module tt_um_brukstus_tdc_with_spi (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire \coarse_result[0] ;
 wire \coarse_result[10] ;
 wire \coarse_result[11] ;
 wire \coarse_result[12] ;
 wire \coarse_result[13] ;
 wire \coarse_result[14] ;
 wire \coarse_result[15] ;
 wire \coarse_result[16] ;
 wire \coarse_result[17] ;
 wire \coarse_result[18] ;
 wire \coarse_result[19] ;
 wire \coarse_result[1] ;
 wire \coarse_result[20] ;
 wire \coarse_result[21] ;
 wire \coarse_result[22] ;
 wire \coarse_result[23] ;
 wire \coarse_result[24] ;
 wire \coarse_result[25] ;
 wire \coarse_result[26] ;
 wire \coarse_result[27] ;
 wire \coarse_result[28] ;
 wire \coarse_result[29] ;
 wire \coarse_result[2] ;
 wire \coarse_result[30] ;
 wire \coarse_result[31] ;
 wire \coarse_result[3] ;
 wire \coarse_result[4] ;
 wire \coarse_result[5] ;
 wire \coarse_result[6] ;
 wire \coarse_result[7] ;
 wire \coarse_result[8] ;
 wire \coarse_result[9] ;
 wire \config_regs[0] ;
 wire \config_regs[10] ;
 wire \config_regs[11] ;
 wire \config_regs[12] ;
 wire \config_regs[13] ;
 wire \config_regs[14] ;
 wire \config_regs[15] ;
 wire \config_regs[16] ;
 wire \config_regs[17] ;
 wire \config_regs[18] ;
 wire \config_regs[19] ;
 wire \config_regs[1] ;
 wire \config_regs[20] ;
 wire \config_regs[21] ;
 wire \config_regs[22] ;
 wire \config_regs[23] ;
 wire \config_regs[24] ;
 wire \config_regs[25] ;
 wire \config_regs[26] ;
 wire \config_regs[27] ;
 wire \config_regs[28] ;
 wire \config_regs[29] ;
 wire \config_regs[2] ;
 wire \config_regs[30] ;
 wire \config_regs[31] ;
 wire \config_regs[32] ;
 wire \config_regs[33] ;
 wire \config_regs[34] ;
 wire \config_regs[35] ;
 wire \config_regs[36] ;
 wire \config_regs[37] ;
 wire \config_regs[38] ;
 wire \config_regs[39] ;
 wire \config_regs[3] ;
 wire \config_regs[40] ;
 wire \config_regs[41] ;
 wire \config_regs[42] ;
 wire \config_regs[43] ;
 wire \config_regs[44] ;
 wire \config_regs[45] ;
 wire \config_regs[46] ;
 wire \config_regs[47] ;
 wire \config_regs[48] ;
 wire \config_regs[49] ;
 wire \config_regs[4] ;
 wire \config_regs[50] ;
 wire \config_regs[51] ;
 wire \config_regs[52] ;
 wire \config_regs[53] ;
 wire \config_regs[54] ;
 wire \config_regs[55] ;
 wire \config_regs[56] ;
 wire \config_regs[57] ;
 wire \config_regs[58] ;
 wire \config_regs[59] ;
 wire \config_regs[5] ;
 wire \config_regs[60] ;
 wire \config_regs[61] ;
 wire \config_regs[62] ;
 wire \config_regs[63] ;
 wire \config_regs[6] ;
 wire \config_regs[7] ;
 wire \config_regs[8] ;
 wire \config_regs[9] ;
 wire cpha_sync;
 wire cpol_sync;
 wire \fine_result[0] ;
 wire \fine_result[1] ;
 wire \fine_result[2] ;
 wire \fine_result[3] ;
 wire \fine_result[4] ;
 wire \fine_result[5] ;
 wire \fine_result[6] ;
 wire \fine_result[7] ;
 wire \fine_result[8] ;
 wire spi_clk_sync;
 wire spi_cs_n_sync;
 wire spi_miso;
 wire spi_mosi_sync;
 wire \spi_wrapper_i.reg_addr[0] ;
 wire \spi_wrapper_i.reg_addr[1] ;
 wire \spi_wrapper_i.reg_addr[2] ;
 wire \spi_wrapper_i.reg_addr[3] ;
 wire \spi_wrapper_i.reg_data_o[0] ;
 wire \spi_wrapper_i.reg_data_o[1] ;
 wire \spi_wrapper_i.reg_data_o[2] ;
 wire \spi_wrapper_i.reg_data_o[3] ;
 wire \spi_wrapper_i.reg_data_o[4] ;
 wire \spi_wrapper_i.reg_data_o[5] ;
 wire \spi_wrapper_i.reg_data_o[6] ;
 wire \spi_wrapper_i.reg_data_o[7] ;
 wire \spi_wrapper_i.reg_data_o_vld ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.reg_rw ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[6] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[7] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ;
 wire \spi_wrapper_i.spi_reg_inst.state[0] ;
 wire \spi_wrapper_i.spi_reg_inst.state[1] ;
 wire \spi_wrapper_i.spi_reg_inst.state[2] ;
 wire \spi_wrapper_i.spi_reg_inst.state[3] ;
 wire \spi_wrapper_i.spi_reg_inst.state[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[6] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ;
 wire \synchronizer_spi_clk_inst.data_sync[1] ;
 wire \synchronizer_spi_cs_n_inst.data_sync[1] ;
 wire \synchronizer_spi_mode_cpha.data_sync[1] ;
 wire \synchronizer_spi_mode_cpol.data_sync[1] ;
 wire \synchronizer_spi_mosi_inst.data_sync[1] ;
 wire \tdc_inst.busy ;
 wire \tdc_inst.coarse_count[0] ;
 wire \tdc_inst.coarse_count[10] ;
 wire \tdc_inst.coarse_count[11] ;
 wire \tdc_inst.coarse_count[12] ;
 wire \tdc_inst.coarse_count[13] ;
 wire \tdc_inst.coarse_count[14] ;
 wire \tdc_inst.coarse_count[15] ;
 wire \tdc_inst.coarse_count[16] ;
 wire \tdc_inst.coarse_count[17] ;
 wire \tdc_inst.coarse_count[18] ;
 wire \tdc_inst.coarse_count[19] ;
 wire \tdc_inst.coarse_count[1] ;
 wire \tdc_inst.coarse_count[20] ;
 wire \tdc_inst.coarse_count[21] ;
 wire \tdc_inst.coarse_count[22] ;
 wire \tdc_inst.coarse_count[23] ;
 wire \tdc_inst.coarse_count[24] ;
 wire \tdc_inst.coarse_count[25] ;
 wire \tdc_inst.coarse_count[26] ;
 wire \tdc_inst.coarse_count[27] ;
 wire \tdc_inst.coarse_count[28] ;
 wire \tdc_inst.coarse_count[29] ;
 wire \tdc_inst.coarse_count[2] ;
 wire \tdc_inst.coarse_count[30] ;
 wire \tdc_inst.coarse_count[31] ;
 wire \tdc_inst.coarse_count[3] ;
 wire \tdc_inst.coarse_count[4] ;
 wire \tdc_inst.coarse_count[5] ;
 wire \tdc_inst.coarse_count[6] ;
 wire \tdc_inst.coarse_count[7] ;
 wire \tdc_inst.coarse_count[8] ;
 wire \tdc_inst.coarse_count[9] ;
 wire \tdc_inst.fine_another_counter[0] ;
 wire \tdc_inst.fine_another_counter[1] ;
 wire \tdc_inst.fine_another_counter[2] ;
 wire \tdc_inst.fine_another_counter[3] ;
 wire \tdc_inst.fine_another_counter[4] ;
 wire \tdc_inst.fine_another_counter[5] ;
 wire \tdc_inst.fine_another_counter[6] ;
 wire \tdc_inst.fine_another_counter[7] ;
 wire \tdc_inst.fine_another_counter[8] ;
 wire \tdc_inst.fine_procedure_counter[0] ;
 wire \tdc_inst.fine_procedure_counter[1] ;
 wire \tdc_inst.fine_procedure_counter[2] ;
 wire \tdc_inst.fine_procedure_counter[3] ;
 wire \tdc_inst.fine_procedure_counter[4] ;
 wire \tdc_inst.fine_procedure_counter[5] ;
 wire \tdc_inst.fine_procedure_counter[6] ;
 wire \tdc_inst.fine_procedure_counter[7] ;
 wire \tdc_inst.fine_procedure_counter[8] ;
 wire \tdc_inst.fine_start_counter[0] ;
 wire \tdc_inst.fine_start_counter[1] ;
 wire \tdc_inst.fine_start_counter[2] ;
 wire \tdc_inst.fine_start_counter[3] ;
 wire \tdc_inst.fine_start_counter[4] ;
 wire \tdc_inst.fine_start_counter[5] ;
 wire \tdc_inst.fine_start_counter[6] ;
 wire \tdc_inst.fine_start_counter[7] ;
 wire \tdc_inst.fine_start_counter[8] ;
 wire \tdc_inst.fine_stop_counter[0] ;
 wire \tdc_inst.fine_stop_counter[1] ;
 wire \tdc_inst.fine_stop_counter[2] ;
 wire \tdc_inst.fine_stop_counter[3] ;
 wire \tdc_inst.fine_stop_counter[4] ;
 wire \tdc_inst.fine_stop_counter[5] ;
 wire \tdc_inst.fine_stop_counter[6] ;
 wire \tdc_inst.fine_stop_counter[7] ;
 wire \tdc_inst.fine_stop_counter[8] ;
 wire \tdc_inst.positions_sum[4] ;
 wire \tdc_inst.positions_sum[5] ;
 wire \tdc_inst.positions_sum[6] ;
 wire \tdc_inst.positions_sum[7] ;
 wire \tdc_inst.positions_sum[8] ;
 wire \tdc_inst.reset_internal_logic ;
 wire \tdc_inst.start_count_debug[0] ;
 wire \tdc_inst.start_count_debug[100] ;
 wire \tdc_inst.start_count_debug[101] ;
 wire \tdc_inst.start_count_debug[102] ;
 wire \tdc_inst.start_count_debug[103] ;
 wire \tdc_inst.start_count_debug[104] ;
 wire \tdc_inst.start_count_debug[105] ;
 wire \tdc_inst.start_count_debug[106] ;
 wire \tdc_inst.start_count_debug[107] ;
 wire \tdc_inst.start_count_debug[108] ;
 wire \tdc_inst.start_count_debug[109] ;
 wire \tdc_inst.start_count_debug[10] ;
 wire \tdc_inst.start_count_debug[110] ;
 wire \tdc_inst.start_count_debug[111] ;
 wire \tdc_inst.start_count_debug[112] ;
 wire \tdc_inst.start_count_debug[113] ;
 wire \tdc_inst.start_count_debug[114] ;
 wire \tdc_inst.start_count_debug[115] ;
 wire \tdc_inst.start_count_debug[116] ;
 wire \tdc_inst.start_count_debug[117] ;
 wire \tdc_inst.start_count_debug[118] ;
 wire \tdc_inst.start_count_debug[119] ;
 wire \tdc_inst.start_count_debug[11] ;
 wire \tdc_inst.start_count_debug[120] ;
 wire \tdc_inst.start_count_debug[121] ;
 wire \tdc_inst.start_count_debug[122] ;
 wire \tdc_inst.start_count_debug[123] ;
 wire \tdc_inst.start_count_debug[124] ;
 wire \tdc_inst.start_count_debug[125] ;
 wire \tdc_inst.start_count_debug[126] ;
 wire \tdc_inst.start_count_debug[127] ;
 wire \tdc_inst.start_count_debug[128] ;
 wire \tdc_inst.start_count_debug[129] ;
 wire \tdc_inst.start_count_debug[12] ;
 wire \tdc_inst.start_count_debug[130] ;
 wire \tdc_inst.start_count_debug[131] ;
 wire \tdc_inst.start_count_debug[132] ;
 wire \tdc_inst.start_count_debug[133] ;
 wire \tdc_inst.start_count_debug[134] ;
 wire \tdc_inst.start_count_debug[135] ;
 wire \tdc_inst.start_count_debug[136] ;
 wire \tdc_inst.start_count_debug[137] ;
 wire \tdc_inst.start_count_debug[138] ;
 wire \tdc_inst.start_count_debug[139] ;
 wire \tdc_inst.start_count_debug[13] ;
 wire \tdc_inst.start_count_debug[140] ;
 wire \tdc_inst.start_count_debug[141] ;
 wire \tdc_inst.start_count_debug[142] ;
 wire \tdc_inst.start_count_debug[14] ;
 wire \tdc_inst.start_count_debug[15] ;
 wire \tdc_inst.start_count_debug[16] ;
 wire \tdc_inst.start_count_debug[17] ;
 wire \tdc_inst.start_count_debug[18] ;
 wire \tdc_inst.start_count_debug[19] ;
 wire \tdc_inst.start_count_debug[1] ;
 wire \tdc_inst.start_count_debug[20] ;
 wire \tdc_inst.start_count_debug[21] ;
 wire \tdc_inst.start_count_debug[22] ;
 wire \tdc_inst.start_count_debug[23] ;
 wire \tdc_inst.start_count_debug[24] ;
 wire \tdc_inst.start_count_debug[25] ;
 wire \tdc_inst.start_count_debug[26] ;
 wire \tdc_inst.start_count_debug[27] ;
 wire \tdc_inst.start_count_debug[28] ;
 wire \tdc_inst.start_count_debug[29] ;
 wire \tdc_inst.start_count_debug[2] ;
 wire \tdc_inst.start_count_debug[30] ;
 wire \tdc_inst.start_count_debug[31] ;
 wire \tdc_inst.start_count_debug[32] ;
 wire \tdc_inst.start_count_debug[33] ;
 wire \tdc_inst.start_count_debug[34] ;
 wire \tdc_inst.start_count_debug[35] ;
 wire \tdc_inst.start_count_debug[36] ;
 wire \tdc_inst.start_count_debug[37] ;
 wire \tdc_inst.start_count_debug[38] ;
 wire \tdc_inst.start_count_debug[39] ;
 wire \tdc_inst.start_count_debug[3] ;
 wire \tdc_inst.start_count_debug[40] ;
 wire \tdc_inst.start_count_debug[41] ;
 wire \tdc_inst.start_count_debug[42] ;
 wire \tdc_inst.start_count_debug[43] ;
 wire \tdc_inst.start_count_debug[44] ;
 wire \tdc_inst.start_count_debug[45] ;
 wire \tdc_inst.start_count_debug[46] ;
 wire \tdc_inst.start_count_debug[47] ;
 wire \tdc_inst.start_count_debug[48] ;
 wire \tdc_inst.start_count_debug[49] ;
 wire \tdc_inst.start_count_debug[4] ;
 wire \tdc_inst.start_count_debug[50] ;
 wire \tdc_inst.start_count_debug[51] ;
 wire \tdc_inst.start_count_debug[52] ;
 wire \tdc_inst.start_count_debug[53] ;
 wire \tdc_inst.start_count_debug[54] ;
 wire \tdc_inst.start_count_debug[55] ;
 wire \tdc_inst.start_count_debug[56] ;
 wire \tdc_inst.start_count_debug[57] ;
 wire \tdc_inst.start_count_debug[58] ;
 wire \tdc_inst.start_count_debug[59] ;
 wire \tdc_inst.start_count_debug[5] ;
 wire \tdc_inst.start_count_debug[60] ;
 wire \tdc_inst.start_count_debug[61] ;
 wire \tdc_inst.start_count_debug[62] ;
 wire \tdc_inst.start_count_debug[63] ;
 wire \tdc_inst.start_count_debug[64] ;
 wire \tdc_inst.start_count_debug[65] ;
 wire \tdc_inst.start_count_debug[66] ;
 wire \tdc_inst.start_count_debug[67] ;
 wire \tdc_inst.start_count_debug[68] ;
 wire \tdc_inst.start_count_debug[69] ;
 wire \tdc_inst.start_count_debug[6] ;
 wire \tdc_inst.start_count_debug[70] ;
 wire \tdc_inst.start_count_debug[71] ;
 wire \tdc_inst.start_count_debug[72] ;
 wire \tdc_inst.start_count_debug[73] ;
 wire \tdc_inst.start_count_debug[74] ;
 wire \tdc_inst.start_count_debug[75] ;
 wire \tdc_inst.start_count_debug[76] ;
 wire \tdc_inst.start_count_debug[77] ;
 wire \tdc_inst.start_count_debug[78] ;
 wire \tdc_inst.start_count_debug[79] ;
 wire \tdc_inst.start_count_debug[7] ;
 wire \tdc_inst.start_count_debug[80] ;
 wire \tdc_inst.start_count_debug[81] ;
 wire \tdc_inst.start_count_debug[82] ;
 wire \tdc_inst.start_count_debug[83] ;
 wire \tdc_inst.start_count_debug[84] ;
 wire \tdc_inst.start_count_debug[85] ;
 wire \tdc_inst.start_count_debug[86] ;
 wire \tdc_inst.start_count_debug[87] ;
 wire \tdc_inst.start_count_debug[88] ;
 wire \tdc_inst.start_count_debug[89] ;
 wire \tdc_inst.start_count_debug[8] ;
 wire \tdc_inst.start_count_debug[90] ;
 wire \tdc_inst.start_count_debug[91] ;
 wire \tdc_inst.start_count_debug[92] ;
 wire \tdc_inst.start_count_debug[93] ;
 wire \tdc_inst.start_count_debug[94] ;
 wire \tdc_inst.start_count_debug[95] ;
 wire \tdc_inst.start_count_debug[96] ;
 wire \tdc_inst.start_count_debug[97] ;
 wire \tdc_inst.start_count_debug[98] ;
 wire \tdc_inst.start_count_debug[99] ;
 wire \tdc_inst.start_count_debug[9] ;
 wire \tdc_inst.start_signal_activated ;
 wire \tdc_inst.start_signal_sampling_clock_level ;
 wire \tdc_inst.stop_count_debug[0] ;
 wire \tdc_inst.stop_count_debug[100] ;
 wire \tdc_inst.stop_count_debug[101] ;
 wire \tdc_inst.stop_count_debug[102] ;
 wire \tdc_inst.stop_count_debug[103] ;
 wire \tdc_inst.stop_count_debug[104] ;
 wire \tdc_inst.stop_count_debug[105] ;
 wire \tdc_inst.stop_count_debug[106] ;
 wire \tdc_inst.stop_count_debug[107] ;
 wire \tdc_inst.stop_count_debug[108] ;
 wire \tdc_inst.stop_count_debug[109] ;
 wire \tdc_inst.stop_count_debug[10] ;
 wire \tdc_inst.stop_count_debug[110] ;
 wire \tdc_inst.stop_count_debug[111] ;
 wire \tdc_inst.stop_count_debug[112] ;
 wire \tdc_inst.stop_count_debug[113] ;
 wire \tdc_inst.stop_count_debug[114] ;
 wire \tdc_inst.stop_count_debug[115] ;
 wire \tdc_inst.stop_count_debug[116] ;
 wire \tdc_inst.stop_count_debug[117] ;
 wire \tdc_inst.stop_count_debug[118] ;
 wire \tdc_inst.stop_count_debug[119] ;
 wire \tdc_inst.stop_count_debug[11] ;
 wire \tdc_inst.stop_count_debug[120] ;
 wire \tdc_inst.stop_count_debug[121] ;
 wire \tdc_inst.stop_count_debug[122] ;
 wire \tdc_inst.stop_count_debug[123] ;
 wire \tdc_inst.stop_count_debug[124] ;
 wire \tdc_inst.stop_count_debug[125] ;
 wire \tdc_inst.stop_count_debug[126] ;
 wire \tdc_inst.stop_count_debug[127] ;
 wire \tdc_inst.stop_count_debug[128] ;
 wire \tdc_inst.stop_count_debug[129] ;
 wire \tdc_inst.stop_count_debug[12] ;
 wire \tdc_inst.stop_count_debug[130] ;
 wire \tdc_inst.stop_count_debug[131] ;
 wire \tdc_inst.stop_count_debug[132] ;
 wire \tdc_inst.stop_count_debug[133] ;
 wire \tdc_inst.stop_count_debug[134] ;
 wire \tdc_inst.stop_count_debug[135] ;
 wire \tdc_inst.stop_count_debug[136] ;
 wire \tdc_inst.stop_count_debug[137] ;
 wire \tdc_inst.stop_count_debug[138] ;
 wire \tdc_inst.stop_count_debug[139] ;
 wire \tdc_inst.stop_count_debug[13] ;
 wire \tdc_inst.stop_count_debug[140] ;
 wire \tdc_inst.stop_count_debug[141] ;
 wire \tdc_inst.stop_count_debug[142] ;
 wire \tdc_inst.stop_count_debug[14] ;
 wire \tdc_inst.stop_count_debug[15] ;
 wire \tdc_inst.stop_count_debug[16] ;
 wire \tdc_inst.stop_count_debug[17] ;
 wire \tdc_inst.stop_count_debug[18] ;
 wire \tdc_inst.stop_count_debug[19] ;
 wire \tdc_inst.stop_count_debug[1] ;
 wire \tdc_inst.stop_count_debug[20] ;
 wire \tdc_inst.stop_count_debug[21] ;
 wire \tdc_inst.stop_count_debug[22] ;
 wire \tdc_inst.stop_count_debug[23] ;
 wire \tdc_inst.stop_count_debug[24] ;
 wire \tdc_inst.stop_count_debug[25] ;
 wire \tdc_inst.stop_count_debug[26] ;
 wire \tdc_inst.stop_count_debug[27] ;
 wire \tdc_inst.stop_count_debug[28] ;
 wire \tdc_inst.stop_count_debug[29] ;
 wire \tdc_inst.stop_count_debug[2] ;
 wire \tdc_inst.stop_count_debug[30] ;
 wire \tdc_inst.stop_count_debug[31] ;
 wire \tdc_inst.stop_count_debug[32] ;
 wire \tdc_inst.stop_count_debug[33] ;
 wire \tdc_inst.stop_count_debug[34] ;
 wire \tdc_inst.stop_count_debug[35] ;
 wire \tdc_inst.stop_count_debug[36] ;
 wire \tdc_inst.stop_count_debug[37] ;
 wire \tdc_inst.stop_count_debug[38] ;
 wire \tdc_inst.stop_count_debug[39] ;
 wire \tdc_inst.stop_count_debug[3] ;
 wire \tdc_inst.stop_count_debug[40] ;
 wire \tdc_inst.stop_count_debug[41] ;
 wire \tdc_inst.stop_count_debug[42] ;
 wire \tdc_inst.stop_count_debug[43] ;
 wire \tdc_inst.stop_count_debug[44] ;
 wire \tdc_inst.stop_count_debug[45] ;
 wire \tdc_inst.stop_count_debug[46] ;
 wire \tdc_inst.stop_count_debug[47] ;
 wire \tdc_inst.stop_count_debug[48] ;
 wire \tdc_inst.stop_count_debug[49] ;
 wire \tdc_inst.stop_count_debug[4] ;
 wire \tdc_inst.stop_count_debug[50] ;
 wire \tdc_inst.stop_count_debug[51] ;
 wire \tdc_inst.stop_count_debug[52] ;
 wire \tdc_inst.stop_count_debug[53] ;
 wire \tdc_inst.stop_count_debug[54] ;
 wire \tdc_inst.stop_count_debug[55] ;
 wire \tdc_inst.stop_count_debug[56] ;
 wire \tdc_inst.stop_count_debug[57] ;
 wire \tdc_inst.stop_count_debug[58] ;
 wire \tdc_inst.stop_count_debug[59] ;
 wire \tdc_inst.stop_count_debug[5] ;
 wire \tdc_inst.stop_count_debug[60] ;
 wire \tdc_inst.stop_count_debug[61] ;
 wire \tdc_inst.stop_count_debug[62] ;
 wire \tdc_inst.stop_count_debug[63] ;
 wire \tdc_inst.stop_count_debug[64] ;
 wire \tdc_inst.stop_count_debug[65] ;
 wire \tdc_inst.stop_count_debug[66] ;
 wire \tdc_inst.stop_count_debug[67] ;
 wire \tdc_inst.stop_count_debug[68] ;
 wire \tdc_inst.stop_count_debug[69] ;
 wire \tdc_inst.stop_count_debug[6] ;
 wire \tdc_inst.stop_count_debug[70] ;
 wire \tdc_inst.stop_count_debug[71] ;
 wire \tdc_inst.stop_count_debug[72] ;
 wire \tdc_inst.stop_count_debug[73] ;
 wire \tdc_inst.stop_count_debug[74] ;
 wire \tdc_inst.stop_count_debug[75] ;
 wire \tdc_inst.stop_count_debug[76] ;
 wire \tdc_inst.stop_count_debug[77] ;
 wire \tdc_inst.stop_count_debug[78] ;
 wire \tdc_inst.stop_count_debug[79] ;
 wire \tdc_inst.stop_count_debug[7] ;
 wire \tdc_inst.stop_count_debug[80] ;
 wire \tdc_inst.stop_count_debug[81] ;
 wire \tdc_inst.stop_count_debug[82] ;
 wire \tdc_inst.stop_count_debug[83] ;
 wire \tdc_inst.stop_count_debug[84] ;
 wire \tdc_inst.stop_count_debug[85] ;
 wire \tdc_inst.stop_count_debug[86] ;
 wire \tdc_inst.stop_count_debug[87] ;
 wire \tdc_inst.stop_count_debug[88] ;
 wire \tdc_inst.stop_count_debug[89] ;
 wire \tdc_inst.stop_count_debug[8] ;
 wire \tdc_inst.stop_count_debug[90] ;
 wire \tdc_inst.stop_count_debug[91] ;
 wire \tdc_inst.stop_count_debug[92] ;
 wire \tdc_inst.stop_count_debug[93] ;
 wire \tdc_inst.stop_count_debug[94] ;
 wire \tdc_inst.stop_count_debug[95] ;
 wire \tdc_inst.stop_count_debug[96] ;
 wire \tdc_inst.stop_count_debug[97] ;
 wire \tdc_inst.stop_count_debug[98] ;
 wire \tdc_inst.stop_count_debug[99] ;
 wire \tdc_inst.stop_count_debug[9] ;
 wire \tdc_inst.stop_signal_activated ;
 wire \tdc_inst.stop_signal_sampling_clock_level ;
 wire \tdc_inst.tdc_xor_result[0] ;
 wire \tdc_inst.tdc_xor_result[100] ;
 wire \tdc_inst.tdc_xor_result[101] ;
 wire \tdc_inst.tdc_xor_result[102] ;
 wire \tdc_inst.tdc_xor_result[103] ;
 wire \tdc_inst.tdc_xor_result[104] ;
 wire \tdc_inst.tdc_xor_result[105] ;
 wire \tdc_inst.tdc_xor_result[106] ;
 wire \tdc_inst.tdc_xor_result[107] ;
 wire \tdc_inst.tdc_xor_result[108] ;
 wire \tdc_inst.tdc_xor_result[109] ;
 wire \tdc_inst.tdc_xor_result[10] ;
 wire \tdc_inst.tdc_xor_result[110] ;
 wire \tdc_inst.tdc_xor_result[111] ;
 wire \tdc_inst.tdc_xor_result[112] ;
 wire \tdc_inst.tdc_xor_result[113] ;
 wire \tdc_inst.tdc_xor_result[114] ;
 wire \tdc_inst.tdc_xor_result[115] ;
 wire \tdc_inst.tdc_xor_result[116] ;
 wire \tdc_inst.tdc_xor_result[117] ;
 wire \tdc_inst.tdc_xor_result[118] ;
 wire \tdc_inst.tdc_xor_result[119] ;
 wire \tdc_inst.tdc_xor_result[11] ;
 wire \tdc_inst.tdc_xor_result[120] ;
 wire \tdc_inst.tdc_xor_result[121] ;
 wire \tdc_inst.tdc_xor_result[122] ;
 wire \tdc_inst.tdc_xor_result[123] ;
 wire \tdc_inst.tdc_xor_result[124] ;
 wire \tdc_inst.tdc_xor_result[125] ;
 wire \tdc_inst.tdc_xor_result[126] ;
 wire \tdc_inst.tdc_xor_result[127] ;
 wire \tdc_inst.tdc_xor_result[128] ;
 wire \tdc_inst.tdc_xor_result[129] ;
 wire \tdc_inst.tdc_xor_result[12] ;
 wire \tdc_inst.tdc_xor_result[130] ;
 wire \tdc_inst.tdc_xor_result[131] ;
 wire \tdc_inst.tdc_xor_result[132] ;
 wire \tdc_inst.tdc_xor_result[133] ;
 wire \tdc_inst.tdc_xor_result[134] ;
 wire \tdc_inst.tdc_xor_result[135] ;
 wire \tdc_inst.tdc_xor_result[136] ;
 wire \tdc_inst.tdc_xor_result[137] ;
 wire \tdc_inst.tdc_xor_result[138] ;
 wire \tdc_inst.tdc_xor_result[139] ;
 wire \tdc_inst.tdc_xor_result[13] ;
 wire \tdc_inst.tdc_xor_result[140] ;
 wire \tdc_inst.tdc_xor_result[141] ;
 wire \tdc_inst.tdc_xor_result[142] ;
 wire \tdc_inst.tdc_xor_result[14] ;
 wire \tdc_inst.tdc_xor_result[15] ;
 wire \tdc_inst.tdc_xor_result[16] ;
 wire \tdc_inst.tdc_xor_result[17] ;
 wire \tdc_inst.tdc_xor_result[18] ;
 wire \tdc_inst.tdc_xor_result[19] ;
 wire \tdc_inst.tdc_xor_result[1] ;
 wire \tdc_inst.tdc_xor_result[20] ;
 wire \tdc_inst.tdc_xor_result[21] ;
 wire \tdc_inst.tdc_xor_result[22] ;
 wire \tdc_inst.tdc_xor_result[23] ;
 wire \tdc_inst.tdc_xor_result[24] ;
 wire \tdc_inst.tdc_xor_result[25] ;
 wire \tdc_inst.tdc_xor_result[26] ;
 wire \tdc_inst.tdc_xor_result[27] ;
 wire \tdc_inst.tdc_xor_result[28] ;
 wire \tdc_inst.tdc_xor_result[29] ;
 wire \tdc_inst.tdc_xor_result[2] ;
 wire \tdc_inst.tdc_xor_result[30] ;
 wire \tdc_inst.tdc_xor_result[31] ;
 wire \tdc_inst.tdc_xor_result[32] ;
 wire \tdc_inst.tdc_xor_result[33] ;
 wire \tdc_inst.tdc_xor_result[34] ;
 wire \tdc_inst.tdc_xor_result[35] ;
 wire \tdc_inst.tdc_xor_result[36] ;
 wire \tdc_inst.tdc_xor_result[37] ;
 wire \tdc_inst.tdc_xor_result[38] ;
 wire \tdc_inst.tdc_xor_result[39] ;
 wire \tdc_inst.tdc_xor_result[3] ;
 wire \tdc_inst.tdc_xor_result[40] ;
 wire \tdc_inst.tdc_xor_result[41] ;
 wire \tdc_inst.tdc_xor_result[42] ;
 wire \tdc_inst.tdc_xor_result[43] ;
 wire \tdc_inst.tdc_xor_result[44] ;
 wire \tdc_inst.tdc_xor_result[45] ;
 wire \tdc_inst.tdc_xor_result[46] ;
 wire \tdc_inst.tdc_xor_result[47] ;
 wire \tdc_inst.tdc_xor_result[48] ;
 wire \tdc_inst.tdc_xor_result[49] ;
 wire \tdc_inst.tdc_xor_result[4] ;
 wire \tdc_inst.tdc_xor_result[50] ;
 wire \tdc_inst.tdc_xor_result[51] ;
 wire \tdc_inst.tdc_xor_result[52] ;
 wire \tdc_inst.tdc_xor_result[53] ;
 wire \tdc_inst.tdc_xor_result[54] ;
 wire \tdc_inst.tdc_xor_result[55] ;
 wire \tdc_inst.tdc_xor_result[56] ;
 wire \tdc_inst.tdc_xor_result[57] ;
 wire \tdc_inst.tdc_xor_result[58] ;
 wire \tdc_inst.tdc_xor_result[59] ;
 wire \tdc_inst.tdc_xor_result[5] ;
 wire \tdc_inst.tdc_xor_result[60] ;
 wire \tdc_inst.tdc_xor_result[61] ;
 wire \tdc_inst.tdc_xor_result[62] ;
 wire \tdc_inst.tdc_xor_result[63] ;
 wire \tdc_inst.tdc_xor_result[64] ;
 wire \tdc_inst.tdc_xor_result[65] ;
 wire \tdc_inst.tdc_xor_result[66] ;
 wire \tdc_inst.tdc_xor_result[67] ;
 wire \tdc_inst.tdc_xor_result[68] ;
 wire \tdc_inst.tdc_xor_result[69] ;
 wire \tdc_inst.tdc_xor_result[6] ;
 wire \tdc_inst.tdc_xor_result[70] ;
 wire \tdc_inst.tdc_xor_result[71] ;
 wire \tdc_inst.tdc_xor_result[72] ;
 wire \tdc_inst.tdc_xor_result[73] ;
 wire \tdc_inst.tdc_xor_result[74] ;
 wire \tdc_inst.tdc_xor_result[75] ;
 wire \tdc_inst.tdc_xor_result[76] ;
 wire \tdc_inst.tdc_xor_result[77] ;
 wire \tdc_inst.tdc_xor_result[78] ;
 wire \tdc_inst.tdc_xor_result[79] ;
 wire \tdc_inst.tdc_xor_result[7] ;
 wire \tdc_inst.tdc_xor_result[80] ;
 wire \tdc_inst.tdc_xor_result[81] ;
 wire \tdc_inst.tdc_xor_result[82] ;
 wire \tdc_inst.tdc_xor_result[83] ;
 wire \tdc_inst.tdc_xor_result[84] ;
 wire \tdc_inst.tdc_xor_result[85] ;
 wire \tdc_inst.tdc_xor_result[86] ;
 wire \tdc_inst.tdc_xor_result[87] ;
 wire \tdc_inst.tdc_xor_result[88] ;
 wire \tdc_inst.tdc_xor_result[89] ;
 wire \tdc_inst.tdc_xor_result[8] ;
 wire \tdc_inst.tdc_xor_result[90] ;
 wire \tdc_inst.tdc_xor_result[91] ;
 wire \tdc_inst.tdc_xor_result[92] ;
 wire \tdc_inst.tdc_xor_result[93] ;
 wire \tdc_inst.tdc_xor_result[94] ;
 wire \tdc_inst.tdc_xor_result[95] ;
 wire \tdc_inst.tdc_xor_result[96] ;
 wire \tdc_inst.tdc_xor_result[97] ;
 wire \tdc_inst.tdc_xor_result[98] ;
 wire \tdc_inst.tdc_xor_result[99] ;
 wire \tdc_inst.tdc_xor_result[9] ;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_leaf_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;

 sg13g2_a22oi_1 _2770_ (.Y(_1422_),
    .B1(net958),
    .B2(net644),
    .A2(net961),
    .A1(\tdc_inst.coarse_count[25] ));
 sg13g2_inv_1 _2771_ (.Y(_0620_),
    .A(_1422_));
 sg13g2_nor2b_1 _2772_ (.A(_0042_),
    .B_N(_1392_),
    .Y(_1423_));
 sg13g2_o21ai_1 _2773_ (.B1(net961),
    .Y(_1424_),
    .A1(\tdc_inst.coarse_count[26] ),
    .A2(_1423_));
 sg13g2_o21ai_1 _2774_ (.B1(_1424_),
    .Y(_0621_),
    .A1(_0716_),
    .A2(_1380_));
 sg13g2_a22oi_1 _2775_ (.Y(_1425_),
    .B1(net958),
    .B2(net567),
    .A2(net964),
    .A1(\tdc_inst.coarse_count[27] ));
 sg13g2_inv_1 _2776_ (.Y(_0622_),
    .A(_1425_));
 sg13g2_a22oi_1 _2777_ (.Y(_1426_),
    .B1(net958),
    .B2(net586),
    .A2(net960),
    .A1(\tdc_inst.coarse_count[28] ));
 sg13g2_inv_1 _2778_ (.Y(_0623_),
    .A(_1426_));
 sg13g2_a22oi_1 _2779_ (.Y(_1427_),
    .B1(net958),
    .B2(net881),
    .A2(net960),
    .A1(\tdc_inst.coarse_count[29] ));
 sg13g2_inv_1 _2780_ (.Y(_0624_),
    .A(_1427_));
 sg13g2_nor2b_1 _2781_ (.A(_0043_),
    .B_N(_1392_),
    .Y(_1428_));
 sg13g2_o21ai_1 _2782_ (.B1(net960),
    .Y(_1429_),
    .A1(\tdc_inst.coarse_count[30] ),
    .A2(_1428_));
 sg13g2_o21ai_1 _2783_ (.B1(_1429_),
    .Y(_0625_),
    .A1(_0715_),
    .A2(_1380_));
 sg13g2_a22oi_1 _2784_ (.Y(_1430_),
    .B1(net958),
    .B2(net573),
    .A2(net960),
    .A1(\tdc_inst.coarse_count[31] ));
 sg13g2_inv_1 _2785_ (.Y(_0626_),
    .A(_1430_));
 sg13g2_mux2_1 _2786_ (.A0(\tdc_inst.start_signal_sampling_clock_level ),
    .A1(net1235),
    .S(net1215),
    .X(_0627_));
 sg13g2_a21o_1 _2787_ (.A2(net1159),
    .A1(net1339),
    .B1(_0919_),
    .X(_0628_));
 sg13g2_a21o_1 _2788_ (.A2(net1158),
    .A1(net1377),
    .B1(_0774_),
    .X(_0629_));
 sg13g2_a21o_1 _2789_ (.A2(net1158),
    .A1(net1318),
    .B1(_1063_),
    .X(_0630_));
 sg13g2_a21oi_1 _2790_ (.A1(net1209),
    .A2(_1366_),
    .Y(_1431_),
    .B1(net1749));
 sg13g2_and2_1 _2791_ (.A(net1209),
    .B(net1749),
    .X(_1432_));
 sg13g2_nor3_1 _2792_ (.A(net1228),
    .B(net1750),
    .C(_1432_),
    .Y(_0631_));
 sg13g2_and2_1 _2793_ (.A(net1787),
    .B(_1432_),
    .X(_1433_));
 sg13g2_o21ai_1 _2794_ (.B1(_1379_),
    .Y(_1434_),
    .A1(net1787),
    .A2(_1432_));
 sg13g2_nor2_1 _2795_ (.A(_1433_),
    .B(_1434_),
    .Y(_0632_));
 sg13g2_and2_1 _2796_ (.A(net1772),
    .B(_1433_),
    .X(_1435_));
 sg13g2_nor2_1 _2797_ (.A(net1772),
    .B(_1433_),
    .Y(_1436_));
 sg13g2_nor3_1 _2798_ (.A(_1380_),
    .B(_1435_),
    .C(net1773),
    .Y(_0633_));
 sg13g2_nor2_1 _2799_ (.A(net1770),
    .B(_1435_),
    .Y(_1437_));
 sg13g2_and2_1 _2800_ (.A(net1770),
    .B(_1435_),
    .X(_1438_));
 sg13g2_nor3_1 _2801_ (.A(_1380_),
    .B(net1771),
    .C(_1438_),
    .Y(_0634_));
 sg13g2_and2_2 _2802_ (.A(net1210),
    .B(_1369_),
    .X(_1439_));
 sg13g2_nand4_1 _2803_ (.B(\tdc_inst.fine_procedure_counter[2] ),
    .C(\tdc_inst.fine_procedure_counter[1] ),
    .A(\tdc_inst.fine_procedure_counter[3] ),
    .Y(_1440_),
    .D(net1749));
 sg13g2_xor2_1 _2804_ (.B(_1440_),
    .A(net1755),
    .X(_1441_));
 sg13g2_a22oi_1 _2805_ (.Y(_1442_),
    .B1(_1439_),
    .B2(net1756),
    .A2(\tdc_inst.fine_procedure_counter[4] ),
    .A1(_0712_));
 sg13g2_nor2_1 _2806_ (.A(net1228),
    .B(net1757),
    .Y(_0635_));
 sg13g2_nand3_1 _2807_ (.B(\tdc_inst.fine_procedure_counter[4] ),
    .C(_1438_),
    .A(net1801),
    .Y(_1443_));
 sg13g2_a21o_1 _2808_ (.A2(_1438_),
    .A1(\tdc_inst.fine_procedure_counter[4] ),
    .B1(net1801),
    .X(_1444_));
 sg13g2_and3_1 _2809_ (.X(_0636_),
    .A(_1379_),
    .B(_1443_),
    .C(net1802));
 sg13g2_o21ai_1 _2810_ (.B1(net959),
    .Y(_1445_),
    .A1(_0714_),
    .A2(_1443_));
 sg13g2_a21oi_1 _2811_ (.A1(_0714_),
    .A2(_1443_),
    .Y(_0637_),
    .B1(_1445_));
 sg13g2_o21ai_1 _2812_ (.B1(_0713_),
    .Y(_1446_),
    .A1(_0714_),
    .A2(_1443_));
 sg13g2_and2_1 _2813_ (.A(net959),
    .B(net1800),
    .X(_0638_));
 sg13g2_a22oi_1 _2814_ (.Y(_1447_),
    .B1(_0728_),
    .B2(_1439_),
    .A2(\tdc_inst.fine_procedure_counter[8] ),
    .A1(net1208));
 sg13g2_nor2_1 _2815_ (.A(_0729_),
    .B(net597),
    .Y(_0639_));
 sg13g2_nand2_1 _2816_ (.Y(_1448_),
    .A(\tdc_inst.fine_another_counter[0] ),
    .B(net1766));
 sg13g2_nand2_1 _2817_ (.Y(_1449_),
    .A(_0032_),
    .B(_1448_));
 sg13g2_nand3b_1 _2818_ (.B(\tdc_inst.tdc_xor_result[0] ),
    .C(\tdc_inst.fine_another_counter[0] ),
    .Y(_1450_),
    .A_N(_0032_));
 sg13g2_nand3_1 _2819_ (.B(_1449_),
    .C(_1450_),
    .A(net1119),
    .Y(_1451_));
 sg13g2_or3_1 _2820_ (.A(\tdc_inst.positions_sum[6] ),
    .B(\tdc_inst.positions_sum[5] ),
    .C(\tdc_inst.positions_sum[4] ),
    .X(_1452_));
 sg13g2_a21oi_2 _2821_ (.B1(\tdc_inst.positions_sum[8] ),
    .Y(_1453_),
    .A2(_1452_),
    .A1(\tdc_inst.positions_sum[7] ));
 sg13g2_nand3b_1 _2822_ (.B(_0768_),
    .C(_0918_),
    .Y(_1454_),
    .A_N(\tdc_inst.fine_procedure_counter[8] ));
 sg13g2_nor3_2 _2823_ (.A(_1368_),
    .B(_1453_),
    .C(_1454_),
    .Y(_1455_));
 sg13g2_and2_1 _2824_ (.A(net1209),
    .B(_1455_),
    .X(_1456_));
 sg13g2_nand2_1 _2825_ (.Y(_1457_),
    .A(net1209),
    .B(_1455_));
 sg13g2_or3_2 _2826_ (.A(_1368_),
    .B(_1453_),
    .C(_1454_),
    .X(_1458_));
 sg13g2_nand2_1 _2827_ (.Y(_1459_),
    .A(_1451_),
    .B(_1457_));
 sg13g2_or2_1 _2828_ (.X(_1460_),
    .B(\tdc_inst.fine_another_counter[1] ),
    .A(\tdc_inst.fine_another_counter[0] ));
 sg13g2_nand2_2 _2829_ (.Y(_1461_),
    .A(\tdc_inst.fine_another_counter[0] ),
    .B(\tdc_inst.fine_another_counter[1] ));
 sg13g2_nand3_1 _2830_ (.B(_1460_),
    .C(_1461_),
    .A(_1455_),
    .Y(_1462_));
 sg13g2_a22oi_1 _2831_ (.Y(_1463_),
    .B1(_1459_),
    .B2(_1462_),
    .A2(net1778),
    .A1(net1208));
 sg13g2_nor2_1 _2832_ (.A(net1229),
    .B(net1779),
    .Y(_0640_));
 sg13g2_nor2_1 _2833_ (.A(_0033_),
    .B(_1450_),
    .Y(_1464_));
 sg13g2_xor2_1 _2834_ (.B(_1450_),
    .A(_0033_),
    .X(_1465_));
 sg13g2_a21oi_1 _2835_ (.A1(net1119),
    .A2(_1465_),
    .Y(_1466_),
    .B1(_1456_));
 sg13g2_nor2_1 _2836_ (.A(_0033_),
    .B(_1461_),
    .Y(_1467_));
 sg13g2_nand2b_1 _2837_ (.Y(_1468_),
    .B(_1455_),
    .A_N(_1467_));
 sg13g2_a21oi_1 _2838_ (.A1(_0033_),
    .A2(_1461_),
    .Y(_1469_),
    .B1(_1468_));
 sg13g2_nor2_1 _2839_ (.A(_1466_),
    .B(_1469_),
    .Y(_1470_));
 sg13g2_a21oi_1 _2840_ (.A1(net1208),
    .A2(net1764),
    .Y(_1471_),
    .B1(_1470_));
 sg13g2_nor2_1 _2841_ (.A(net1229),
    .B(net1765),
    .Y(_0641_));
 sg13g2_nand2_2 _2842_ (.Y(_1472_),
    .A(net1209),
    .B(_1458_));
 sg13g2_inv_1 _2843_ (.Y(_1473_),
    .A(_1472_));
 sg13g2_nand2_2 _2844_ (.Y(_1474_),
    .A(net1119),
    .B(_1458_));
 sg13g2_nor2_1 _2845_ (.A(_1464_),
    .B(_1474_),
    .Y(_1475_));
 sg13g2_a21oi_1 _2846_ (.A1(_1456_),
    .A2(_1467_),
    .Y(_1476_),
    .B1(_1475_));
 sg13g2_nand3_1 _2847_ (.B(_1458_),
    .C(_1464_),
    .A(net1119),
    .Y(_1477_));
 sg13g2_o21ai_1 _2848_ (.B1(_1477_),
    .Y(_1478_),
    .A1(_1457_),
    .A2(_1467_));
 sg13g2_a22oi_1 _2849_ (.Y(_1479_),
    .B1(net1725),
    .B2(_1478_),
    .A2(\tdc_inst.fine_another_counter[3] ),
    .A1(net1208));
 sg13g2_o21ai_1 _2850_ (.B1(_1479_),
    .Y(_1480_),
    .A1(net1725),
    .A2(_1476_));
 sg13g2_and2_1 _2851_ (.A(net1237),
    .B(net1726),
    .X(_0642_));
 sg13g2_nand2_1 _2852_ (.Y(_1481_),
    .A(\tdc_inst.fine_another_counter[3] ),
    .B(\tdc_inst.fine_another_counter[2] ));
 sg13g2_nor2_1 _2853_ (.A(_1450_),
    .B(_1481_),
    .Y(_1482_));
 sg13g2_xor2_1 _2854_ (.B(_1482_),
    .A(_0035_),
    .X(_1483_));
 sg13g2_nor2_1 _2855_ (.A(_1474_),
    .B(_1483_),
    .Y(_1484_));
 sg13g2_nor2_1 _2856_ (.A(_1461_),
    .B(_1481_),
    .Y(_1485_));
 sg13g2_xor2_1 _2857_ (.B(_1485_),
    .A(_0035_),
    .X(_1486_));
 sg13g2_a221oi_1 _2858_ (.B2(_1486_),
    .C1(_1484_),
    .B1(_1456_),
    .A1(net1208),
    .Y(_1487_),
    .A2(net1807));
 sg13g2_nor2_1 _2859_ (.A(net1229),
    .B(net1808),
    .Y(_0643_));
 sg13g2_nor4_1 _2860_ (.A(net1208),
    .B(_0035_),
    .C(_1461_),
    .D(_1481_),
    .Y(_1488_));
 sg13g2_xor2_1 _2861_ (.B(_1488_),
    .A(net1805),
    .X(_1489_));
 sg13g2_nand3_1 _2862_ (.B(\tdc_inst.fine_another_counter[4] ),
    .C(_1482_),
    .A(\tdc_inst.fine_another_counter[5] ),
    .Y(_1490_));
 sg13g2_inv_1 _2863_ (.Y(_1491_),
    .A(_1490_));
 sg13g2_a21oi_1 _2864_ (.A1(\tdc_inst.fine_another_counter[4] ),
    .A2(_1482_),
    .Y(_1492_),
    .B1(net1805));
 sg13g2_nor3_1 _2865_ (.A(_1474_),
    .B(_1491_),
    .C(net1806),
    .Y(_1493_));
 sg13g2_a21oi_1 _2866_ (.A1(_1472_),
    .A2(_1489_),
    .Y(_1494_),
    .B1(_1493_));
 sg13g2_nor2_1 _2867_ (.A(net1229),
    .B(_1494_),
    .Y(_0644_));
 sg13g2_a21o_1 _2868_ (.A2(_1485_),
    .A1(\tdc_inst.fine_another_counter[4] ),
    .B1(\tdc_inst.fine_another_counter[5] ),
    .X(_1495_));
 sg13g2_nand2_1 _2869_ (.Y(_1496_),
    .A(net1209),
    .B(_1495_));
 sg13g2_xnor2_1 _2870_ (.Y(_1497_),
    .A(\tdc_inst.fine_another_counter[6] ),
    .B(_1496_));
 sg13g2_nand2b_1 _2871_ (.Y(_1498_),
    .B(_0735_),
    .A_N(_1490_));
 sg13g2_a21oi_1 _2872_ (.A1(net1546),
    .A2(_1490_),
    .Y(_1499_),
    .B1(_1474_));
 sg13g2_a22oi_1 _2873_ (.Y(_1500_),
    .B1(_1498_),
    .B2(net1547),
    .A2(_1497_),
    .A1(_1472_));
 sg13g2_nor2_1 _2874_ (.A(net1229),
    .B(net1548),
    .Y(_0645_));
 sg13g2_xnor2_1 _2875_ (.Y(_1501_),
    .A(_0037_),
    .B(_1498_));
 sg13g2_nor2_1 _2876_ (.A(_1474_),
    .B(_1501_),
    .Y(_1502_));
 sg13g2_nor2_1 _2877_ (.A(_0735_),
    .B(_1495_),
    .Y(_1503_));
 sg13g2_xor2_1 _2878_ (.B(_1503_),
    .A(_0037_),
    .X(_1504_));
 sg13g2_a221oi_1 _2879_ (.B2(_1504_),
    .C1(_1502_),
    .B1(_1456_),
    .A1(net1208),
    .Y(_1505_),
    .A2(net1803));
 sg13g2_nor2_1 _2880_ (.A(net1229),
    .B(net1804),
    .Y(_0646_));
 sg13g2_and3_1 _2881_ (.X(_1506_),
    .A(\tdc_inst.fine_another_counter[7] ),
    .B(\tdc_inst.fine_another_counter[6] ),
    .C(_1491_));
 sg13g2_xnor2_1 _2882_ (.Y(_1507_),
    .A(_0038_),
    .B(_1506_));
 sg13g2_nand3_1 _2883_ (.B(_1458_),
    .C(_1507_),
    .A(_0769_),
    .Y(_1508_));
 sg13g2_or3_1 _2884_ (.A(\tdc_inst.fine_another_counter[7] ),
    .B(\tdc_inst.fine_another_counter[6] ),
    .C(_1495_),
    .X(_1509_));
 sg13g2_or2_1 _2885_ (.X(_1510_),
    .B(_1509_),
    .A(_0038_));
 sg13g2_a21oi_1 _2886_ (.A1(_0038_),
    .A2(_1509_),
    .Y(_1511_),
    .B1(_1458_));
 sg13g2_a21oi_1 _2887_ (.A1(_1510_),
    .A2(_1511_),
    .Y(_1512_),
    .B1(net1208));
 sg13g2_o21ai_1 _2888_ (.B1(net1237),
    .Y(_1513_),
    .A1(net1776),
    .A2(net1209));
 sg13g2_a21oi_1 _2889_ (.A1(_1508_),
    .A2(_1512_),
    .Y(_0647_),
    .B1(_1513_));
 sg13g2_a21oi_1 _2890_ (.A1(\tdc_inst.start_count_debug[0] ),
    .A2(_0770_),
    .Y(_1514_),
    .B1(net1634));
 sg13g2_nand3_1 _2891_ (.B(\tdc_inst.start_count_debug[0] ),
    .C(_0770_),
    .A(net1634),
    .Y(_1515_));
 sg13g2_nand2_1 _2892_ (.Y(_1516_),
    .A(net1238),
    .B(_1515_));
 sg13g2_nor2_1 _2893_ (.A(net1635),
    .B(_1516_),
    .Y(_0648_));
 sg13g2_nor2b_1 _2894_ (.A(net1746),
    .B_N(_1515_),
    .Y(_1517_));
 sg13g2_and4_2 _2895_ (.A(net1746),
    .B(net1634),
    .C(\tdc_inst.start_count_debug[0] ),
    .D(net1119),
    .X(_1518_));
 sg13g2_nor3_1 _2896_ (.A(_0729_),
    .B(net1747),
    .C(_1518_),
    .Y(_0649_));
 sg13g2_xnor2_1 _2897_ (.Y(_1519_),
    .A(net1788),
    .B(_1518_));
 sg13g2_nor2_1 _2898_ (.A(net1228),
    .B(net1789),
    .Y(_0650_));
 sg13g2_a21oi_1 _2899_ (.A1(\tdc_inst.fine_start_counter[2] ),
    .A2(_1518_),
    .Y(_1520_),
    .B1(net1706));
 sg13g2_nand3_1 _2900_ (.B(\tdc_inst.fine_start_counter[2] ),
    .C(_1518_),
    .A(net1706),
    .Y(_1521_));
 sg13g2_nand2_1 _2901_ (.Y(_1522_),
    .A(net1238),
    .B(_1521_));
 sg13g2_nor2_1 _2902_ (.A(net1707),
    .B(_1522_),
    .Y(_0651_));
 sg13g2_nor2b_1 _2903_ (.A(net1751),
    .B_N(_1521_),
    .Y(_1523_));
 sg13g2_and4_2 _2904_ (.A(net1751),
    .B(\tdc_inst.fine_start_counter[3] ),
    .C(\tdc_inst.fine_start_counter[2] ),
    .D(_1518_),
    .X(_1524_));
 sg13g2_nor3_1 _2905_ (.A(net1228),
    .B(net1752),
    .C(_1524_),
    .Y(_0652_));
 sg13g2_xnor2_1 _2906_ (.Y(_1525_),
    .A(net1790),
    .B(_1524_));
 sg13g2_nor2_1 _2907_ (.A(net1228),
    .B(net1791),
    .Y(_0653_));
 sg13g2_a21oi_1 _2908_ (.A1(\tdc_inst.fine_start_counter[5] ),
    .A2(_1524_),
    .Y(_1526_),
    .B1(net1737));
 sg13g2_nand3_1 _2909_ (.B(net1790),
    .C(_1524_),
    .A(net1737),
    .Y(_1527_));
 sg13g2_nand2_1 _2910_ (.Y(_1528_),
    .A(net1236),
    .B(_1527_));
 sg13g2_nor2_1 _2911_ (.A(net1738),
    .B(_1528_),
    .Y(_0654_));
 sg13g2_nand2b_1 _2912_ (.Y(_1529_),
    .B(_1527_),
    .A_N(net1793));
 sg13g2_nand4_1 _2913_ (.B(net1737),
    .C(\tdc_inst.fine_start_counter[5] ),
    .A(net1793),
    .Y(_1530_),
    .D(_1524_));
 sg13g2_and3_1 _2914_ (.X(_0655_),
    .A(net1236),
    .B(_1529_),
    .C(_1530_));
 sg13g2_o21ai_1 _2915_ (.B1(net1236),
    .Y(_1531_),
    .A1(_0710_),
    .A2(_1530_));
 sg13g2_a21oi_1 _2916_ (.A1(_0710_),
    .A2(_1530_),
    .Y(_0656_),
    .B1(_1531_));
 sg13g2_a21oi_1 _2917_ (.A1(\tdc_inst.stop_count_debug[0] ),
    .A2(net1119),
    .Y(_1532_),
    .B1(net1427));
 sg13g2_nand3_1 _2918_ (.B(\tdc_inst.stop_count_debug[0] ),
    .C(net1119),
    .A(net1427),
    .Y(_1533_));
 sg13g2_nand2_1 _2919_ (.Y(_1534_),
    .A(net1238),
    .B(_1533_));
 sg13g2_nor2_1 _2920_ (.A(net1428),
    .B(_1534_),
    .Y(_0657_));
 sg13g2_nor2b_1 _2921_ (.A(net1709),
    .B_N(_1533_),
    .Y(_1535_));
 sg13g2_and4_2 _2922_ (.A(net1709),
    .B(net1427),
    .C(\tdc_inst.stop_count_debug[0] ),
    .D(net1119),
    .X(_1536_));
 sg13g2_nor3_1 _2923_ (.A(net1228),
    .B(net1710),
    .C(_1536_),
    .Y(_0658_));
 sg13g2_xnor2_1 _2924_ (.Y(_1537_),
    .A(net1785),
    .B(_1536_));
 sg13g2_nor2_1 _2925_ (.A(net1228),
    .B(net1786),
    .Y(_0659_));
 sg13g2_a21oi_1 _2926_ (.A1(\tdc_inst.fine_stop_counter[2] ),
    .A2(_1536_),
    .Y(_1538_),
    .B1(net1688));
 sg13g2_nand3_1 _2927_ (.B(net1810),
    .C(_1536_),
    .A(net1688),
    .Y(_1539_));
 sg13g2_nand2_1 _2928_ (.Y(_1540_),
    .A(net1236),
    .B(_1539_));
 sg13g2_nor2_1 _2929_ (.A(net1689),
    .B(_1540_),
    .Y(_0660_));
 sg13g2_nor2b_1 _2930_ (.A(net1762),
    .B_N(_1539_),
    .Y(_1541_));
 sg13g2_and4_2 _2931_ (.A(net1762),
    .B(net1688),
    .C(\tdc_inst.fine_stop_counter[2] ),
    .D(_1536_),
    .X(_1542_));
 sg13g2_nor3_1 _2932_ (.A(net1228),
    .B(net1763),
    .C(_1542_),
    .Y(_0661_));
 sg13g2_xnor2_1 _2933_ (.Y(_1543_),
    .A(net1798),
    .B(_1542_));
 sg13g2_nor2_1 _2934_ (.A(net1229),
    .B(_1543_),
    .Y(_0662_));
 sg13g2_a21oi_1 _2935_ (.A1(\tdc_inst.fine_stop_counter[5] ),
    .A2(_1542_),
    .Y(_1544_),
    .B1(net1758));
 sg13g2_nand3_1 _2936_ (.B(net1811),
    .C(_1542_),
    .A(net1758),
    .Y(_1545_));
 sg13g2_nand2_1 _2937_ (.Y(_1546_),
    .A(net1236),
    .B(_1545_));
 sg13g2_nor2_1 _2938_ (.A(net1759),
    .B(_1546_),
    .Y(_0663_));
 sg13g2_nand2b_1 _2939_ (.Y(_1547_),
    .B(_1545_),
    .A_N(net1795));
 sg13g2_nand4_1 _2940_ (.B(\tdc_inst.fine_stop_counter[6] ),
    .C(\tdc_inst.fine_stop_counter[5] ),
    .A(net1795),
    .Y(_1548_),
    .D(_1542_));
 sg13g2_and3_1 _2941_ (.X(_0664_),
    .A(net1236),
    .B(net1796),
    .C(_1548_));
 sg13g2_o21ai_1 _2942_ (.B1(net1236),
    .Y(_1549_),
    .A1(_0708_),
    .A2(_1548_));
 sg13g2_a21oi_1 _2943_ (.A1(_0708_),
    .A2(_1548_),
    .Y(_0665_),
    .B1(_1549_));
 sg13g2_mux2_1 _2944_ (.A0(net604),
    .A1(net632),
    .S(net1262),
    .X(_0666_));
 sg13g2_o21ai_1 _2945_ (.B1(net1237),
    .Y(_1550_),
    .A1(_0004_),
    .A2(_1439_));
 sg13g2_a21oi_1 _2946_ (.A1(_0707_),
    .A2(_1439_),
    .Y(_0667_),
    .B1(_1550_));
 sg13g2_nor2_1 _2947_ (.A(net843),
    .B(net1067),
    .Y(_1551_));
 sg13g2_nand2_1 _2948_ (.Y(_1552_),
    .A(\tdc_inst.fine_stop_counter[4] ),
    .B(\tdc_inst.fine_start_counter[4] ));
 sg13g2_xor2_1 _2949_ (.B(\tdc_inst.fine_start_counter[4] ),
    .A(\tdc_inst.fine_stop_counter[4] ),
    .X(_1553_));
 sg13g2_nor2_1 _2950_ (.A(\tdc_inst.fine_stop_counter[2] ),
    .B(\tdc_inst.fine_start_counter[2] ),
    .Y(_1554_));
 sg13g2_nor2_1 _2951_ (.A(\tdc_inst.fine_stop_counter[1] ),
    .B(\tdc_inst.fine_start_counter[1] ),
    .Y(_1555_));
 sg13g2_a22oi_1 _2952_ (.Y(_1556_),
    .B1(\tdc_inst.fine_start_counter[0] ),
    .B2(\tdc_inst.fine_stop_counter[0] ),
    .A2(\tdc_inst.fine_start_counter[1] ),
    .A1(\tdc_inst.fine_stop_counter[1] ));
 sg13g2_or3_1 _2953_ (.A(_1554_),
    .B(_1555_),
    .C(_1556_),
    .X(_1557_));
 sg13g2_a22oi_1 _2954_ (.Y(_1558_),
    .B1(\tdc_inst.fine_start_counter[2] ),
    .B2(\tdc_inst.fine_stop_counter[2] ),
    .A2(\tdc_inst.fine_start_counter[3] ),
    .A1(\tdc_inst.fine_stop_counter[3] ));
 sg13g2_a22oi_1 _2955_ (.Y(_1559_),
    .B1(_1557_),
    .B2(_1558_),
    .A2(_0711_),
    .A1(_0709_));
 sg13g2_nand2_1 _2956_ (.Y(_1560_),
    .A(_1553_),
    .B(_1559_));
 sg13g2_xnor2_1 _2957_ (.Y(_1561_),
    .A(_1553_),
    .B(_1559_));
 sg13g2_a21oi_1 _2958_ (.A1(net1067),
    .A2(_1561_),
    .Y(_0668_),
    .B1(_1551_));
 sg13g2_nor2_1 _2959_ (.A(net936),
    .B(net1056),
    .Y(_1562_));
 sg13g2_nand2_1 _2960_ (.Y(_1563_),
    .A(\tdc_inst.fine_stop_counter[5] ),
    .B(\tdc_inst.fine_start_counter[5] ));
 sg13g2_nor2_1 _2961_ (.A(\tdc_inst.fine_stop_counter[5] ),
    .B(\tdc_inst.fine_start_counter[5] ),
    .Y(_1564_));
 sg13g2_xor2_1 _2962_ (.B(\tdc_inst.fine_start_counter[5] ),
    .A(\tdc_inst.fine_stop_counter[5] ),
    .X(_1565_));
 sg13g2_nand2_1 _2963_ (.Y(_1566_),
    .A(_1552_),
    .B(_1560_));
 sg13g2_xnor2_1 _2964_ (.Y(_1567_),
    .A(_1565_),
    .B(_1566_));
 sg13g2_a21oi_1 _2965_ (.A1(net1056),
    .A2(_1567_),
    .Y(_0669_),
    .B1(_1562_));
 sg13g2_nand2_1 _2966_ (.Y(_1568_),
    .A(\tdc_inst.fine_stop_counter[6] ),
    .B(\tdc_inst.fine_start_counter[6] ));
 sg13g2_xor2_1 _2967_ (.B(\tdc_inst.fine_start_counter[6] ),
    .A(\tdc_inst.fine_stop_counter[6] ),
    .X(_1569_));
 sg13g2_o21ai_1 _2968_ (.B1(_1563_),
    .Y(_1570_),
    .A1(_1552_),
    .A2(_1564_));
 sg13g2_nand3b_1 _2969_ (.B(_1553_),
    .C(_1563_),
    .Y(_1571_),
    .A_N(_1564_));
 sg13g2_a221oi_1 _2970_ (.B2(_1558_),
    .C1(_1571_),
    .B1(_1557_),
    .A1(_0709_),
    .Y(_1572_),
    .A2(_0711_));
 sg13g2_o21ai_1 _2971_ (.B1(_1569_),
    .Y(_1573_),
    .A1(_1570_),
    .A2(_1572_));
 sg13g2_or3_1 _2972_ (.A(_1569_),
    .B(_1570_),
    .C(_1572_),
    .X(_1574_));
 sg13g2_nand3_1 _2973_ (.B(_1573_),
    .C(_1574_),
    .A(net1057),
    .Y(_1575_));
 sg13g2_o21ai_1 _2974_ (.B1(_1575_),
    .Y(_0670_),
    .A1(_0732_),
    .A2(net1057));
 sg13g2_xnor2_1 _2975_ (.Y(_1576_),
    .A(\tdc_inst.fine_stop_counter[7] ),
    .B(\tdc_inst.fine_start_counter[7] ));
 sg13g2_and3_1 _2976_ (.X(_1577_),
    .A(_1568_),
    .B(_1573_),
    .C(_1576_));
 sg13g2_a21oi_1 _2977_ (.A1(_1568_),
    .A2(_1573_),
    .Y(_1578_),
    .B1(_1576_));
 sg13g2_nor2_1 _2978_ (.A(_1577_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_mux2_1 _2979_ (.A0(net1657),
    .A1(_1579_),
    .S(net1057),
    .X(_0671_));
 sg13g2_nor2_1 _2980_ (.A(net1624),
    .B(net1070),
    .Y(_1580_));
 sg13g2_a21oi_1 _2981_ (.A1(\tdc_inst.fine_stop_counter[7] ),
    .A2(\tdc_inst.fine_start_counter[7] ),
    .Y(_1581_),
    .B1(_1578_));
 sg13g2_xnor2_1 _2982_ (.Y(_1582_),
    .A(\tdc_inst.fine_stop_counter[8] ),
    .B(net1537));
 sg13g2_xnor2_1 _2983_ (.Y(_1583_),
    .A(_1581_),
    .B(_1582_));
 sg13g2_a21oi_1 _2984_ (.A1(net1057),
    .A2(_1583_),
    .Y(_0672_),
    .B1(_1580_));
 sg13g2_xor2_1 _2985_ (.B(\tdc_inst.start_signal_activated ),
    .A(net1210),
    .X(_1584_));
 sg13g2_nand2_1 _2986_ (.Y(_1585_),
    .A(_0044_),
    .B(_1584_));
 sg13g2_o21ai_1 _2987_ (.B1(_1585_),
    .Y(_0673_),
    .A1(_0720_),
    .A2(_1584_));
 sg13g2_nand3_1 _2988_ (.B(\tdc_inst.coarse_count[1] ),
    .C(_1584_),
    .A(\tdc_inst.coarse_count[0] ),
    .Y(_1586_));
 sg13g2_a21o_1 _2989_ (.A2(_1584_),
    .A1(\tdc_inst.coarse_count[0] ),
    .B1(\tdc_inst.coarse_count[1] ),
    .X(_1587_));
 sg13g2_and2_1 _2990_ (.A(_1586_),
    .B(_1587_),
    .X(_0674_));
 sg13g2_and4_2 _2991_ (.A(\tdc_inst.coarse_count[0] ),
    .B(\tdc_inst.coarse_count[1] ),
    .C(\tdc_inst.coarse_count[2] ),
    .D(_1584_),
    .X(_1588_));
 sg13g2_xnor2_1 _2992_ (.Y(_0675_),
    .A(\tdc_inst.coarse_count[2] ),
    .B(_1586_));
 sg13g2_and2_1 _2993_ (.A(\tdc_inst.coarse_count[3] ),
    .B(_1588_),
    .X(_1589_));
 sg13g2_xor2_1 _2994_ (.B(_1588_),
    .A(\tdc_inst.coarse_count[3] ),
    .X(_0676_));
 sg13g2_xor2_1 _2995_ (.B(_1589_),
    .A(\tdc_inst.coarse_count[4] ),
    .X(_0677_));
 sg13g2_and4_2 _2996_ (.A(\tdc_inst.coarse_count[3] ),
    .B(\tdc_inst.coarse_count[5] ),
    .C(\tdc_inst.coarse_count[4] ),
    .D(_1588_),
    .X(_1590_));
 sg13g2_a21oi_1 _2997_ (.A1(\tdc_inst.coarse_count[4] ),
    .A2(_1589_),
    .Y(_1591_),
    .B1(\tdc_inst.coarse_count[5] ));
 sg13g2_nor2_1 _2998_ (.A(_1590_),
    .B(_1591_),
    .Y(_0678_));
 sg13g2_and2_1 _2999_ (.A(\tdc_inst.coarse_count[6] ),
    .B(_1590_),
    .X(_1592_));
 sg13g2_xor2_1 _3000_ (.B(_1590_),
    .A(\tdc_inst.coarse_count[6] ),
    .X(_0679_));
 sg13g2_xor2_1 _3001_ (.B(_1592_),
    .A(\tdc_inst.coarse_count[7] ),
    .X(_0680_));
 sg13g2_nand3_1 _3002_ (.B(\tdc_inst.coarse_count[8] ),
    .C(_1592_),
    .A(\tdc_inst.coarse_count[7] ),
    .Y(_1593_));
 sg13g2_a21o_1 _3003_ (.A2(_1592_),
    .A1(\tdc_inst.coarse_count[7] ),
    .B1(\tdc_inst.coarse_count[8] ),
    .X(_1594_));
 sg13g2_and2_1 _3004_ (.A(_1593_),
    .B(_1594_),
    .X(_0681_));
 sg13g2_and2_1 _3005_ (.A(\tdc_inst.coarse_count[9] ),
    .B(\tdc_inst.coarse_count[8] ),
    .X(_1595_));
 sg13g2_and3_1 _3006_ (.X(_1596_),
    .A(\tdc_inst.coarse_count[7] ),
    .B(_1592_),
    .C(_1595_));
 sg13g2_nand4_1 _3007_ (.B(\tdc_inst.coarse_count[6] ),
    .C(_1590_),
    .A(\tdc_inst.coarse_count[7] ),
    .Y(_1597_),
    .D(_1595_));
 sg13g2_a21oi_1 _3008_ (.A1(_0736_),
    .A2(_1593_),
    .Y(_0682_),
    .B1(_1596_));
 sg13g2_and2_1 _3009_ (.A(\tdc_inst.coarse_count[10] ),
    .B(_1596_),
    .X(_1598_));
 sg13g2_xnor2_1 _3010_ (.Y(_0683_),
    .A(\tdc_inst.coarse_count[10] ),
    .B(_1597_));
 sg13g2_xor2_1 _3011_ (.B(_1598_),
    .A(\tdc_inst.coarse_count[11] ),
    .X(_0684_));
 sg13g2_a21oi_1 _3012_ (.A1(\tdc_inst.coarse_count[11] ),
    .A2(_1598_),
    .Y(_1599_),
    .B1(\tdc_inst.coarse_count[12] ));
 sg13g2_nand3_1 _3013_ (.B(\tdc_inst.coarse_count[12] ),
    .C(_1598_),
    .A(\tdc_inst.coarse_count[11] ),
    .Y(_1600_));
 sg13g2_nor2b_1 _3014_ (.A(_1599_),
    .B_N(_1600_),
    .Y(_0685_));
 sg13g2_xnor2_1 _3015_ (.Y(_0686_),
    .A(\tdc_inst.coarse_count[13] ),
    .B(_1600_));
 sg13g2_nand4_1 _3016_ (.B(\tdc_inst.coarse_count[10] ),
    .C(\tdc_inst.coarse_count[13] ),
    .A(\tdc_inst.coarse_count[11] ),
    .Y(_1601_),
    .D(\tdc_inst.coarse_count[12] ));
 sg13g2_nor2_1 _3017_ (.A(_1597_),
    .B(_1601_),
    .Y(_1602_));
 sg13g2_xor2_1 _3018_ (.B(_1602_),
    .A(\tdc_inst.coarse_count[14] ),
    .X(_0687_));
 sg13g2_nor3_1 _3019_ (.A(_0039_),
    .B(_1597_),
    .C(_1601_),
    .Y(_1603_));
 sg13g2_xor2_1 _3020_ (.B(_1603_),
    .A(\tdc_inst.coarse_count[15] ),
    .X(_0688_));
 sg13g2_nand3_1 _3021_ (.B(\tdc_inst.coarse_count[14] ),
    .C(\tdc_inst.coarse_count[16] ),
    .A(\tdc_inst.coarse_count[15] ),
    .Y(_1604_));
 sg13g2_nor3_2 _3022_ (.A(_1597_),
    .B(_1601_),
    .C(_1604_),
    .Y(_1605_));
 sg13g2_nand3_1 _3023_ (.B(\tdc_inst.coarse_count[14] ),
    .C(_1602_),
    .A(\tdc_inst.coarse_count[15] ),
    .Y(_1606_));
 sg13g2_a21oi_1 _3024_ (.A1(_0737_),
    .A2(_1606_),
    .Y(_0689_),
    .B1(_1605_));
 sg13g2_nand2_1 _3025_ (.Y(_1607_),
    .A(\tdc_inst.coarse_count[17] ),
    .B(_1605_));
 sg13g2_xor2_1 _3026_ (.B(_1605_),
    .A(\tdc_inst.coarse_count[17] ),
    .X(_0690_));
 sg13g2_xnor2_1 _3027_ (.Y(_0691_),
    .A(\tdc_inst.coarse_count[18] ),
    .B(_1607_));
 sg13g2_nor2_1 _3028_ (.A(_0040_),
    .B(_1607_),
    .Y(_1608_));
 sg13g2_xor2_1 _3029_ (.B(_1608_),
    .A(\tdc_inst.coarse_count[19] ),
    .X(_0692_));
 sg13g2_nand3_1 _3030_ (.B(\tdc_inst.coarse_count[19] ),
    .C(\tdc_inst.coarse_count[18] ),
    .A(\tdc_inst.coarse_count[17] ),
    .Y(_1609_));
 sg13g2_nor4_2 _3031_ (.A(_1597_),
    .B(_1601_),
    .C(_1604_),
    .Y(_1610_),
    .D(_1609_));
 sg13g2_and2_1 _3032_ (.A(\tdc_inst.coarse_count[20] ),
    .B(_1610_),
    .X(_1611_));
 sg13g2_xor2_1 _3033_ (.B(_1610_),
    .A(\tdc_inst.coarse_count[20] ),
    .X(_0693_));
 sg13g2_nand3_1 _3034_ (.B(\tdc_inst.coarse_count[20] ),
    .C(_1610_),
    .A(\tdc_inst.coarse_count[21] ),
    .Y(_1612_));
 sg13g2_xor2_1 _3035_ (.B(_1611_),
    .A(\tdc_inst.coarse_count[21] ),
    .X(_0694_));
 sg13g2_xnor2_1 _3036_ (.Y(_0695_),
    .A(\tdc_inst.coarse_count[22] ),
    .B(_1612_));
 sg13g2_nor2_1 _3037_ (.A(_0041_),
    .B(_1612_),
    .Y(_1613_));
 sg13g2_xor2_1 _3038_ (.B(_1613_),
    .A(\tdc_inst.coarse_count[23] ),
    .X(_0696_));
 sg13g2_and3_1 _3039_ (.X(_1614_),
    .A(\tdc_inst.coarse_count[21] ),
    .B(\tdc_inst.coarse_count[23] ),
    .C(\tdc_inst.coarse_count[22] ));
 sg13g2_and4_2 _3040_ (.A(\tdc_inst.coarse_count[20] ),
    .B(\tdc_inst.coarse_count[24] ),
    .C(_1610_),
    .D(_1614_),
    .X(_1615_));
 sg13g2_nand4_1 _3041_ (.B(\tdc_inst.coarse_count[24] ),
    .C(_1610_),
    .A(\tdc_inst.coarse_count[20] ),
    .Y(_1616_),
    .D(_1614_));
 sg13g2_a21oi_1 _3042_ (.A1(_1611_),
    .A2(_1614_),
    .Y(_1617_),
    .B1(\tdc_inst.coarse_count[24] ));
 sg13g2_nor2_1 _3043_ (.A(_1615_),
    .B(_1617_),
    .Y(_0697_));
 sg13g2_nand2_1 _3044_ (.Y(_1618_),
    .A(\tdc_inst.coarse_count[25] ),
    .B(_1615_));
 sg13g2_xnor2_1 _3045_ (.Y(_0698_),
    .A(_0738_),
    .B(_1615_));
 sg13g2_xnor2_1 _3046_ (.Y(_0699_),
    .A(\tdc_inst.coarse_count[26] ),
    .B(_1618_));
 sg13g2_nor3_1 _3047_ (.A(_0738_),
    .B(_0042_),
    .C(_1616_),
    .Y(_1619_));
 sg13g2_xor2_1 _3048_ (.B(_1619_),
    .A(\tdc_inst.coarse_count[27] ),
    .X(_0700_));
 sg13g2_nand3_1 _3049_ (.B(\tdc_inst.coarse_count[27] ),
    .C(\tdc_inst.coarse_count[26] ),
    .A(\tdc_inst.coarse_count[25] ),
    .Y(_1620_));
 sg13g2_inv_1 _3050_ (.Y(_1621_),
    .A(_1620_));
 sg13g2_nand2_1 _3051_ (.Y(_1622_),
    .A(_1615_),
    .B(_1621_));
 sg13g2_nand3_1 _3052_ (.B(_1615_),
    .C(_1621_),
    .A(\tdc_inst.coarse_count[28] ),
    .Y(_1623_));
 sg13g2_xnor2_1 _3053_ (.Y(_0701_),
    .A(\tdc_inst.coarse_count[28] ),
    .B(_1622_));
 sg13g2_nand2_1 _3054_ (.Y(_1624_),
    .A(\tdc_inst.coarse_count[29] ),
    .B(\tdc_inst.coarse_count[28] ));
 sg13g2_nor3_1 _3055_ (.A(_1616_),
    .B(_1620_),
    .C(_1624_),
    .Y(_1625_));
 sg13g2_a21oi_1 _3056_ (.A1(_0739_),
    .A2(_1623_),
    .Y(_0702_),
    .B1(_1625_));
 sg13g2_xor2_1 _3057_ (.B(_1625_),
    .A(\tdc_inst.coarse_count[30] ),
    .X(_0703_));
 sg13g2_nor4_1 _3058_ (.A(_0043_),
    .B(_1616_),
    .C(_1620_),
    .D(_1624_),
    .Y(_1626_));
 sg13g2_xor2_1 _3059_ (.B(_1626_),
    .A(\tdc_inst.coarse_count[31] ),
    .X(_0704_));
 sg13g2_mux2_1 _3060_ (.A0(\tdc_inst.stop_signal_sampling_clock_level ),
    .A1(net1235),
    .S(net1215),
    .X(_0705_));
 sg13g2_a21oi_1 _3061_ (.A1(net1766),
    .A2(_1473_),
    .Y(_1627_),
    .B1(\tdc_inst.fine_another_counter[0] ));
 sg13g2_a21oi_1 _3062_ (.A1(_0769_),
    .A2(_1448_),
    .Y(_1628_),
    .B1(_1472_));
 sg13g2_nor3_1 _3063_ (.A(net1229),
    .B(net1767),
    .C(_1628_),
    .Y(_0706_));
 sg13g2_inv_1 _3064_ (.Y(_0707_),
    .A(net1215));
 sg13g2_inv_1 _3065_ (.Y(_0708_),
    .A(net1712));
 sg13g2_inv_1 _3066_ (.Y(_0709_),
    .A(\tdc_inst.fine_stop_counter[3] ));
 sg13g2_inv_1 _3067_ (.Y(_0710_),
    .A(net1537));
 sg13g2_inv_1 _3068_ (.Y(_0711_),
    .A(\tdc_inst.fine_start_counter[3] ));
 sg13g2_inv_1 _3069_ (.Y(_0712_),
    .A(net1210));
 sg13g2_inv_1 _3070_ (.Y(_0713_),
    .A(net1799));
 sg13g2_inv_1 _3071_ (.Y(_0714_),
    .A(net1774));
 sg13g2_inv_1 _3072_ (.Y(_0715_),
    .A(net770));
 sg13g2_inv_1 _3073_ (.Y(_0716_),
    .A(net1295));
 sg13g2_inv_1 _3074_ (.Y(_0717_),
    .A(net935));
 sg13g2_inv_1 _3075_ (.Y(_0718_),
    .A(net810));
 sg13g2_inv_1 _3076_ (.Y(_0719_),
    .A(net1274));
 sg13g2_inv_1 _3077_ (.Y(_0720_),
    .A(\tdc_inst.coarse_count[0] ));
 sg13g2_inv_1 _3078_ (.Y(_0721_),
    .A(net661));
 sg13g2_inv_1 _3079_ (.Y(_0722_),
    .A(net1259));
 sg13g2_inv_1 _3080_ (.Y(_0723_),
    .A(net1627));
 sg13g2_inv_1 _3081_ (.Y(_0724_),
    .A(net1769));
 sg13g2_inv_1 _3082_ (.Y(_0725_),
    .A(net1792));
 sg13g2_inv_1 _3083_ (.Y(_0726_),
    .A(net1780));
 sg13g2_inv_1 _3084_ (.Y(_0727_),
    .A(net555));
 sg13g2_inv_1 _3085_ (.Y(_0728_),
    .A(net596));
 sg13g2_inv_2 _3086_ (.Y(_0729_),
    .A(net1236));
 sg13g2_inv_1 _3087_ (.Y(_0730_),
    .A(net1227));
 sg13g2_inv_1 _3088_ (.Y(_0731_),
    .A(net1226));
 sg13g2_inv_1 _3089_ (.Y(_0732_),
    .A(net730));
 sg13g2_inv_1 _3090_ (.Y(_0733_),
    .A(_0010_));
 sg13g2_inv_2 _3091_ (.Y(_0734_),
    .A(net1224));
 sg13g2_inv_1 _3092_ (.Y(_0735_),
    .A(net1546));
 sg13g2_inv_1 _3093_ (.Y(_0736_),
    .A(\tdc_inst.coarse_count[9] ));
 sg13g2_inv_1 _3094_ (.Y(_0737_),
    .A(\tdc_inst.coarse_count[16] ));
 sg13g2_inv_1 _3095_ (.Y(_0738_),
    .A(\tdc_inst.coarse_count[25] ));
 sg13g2_inv_1 _3096_ (.Y(_0739_),
    .A(\tdc_inst.coarse_count[29] ));
 sg13g2_nor3_2 _3097_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .B(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ),
    .C(net1784),
    .Y(_0740_));
 sg13g2_nand2b_1 _3098_ (.Y(_0741_),
    .B(net1405),
    .A_N(_0740_));
 sg13g2_nor4_2 _3099_ (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ),
    .B(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .C(_0726_),
    .Y(_0742_),
    .D(net1794));
 sg13g2_nor2_1 _3100_ (.A(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .B(\spi_wrapper_i.spi_reg_inst.state[4] ),
    .Y(_0743_));
 sg13g2_o21ai_1 _3101_ (.B1(_0741_),
    .Y(_0744_),
    .A1(_0742_),
    .A2(_0743_));
 sg13g2_nor2b_1 _3102_ (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .B_N(spi_cs_n_sync),
    .Y(_0745_));
 sg13g2_nand3_1 _3103_ (.B(_0744_),
    .C(_0745_),
    .A(net1259),
    .Y(_0746_));
 sg13g2_nand3_1 _3104_ (.B(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .C(_0740_),
    .A(net1262),
    .Y(_0747_));
 sg13g2_nand4_1 _3105_ (.B(net1809),
    .C(net1405),
    .A(net1259),
    .Y(_0748_),
    .D(_0740_));
 sg13g2_and2_1 _3106_ (.A(net1260),
    .B(net1699),
    .X(_0749_));
 sg13g2_nand2_2 _3107_ (.Y(_0750_),
    .A(net1475),
    .B(_0749_));
 sg13g2_nor2b_2 _3108_ (.A(spi_cs_n_sync),
    .B_N(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .Y(_0751_));
 sg13g2_nand2_1 _3109_ (.Y(_0752_),
    .A(net1259),
    .B(_0751_));
 sg13g2_nand2_1 _3110_ (.Y(_0753_),
    .A(net555),
    .B(_0752_));
 sg13g2_and4_1 _3111_ (.A(_0746_),
    .B(_0748_),
    .C(net1042),
    .D(_0753_),
    .X(_0046_));
 sg13g2_nand2_1 _3112_ (.Y(_0754_),
    .A(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .B(_0740_));
 sg13g2_nor2_2 _3113_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_nand3b_1 _3114_ (.B(net1405),
    .C(_0740_),
    .Y(_0756_),
    .A_N(net1812));
 sg13g2_nor2_1 _3115_ (.A(net1259),
    .B(net1405),
    .Y(_0757_));
 sg13g2_o21ai_1 _3116_ (.B1(net1259),
    .Y(_0758_),
    .A1(_0741_),
    .A2(_0745_));
 sg13g2_a21oi_1 _3117_ (.A1(_0721_),
    .A2(net1627),
    .Y(_0759_),
    .B1(_0758_));
 sg13g2_o21ai_1 _3118_ (.B1(net1133),
    .Y(_0000_),
    .A1(_0757_),
    .A2(_0759_));
 sg13g2_nand2_1 _3119_ (.Y(_0760_),
    .A(net1613),
    .B(_0749_));
 sg13g2_o21ai_1 _3120_ (.B1(_0760_),
    .Y(_0001_),
    .A1(net1260),
    .A2(_0723_));
 sg13g2_o21ai_1 _3121_ (.B1(net1259),
    .Y(_0761_),
    .A1(_0742_),
    .A2(_0745_));
 sg13g2_nand2_1 _3122_ (.Y(_0762_),
    .A(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .B(_0761_));
 sg13g2_o21ai_1 _3123_ (.B1(_0762_),
    .Y(_0002_),
    .A1(_0727_),
    .A2(_0752_));
 sg13g2_nand2_1 _3124_ (.Y(_0763_),
    .A(\spi_wrapper_i.spi_reg_inst.state[4] ),
    .B(_0761_));
 sg13g2_nand3_1 _3125_ (.B(net1260),
    .C(\spi_wrapper_i.spi_reg_inst.state[2] ),
    .A(net661),
    .Y(_0764_));
 sg13g2_nand2_1 _3126_ (.Y(_0003_),
    .A(_0763_),
    .B(net662));
 sg13g2_or2_1 _3127_ (.X(\tdc_inst.busy ),
    .B(\tdc_inst.start_signal_activated ),
    .A(net1210));
 sg13g2_nor2_1 _3128_ (.A(\tdc_inst.fine_procedure_counter[6] ),
    .B(\tdc_inst.fine_procedure_counter[5] ),
    .Y(_0765_));
 sg13g2_nor4_2 _3129_ (.A(\tdc_inst.fine_procedure_counter[6] ),
    .B(\tdc_inst.fine_procedure_counter[5] ),
    .C(\tdc_inst.fine_procedure_counter[3] ),
    .Y(_0766_),
    .D(\tdc_inst.fine_procedure_counter[2] ));
 sg13g2_nor2_1 _3130_ (.A(\tdc_inst.fine_procedure_counter[7] ),
    .B(\tdc_inst.fine_procedure_counter[4] ),
    .Y(_0767_));
 sg13g2_nor2_1 _3131_ (.A(\tdc_inst.fine_procedure_counter[1] ),
    .B(\tdc_inst.fine_procedure_counter[0] ),
    .Y(_0768_));
 sg13g2_nand4_1 _3132_ (.B(_0766_),
    .C(_0767_),
    .A(_0006_),
    .Y(_0769_),
    .D(_0768_));
 sg13g2_and2_1 _3133_ (.A(net1209),
    .B(_0769_),
    .X(_0770_));
 sg13g2_nand2_1 _3134_ (.Y(_0771_),
    .A(net1210),
    .B(net1244));
 sg13g2_nor2b_1 _3135_ (.A(net1159),
    .B_N(_0769_),
    .Y(_0772_));
 sg13g2_nor2_2 _3136_ (.A(_0769_),
    .B(net1159),
    .Y(_0773_));
 sg13g2_and2_1 _3137_ (.A(\tdc_inst.start_signal_sampling_clock_level ),
    .B(_0773_),
    .X(_0774_));
 sg13g2_nand2_1 _3138_ (.Y(_0775_),
    .A(\tdc_inst.start_signal_sampling_clock_level ),
    .B(_0773_));
 sg13g2_a22oi_1 _3139_ (.Y(_0776_),
    .B1(net1071),
    .B2(net1741),
    .A2(net1158),
    .A1(\tdc_inst.start_count_debug[0] ));
 sg13g2_nand2_1 _3140_ (.Y(_0047_),
    .A(net1016),
    .B(net1742));
 sg13g2_a22oi_1 _3141_ (.Y(_0777_),
    .B1(net1071),
    .B2(net897),
    .A2(net1158),
    .A1(\tdc_inst.start_count_debug[1] ));
 sg13g2_nand2_1 _3142_ (.Y(_0048_),
    .A(net1016),
    .B(net898));
 sg13g2_a22oi_1 _3143_ (.Y(_0778_),
    .B1(net1095),
    .B2(net1582),
    .A2(net1184),
    .A1(net897));
 sg13g2_nand2_1 _3144_ (.Y(_0049_),
    .A(net1016),
    .B(_0778_));
 sg13g2_a22oi_1 _3145_ (.Y(_0779_),
    .B1(net1095),
    .B2(net580),
    .A2(net1184),
    .A1(\tdc_inst.start_count_debug[3] ));
 sg13g2_nand2_1 _3146_ (.Y(_0050_),
    .A(net1016),
    .B(net581));
 sg13g2_a22oi_1 _3147_ (.Y(_0780_),
    .B1(net1095),
    .B2(net1704),
    .A2(net1184),
    .A1(net580));
 sg13g2_nand2_1 _3148_ (.Y(_0051_),
    .A(net1016),
    .B(_0780_));
 sg13g2_a22oi_1 _3149_ (.Y(_0781_),
    .B1(net1096),
    .B2(net1631),
    .A2(net1185),
    .A1(\tdc_inst.start_count_debug[5] ));
 sg13g2_nand2_1 _3150_ (.Y(_0052_),
    .A(net1016),
    .B(net1632));
 sg13g2_a22oi_1 _3151_ (.Y(_0782_),
    .B1(net1096),
    .B2(net1373),
    .A2(net1185),
    .A1(\tdc_inst.start_count_debug[6] ));
 sg13g2_nand2_1 _3152_ (.Y(_0053_),
    .A(net1021),
    .B(net1374));
 sg13g2_a22oi_1 _3153_ (.Y(_0783_),
    .B1(net1095),
    .B2(net1587),
    .A2(net1184),
    .A1(net1373));
 sg13g2_nand2_1 _3154_ (.Y(_0054_),
    .A(net1019),
    .B(_0783_));
 sg13g2_a22oi_1 _3155_ (.Y(_0784_),
    .B1(net1096),
    .B2(net624),
    .A2(net1185),
    .A1(\tdc_inst.start_count_debug[8] ));
 sg13g2_nand2_1 _3156_ (.Y(_0055_),
    .A(net1017),
    .B(net625));
 sg13g2_a22oi_1 _3157_ (.Y(_0785_),
    .B1(net1096),
    .B2(net1555),
    .A2(net1185),
    .A1(net624));
 sg13g2_nand2_1 _3158_ (.Y(_0056_),
    .A(net1017),
    .B(_0785_));
 sg13g2_a22oi_1 _3159_ (.Y(_0786_),
    .B1(net1095),
    .B2(net808),
    .A2(net1184),
    .A1(\tdc_inst.start_count_debug[10] ));
 sg13g2_nand2_1 _3160_ (.Y(_0057_),
    .A(net1017),
    .B(net809));
 sg13g2_a22oi_1 _3161_ (.Y(_0787_),
    .B1(net1095),
    .B2(net1703),
    .A2(net1184),
    .A1(net808));
 sg13g2_nand2_1 _3162_ (.Y(_0058_),
    .A(net1017),
    .B(_0787_));
 sg13g2_a22oi_1 _3163_ (.Y(_0788_),
    .B1(net1098),
    .B2(net949),
    .A2(net1187),
    .A1(\tdc_inst.start_count_debug[12] ));
 sg13g2_nand2_1 _3164_ (.Y(_0059_),
    .A(net1017),
    .B(net950));
 sg13g2_a22oi_1 _3165_ (.Y(_0789_),
    .B1(net1098),
    .B2(net1300),
    .A2(net1187),
    .A1(net949));
 sg13g2_nand2_1 _3166_ (.Y(_0060_),
    .A(net1017),
    .B(_0789_));
 sg13g2_a22oi_1 _3167_ (.Y(_0790_),
    .B1(net1098),
    .B2(net786),
    .A2(net1187),
    .A1(\tdc_inst.start_count_debug[14] ));
 sg13g2_nand2_1 _3168_ (.Y(_0061_),
    .A(net1017),
    .B(net787));
 sg13g2_a22oi_1 _3169_ (.Y(_0791_),
    .B1(net1098),
    .B2(net1693),
    .A2(net1187),
    .A1(net786));
 sg13g2_nand2_1 _3170_ (.Y(_0062_),
    .A(net1018),
    .B(_0791_));
 sg13g2_a22oi_1 _3171_ (.Y(_0792_),
    .B1(net1103),
    .B2(net945),
    .A2(net1192),
    .A1(\tdc_inst.start_count_debug[16] ));
 sg13g2_nand2_1 _3172_ (.Y(_0063_),
    .A(net1023),
    .B(net946));
 sg13g2_a22oi_1 _3173_ (.Y(_0793_),
    .B1(net1103),
    .B2(net1605),
    .A2(net1192),
    .A1(net945));
 sg13g2_nand2_1 _3174_ (.Y(_0064_),
    .A(net1023),
    .B(_0793_));
 sg13g2_a22oi_1 _3175_ (.Y(_0794_),
    .B1(net1105),
    .B2(net1533),
    .A2(net1194),
    .A1(\tdc_inst.start_count_debug[18] ));
 sg13g2_nand2_1 _3176_ (.Y(_0065_),
    .A(net1024),
    .B(net1534));
 sg13g2_a22oi_1 _3177_ (.Y(_0795_),
    .B1(net1106),
    .B2(net1375),
    .A2(net1195),
    .A1(\tdc_inst.start_count_debug[19] ));
 sg13g2_nand2_1 _3178_ (.Y(_0066_),
    .A(net1027),
    .B(net1376));
 sg13g2_a22oi_1 _3179_ (.Y(_0796_),
    .B1(net1106),
    .B2(net1515),
    .A2(net1195),
    .A1(net1375));
 sg13g2_nand2_1 _3180_ (.Y(_0067_),
    .A(net1027),
    .B(_0796_));
 sg13g2_a22oi_1 _3181_ (.Y(_0797_),
    .B1(net1108),
    .B2(net1473),
    .A2(net1197),
    .A1(\tdc_inst.start_count_debug[21] ));
 sg13g2_nand2_1 _3182_ (.Y(_0068_),
    .A(net1030),
    .B(net1474));
 sg13g2_a22oi_1 _3183_ (.Y(_0798_),
    .B1(net1108),
    .B2(net1419),
    .A2(net1197),
    .A1(\tdc_inst.start_count_debug[22] ));
 sg13g2_nand2_1 _3184_ (.Y(_0069_),
    .A(net1030),
    .B(net1420));
 sg13g2_a22oi_1 _3185_ (.Y(_0799_),
    .B1(net1108),
    .B2(net1513),
    .A2(net1195),
    .A1(net1419));
 sg13g2_nand2_1 _3186_ (.Y(_0070_),
    .A(net1030),
    .B(_0799_));
 sg13g2_a22oi_1 _3187_ (.Y(_0800_),
    .B1(net1106),
    .B2(net1584),
    .A2(net1195),
    .A1(net1513));
 sg13g2_nand2_1 _3188_ (.Y(_0071_),
    .A(net1027),
    .B(_0800_));
 sg13g2_a22oi_1 _3189_ (.Y(_0801_),
    .B1(net1106),
    .B2(net612),
    .A2(net1195),
    .A1(\tdc_inst.start_count_debug[25] ));
 sg13g2_nand2_1 _3190_ (.Y(_0072_),
    .A(net1027),
    .B(net613));
 sg13g2_a22oi_1 _3191_ (.Y(_0802_),
    .B1(net1106),
    .B2(net692),
    .A2(net1197),
    .A1(net612));
 sg13g2_nand2_1 _3192_ (.Y(_0073_),
    .A(net1027),
    .B(_0802_));
 sg13g2_a22oi_1 _3193_ (.Y(_0803_),
    .B1(net1106),
    .B2(net1535),
    .A2(net1195),
    .A1(net692));
 sg13g2_nand2_1 _3194_ (.Y(_0074_),
    .A(net1027),
    .B(_0803_));
 sg13g2_a22oi_1 _3195_ (.Y(_0804_),
    .B1(net1106),
    .B2(net798),
    .A2(net1195),
    .A1(\tdc_inst.start_count_debug[28] ));
 sg13g2_nand2_1 _3196_ (.Y(_0075_),
    .A(net1029),
    .B(net799));
 sg13g2_a22oi_1 _3197_ (.Y(_0805_),
    .B1(net1106),
    .B2(net1670),
    .A2(net1195),
    .A1(net798));
 sg13g2_nand2_1 _3198_ (.Y(_0076_),
    .A(net1029),
    .B(_0805_));
 sg13g2_a22oi_1 _3199_ (.Y(_0806_),
    .B1(net1103),
    .B2(net745),
    .A2(net1192),
    .A1(\tdc_inst.start_count_debug[30] ));
 sg13g2_nand2_1 _3200_ (.Y(_0077_),
    .A(net1027),
    .B(net746));
 sg13g2_a22oi_1 _3201_ (.Y(_0807_),
    .B1(net1103),
    .B2(net1491),
    .A2(net1192),
    .A1(net745));
 sg13g2_nand2_1 _3202_ (.Y(_0078_),
    .A(net1027),
    .B(_0807_));
 sg13g2_a22oi_1 _3203_ (.Y(_0808_),
    .B1(net1103),
    .B2(net941),
    .A2(net1192),
    .A1(\tdc_inst.start_count_debug[32] ));
 sg13g2_nand2_1 _3204_ (.Y(_0079_),
    .A(net1024),
    .B(net942));
 sg13g2_a22oi_1 _3205_ (.Y(_0809_),
    .B1(net1105),
    .B2(net1502),
    .A2(net1194),
    .A1(net941));
 sg13g2_nand2_1 _3206_ (.Y(_0080_),
    .A(net1024),
    .B(_0809_));
 sg13g2_a22oi_1 _3207_ (.Y(_0810_),
    .B1(net1089),
    .B2(net1399),
    .A2(net1178),
    .A1(\tdc_inst.start_count_debug[34] ));
 sg13g2_nand2_1 _3208_ (.Y(_0081_),
    .A(net1024),
    .B(net1400));
 sg13g2_a22oi_1 _3209_ (.Y(_0811_),
    .B1(net1089),
    .B2(net1597),
    .A2(net1178),
    .A1(net1399));
 sg13g2_nand2_1 _3210_ (.Y(_0082_),
    .A(net1024),
    .B(_0811_));
 sg13g2_a22oi_1 _3211_ (.Y(_0812_),
    .B1(net1089),
    .B2(net1701),
    .A2(net1178),
    .A1(net1597));
 sg13g2_nand2_1 _3212_ (.Y(_0083_),
    .A(net1023),
    .B(_0812_));
 sg13g2_a22oi_1 _3213_ (.Y(_0813_),
    .B1(net1099),
    .B2(net628),
    .A2(net1188),
    .A1(\tdc_inst.start_count_debug[37] ));
 sg13g2_nand2_1 _3214_ (.Y(_0084_),
    .A(net1023),
    .B(net629));
 sg13g2_a22oi_1 _3215_ (.Y(_0814_),
    .B1(net1098),
    .B2(net1721),
    .A2(net1187),
    .A1(net628));
 sg13g2_nand2_1 _3216_ (.Y(_0085_),
    .A(net1018),
    .B(_0814_));
 sg13g2_a22oi_1 _3217_ (.Y(_0815_),
    .B1(net1099),
    .B2(net764),
    .A2(net1188),
    .A1(\tdc_inst.start_count_debug[39] ));
 sg13g2_nand2_1 _3218_ (.Y(_0086_),
    .A(net1018),
    .B(net765));
 sg13g2_a22oi_1 _3219_ (.Y(_0816_),
    .B1(net1099),
    .B2(net1390),
    .A2(net1188),
    .A1(net764));
 sg13g2_nand2_1 _3220_ (.Y(_0087_),
    .A(net1018),
    .B(_0816_));
 sg13g2_a22oi_1 _3221_ (.Y(_0817_),
    .B1(net1098),
    .B2(net1411),
    .A2(net1187),
    .A1(net1390));
 sg13g2_nand2_1 _3222_ (.Y(_0088_),
    .A(net1017),
    .B(_0817_));
 sg13g2_a22oi_1 _3223_ (.Y(_0818_),
    .B1(net1098),
    .B2(net1452),
    .A2(net1187),
    .A1(net1411));
 sg13g2_nand2_1 _3224_ (.Y(_0089_),
    .A(net1019),
    .B(_0818_));
 sg13g2_a22oi_1 _3225_ (.Y(_0819_),
    .B1(net1098),
    .B2(net1681),
    .A2(net1187),
    .A1(net1452));
 sg13g2_nand2_1 _3226_ (.Y(_0090_),
    .A(net1023),
    .B(_0819_));
 sg13g2_a22oi_1 _3227_ (.Y(_0820_),
    .B1(net1103),
    .B2(net951),
    .A2(net1192),
    .A1(\tdc_inst.start_count_debug[44] ));
 sg13g2_nand2_1 _3228_ (.Y(_0091_),
    .A(net1023),
    .B(net952));
 sg13g2_a22oi_1 _3229_ (.Y(_0821_),
    .B1(net1103),
    .B2(net1397),
    .A2(net1192),
    .A1(net951));
 sg13g2_nand2_1 _3230_ (.Y(_0092_),
    .A(net1023),
    .B(_0821_));
 sg13g2_a22oi_1 _3231_ (.Y(_0822_),
    .B1(net1103),
    .B2(net1642),
    .A2(net1192),
    .A1(net1397));
 sg13g2_nand2_1 _3232_ (.Y(_0093_),
    .A(net1023),
    .B(_0822_));
 sg13g2_a22oi_1 _3233_ (.Y(_0823_),
    .B1(net1105),
    .B2(net639),
    .A2(net1194),
    .A1(\tdc_inst.start_count_debug[47] ));
 sg13g2_nand2_1 _3234_ (.Y(_0094_),
    .A(net1025),
    .B(net640));
 sg13g2_a22oi_1 _3235_ (.Y(_0824_),
    .B1(net1104),
    .B2(net1488),
    .A2(net1193),
    .A1(net639));
 sg13g2_nand2_1 _3236_ (.Y(_0095_),
    .A(net1025),
    .B(_0824_));
 sg13g2_a22oi_1 _3237_ (.Y(_0825_),
    .B1(net1105),
    .B2(net1604),
    .A2(net1194),
    .A1(net1488));
 sg13g2_nand2_1 _3238_ (.Y(_0096_),
    .A(net1025),
    .B(_0825_));
 sg13g2_a22oi_1 _3239_ (.Y(_0826_),
    .B1(net1104),
    .B2(net1443),
    .A2(net1193),
    .A1(\tdc_inst.start_count_debug[50] ));
 sg13g2_nand2_1 _3240_ (.Y(_0097_),
    .A(net1029),
    .B(net1444));
 sg13g2_a22oi_1 _3241_ (.Y(_0827_),
    .B1(net1104),
    .B2(net947),
    .A2(net1193),
    .A1(\tdc_inst.start_count_debug[51] ));
 sg13g2_nand2_1 _3242_ (.Y(_0098_),
    .A(net1029),
    .B(net948));
 sg13g2_a22oi_1 _3243_ (.Y(_0828_),
    .B1(net1104),
    .B2(net1677),
    .A2(net1193),
    .A1(net947));
 sg13g2_nand2_1 _3244_ (.Y(_0099_),
    .A(net1029),
    .B(_0828_));
 sg13g2_a22oi_1 _3245_ (.Y(_0829_),
    .B1(net1111),
    .B2(net1264),
    .A2(net1200),
    .A1(\tdc_inst.start_count_debug[53] ));
 sg13g2_nand2_1 _3246_ (.Y(_0100_),
    .A(net1035),
    .B(net1265));
 sg13g2_a22oi_1 _3247_ (.Y(_0830_),
    .B1(net1111),
    .B2(net1730),
    .A2(net1200),
    .A1(net1264));
 sg13g2_nand2_1 _3248_ (.Y(_0101_),
    .A(net1035),
    .B(_0830_));
 sg13g2_a22oi_1 _3249_ (.Y(_0831_),
    .B1(net1111),
    .B2(net887),
    .A2(net1200),
    .A1(\tdc_inst.start_count_debug[55] ));
 sg13g2_nand2_1 _3250_ (.Y(_0102_),
    .A(net1035),
    .B(net888));
 sg13g2_a22oi_1 _3251_ (.Y(_0832_),
    .B1(net1111),
    .B2(net594),
    .A2(net1200),
    .A1(\tdc_inst.start_count_debug[56] ));
 sg13g2_nand2_1 _3252_ (.Y(_0103_),
    .A(net1035),
    .B(net595));
 sg13g2_a22oi_1 _3253_ (.Y(_0833_),
    .B1(net1107),
    .B2(net783),
    .A2(net1196),
    .A1(net594));
 sg13g2_nand2_1 _3254_ (.Y(_0104_),
    .A(net1036),
    .B(_0833_));
 sg13g2_a22oi_1 _3255_ (.Y(_0834_),
    .B1(net1107),
    .B2(net1389),
    .A2(net1196),
    .A1(net783));
 sg13g2_nand2_1 _3256_ (.Y(_0105_),
    .A(net1029),
    .B(_0834_));
 sg13g2_a22oi_1 _3257_ (.Y(_0835_),
    .B1(net1107),
    .B2(net839),
    .A2(net1196),
    .A1(\tdc_inst.start_count_debug[59] ));
 sg13g2_nand2_1 _3258_ (.Y(_0106_),
    .A(net1028),
    .B(net840));
 sg13g2_a22oi_1 _3259_ (.Y(_0836_),
    .B1(net1107),
    .B2(net1340),
    .A2(net1196),
    .A1(net839));
 sg13g2_nand2_1 _3260_ (.Y(_0107_),
    .A(net1028),
    .B(_0836_));
 sg13g2_a22oi_1 _3261_ (.Y(_0837_),
    .B1(net1107),
    .B2(net823),
    .A2(net1196),
    .A1(\tdc_inst.start_count_debug[61] ));
 sg13g2_nand2_1 _3262_ (.Y(_0108_),
    .A(net1028),
    .B(net824));
 sg13g2_a22oi_1 _3263_ (.Y(_0838_),
    .B1(net1107),
    .B2(net768),
    .A2(net1196),
    .A1(\tdc_inst.start_count_debug[62] ));
 sg13g2_nand2_1 _3264_ (.Y(_0109_),
    .A(net1028),
    .B(net769));
 sg13g2_a22oi_1 _3265_ (.Y(_0839_),
    .B1(net1107),
    .B2(net1476),
    .A2(net1197),
    .A1(net768));
 sg13g2_nand2_1 _3266_ (.Y(_0110_),
    .A(net1028),
    .B(_0839_));
 sg13g2_a22oi_1 _3267_ (.Y(_0840_),
    .B1(net1108),
    .B2(net1279),
    .A2(net1196),
    .A1(\tdc_inst.start_count_debug[64] ));
 sg13g2_nand2_1 _3268_ (.Y(_0111_),
    .A(net1028),
    .B(net1280));
 sg13g2_a22oi_1 _3269_ (.Y(_0841_),
    .B1(net1108),
    .B2(net1408),
    .A2(net1197),
    .A1(net1279));
 sg13g2_nand2_1 _3270_ (.Y(_0112_),
    .A(net1028),
    .B(_0841_));
 sg13g2_a22oi_1 _3271_ (.Y(_0842_),
    .B1(net1107),
    .B2(net1716),
    .A2(net1196),
    .A1(net1408));
 sg13g2_nand2_1 _3272_ (.Y(_0113_),
    .A(net1028),
    .B(_0842_));
 sg13g2_a22oi_1 _3273_ (.Y(_0843_),
    .B1(net1112),
    .B2(net1358),
    .A2(net1201),
    .A1(\tdc_inst.start_count_debug[67] ));
 sg13g2_nand2_1 _3274_ (.Y(_0114_),
    .A(net1036),
    .B(net1359));
 sg13g2_a22oi_1 _3275_ (.Y(_0844_),
    .B1(net1112),
    .B2(net802),
    .A2(net1201),
    .A1(\tdc_inst.start_count_debug[68] ));
 sg13g2_nand2_1 _3276_ (.Y(_0115_),
    .A(net1036),
    .B(net803));
 sg13g2_a22oi_1 _3277_ (.Y(_0845_),
    .B1(net1112),
    .B2(net784),
    .A2(net1201),
    .A1(\tdc_inst.start_count_debug[69] ));
 sg13g2_nand2_1 _3278_ (.Y(_0116_),
    .A(net1036),
    .B(net785));
 sg13g2_a22oi_1 _3279_ (.Y(_0846_),
    .B1(net1111),
    .B2(net1679),
    .A2(net1200),
    .A1(net784));
 sg13g2_nand2_1 _3280_ (.Y(_0117_),
    .A(net1036),
    .B(_0846_));
 sg13g2_a22oi_1 _3281_ (.Y(_0847_),
    .B1(net1112),
    .B2(net1293),
    .A2(net1201),
    .A1(\tdc_inst.start_count_debug[71] ));
 sg13g2_nand2_1 _3282_ (.Y(_0118_),
    .A(net1036),
    .B(net1294));
 sg13g2_a22oi_1 _3283_ (.Y(_0848_),
    .B1(net1112),
    .B2(net917),
    .A2(net1201),
    .A1(\tdc_inst.start_count_debug[72] ));
 sg13g2_nand2_1 _3284_ (.Y(_0119_),
    .A(net1036),
    .B(net918));
 sg13g2_a22oi_1 _3285_ (.Y(_0849_),
    .B1(net1114),
    .B2(net1278),
    .A2(net1203),
    .A1(net917));
 sg13g2_nand2_1 _3286_ (.Y(_0120_),
    .A(net1037),
    .B(_0849_));
 sg13g2_a22oi_1 _3287_ (.Y(_0850_),
    .B1(net1114),
    .B2(net652),
    .A2(net1203),
    .A1(\tdc_inst.start_count_debug[74] ));
 sg13g2_nand2_1 _3288_ (.Y(_0121_),
    .A(net1037),
    .B(net653));
 sg13g2_a22oi_1 _3289_ (.Y(_0851_),
    .B1(net1114),
    .B2(net1579),
    .A2(net1202),
    .A1(net652));
 sg13g2_nand2_1 _3290_ (.Y(_0122_),
    .A(net1037),
    .B(_0851_));
 sg13g2_a22oi_1 _3291_ (.Y(_0852_),
    .B1(net1114),
    .B2(net1345),
    .A2(net1203),
    .A1(\tdc_inst.start_count_debug[76] ));
 sg13g2_nand2_1 _3292_ (.Y(_0123_),
    .A(net1037),
    .B(net1346));
 sg13g2_a22oi_1 _3293_ (.Y(_0853_),
    .B1(net1113),
    .B2(net1396),
    .A2(net1203),
    .A1(net1345));
 sg13g2_nand2_1 _3294_ (.Y(_0124_),
    .A(net1038),
    .B(_0853_));
 sg13g2_a22oi_1 _3295_ (.Y(_0854_),
    .B1(net1114),
    .B2(net1496),
    .A2(net1203),
    .A1(net1396));
 sg13g2_nand2_1 _3296_ (.Y(_0125_),
    .A(net1037),
    .B(_0854_));
 sg13g2_a22oi_1 _3297_ (.Y(_0855_),
    .B1(net1114),
    .B2(net1690),
    .A2(net1203),
    .A1(net1496));
 sg13g2_nand2_1 _3298_ (.Y(_0126_),
    .A(net1038),
    .B(_0855_));
 sg13g2_a22oi_1 _3299_ (.Y(_0856_),
    .B1(net1113),
    .B2(net735),
    .A2(net1202),
    .A1(\tdc_inst.start_count_debug[80] ));
 sg13g2_nand2_1 _3300_ (.Y(_0127_),
    .A(net1038),
    .B(net736));
 sg13g2_a22oi_1 _3301_ (.Y(_0857_),
    .B1(net1109),
    .B2(net563),
    .A2(net1198),
    .A1(\tdc_inst.start_count_debug[81] ));
 sg13g2_nand2_1 _3302_ (.Y(_0128_),
    .A(net1038),
    .B(net564));
 sg13g2_a22oi_1 _3303_ (.Y(_0858_),
    .B1(net1109),
    .B2(net1466),
    .A2(net1198),
    .A1(net563));
 sg13g2_nand2_1 _3304_ (.Y(_0129_),
    .A(net1032),
    .B(_0858_));
 sg13g2_a22oi_1 _3305_ (.Y(_0859_),
    .B1(net1116),
    .B2(net1745),
    .A2(net1205),
    .A1(net1466));
 sg13g2_nand2_1 _3306_ (.Y(_0130_),
    .A(net1032),
    .B(_0859_));
 sg13g2_a22oi_1 _3307_ (.Y(_0860_),
    .B1(net1109),
    .B2(net915),
    .A2(net1198),
    .A1(\tdc_inst.start_count_debug[84] ));
 sg13g2_nand2_1 _3308_ (.Y(_0131_),
    .A(net1032),
    .B(net916));
 sg13g2_a22oi_1 _3309_ (.Y(_0861_),
    .B1(net1109),
    .B2(net1719),
    .A2(net1198),
    .A1(net915));
 sg13g2_nand2_1 _3310_ (.Y(_0132_),
    .A(net1033),
    .B(_0861_));
 sg13g2_a22oi_1 _3311_ (.Y(_0862_),
    .B1(net1109),
    .B2(net1349),
    .A2(net1198),
    .A1(\tdc_inst.start_count_debug[86] ));
 sg13g2_nand2_1 _3312_ (.Y(_0133_),
    .A(net1032),
    .B(net1350));
 sg13g2_a22oi_1 _3313_ (.Y(_0863_),
    .B1(net1116),
    .B2(net1484),
    .A2(net1205),
    .A1(net1349));
 sg13g2_nand2_1 _3314_ (.Y(_0134_),
    .A(net1032),
    .B(_0863_));
 sg13g2_a22oi_1 _3315_ (.Y(_0864_),
    .B1(net1116),
    .B2(net1648),
    .A2(net1198),
    .A1(net1484));
 sg13g2_nand2_1 _3316_ (.Y(_0135_),
    .A(net1032),
    .B(_0864_));
 sg13g2_a22oi_1 _3317_ (.Y(_0865_),
    .B1(net1113),
    .B2(net953),
    .A2(net1202),
    .A1(\tdc_inst.start_count_debug[89] ));
 sg13g2_nand2_1 _3318_ (.Y(_0136_),
    .A(net1038),
    .B(net954));
 sg13g2_a22oi_1 _3319_ (.Y(_0866_),
    .B1(net1113),
    .B2(net1461),
    .A2(net1202),
    .A1(net953));
 sg13g2_nand2_1 _3320_ (.Y(_0137_),
    .A(net1038),
    .B(_0866_));
 sg13g2_a22oi_1 _3321_ (.Y(_0867_),
    .B1(net1113),
    .B2(net680),
    .A2(net1202),
    .A1(\tdc_inst.start_count_debug[91] ));
 sg13g2_nand2_1 _3322_ (.Y(_0138_),
    .A(net1038),
    .B(net681));
 sg13g2_a22oi_1 _3323_ (.Y(_0868_),
    .B1(net1113),
    .B2(net1336),
    .A2(net1202),
    .A1(net680));
 sg13g2_nand2_1 _3324_ (.Y(_0139_),
    .A(net1037),
    .B(_0868_));
 sg13g2_a22oi_1 _3325_ (.Y(_0869_),
    .B1(net1113),
    .B2(net1623),
    .A2(net1202),
    .A1(net1336));
 sg13g2_nand2_1 _3326_ (.Y(_0140_),
    .A(net1037),
    .B(_0869_));
 sg13g2_a22oi_1 _3327_ (.Y(_0870_),
    .B1(net1113),
    .B2(net741),
    .A2(net1202),
    .A1(\tdc_inst.start_count_debug[94] ));
 sg13g2_nand2_1 _3328_ (.Y(_0141_),
    .A(net1037),
    .B(net742));
 sg13g2_a22oi_1 _3329_ (.Y(_0871_),
    .B1(net1111),
    .B2(net1714),
    .A2(net1200),
    .A1(net741));
 sg13g2_nand2_1 _3330_ (.Y(_0142_),
    .A(net1035),
    .B(_0871_));
 sg13g2_a22oi_1 _3331_ (.Y(_0872_),
    .B1(net1111),
    .B2(net771),
    .A2(net1200),
    .A1(\tdc_inst.start_count_debug[96] ));
 sg13g2_nand2_1 _3332_ (.Y(_0143_),
    .A(net1035),
    .B(net772));
 sg13g2_a22oi_1 _3333_ (.Y(_0873_),
    .B1(net1111),
    .B2(net694),
    .A2(net1200),
    .A1(\tdc_inst.start_count_debug[97] ));
 sg13g2_nand2_1 _3334_ (.Y(_0144_),
    .A(net1035),
    .B(net695));
 sg13g2_a22oi_1 _3335_ (.Y(_0874_),
    .B1(net1110),
    .B2(net919),
    .A2(net1199),
    .A1(net694));
 sg13g2_nand2_1 _3336_ (.Y(_0145_),
    .A(net1035),
    .B(_0874_));
 sg13g2_a22oi_1 _3337_ (.Y(_0875_),
    .B1(net1109),
    .B2(net1691),
    .A2(net1205),
    .A1(net919));
 sg13g2_nand2_1 _3338_ (.Y(_0146_),
    .A(net1032),
    .B(_0875_));
 sg13g2_a22oi_1 _3339_ (.Y(_0876_),
    .B1(net1110),
    .B2(net578),
    .A2(net1199),
    .A1(\tdc_inst.start_count_debug[100] ));
 sg13g2_nand2_1 _3340_ (.Y(_0147_),
    .A(net1032),
    .B(net579));
 sg13g2_a22oi_1 _3341_ (.Y(_0877_),
    .B1(net1110),
    .B2(net848),
    .A2(net1199),
    .A1(net578));
 sg13g2_nand2_1 _3342_ (.Y(_0148_),
    .A(net1034),
    .B(_0877_));
 sg13g2_a22oi_1 _3343_ (.Y(_0878_),
    .B1(net1110),
    .B2(net1495),
    .A2(net1199),
    .A1(net848));
 sg13g2_nand2_1 _3344_ (.Y(_0149_),
    .A(net1031),
    .B(_0878_));
 sg13g2_a22oi_1 _3345_ (.Y(_0879_),
    .B1(net1110),
    .B2(net1499),
    .A2(net1199),
    .A1(net1495));
 sg13g2_nand2_1 _3346_ (.Y(_0150_),
    .A(net1034),
    .B(_0879_));
 sg13g2_a22oi_1 _3347_ (.Y(_0880_),
    .B1(net1110),
    .B2(net905),
    .A2(net1199),
    .A1(\tdc_inst.start_count_debug[104] ));
 sg13g2_nand2_1 _3348_ (.Y(_0151_),
    .A(net1031),
    .B(net906));
 sg13g2_a22oi_1 _3349_ (.Y(_0881_),
    .B1(net1110),
    .B2(net1685),
    .A2(net1199),
    .A1(net905));
 sg13g2_nand2_1 _3350_ (.Y(_0152_),
    .A(net1034),
    .B(_0881_));
 sg13g2_a22oi_1 _3351_ (.Y(_0882_),
    .B1(net1104),
    .B2(net1519),
    .A2(net1193),
    .A1(\tdc_inst.start_count_debug[106] ));
 sg13g2_nand2_1 _3352_ (.Y(_0153_),
    .A(net1026),
    .B(net1520));
 sg13g2_a22oi_1 _3353_ (.Y(_0883_),
    .B1(net1104),
    .B2(net1459),
    .A2(net1193),
    .A1(\tdc_inst.start_count_debug[107] ));
 sg13g2_nand2_1 _3354_ (.Y(_0154_),
    .A(net1025),
    .B(net1460));
 sg13g2_a22oi_1 _3355_ (.Y(_0884_),
    .B1(net1104),
    .B2(net1385),
    .A2(net1193),
    .A1(\tdc_inst.start_count_debug[108] ));
 sg13g2_nand2_1 _3356_ (.Y(_0155_),
    .A(net1025),
    .B(net1386));
 sg13g2_a22oi_1 _3357_ (.Y(_0885_),
    .B1(net1104),
    .B2(net1740),
    .A2(net1193),
    .A1(net1385));
 sg13g2_nand2_1 _3358_ (.Y(_0156_),
    .A(net1025),
    .B(_0885_));
 sg13g2_a22oi_1 _3359_ (.Y(_0886_),
    .B1(net1100),
    .B2(net1412),
    .A2(net1189),
    .A1(\tdc_inst.start_count_debug[110] ));
 sg13g2_nand2_1 _3360_ (.Y(_0157_),
    .A(net1025),
    .B(net1413));
 sg13g2_a22oi_1 _3361_ (.Y(_0887_),
    .B1(net1100),
    .B2(net1417),
    .A2(net1189),
    .A1(net1412));
 sg13g2_nand2_1 _3362_ (.Y(_0158_),
    .A(net1020),
    .B(_0887_));
 sg13g2_a22oi_1 _3363_ (.Y(_0888_),
    .B1(net1099),
    .B2(net1531),
    .A2(net1188),
    .A1(net1417));
 sg13g2_nand2_1 _3364_ (.Y(_0159_),
    .A(net1019),
    .B(_0888_));
 sg13g2_a22oi_1 _3365_ (.Y(_0889_),
    .B1(net1100),
    .B2(net1321),
    .A2(net1189),
    .A1(\tdc_inst.start_count_debug[113] ));
 sg13g2_nand2_1 _3366_ (.Y(_0160_),
    .A(net1025),
    .B(net1322));
 sg13g2_a22oi_1 _3367_ (.Y(_0890_),
    .B1(net1101),
    .B2(net600),
    .A2(net1190),
    .A1(\tdc_inst.start_count_debug[114] ));
 sg13g2_nand2_1 _3368_ (.Y(_0161_),
    .A(net1031),
    .B(net601));
 sg13g2_a22oi_1 _3369_ (.Y(_0891_),
    .B1(net1101),
    .B2(net1733),
    .A2(net1190),
    .A1(net600));
 sg13g2_nand2_1 _3370_ (.Y(_0162_),
    .A(net1031),
    .B(_0891_));
 sg13g2_a22oi_1 _3371_ (.Y(_0892_),
    .B1(net1101),
    .B2(net1453),
    .A2(net1190),
    .A1(\tdc_inst.start_count_debug[116] ));
 sg13g2_nand2_1 _3372_ (.Y(_0163_),
    .A(net1031),
    .B(net1454));
 sg13g2_a22oi_1 _3373_ (.Y(_0893_),
    .B1(net1101),
    .B2(net633),
    .A2(net1190),
    .A1(\tdc_inst.start_count_debug[117] ));
 sg13g2_nand2_1 _3374_ (.Y(_0164_),
    .A(net1031),
    .B(net634));
 sg13g2_a22oi_1 _3375_ (.Y(_0894_),
    .B1(net1101),
    .B2(net1743),
    .A2(net1190),
    .A1(net633));
 sg13g2_nand2_1 _3376_ (.Y(_0165_),
    .A(net1031),
    .B(_0894_));
 sg13g2_a22oi_1 _3377_ (.Y(_0895_),
    .B1(net1109),
    .B2(net568),
    .A2(net1198),
    .A1(\tdc_inst.start_count_debug[119] ));
 sg13g2_nand2_1 _3378_ (.Y(_0166_),
    .A(net1031),
    .B(net569));
 sg13g2_a22oi_1 _3379_ (.Y(_0896_),
    .B1(net1109),
    .B2(net1734),
    .A2(net1198),
    .A1(net568));
 sg13g2_nand2_1 _3380_ (.Y(_0167_),
    .A(net1033),
    .B(_0896_));
 sg13g2_a22oi_1 _3381_ (.Y(_0897_),
    .B1(net1102),
    .B2(net1556),
    .A2(net1191),
    .A1(\tdc_inst.start_count_debug[121] ));
 sg13g2_nand2_1 _3382_ (.Y(_0168_),
    .A(net1033),
    .B(net1557));
 sg13g2_a22oi_1 _3383_ (.Y(_0898_),
    .B1(net1102),
    .B2(net1671),
    .A2(net1191),
    .A1(net1556));
 sg13g2_nand2_1 _3384_ (.Y(_0169_),
    .A(net1033),
    .B(_0898_));
 sg13g2_a22oi_1 _3385_ (.Y(_0899_),
    .B1(net1102),
    .B2(net760),
    .A2(net1191),
    .A1(\tdc_inst.start_count_debug[123] ));
 sg13g2_nand2_1 _3386_ (.Y(_0170_),
    .A(net1033),
    .B(net761));
 sg13g2_a22oi_1 _3387_ (.Y(_0900_),
    .B1(net1102),
    .B2(net832),
    .A2(net1191),
    .A1(net760));
 sg13g2_nand2_1 _3388_ (.Y(_0171_),
    .A(net1022),
    .B(_0900_));
 sg13g2_a22oi_1 _3389_ (.Y(_0901_),
    .B1(net1102),
    .B2(net1392),
    .A2(net1191),
    .A1(net832));
 sg13g2_nand2_1 _3390_ (.Y(_0172_),
    .A(net1022),
    .B(_0901_));
 sg13g2_a22oi_1 _3391_ (.Y(_0902_),
    .B1(net1102),
    .B2(net790),
    .A2(net1191),
    .A1(\tdc_inst.start_count_debug[126] ));
 sg13g2_nand2_1 _3392_ (.Y(_0173_),
    .A(net1022),
    .B(net791));
 sg13g2_a22oi_1 _3393_ (.Y(_0903_),
    .B1(net1102),
    .B2(net1479),
    .A2(net1191),
    .A1(net790));
 sg13g2_nand2_1 _3394_ (.Y(_0174_),
    .A(net1022),
    .B(_0903_));
 sg13g2_a22oi_1 _3395_ (.Y(_0904_),
    .B1(net1102),
    .B2(net1433),
    .A2(net1191),
    .A1(\tdc_inst.start_count_debug[128] ));
 sg13g2_nand2_1 _3396_ (.Y(_0175_),
    .A(net1040),
    .B(net1434));
 sg13g2_a22oi_1 _3397_ (.Y(_0905_),
    .B1(net1101),
    .B2(net1403),
    .A2(net1190),
    .A1(\tdc_inst.start_count_debug[129] ));
 sg13g2_nand2_1 _3398_ (.Y(_0176_),
    .A(net1022),
    .B(net1404));
 sg13g2_a22oi_1 _3399_ (.Y(_0906_),
    .B1(net1101),
    .B2(net1647),
    .A2(net1190),
    .A1(net1403));
 sg13g2_nand2_1 _3400_ (.Y(_0177_),
    .A(net1022),
    .B(_0906_));
 sg13g2_a22oi_1 _3401_ (.Y(_0907_),
    .B1(net1101),
    .B2(net1682),
    .A2(net1190),
    .A1(net1647));
 sg13g2_nand2_1 _3402_ (.Y(_0178_),
    .A(net1022),
    .B(_0907_));
 sg13g2_a22oi_1 _3403_ (.Y(_0908_),
    .B1(net1099),
    .B2(net939),
    .A2(net1188),
    .A1(\tdc_inst.start_count_debug[132] ));
 sg13g2_nand2_1 _3404_ (.Y(_0179_),
    .A(net1019),
    .B(net940));
 sg13g2_a22oi_1 _3405_ (.Y(_0909_),
    .B1(net1099),
    .B2(net856),
    .A2(net1188),
    .A1(\tdc_inst.start_count_debug[133] ));
 sg13g2_nand2_1 _3406_ (.Y(_0180_),
    .A(net1019),
    .B(net857));
 sg13g2_a22oi_1 _3407_ (.Y(_0910_),
    .B1(net1099),
    .B2(net1514),
    .A2(net1188),
    .A1(net856));
 sg13g2_nand2_1 _3408_ (.Y(_0181_),
    .A(net1019),
    .B(_0910_));
 sg13g2_a22oi_1 _3409_ (.Y(_0911_),
    .B1(net1097),
    .B2(net925),
    .A2(net1186),
    .A1(\tdc_inst.start_count_debug[135] ));
 sg13g2_nand2_1 _3410_ (.Y(_0182_),
    .A(net1019),
    .B(net926));
 sg13g2_a22oi_1 _3411_ (.Y(_0912_),
    .B1(net1097),
    .B2(net827),
    .A2(net1186),
    .A1(\tdc_inst.start_count_debug[136] ));
 sg13g2_nand2_1 _3412_ (.Y(_0183_),
    .A(net1019),
    .B(net828));
 sg13g2_a22oi_1 _3413_ (.Y(_0913_),
    .B1(net1097),
    .B2(net1323),
    .A2(net1186),
    .A1(net827));
 sg13g2_nand2_1 _3414_ (.Y(_0184_),
    .A(net1016),
    .B(_0913_));
 sg13g2_a22oi_1 _3415_ (.Y(_0914_),
    .B1(net1097),
    .B2(net1431),
    .A2(net1186),
    .A1(net1323));
 sg13g2_nand2_1 _3416_ (.Y(_0185_),
    .A(net1016),
    .B(_0914_));
 sg13g2_a22oi_1 _3417_ (.Y(_0915_),
    .B1(net1097),
    .B2(net1643),
    .A2(net1186),
    .A1(net1431));
 sg13g2_nand2_1 _3418_ (.Y(_0186_),
    .A(net1021),
    .B(_0915_));
 sg13g2_a22oi_1 _3419_ (.Y(_0916_),
    .B1(net1071),
    .B2(net1275),
    .A2(net1159),
    .A1(\tdc_inst.start_count_debug[140] ));
 sg13g2_nand2_1 _3420_ (.Y(_0187_),
    .A(net1021),
    .B(net1276));
 sg13g2_a221oi_1 _3421_ (.B2(net1377),
    .C1(_0774_),
    .B1(net1071),
    .A1(net1275),
    .Y(_0917_),
    .A2(net1159));
 sg13g2_inv_1 _3422_ (.Y(_0188_),
    .A(_0917_));
 sg13g2_xor2_1 _3423_ (.B(\tdc_inst.start_signal_sampling_clock_level ),
    .A(\tdc_inst.stop_signal_sampling_clock_level ),
    .X(_0918_));
 sg13g2_and2_1 _3424_ (.A(_0773_),
    .B(_0918_),
    .X(_0919_));
 sg13g2_nand2_1 _3425_ (.Y(_0920_),
    .A(_0773_),
    .B(_0918_));
 sg13g2_a22oi_1 _3426_ (.Y(_0921_),
    .B1(net1070),
    .B2(net1364),
    .A2(net1160),
    .A1(\tdc_inst.tdc_xor_result[0] ));
 sg13g2_nand2_1 _3427_ (.Y(_0189_),
    .A(net1003),
    .B(net1365));
 sg13g2_a22oi_1 _3428_ (.Y(_0922_),
    .B1(net1070),
    .B2(net1536),
    .A2(net1160),
    .A1(net1364));
 sg13g2_nand2_1 _3429_ (.Y(_0190_),
    .A(net1001),
    .B(_0922_));
 sg13g2_a22oi_1 _3430_ (.Y(_0923_),
    .B1(net1070),
    .B2(net1492),
    .A2(net1160),
    .A1(\tdc_inst.tdc_xor_result[2] ));
 sg13g2_nand2_1 _3431_ (.Y(_0191_),
    .A(net1001),
    .B(net1493));
 sg13g2_a22oi_1 _3432_ (.Y(_0924_),
    .B1(net1070),
    .B2(net1314),
    .A2(net1160),
    .A1(\tdc_inst.tdc_xor_result[3] ));
 sg13g2_nand2_1 _3433_ (.Y(_0192_),
    .A(net1000),
    .B(net1315));
 sg13g2_a22oi_1 _3434_ (.Y(_0925_),
    .B1(net1070),
    .B2(net1628),
    .A2(net1160),
    .A1(net1314));
 sg13g2_nand2_1 _3435_ (.Y(_0193_),
    .A(net1000),
    .B(_0925_));
 sg13g2_a22oi_1 _3436_ (.Y(_0926_),
    .B1(net1070),
    .B2(net1571),
    .A2(net1160),
    .A1(\tdc_inst.tdc_xor_result[5] ));
 sg13g2_nand2_1 _3437_ (.Y(_0194_),
    .A(net1000),
    .B(net1572));
 sg13g2_a22oi_1 _3438_ (.Y(_0927_),
    .B1(net1070),
    .B2(net1268),
    .A2(net1160),
    .A1(\tdc_inst.tdc_xor_result[6] ));
 sg13g2_nand2_1 _3439_ (.Y(_0195_),
    .A(net1000),
    .B(net1269));
 sg13g2_a22oi_1 _3440_ (.Y(_0928_),
    .B1(net1055),
    .B2(net1598),
    .A2(net1145),
    .A1(net1268));
 sg13g2_nand2_1 _3441_ (.Y(_0196_),
    .A(net1000),
    .B(_0928_));
 sg13g2_a22oi_1 _3442_ (.Y(_0929_),
    .B1(net1055),
    .B2(net1308),
    .A2(net1145),
    .A1(\tdc_inst.tdc_xor_result[8] ));
 sg13g2_nand2_1 _3443_ (.Y(_0197_),
    .A(net1000),
    .B(net1309));
 sg13g2_a22oi_1 _3444_ (.Y(_0930_),
    .B1(net1055),
    .B2(net1494),
    .A2(net1145),
    .A1(net1308));
 sg13g2_nand2_1 _3445_ (.Y(_0198_),
    .A(net1000),
    .B(_0930_));
 sg13g2_a22oi_1 _3446_ (.Y(_0931_),
    .B1(net1055),
    .B2(net1298),
    .A2(net1145),
    .A1(\tdc_inst.tdc_xor_result[10] ));
 sg13g2_nand2_1 _3447_ (.Y(_0199_),
    .A(net1000),
    .B(net1299));
 sg13g2_a22oi_1 _3448_ (.Y(_0932_),
    .B1(net1055),
    .B2(net1398),
    .A2(net1145),
    .A1(net1298));
 sg13g2_nand2_1 _3449_ (.Y(_0200_),
    .A(net998),
    .B(_0932_));
 sg13g2_a22oi_1 _3450_ (.Y(_0933_),
    .B1(net1053),
    .B2(net1285),
    .A2(net1143),
    .A1(\tdc_inst.tdc_xor_result[12] ));
 sg13g2_nand2_1 _3451_ (.Y(_0201_),
    .A(net998),
    .B(net1286));
 sg13g2_a22oi_1 _3452_ (.Y(_0934_),
    .B1(net1053),
    .B2(net1577),
    .A2(net1143),
    .A1(net1285));
 sg13g2_nand2_1 _3453_ (.Y(_0202_),
    .A(net998),
    .B(_0934_));
 sg13g2_a22oi_1 _3454_ (.Y(_0935_),
    .B1(net1053),
    .B2(net821),
    .A2(net1143),
    .A1(\tdc_inst.tdc_xor_result[14] ));
 sg13g2_nand2_1 _3455_ (.Y(_0203_),
    .A(net998),
    .B(net822));
 sg13g2_a22oi_1 _3456_ (.Y(_0936_),
    .B1(net1053),
    .B2(net1569),
    .A2(net1143),
    .A1(net821));
 sg13g2_nand2_1 _3457_ (.Y(_0204_),
    .A(net998),
    .B(_0936_));
 sg13g2_a22oi_1 _3458_ (.Y(_0937_),
    .B1(net1053),
    .B2(net622),
    .A2(net1143),
    .A1(\tdc_inst.tdc_xor_result[16] ));
 sg13g2_nand2_1 _3459_ (.Y(_0205_),
    .A(net998),
    .B(net623));
 sg13g2_a22oi_1 _3460_ (.Y(_0938_),
    .B1(net1053),
    .B2(net1680),
    .A2(net1143),
    .A1(net622));
 sg13g2_nand2_1 _3461_ (.Y(_0206_),
    .A(net993),
    .B(_0938_));
 sg13g2_a22oi_1 _3462_ (.Y(_0939_),
    .B1(net1047),
    .B2(net1591),
    .A2(net1137),
    .A1(\tdc_inst.tdc_xor_result[18] ));
 sg13g2_nand2_1 _3463_ (.Y(_0207_),
    .A(net993),
    .B(net1592));
 sg13g2_a22oi_1 _3464_ (.Y(_0940_),
    .B1(net1047),
    .B2(net702),
    .A2(net1137),
    .A1(\tdc_inst.tdc_xor_result[19] ));
 sg13g2_nand2_1 _3465_ (.Y(_0208_),
    .A(net993),
    .B(net703));
 sg13g2_a22oi_1 _3466_ (.Y(_0941_),
    .B1(net1047),
    .B2(net1705),
    .A2(net1137),
    .A1(net702));
 sg13g2_nand2_1 _3467_ (.Y(_0209_),
    .A(net993),
    .B(_0941_));
 sg13g2_a22oi_1 _3468_ (.Y(_0942_),
    .B1(net1047),
    .B2(net1471),
    .A2(net1137),
    .A1(\tdc_inst.tdc_xor_result[21] ));
 sg13g2_nand2_1 _3469_ (.Y(_0210_),
    .A(net993),
    .B(net1472));
 sg13g2_a22oi_1 _3470_ (.Y(_0943_),
    .B1(net1047),
    .B2(net667),
    .A2(net1137),
    .A1(\tdc_inst.tdc_xor_result[22] ));
 sg13g2_nand2_1 _3471_ (.Y(_0211_),
    .A(net993),
    .B(net668));
 sg13g2_a22oi_1 _3472_ (.Y(_0944_),
    .B1(net1047),
    .B2(net1608),
    .A2(net1137),
    .A1(net667));
 sg13g2_nand2_1 _3473_ (.Y(_0212_),
    .A(net993),
    .B(_0944_));
 sg13g2_a22oi_1 _3474_ (.Y(_0945_),
    .B1(net1045),
    .B2(net1529),
    .A2(net1135),
    .A1(\tdc_inst.tdc_xor_result[24] ));
 sg13g2_nand2_1 _3475_ (.Y(_0213_),
    .A(net991),
    .B(net1530));
 sg13g2_a22oi_1 _3476_ (.Y(_0946_),
    .B1(net1045),
    .B2(net1272),
    .A2(net1135),
    .A1(\tdc_inst.tdc_xor_result[25] ));
 sg13g2_nand2_1 _3477_ (.Y(_0214_),
    .A(net991),
    .B(net1273));
 sg13g2_a22oi_1 _3478_ (.Y(_0947_),
    .B1(net1045),
    .B2(net866),
    .A2(net1135),
    .A1(\tdc_inst.tdc_xor_result[26] ));
 sg13g2_nand2_1 _3479_ (.Y(_0215_),
    .A(net991),
    .B(net867));
 sg13g2_a22oi_1 _3480_ (.Y(_0948_),
    .B1(net1045),
    .B2(net673),
    .A2(net1135),
    .A1(\tdc_inst.tdc_xor_result[27] ));
 sg13g2_nand2_1 _3481_ (.Y(_0216_),
    .A(net991),
    .B(net674));
 sg13g2_a22oi_1 _3482_ (.Y(_0949_),
    .B1(net1045),
    .B2(net904),
    .A2(net1135),
    .A1(net673));
 sg13g2_nand2_1 _3483_ (.Y(_0217_),
    .A(net991),
    .B(_0949_));
 sg13g2_a22oi_1 _3484_ (.Y(_0950_),
    .B1(net1045),
    .B2(net1609),
    .A2(net1135),
    .A1(net904));
 sg13g2_nand2_1 _3485_ (.Y(_0218_),
    .A(net991),
    .B(_0950_));
 sg13g2_a22oi_1 _3486_ (.Y(_0951_),
    .B1(net1045),
    .B2(net1644),
    .A2(net1135),
    .A1(net1609));
 sg13g2_nand2_1 _3487_ (.Y(_0219_),
    .A(net991),
    .B(_0951_));
 sg13g2_a22oi_1 _3488_ (.Y(_0952_),
    .B1(net1045),
    .B2(net829),
    .A2(net1135),
    .A1(\tdc_inst.tdc_xor_result[31] ));
 sg13g2_nand2_1 _3489_ (.Y(_0220_),
    .A(net992),
    .B(net830));
 sg13g2_a22oi_1 _3490_ (.Y(_0953_),
    .B1(net1046),
    .B2(net911),
    .A2(net1136),
    .A1(net829));
 sg13g2_nand2_1 _3491_ (.Y(_0221_),
    .A(net992),
    .B(_0953_));
 sg13g2_a22oi_1 _3492_ (.Y(_0954_),
    .B1(net1046),
    .B2(net1633),
    .A2(net1136),
    .A1(net911));
 sg13g2_nand2_1 _3493_ (.Y(_0222_),
    .A(net991),
    .B(_0954_));
 sg13g2_a22oi_1 _3494_ (.Y(_0955_),
    .B1(net1050),
    .B2(net1618),
    .A2(net1140),
    .A1(\tdc_inst.tdc_xor_result[34] ));
 sg13g2_nand2_1 _3495_ (.Y(_0223_),
    .A(net995),
    .B(net1619));
 sg13g2_a22oi_1 _3496_ (.Y(_0956_),
    .B1(net1050),
    .B2(net885),
    .A2(net1140),
    .A1(\tdc_inst.tdc_xor_result[35] ));
 sg13g2_nand2_1 _3497_ (.Y(_0224_),
    .A(net995),
    .B(net886));
 sg13g2_a22oi_1 _3498_ (.Y(_0957_),
    .B1(net1050),
    .B2(net1637),
    .A2(net1140),
    .A1(net885));
 sg13g2_nand2_1 _3499_ (.Y(_0225_),
    .A(net995),
    .B(_0957_));
 sg13g2_a22oi_1 _3500_ (.Y(_0958_),
    .B1(net1050),
    .B2(net1505),
    .A2(net1140),
    .A1(\tdc_inst.tdc_xor_result[37] ));
 sg13g2_nand2_1 _3501_ (.Y(_0226_),
    .A(net995),
    .B(net1506));
 sg13g2_a22oi_1 _3502_ (.Y(_0959_),
    .B1(net1051),
    .B2(net899),
    .A2(net1141),
    .A1(\tdc_inst.tdc_xor_result[38] ));
 sg13g2_nand2_1 _3503_ (.Y(_0227_),
    .A(net1004),
    .B(net900));
 sg13g2_a22oi_1 _3504_ (.Y(_0960_),
    .B1(net1059),
    .B2(net1501),
    .A2(net1148),
    .A1(net899));
 sg13g2_nand2_1 _3505_ (.Y(_0228_),
    .A(net1004),
    .B(_0960_));
 sg13g2_a22oi_1 _3506_ (.Y(_0961_),
    .B1(net1059),
    .B2(net1594),
    .A2(net1148),
    .A1(net1501));
 sg13g2_nand2_1 _3507_ (.Y(_0229_),
    .A(net1004),
    .B(_0961_));
 sg13g2_a22oi_1 _3508_ (.Y(_0962_),
    .B1(net1059),
    .B2(net1668),
    .A2(net1148),
    .A1(net1594));
 sg13g2_nand2_1 _3509_ (.Y(_0230_),
    .A(net1004),
    .B(_0962_));
 sg13g2_a22oi_1 _3510_ (.Y(_0963_),
    .B1(net1059),
    .B2(net1327),
    .A2(net1148),
    .A1(\tdc_inst.tdc_xor_result[42] ));
 sg13g2_nand2_1 _3511_ (.Y(_0231_),
    .A(net1007),
    .B(net1328));
 sg13g2_a22oi_1 _3512_ (.Y(_0964_),
    .B1(net1059),
    .B2(net1646),
    .A2(net1148),
    .A1(net1327));
 sg13g2_nand2_1 _3513_ (.Y(_0232_),
    .A(net1007),
    .B(_0964_));
 sg13g2_a22oi_1 _3514_ (.Y(_0965_),
    .B1(net1063),
    .B2(net1729),
    .A2(net1152),
    .A1(net1646));
 sg13g2_nand2_1 _3515_ (.Y(_0233_),
    .A(net1007),
    .B(_0965_));
 sg13g2_a22oi_1 _3516_ (.Y(_0966_),
    .B1(net1063),
    .B2(net1312),
    .A2(net1152),
    .A1(\tdc_inst.tdc_xor_result[45] ));
 sg13g2_nand2_1 _3517_ (.Y(_0234_),
    .A(net1007),
    .B(net1313));
 sg13g2_a22oi_1 _3518_ (.Y(_0967_),
    .B1(net1063),
    .B2(net1430),
    .A2(net1152),
    .A1(net1312));
 sg13g2_nand2_1 _3519_ (.Y(_0235_),
    .A(net1007),
    .B(_0967_));
 sg13g2_a22oi_1 _3520_ (.Y(_0968_),
    .B1(net1063),
    .B2(net1566),
    .A2(net1152),
    .A1(net1430));
 sg13g2_nand2_1 _3521_ (.Y(_0236_),
    .A(net1008),
    .B(_0968_));
 sg13g2_a22oi_1 _3522_ (.Y(_0969_),
    .B1(net1063),
    .B2(net775),
    .A2(net1152),
    .A1(\tdc_inst.tdc_xor_result[48] ));
 sg13g2_nand2_1 _3523_ (.Y(_0237_),
    .A(net1008),
    .B(net776));
 sg13g2_a22oi_1 _3524_ (.Y(_0970_),
    .B1(net1062),
    .B2(net637),
    .A2(net1151),
    .A1(\tdc_inst.tdc_xor_result[49] ));
 sg13g2_nand2_1 _3525_ (.Y(_0238_),
    .A(net1009),
    .B(net638));
 sg13g2_a22oi_1 _3526_ (.Y(_0971_),
    .B1(net1062),
    .B2(net1655),
    .A2(net1151),
    .A1(net637));
 sg13g2_nand2_1 _3527_ (.Y(_0239_),
    .A(net1009),
    .B(_0971_));
 sg13g2_a22oi_1 _3528_ (.Y(_0972_),
    .B1(net1060),
    .B2(net688),
    .A2(net1149),
    .A1(\tdc_inst.tdc_xor_result[51] ));
 sg13g2_nand2_1 _3529_ (.Y(_0240_),
    .A(net1009),
    .B(net689));
 sg13g2_a22oi_1 _3530_ (.Y(_0973_),
    .B1(net1060),
    .B2(net1316),
    .A2(net1149),
    .A1(net688));
 sg13g2_nand2_1 _3531_ (.Y(_0241_),
    .A(net1009),
    .B(_0973_));
 sg13g2_a22oi_1 _3532_ (.Y(_0974_),
    .B1(net1060),
    .B2(net1449),
    .A2(net1149),
    .A1(net1316));
 sg13g2_nand2_1 _3533_ (.Y(_0242_),
    .A(net1005),
    .B(_0974_));
 sg13g2_a22oi_1 _3534_ (.Y(_0975_),
    .B1(net1060),
    .B2(net1324),
    .A2(net1149),
    .A1(\tdc_inst.tdc_xor_result[54] ));
 sg13g2_nand2_1 _3535_ (.Y(_0243_),
    .A(net1005),
    .B(net1325));
 sg13g2_a22oi_1 _3536_ (.Y(_0976_),
    .B1(net1060),
    .B2(net1482),
    .A2(net1149),
    .A1(net1324));
 sg13g2_nand2_1 _3537_ (.Y(_0244_),
    .A(net1005),
    .B(_0976_));
 sg13g2_a22oi_1 _3538_ (.Y(_0977_),
    .B1(net1052),
    .B2(net907),
    .A2(net1142),
    .A1(\tdc_inst.tdc_xor_result[56] ));
 sg13g2_nand2_1 _3539_ (.Y(_0245_),
    .A(net1005),
    .B(net908));
 sg13g2_a22oi_1 _3540_ (.Y(_0978_),
    .B1(net1052),
    .B2(net868),
    .A2(net1142),
    .A1(\tdc_inst.tdc_xor_result[57] ));
 sg13g2_nand2_1 _3541_ (.Y(_0246_),
    .A(net996),
    .B(net869));
 sg13g2_a22oi_1 _3542_ (.Y(_0979_),
    .B1(net1052),
    .B2(net1573),
    .A2(net1142),
    .A1(net868));
 sg13g2_nand2_1 _3543_ (.Y(_0247_),
    .A(net997),
    .B(_0979_));
 sg13g2_a22oi_1 _3544_ (.Y(_0980_),
    .B1(net1052),
    .B2(net1610),
    .A2(net1142),
    .A1(net1573));
 sg13g2_nand2_1 _3545_ (.Y(_0248_),
    .A(net997),
    .B(_0980_));
 sg13g2_a22oi_1 _3546_ (.Y(_0981_),
    .B1(net1052),
    .B2(net671),
    .A2(net1142),
    .A1(\tdc_inst.tdc_xor_result[60] ));
 sg13g2_nand2_1 _3547_ (.Y(_0249_),
    .A(net997),
    .B(net672));
 sg13g2_a22oi_1 _3548_ (.Y(_0982_),
    .B1(net1052),
    .B2(net1731),
    .A2(net1142),
    .A1(net671));
 sg13g2_nand2_1 _3549_ (.Y(_0250_),
    .A(net1005),
    .B(_0982_));
 sg13g2_a22oi_1 _3550_ (.Y(_0983_),
    .B1(net1060),
    .B2(net1511),
    .A2(net1149),
    .A1(\tdc_inst.tdc_xor_result[62] ));
 sg13g2_nand2_1 _3551_ (.Y(_0251_),
    .A(net1005),
    .B(net1512));
 sg13g2_a22oi_1 _3552_ (.Y(_0984_),
    .B1(net1060),
    .B2(net1659),
    .A2(net1149),
    .A1(net1511));
 sg13g2_nand2_1 _3553_ (.Y(_0252_),
    .A(net1005),
    .B(_0984_));
 sg13g2_a22oi_1 _3554_ (.Y(_0985_),
    .B1(net1061),
    .B2(net1552),
    .A2(net1150),
    .A1(\tdc_inst.tdc_xor_result[64] ));
 sg13g2_nand2_1 _3555_ (.Y(_0253_),
    .A(net1006),
    .B(net1553));
 sg13g2_a22oi_1 _3556_ (.Y(_0986_),
    .B1(net1061),
    .B2(net748),
    .A2(net1150),
    .A1(\tdc_inst.tdc_xor_result[65] ));
 sg13g2_nand2_1 _3557_ (.Y(_0254_),
    .A(net1005),
    .B(net749));
 sg13g2_a22oi_1 _3558_ (.Y(_0987_),
    .B1(net1060),
    .B2(net1586),
    .A2(net1149),
    .A1(net748));
 sg13g2_nand2_1 _3559_ (.Y(_0255_),
    .A(net1009),
    .B(_0987_));
 sg13g2_a22oi_1 _3560_ (.Y(_0988_),
    .B1(net1062),
    .B2(net1517),
    .A2(net1151),
    .A1(\tdc_inst.tdc_xor_result[67] ));
 sg13g2_nand2_1 _3561_ (.Y(_0256_),
    .A(net1009),
    .B(net1518));
 sg13g2_a22oi_1 _3562_ (.Y(_0989_),
    .B1(net1062),
    .B2(net1394),
    .A2(net1151),
    .A1(\tdc_inst.tdc_xor_result[68] ));
 sg13g2_nand2_1 _3563_ (.Y(_0257_),
    .A(net1009),
    .B(net1395));
 sg13g2_a22oi_1 _3564_ (.Y(_0990_),
    .B1(net1066),
    .B2(net806),
    .A2(net1155),
    .A1(\tdc_inst.tdc_xor_result[69] ));
 sg13g2_nand2_1 _3565_ (.Y(_0258_),
    .A(net1010),
    .B(net807));
 sg13g2_a22oi_1 _3566_ (.Y(_0991_),
    .B1(net1066),
    .B2(net1715),
    .A2(net1155),
    .A1(net806));
 sg13g2_nand2_1 _3567_ (.Y(_0259_),
    .A(net1010),
    .B(_0991_));
 sg13g2_a22oi_1 _3568_ (.Y(_0992_),
    .B1(net1062),
    .B2(net642),
    .A2(net1151),
    .A1(\tdc_inst.tdc_xor_result[71] ));
 sg13g2_nand2_1 _3569_ (.Y(_0260_),
    .A(net1010),
    .B(net643));
 sg13g2_a22oi_1 _3570_ (.Y(_0993_),
    .B1(net1062),
    .B2(net1672),
    .A2(net1151),
    .A1(net642));
 sg13g2_nand2_1 _3571_ (.Y(_0261_),
    .A(net1010),
    .B(_0993_));
 sg13g2_a22oi_1 _3572_ (.Y(_0994_),
    .B1(net1062),
    .B2(net716),
    .A2(net1151),
    .A1(\tdc_inst.tdc_xor_result[73] ));
 sg13g2_nand2_1 _3573_ (.Y(_0262_),
    .A(net1010),
    .B(net717));
 sg13g2_a22oi_1 _3574_ (.Y(_0995_),
    .B1(net1062),
    .B2(net1697),
    .A2(net1151),
    .A1(net716));
 sg13g2_nand2_1 _3575_ (.Y(_0263_),
    .A(net1009),
    .B(_0995_));
 sg13g2_a22oi_1 _3576_ (.Y(_0996_),
    .B1(net1064),
    .B2(net1497),
    .A2(net1153),
    .A1(\tdc_inst.tdc_xor_result[75] ));
 sg13g2_nand2_1 _3577_ (.Y(_0264_),
    .A(net1010),
    .B(net1498));
 sg13g2_a22oi_1 _3578_ (.Y(_0997_),
    .B1(net1064),
    .B2(net1507),
    .A2(net1153),
    .A1(net1497));
 sg13g2_nand2_1 _3579_ (.Y(_0265_),
    .A(net1008),
    .B(_0997_));
 sg13g2_a22oi_1 _3580_ (.Y(_0998_),
    .B1(net1063),
    .B2(net664),
    .A2(net1152),
    .A1(\tdc_inst.tdc_xor_result[77] ));
 sg13g2_nand2_1 _3581_ (.Y(_0266_),
    .A(net1008),
    .B(net665));
 sg13g2_a22oi_1 _3582_ (.Y(_0999_),
    .B1(net1063),
    .B2(net1462),
    .A2(net1152),
    .A1(net664));
 sg13g2_nand2_1 _3583_ (.Y(_0267_),
    .A(net1007),
    .B(_0999_));
 sg13g2_a22oi_1 _3584_ (.Y(_1000_),
    .B1(net1063),
    .B2(net1588),
    .A2(net1152),
    .A1(net1462));
 sg13g2_nand2_1 _3585_ (.Y(_0268_),
    .A(net1007),
    .B(_1000_));
 sg13g2_a22oi_1 _3586_ (.Y(_1001_),
    .B1(net1061),
    .B2(net1467),
    .A2(net1150),
    .A1(\tdc_inst.tdc_xor_result[80] ));
 sg13g2_nand2_1 _3587_ (.Y(_0269_),
    .A(net1007),
    .B(net1468));
 sg13g2_a22oi_1 _3588_ (.Y(_1002_),
    .B1(net1061),
    .B2(net635),
    .A2(net1150),
    .A1(\tdc_inst.tdc_xor_result[81] ));
 sg13g2_nand2_1 _3589_ (.Y(_0270_),
    .A(net1006),
    .B(net636));
 sg13g2_a22oi_1 _3590_ (.Y(_1003_),
    .B1(net1061),
    .B2(net1656),
    .A2(net1150),
    .A1(net635));
 sg13g2_nand2_1 _3591_ (.Y(_0271_),
    .A(net1004),
    .B(_1003_));
 sg13g2_a22oi_1 _3592_ (.Y(_1004_),
    .B1(net1059),
    .B2(net1291),
    .A2(net1148),
    .A1(\tdc_inst.tdc_xor_result[83] ));
 sg13g2_nand2_1 _3593_ (.Y(_0272_),
    .A(net1006),
    .B(net1292));
 sg13g2_a22oi_1 _3594_ (.Y(_1005_),
    .B1(net1059),
    .B2(net704),
    .A2(net1148),
    .A1(\tdc_inst.tdc_xor_result[84] ));
 sg13g2_nand2_1 _3595_ (.Y(_0273_),
    .A(net1004),
    .B(net705));
 sg13g2_a22oi_1 _3596_ (.Y(_1006_),
    .B1(net1059),
    .B2(net1667),
    .A2(net1148),
    .A1(net704));
 sg13g2_nand2_1 _3597_ (.Y(_0274_),
    .A(net1004),
    .B(_1006_));
 sg13g2_a22oi_1 _3598_ (.Y(_1007_),
    .B1(net1051),
    .B2(net1599),
    .A2(net1141),
    .A1(\tdc_inst.tdc_xor_result[86] ));
 sg13g2_nand2_1 _3599_ (.Y(_0275_),
    .A(net1004),
    .B(net1600));
 sg13g2_a22oi_1 _3600_ (.Y(_1008_),
    .B1(net1051),
    .B2(net645),
    .A2(net1141),
    .A1(\tdc_inst.tdc_xor_result[87] ));
 sg13g2_nand2_1 _3601_ (.Y(_0276_),
    .A(net997),
    .B(net646));
 sg13g2_a22oi_1 _3602_ (.Y(_1009_),
    .B1(net1051),
    .B2(net1675),
    .A2(net1141),
    .A1(net645));
 sg13g2_nand2_1 _3603_ (.Y(_0277_),
    .A(net997),
    .B(_1009_));
 sg13g2_a22oi_1 _3604_ (.Y(_1010_),
    .B1(net1050),
    .B2(net835),
    .A2(net1140),
    .A1(\tdc_inst.tdc_xor_result[89] ));
 sg13g2_nand2_1 _3605_ (.Y(_0278_),
    .A(net997),
    .B(net836));
 sg13g2_a22oi_1 _3606_ (.Y(_1011_),
    .B1(net1050),
    .B2(net1353),
    .A2(net1140),
    .A1(net835));
 sg13g2_nand2_1 _3607_ (.Y(_0279_),
    .A(net995),
    .B(_1011_));
 sg13g2_a22oi_1 _3608_ (.Y(_1012_),
    .B1(net1050),
    .B2(net650),
    .A2(net1140),
    .A1(\tdc_inst.tdc_xor_result[91] ));
 sg13g2_nand2_1 _3609_ (.Y(_0280_),
    .A(net995),
    .B(net651));
 sg13g2_a22oi_1 _3610_ (.Y(_1013_),
    .B1(net1050),
    .B2(net1277),
    .A2(net1140),
    .A1(net650));
 sg13g2_nand2_1 _3611_ (.Y(_0281_),
    .A(net995),
    .B(_1013_));
 sg13g2_a22oi_1 _3612_ (.Y(_1014_),
    .B1(net1046),
    .B2(net1307),
    .A2(net1136),
    .A1(net1277));
 sg13g2_nand2_1 _3613_ (.Y(_0282_),
    .A(net995),
    .B(_1014_));
 sg13g2_a22oi_1 _3614_ (.Y(_1015_),
    .B1(net1046),
    .B2(net1662),
    .A2(net1136),
    .A1(net1307));
 sg13g2_nand2_1 _3615_ (.Y(_0283_),
    .A(net992),
    .B(_1015_));
 sg13g2_a22oi_1 _3616_ (.Y(_1016_),
    .B1(net1046),
    .B2(net882),
    .A2(net1136),
    .A1(\tdc_inst.tdc_xor_result[95] ));
 sg13g2_nand2_1 _3617_ (.Y(_0284_),
    .A(net992),
    .B(net883));
 sg13g2_a22oi_1 _3618_ (.Y(_1017_),
    .B1(net1046),
    .B2(net1521),
    .A2(net1136),
    .A1(net882));
 sg13g2_nand2_1 _3619_ (.Y(_0285_),
    .A(net992),
    .B(_1017_));
 sg13g2_a22oi_1 _3620_ (.Y(_1018_),
    .B1(net1048),
    .B2(net1585),
    .A2(net1138),
    .A1(net1521));
 sg13g2_nand2_1 _3621_ (.Y(_0286_),
    .A(net992),
    .B(_1018_));
 sg13g2_a22oi_1 _3622_ (.Y(_1019_),
    .B1(net1048),
    .B2(net1485),
    .A2(net1138),
    .A1(\tdc_inst.tdc_xor_result[98] ));
 sg13g2_nand2_1 _3623_ (.Y(_0287_),
    .A(net994),
    .B(net1486));
 sg13g2_a22oi_1 _3624_ (.Y(_1020_),
    .B1(net1048),
    .B2(net1447),
    .A2(net1138),
    .A1(\tdc_inst.tdc_xor_result[99] ));
 sg13g2_nand2_1 _3625_ (.Y(_0288_),
    .A(net994),
    .B(net1448));
 sg13g2_a22oi_1 _3626_ (.Y(_1021_),
    .B1(net1048),
    .B2(net1603),
    .A2(net1138),
    .A1(net1447));
 sg13g2_nand2_1 _3627_ (.Y(_0289_),
    .A(net996),
    .B(_1021_));
 sg13g2_a22oi_1 _3628_ (.Y(_1022_),
    .B1(net1048),
    .B2(net1550),
    .A2(net1138),
    .A1(\tdc_inst.tdc_xor_result[101] ));
 sg13g2_nand2_1 _3629_ (.Y(_0290_),
    .A(net996),
    .B(net1551));
 sg13g2_a22oi_1 _3630_ (.Y(_1023_),
    .B1(net1048),
    .B2(net933),
    .A2(net1137),
    .A1(\tdc_inst.tdc_xor_result[102] ));
 sg13g2_nand2_1 _3631_ (.Y(_0291_),
    .A(net996),
    .B(net934));
 sg13g2_a22oi_1 _3632_ (.Y(_1024_),
    .B1(net1047),
    .B2(net1329),
    .A2(net1137),
    .A1(net933));
 sg13g2_nand2_1 _3633_ (.Y(_0292_),
    .A(net996),
    .B(_1024_));
 sg13g2_a22oi_1 _3634_ (.Y(_1025_),
    .B1(net1047),
    .B2(net1371),
    .A2(net1138),
    .A1(net1329));
 sg13g2_nand2_1 _3635_ (.Y(_0293_),
    .A(net994),
    .B(_1025_));
 sg13g2_a22oi_1 _3636_ (.Y(_1026_),
    .B1(net1054),
    .B2(net686),
    .A2(net1144),
    .A1(\tdc_inst.tdc_xor_result[105] ));
 sg13g2_nand2_1 _3637_ (.Y(_0294_),
    .A(net993),
    .B(net687));
 sg13g2_a22oi_1 _3638_ (.Y(_1027_),
    .B1(net1054),
    .B2(net1589),
    .A2(net1144),
    .A1(net686));
 sg13g2_nand2_1 _3639_ (.Y(_0295_),
    .A(net999),
    .B(_1027_));
 sg13g2_a22oi_1 _3640_ (.Y(_1028_),
    .B1(net1054),
    .B2(net648),
    .A2(net1144),
    .A1(\tdc_inst.tdc_xor_result[107] ));
 sg13g2_nand2_1 _3641_ (.Y(_0296_),
    .A(net999),
    .B(net649));
 sg13g2_a22oi_1 _3642_ (.Y(_1029_),
    .B1(net1054),
    .B2(net1391),
    .A2(net1144),
    .A1(net648));
 sg13g2_nand2_1 _3643_ (.Y(_0297_),
    .A(net999),
    .B(_1029_));
 sg13g2_a22oi_1 _3644_ (.Y(_1030_),
    .B1(net1053),
    .B2(net1401),
    .A2(net1143),
    .A1(net1391));
 sg13g2_nand2_1 _3645_ (.Y(_0298_),
    .A(net999),
    .B(_1030_));
 sg13g2_a22oi_1 _3646_ (.Y(_1031_),
    .B1(net1055),
    .B2(net1367),
    .A2(net1145),
    .A1(\tdc_inst.tdc_xor_result[110] ));
 sg13g2_nand2_1 _3647_ (.Y(_0299_),
    .A(net998),
    .B(net1368));
 sg13g2_a22oi_1 _3648_ (.Y(_1032_),
    .B1(net1058),
    .B2(net1337),
    .A2(net1147),
    .A1(\tdc_inst.tdc_xor_result[111] ));
 sg13g2_nand2_1 _3649_ (.Y(_0300_),
    .A(net1001),
    .B(net1338));
 sg13g2_a22oi_1 _3650_ (.Y(_1033_),
    .B1(net1058),
    .B2(net872),
    .A2(net1147),
    .A1(\tdc_inst.tdc_xor_result[112] ));
 sg13g2_nand2_1 _3651_ (.Y(_0301_),
    .A(net1001),
    .B(net873));
 sg13g2_a22oi_1 _3652_ (.Y(_1034_),
    .B1(net1054),
    .B2(net1676),
    .A2(net1144),
    .A1(net872));
 sg13g2_nand2_1 _3653_ (.Y(_0302_),
    .A(net998),
    .B(_1034_));
 sg13g2_a22oi_1 _3654_ (.Y(_1035_),
    .B1(net1053),
    .B2(net889),
    .A2(net1143),
    .A1(\tdc_inst.tdc_xor_result[114] ));
 sg13g2_nand2_1 _3655_ (.Y(_0303_),
    .A(net1003),
    .B(net890));
 sg13g2_a22oi_1 _3656_ (.Y(_1036_),
    .B1(net1056),
    .B2(net870),
    .A2(net1146),
    .A1(\tdc_inst.tdc_xor_result[115] ));
 sg13g2_nand2_1 _3657_ (.Y(_0304_),
    .A(net1003),
    .B(net871));
 sg13g2_a22oi_1 _3658_ (.Y(_1037_),
    .B1(net1056),
    .B2(net1563),
    .A2(net1146),
    .A1(net870));
 sg13g2_nand2_1 _3659_ (.Y(_0305_),
    .A(net1003),
    .B(_1037_));
 sg13g2_a22oi_1 _3660_ (.Y(_1038_),
    .B1(net1056),
    .B2(net1683),
    .A2(net1146),
    .A1(net1563));
 sg13g2_nand2_1 _3661_ (.Y(_0306_),
    .A(net1003),
    .B(_1038_));
 sg13g2_a22oi_1 _3662_ (.Y(_1039_),
    .B1(net1056),
    .B2(net927),
    .A2(net1146),
    .A1(\tdc_inst.tdc_xor_result[118] ));
 sg13g2_nand2_1 _3663_ (.Y(_0307_),
    .A(net1003),
    .B(net928));
 sg13g2_a22oi_1 _3664_ (.Y(_1040_),
    .B1(net1056),
    .B2(net846),
    .A2(net1146),
    .A1(\tdc_inst.tdc_xor_result[119] ));
 sg13g2_nand2_1 _3665_ (.Y(_0308_),
    .A(net996),
    .B(net847));
 sg13g2_a22oi_1 _3666_ (.Y(_1041_),
    .B1(net1057),
    .B2(net1649),
    .A2(net1147),
    .A1(net846));
 sg13g2_nand2_1 _3667_ (.Y(_0309_),
    .A(net996),
    .B(_1041_));
 sg13g2_a22oi_1 _3668_ (.Y(_1042_),
    .B1(net1057),
    .B2(net598),
    .A2(net1146),
    .A1(\tdc_inst.tdc_xor_result[121] ));
 sg13g2_nand2_1 _3669_ (.Y(_0310_),
    .A(net996),
    .B(net599));
 sg13g2_a22oi_1 _3670_ (.Y(_1043_),
    .B1(net1057),
    .B2(net1344),
    .A2(net1146),
    .A1(net598));
 sg13g2_nand2_1 _3671_ (.Y(_0311_),
    .A(net1014),
    .B(_1043_));
 sg13g2_a22oi_1 _3672_ (.Y(_1044_),
    .B1(net1056),
    .B2(net1319),
    .A2(net1146),
    .A1(\tdc_inst.tdc_xor_result[123] ));
 sg13g2_nand2_1 _3673_ (.Y(_0312_),
    .A(net1014),
    .B(net1320));
 sg13g2_a22oi_1 _3674_ (.Y(_1045_),
    .B1(net1067),
    .B2(net1425),
    .A2(net1156),
    .A1(net1319));
 sg13g2_nand2_1 _3675_ (.Y(_0313_),
    .A(net1014),
    .B(_1045_));
 sg13g2_a22oi_1 _3676_ (.Y(_1046_),
    .B1(net1067),
    .B2(net909),
    .A2(net1156),
    .A1(\tdc_inst.tdc_xor_result[125] ));
 sg13g2_nand2_1 _3677_ (.Y(_0314_),
    .A(net1014),
    .B(net910));
 sg13g2_a22oi_1 _3678_ (.Y(_1047_),
    .B1(net1067),
    .B2(net1415),
    .A2(net1156),
    .A1(net909));
 sg13g2_nand2_1 _3679_ (.Y(_0315_),
    .A(net1014),
    .B(_1047_));
 sg13g2_a22oi_1 _3680_ (.Y(_1048_),
    .B1(net1067),
    .B2(net792),
    .A2(net1156),
    .A1(\tdc_inst.tdc_xor_result[127] ));
 sg13g2_nand2_1 _3681_ (.Y(_0316_),
    .A(net1014),
    .B(net793));
 sg13g2_a22oi_1 _3682_ (.Y(_1049_),
    .B1(net1067),
    .B2(net1593),
    .A2(net1156),
    .A1(net792));
 sg13g2_nand2_1 _3683_ (.Y(_0317_),
    .A(net1012),
    .B(_1049_));
 sg13g2_a22oi_1 _3684_ (.Y(_1050_),
    .B1(net1066),
    .B2(net1469),
    .A2(net1155),
    .A1(\tdc_inst.tdc_xor_result[129] ));
 sg13g2_nand2_1 _3685_ (.Y(_0318_),
    .A(net1012),
    .B(net1470));
 sg13g2_a22oi_1 _3686_ (.Y(_1051_),
    .B1(net1066),
    .B2(net756),
    .A2(net1155),
    .A1(\tdc_inst.tdc_xor_result[130] ));
 sg13g2_nand2_1 _3687_ (.Y(_0319_),
    .A(net1012),
    .B(net757));
 sg13g2_a22oi_1 _3688_ (.Y(_1052_),
    .B1(net1066),
    .B2(net1645),
    .A2(net1155),
    .A1(net756));
 sg13g2_nand2_1 _3689_ (.Y(_0320_),
    .A(net1012),
    .B(_1052_));
 sg13g2_a22oi_1 _3690_ (.Y(_1053_),
    .B1(net1066),
    .B2(net1508),
    .A2(net1155),
    .A1(\tdc_inst.tdc_xor_result[132] ));
 sg13g2_nand2_1 _3691_ (.Y(_0321_),
    .A(net1013),
    .B(net1509));
 sg13g2_a22oi_1 _3692_ (.Y(_1054_),
    .B1(net1066),
    .B2(net895),
    .A2(net1155),
    .A1(\tdc_inst.tdc_xor_result[133] ));
 sg13g2_nand2_1 _3693_ (.Y(_0322_),
    .A(net1012),
    .B(net896));
 sg13g2_a22oi_1 _3694_ (.Y(_1055_),
    .B1(net1066),
    .B2(net1595),
    .A2(net1155),
    .A1(net895));
 sg13g2_nand2_1 _3695_ (.Y(_0323_),
    .A(net1012),
    .B(_1055_));
 sg13g2_a22oi_1 _3696_ (.Y(_1056_),
    .B1(net1065),
    .B2(net1362),
    .A2(net1154),
    .A1(\tdc_inst.tdc_xor_result[135] ));
 sg13g2_nand2_1 _3697_ (.Y(_0324_),
    .A(net1012),
    .B(net1363));
 sg13g2_a22oi_1 _3698_ (.Y(_1057_),
    .B1(net1065),
    .B2(net1626),
    .A2(net1154),
    .A1(net1362));
 sg13g2_nand2_1 _3699_ (.Y(_0325_),
    .A(net1012),
    .B(_1057_));
 sg13g2_a22oi_1 _3700_ (.Y(_1058_),
    .B1(net1065),
    .B2(net690),
    .A2(net1154),
    .A1(\tdc_inst.tdc_xor_result[137] ));
 sg13g2_nand2_1 _3701_ (.Y(_0326_),
    .A(net1013),
    .B(net691));
 sg13g2_a22oi_1 _3702_ (.Y(_1059_),
    .B1(net1065),
    .B2(net1393),
    .A2(net1154),
    .A1(net690));
 sg13g2_nand2_1 _3703_ (.Y(_0327_),
    .A(net1013),
    .B(_1059_));
 sg13g2_a22oi_1 _3704_ (.Y(_1060_),
    .B1(net1065),
    .B2(net1702),
    .A2(net1154),
    .A1(net1393));
 sg13g2_nand2_1 _3705_ (.Y(_0328_),
    .A(net1013),
    .B(_1060_));
 sg13g2_a22oi_1 _3706_ (.Y(_1061_),
    .B1(net1071),
    .B2(net1652),
    .A2(net1158),
    .A1(\tdc_inst.tdc_xor_result[140] ));
 sg13g2_nand2_1 _3707_ (.Y(_0329_),
    .A(net1013),
    .B(net1653));
 sg13g2_a221oi_1 _3708_ (.B2(net1339),
    .C1(_0919_),
    .B1(net1071),
    .A1(net1652),
    .Y(_1062_),
    .A2(net1158));
 sg13g2_inv_1 _3709_ (.Y(_0330_),
    .A(_1062_));
 sg13g2_mux2_1 _3710_ (.A0(net878),
    .A1(net5),
    .S(net1262),
    .X(_0331_));
 sg13g2_mux2_1 _3711_ (.A0(net1306),
    .A1(net943),
    .S(net1262),
    .X(_0332_));
 sg13g2_mux2_1 _3712_ (.A0(net943),
    .A1(net6),
    .S(net1262),
    .X(_0333_));
 sg13g2_mux2_1 _3713_ (.A0(net1617),
    .A1(net1306),
    .S(net1262),
    .X(_0334_));
 sg13g2_mux2_1 _3714_ (.A0(net632),
    .A1(net7),
    .S(net1262),
    .X(_0335_));
 sg13g2_mux2_1 _3715_ (.A0(net1541),
    .A1(net1414),
    .S(net1261),
    .X(_0336_));
 sg13g2_mux2_1 _3716_ (.A0(net1414),
    .A1(net1),
    .S(net1261),
    .X(_0337_));
 sg13g2_mux2_1 _3717_ (.A0(net1445),
    .A1(net1317),
    .S(net1261),
    .X(_0338_));
 sg13g2_mux2_1 _3718_ (.A0(net1317),
    .A1(net2),
    .S(net1261),
    .X(_0339_));
 sg13g2_mux2_1 _3719_ (.A0(net1487),
    .A1(net878),
    .S(net1262),
    .X(_0340_));
 sg13g2_and2_1 _3720_ (.A(\tdc_inst.stop_signal_sampling_clock_level ),
    .B(_0773_),
    .X(_1063_));
 sg13g2_nand2_2 _3721_ (.Y(_1064_),
    .A(\tdc_inst.stop_signal_sampling_clock_level ),
    .B(_0773_));
 sg13g2_a22oi_1 _3722_ (.Y(_1065_),
    .B1(net1068),
    .B2(net1615),
    .A2(net1156),
    .A1(\tdc_inst.stop_count_debug[0] ));
 sg13g2_nand2_1 _3723_ (.Y(_0341_),
    .A(net972),
    .B(net1616));
 sg13g2_a22oi_1 _3724_ (.Y(_1066_),
    .B1(net1068),
    .B2(net1351),
    .A2(net1156),
    .A1(\tdc_inst.stop_count_debug[1] ));
 sg13g2_nand2_1 _3725_ (.Y(_0342_),
    .A(net972),
    .B(net1352));
 sg13g2_a22oi_1 _3726_ (.Y(_1067_),
    .B1(net1065),
    .B2(net1654),
    .A2(net1154),
    .A1(net1351));
 sg13g2_nand2_1 _3727_ (.Y(_0343_),
    .A(net972),
    .B(_1067_));
 sg13g2_a22oi_1 _3728_ (.Y(_1068_),
    .B1(net1065),
    .B2(net893),
    .A2(net1154),
    .A1(\tdc_inst.stop_count_debug[3] ));
 sg13g2_nand2_1 _3729_ (.Y(_0344_),
    .A(net972),
    .B(net894));
 sg13g2_a22oi_1 _3730_ (.Y(_1069_),
    .B1(net1065),
    .B2(net1333),
    .A2(net1154),
    .A1(net893));
 sg13g2_nand2_1 _3731_ (.Y(_0345_),
    .A(net973),
    .B(_1069_));
 sg13g2_a22oi_1 _3732_ (.Y(_1070_),
    .B1(net1076),
    .B2(net1458),
    .A2(net1165),
    .A1(net1333));
 sg13g2_nand2_1 _3733_ (.Y(_0346_),
    .A(net973),
    .B(_1070_));
 sg13g2_a22oi_1 _3734_ (.Y(_1071_),
    .B1(net1076),
    .B2(net1570),
    .A2(net1165),
    .A1(net1458));
 sg13g2_nand2_1 _3735_ (.Y(_0347_),
    .A(net973),
    .B(_1071_));
 sg13g2_a22oi_1 _3736_ (.Y(_1072_),
    .B1(net1076),
    .B2(net1477),
    .A2(net1165),
    .A1(\tdc_inst.stop_count_debug[7] ));
 sg13g2_nand2_1 _3737_ (.Y(_0348_),
    .A(net973),
    .B(net1478));
 sg13g2_a22oi_1 _3738_ (.Y(_1073_),
    .B1(net1078),
    .B2(net1578),
    .A2(net1167),
    .A1(net1477));
 sg13g2_nand2_1 _3739_ (.Y(_0349_),
    .A(net973),
    .B(_1073_));
 sg13g2_a22oi_1 _3740_ (.Y(_1074_),
    .B1(net1078),
    .B2(net1522),
    .A2(net1167),
    .A1(\tdc_inst.stop_count_debug[9] ));
 sg13g2_nand2_1 _3741_ (.Y(_0350_),
    .A(net973),
    .B(net1523));
 sg13g2_a22oi_1 _3742_ (.Y(_1075_),
    .B1(net1078),
    .B2(net1564),
    .A2(net1167),
    .A1(net1522));
 sg13g2_nand2_1 _3743_ (.Y(_0351_),
    .A(net973),
    .B(_1075_));
 sg13g2_a22oi_1 _3744_ (.Y(_1076_),
    .B1(net1079),
    .B2(net1561),
    .A2(net1168),
    .A1(\tdc_inst.stop_count_debug[11] ));
 sg13g2_nand2_1 _3745_ (.Y(_0352_),
    .A(net974),
    .B(net1562));
 sg13g2_a22oi_1 _3746_ (.Y(_1077_),
    .B1(net1077),
    .B2(net955),
    .A2(net1166),
    .A1(\tdc_inst.stop_count_debug[12] ));
 sg13g2_nand2_1 _3747_ (.Y(_0353_),
    .A(net974),
    .B(net1263));
 sg13g2_a22oi_1 _3748_ (.Y(_1078_),
    .B1(net1077),
    .B2(net804),
    .A2(net1166),
    .A1(\tdc_inst.stop_count_debug[13] ));
 sg13g2_nand2_1 _3749_ (.Y(_0354_),
    .A(net974),
    .B(net805));
 sg13g2_a22oi_1 _3750_ (.Y(_1079_),
    .B1(net1077),
    .B2(net1724),
    .A2(net1166),
    .A1(net804));
 sg13g2_nand2_1 _3751_ (.Y(_0355_),
    .A(net974),
    .B(_1079_));
 sg13g2_a22oi_1 _3752_ (.Y(_1080_),
    .B1(net1076),
    .B2(net844),
    .A2(net1165),
    .A1(\tdc_inst.stop_count_debug[15] ));
 sg13g2_nand2_1 _3753_ (.Y(_0356_),
    .A(net974),
    .B(net845));
 sg13g2_a22oi_1 _3754_ (.Y(_1081_),
    .B1(net1077),
    .B2(net1284),
    .A2(net1166),
    .A1(net844));
 sg13g2_nand2_1 _3755_ (.Y(_0357_),
    .A(net968),
    .B(_1081_));
 sg13g2_a22oi_1 _3756_ (.Y(_1082_),
    .B1(net1076),
    .B2(net1432),
    .A2(net1165),
    .A1(net1284));
 sg13g2_nand2_1 _3757_ (.Y(_0358_),
    .A(net968),
    .B(_1082_));
 sg13g2_a22oi_1 _3758_ (.Y(_1083_),
    .B1(net1076),
    .B2(net1341),
    .A2(net1165),
    .A1(\tdc_inst.stop_count_debug[18] ));
 sg13g2_nand2_1 _3759_ (.Y(_0359_),
    .A(net973),
    .B(net1342));
 sg13g2_a22oi_1 _3760_ (.Y(_1084_),
    .B1(net1076),
    .B2(net1402),
    .A2(net1165),
    .A1(net1341));
 sg13g2_nand2_1 _3761_ (.Y(_0360_),
    .A(net968),
    .B(_1084_));
 sg13g2_a22oi_1 _3762_ (.Y(_1085_),
    .B1(net1076),
    .B2(net1437),
    .A2(net1165),
    .A1(net1402));
 sg13g2_nand2_1 _3763_ (.Y(_0361_),
    .A(net968),
    .B(_1085_));
 sg13g2_a22oi_1 _3764_ (.Y(_1086_),
    .B1(net1073),
    .B2(net630),
    .A2(net1162),
    .A1(\tdc_inst.stop_count_debug[21] ));
 sg13g2_nand2_1 _3765_ (.Y(_0362_),
    .A(net968),
    .B(net631));
 sg13g2_a22oi_1 _3766_ (.Y(_1087_),
    .B1(net1072),
    .B2(net1754),
    .A2(net1161),
    .A1(net630));
 sg13g2_nand2_1 _3767_ (.Y(_0363_),
    .A(net968),
    .B(_1087_));
 sg13g2_a22oi_1 _3768_ (.Y(_1088_),
    .B1(net1073),
    .B2(net1489),
    .A2(net1162),
    .A1(\tdc_inst.stop_count_debug[23] ));
 sg13g2_nand2_1 _3769_ (.Y(_0364_),
    .A(net968),
    .B(net1490));
 sg13g2_a22oi_1 _3770_ (.Y(_1089_),
    .B1(net1073),
    .B2(net762),
    .A2(net1162),
    .A1(\tdc_inst.stop_count_debug[24] ));
 sg13g2_nand2_1 _3771_ (.Y(_0365_),
    .A(net969),
    .B(net763));
 sg13g2_a22oi_1 _3772_ (.Y(_1090_),
    .B1(net1073),
    .B2(net1366),
    .A2(net1162),
    .A1(net762));
 sg13g2_nand2_1 _3773_ (.Y(_0366_),
    .A(net968),
    .B(_1090_));
 sg13g2_a22oi_1 _3774_ (.Y(_1091_),
    .B1(net1073),
    .B2(net1516),
    .A2(net1162),
    .A1(net1366));
 sg13g2_nand2_1 _3775_ (.Y(_0367_),
    .A(net969),
    .B(_1091_));
 sg13g2_a22oi_1 _3776_ (.Y(_1092_),
    .B1(net1072),
    .B2(net1266),
    .A2(net1161),
    .A1(\tdc_inst.stop_count_debug[27] ));
 sg13g2_nand2_1 _3777_ (.Y(_0368_),
    .A(net969),
    .B(net1267));
 sg13g2_a22oi_1 _3778_ (.Y(_1093_),
    .B1(net1072),
    .B2(net1332),
    .A2(net1161),
    .A1(net1266));
 sg13g2_nand2_1 _3779_ (.Y(_0369_),
    .A(net969),
    .B(_1093_));
 sg13g2_a22oi_1 _3780_ (.Y(_1094_),
    .B1(net1072),
    .B2(net1289),
    .A2(net1161),
    .A1(\tdc_inst.stop_count_debug[29] ));
 sg13g2_nand2_1 _3781_ (.Y(_0370_),
    .A(net969),
    .B(net1290));
 sg13g2_a22oi_1 _3782_ (.Y(_1095_),
    .B1(net1072),
    .B2(net1611),
    .A2(net1161),
    .A1(net1289));
 sg13g2_nand2_1 _3783_ (.Y(_0371_),
    .A(net969),
    .B(_1095_));
 sg13g2_a22oi_1 _3784_ (.Y(_1096_),
    .B1(net1072),
    .B2(net923),
    .A2(net1161),
    .A1(\tdc_inst.stop_count_debug[31] ));
 sg13g2_nand2_1 _3785_ (.Y(_0372_),
    .A(net971),
    .B(net924));
 sg13g2_a22oi_1 _3786_ (.Y(_1097_),
    .B1(net1072),
    .B2(net1303),
    .A2(net1161),
    .A1(net923));
 sg13g2_nand2_1 _3787_ (.Y(_0373_),
    .A(net971),
    .B(_1097_));
 sg13g2_a22oi_1 _3788_ (.Y(_1098_),
    .B1(net1072),
    .B2(net1692),
    .A2(net1161),
    .A1(net1303));
 sg13g2_nand2_1 _3789_ (.Y(_0374_),
    .A(net971),
    .B(_1098_));
 sg13g2_a22oi_1 _3790_ (.Y(_1099_),
    .B1(net1075),
    .B2(net552),
    .A2(net1164),
    .A1(\tdc_inst.stop_count_debug[34] ));
 sg13g2_nand2_1 _3791_ (.Y(_0375_),
    .A(net970),
    .B(net553));
 sg13g2_a22oi_1 _3792_ (.Y(_1100_),
    .B1(net1075),
    .B2(net1661),
    .A2(net1164),
    .A1(net552));
 sg13g2_nand2_1 _3793_ (.Y(_0376_),
    .A(net970),
    .B(_1100_));
 sg13g2_a22oi_1 _3794_ (.Y(_1101_),
    .B1(net1075),
    .B2(net1558),
    .A2(net1164),
    .A1(\tdc_inst.stop_count_debug[36] ));
 sg13g2_nand2_1 _3795_ (.Y(_0377_),
    .A(net970),
    .B(net1559));
 sg13g2_a22oi_1 _3796_ (.Y(_1102_),
    .B1(net1074),
    .B2(net1435),
    .A2(net1163),
    .A1(\tdc_inst.stop_count_debug[37] ));
 sg13g2_nand2_1 _3797_ (.Y(_0378_),
    .A(net977),
    .B(net1436));
 sg13g2_a22oi_1 _3798_ (.Y(_1103_),
    .B1(net1074),
    .B2(net1423),
    .A2(net1163),
    .A1(\tdc_inst.stop_count_debug[38] ));
 sg13g2_nand2_1 _3799_ (.Y(_0379_),
    .A(net970),
    .B(net1424));
 sg13g2_a22oi_1 _3800_ (.Y(_1104_),
    .B1(net1074),
    .B2(net733),
    .A2(net1163),
    .A1(\tdc_inst.stop_count_debug[39] ));
 sg13g2_nand2_1 _3801_ (.Y(_0380_),
    .A(net971),
    .B(net734));
 sg13g2_a22oi_1 _3802_ (.Y(_1105_),
    .B1(net1074),
    .B2(net920),
    .A2(net1163),
    .A1(net733));
 sg13g2_nand2_1 _3803_ (.Y(_0381_),
    .A(net971),
    .B(_1105_));
 sg13g2_a22oi_1 _3804_ (.Y(_1106_),
    .B1(net1074),
    .B2(net1641),
    .A2(net1163),
    .A1(net920));
 sg13g2_nand2_1 _3805_ (.Y(_0382_),
    .A(net971),
    .B(_1106_));
 sg13g2_a22oi_1 _3806_ (.Y(_1107_),
    .B1(net1074),
    .B2(net1542),
    .A2(net1163),
    .A1(\tdc_inst.stop_count_debug[42] ));
 sg13g2_nand2_1 _3807_ (.Y(_0383_),
    .A(net971),
    .B(net1543));
 sg13g2_a22oi_1 _3808_ (.Y(_1108_),
    .B1(net1074),
    .B2(net1684),
    .A2(net1163),
    .A1(net1542));
 sg13g2_nand2_1 _3809_ (.Y(_0384_),
    .A(net978),
    .B(_1108_));
 sg13g2_a22oi_1 _3810_ (.Y(_1109_),
    .B1(net1084),
    .B2(net1621),
    .A2(net1173),
    .A1(\tdc_inst.stop_count_debug[44] ));
 sg13g2_nand2_1 _3811_ (.Y(_0385_),
    .A(net978),
    .B(net1622));
 sg13g2_a22oi_1 _3812_ (.Y(_1110_),
    .B1(net1084),
    .B2(net708),
    .A2(net1173),
    .A1(\tdc_inst.stop_count_debug[45] ));
 sg13g2_nand2_1 _3813_ (.Y(_0386_),
    .A(net978),
    .B(net709));
 sg13g2_a22oi_1 _3814_ (.Y(_1111_),
    .B1(net1084),
    .B2(net1607),
    .A2(net1173),
    .A1(net708));
 sg13g2_nand2_1 _3815_ (.Y(_0387_),
    .A(net979),
    .B(_1111_));
 sg13g2_a22oi_1 _3816_ (.Y(_1112_),
    .B1(net1084),
    .B2(net876),
    .A2(net1173),
    .A1(\tdc_inst.stop_count_debug[47] ));
 sg13g2_nand2_1 _3817_ (.Y(_0388_),
    .A(net978),
    .B(net877));
 sg13g2_a22oi_1 _3818_ (.Y(_1113_),
    .B1(net1084),
    .B2(net1450),
    .A2(net1173),
    .A1(net876));
 sg13g2_nand2_1 _3819_ (.Y(_0389_),
    .A(net978),
    .B(_1113_));
 sg13g2_a22oi_1 _3820_ (.Y(_1114_),
    .B1(net1084),
    .B2(net1590),
    .A2(net1173),
    .A1(net1450));
 sg13g2_nand2_1 _3821_ (.Y(_0390_),
    .A(net981),
    .B(_1114_));
 sg13g2_a22oi_1 _3822_ (.Y(_1115_),
    .B1(net1085),
    .B2(net1421),
    .A2(net1174),
    .A1(\tdc_inst.stop_count_debug[50] ));
 sg13g2_nand2_1 _3823_ (.Y(_0391_),
    .A(net981),
    .B(net1422));
 sg13g2_a22oi_1 _3824_ (.Y(_1116_),
    .B1(net1085),
    .B2(net1576),
    .A2(net1174),
    .A1(net1421));
 sg13g2_nand2_1 _3825_ (.Y(_0392_),
    .A(net981),
    .B(_1116_));
 sg13g2_a22oi_1 _3826_ (.Y(_1117_),
    .B1(net1085),
    .B2(net1567),
    .A2(net1174),
    .A1(\tdc_inst.stop_count_debug[52] ));
 sg13g2_nand2_1 _3827_ (.Y(_0393_),
    .A(net981),
    .B(net1568));
 sg13g2_a22oi_1 _3828_ (.Y(_1118_),
    .B1(net1085),
    .B2(net1525),
    .A2(net1174),
    .A1(\tdc_inst.stop_count_debug[53] ));
 sg13g2_nand2_1 _3829_ (.Y(_0394_),
    .A(net980),
    .B(net1526));
 sg13g2_a22oi_1 _3830_ (.Y(_1119_),
    .B1(net1085),
    .B2(net1296),
    .A2(net1174),
    .A1(\tdc_inst.stop_count_debug[54] ));
 sg13g2_nand2_1 _3831_ (.Y(_0395_),
    .A(net980),
    .B(net1297));
 sg13g2_a22oi_1 _3832_ (.Y(_1120_),
    .B1(net1085),
    .B2(net851),
    .A2(net1174),
    .A1(\tdc_inst.stop_count_debug[55] ));
 sg13g2_nand2_1 _3833_ (.Y(_0396_),
    .A(net980),
    .B(net852));
 sg13g2_a22oi_1 _3834_ (.Y(_1121_),
    .B1(net1085),
    .B2(net1544),
    .A2(net1174),
    .A1(net851));
 sg13g2_nand2_1 _3835_ (.Y(_0397_),
    .A(net980),
    .B(_1121_));
 sg13g2_a22oi_1 _3836_ (.Y(_1122_),
    .B1(net1087),
    .B2(net1387),
    .A2(net1176),
    .A1(\tdc_inst.stop_count_debug[57] ));
 sg13g2_nand2_1 _3837_ (.Y(_0398_),
    .A(net980),
    .B(net1388));
 sg13g2_a22oi_1 _3838_ (.Y(_1123_),
    .B1(net1085),
    .B2(net712),
    .A2(net1174),
    .A1(\tdc_inst.stop_count_debug[58] ));
 sg13g2_nand2_1 _3839_ (.Y(_0399_),
    .A(net980),
    .B(net713));
 sg13g2_a22oi_1 _3840_ (.Y(_1124_),
    .B1(net1087),
    .B2(net1418),
    .A2(net1176),
    .A1(net712));
 sg13g2_nand2_1 _3841_ (.Y(_0400_),
    .A(net981),
    .B(_1124_));
 sg13g2_a22oi_1 _3842_ (.Y(_1125_),
    .B1(net1086),
    .B2(net1658),
    .A2(net1175),
    .A1(net1418));
 sg13g2_nand2_1 _3843_ (.Y(_0401_),
    .A(net980),
    .B(_1125_));
 sg13g2_a22oi_1 _3844_ (.Y(_1126_),
    .B1(net1086),
    .B2(net731),
    .A2(net1175),
    .A1(\tdc_inst.stop_count_debug[61] ));
 sg13g2_nand2_1 _3845_ (.Y(_0402_),
    .A(net980),
    .B(net732));
 sg13g2_a22oi_1 _3846_ (.Y(_1127_),
    .B1(net1087),
    .B2(net831),
    .A2(net1176),
    .A1(net731));
 sg13g2_nand2_1 _3847_ (.Y(_0403_),
    .A(net983),
    .B(_1127_));
 sg13g2_a22oi_1 _3848_ (.Y(_1128_),
    .B1(net1087),
    .B2(net657),
    .A2(net1176),
    .A1(\tdc_inst.stop_count_debug[63] ));
 sg13g2_nand2_1 _3849_ (.Y(_0404_),
    .A(net983),
    .B(net658));
 sg13g2_a22oi_1 _3850_ (.Y(_1129_),
    .B1(net1086),
    .B2(net1602),
    .A2(net1175),
    .A1(net657));
 sg13g2_nand2_1 _3851_ (.Y(_0405_),
    .A(net983),
    .B(_1129_));
 sg13g2_a22oi_1 _3852_ (.Y(_1130_),
    .B1(net1086),
    .B2(net718),
    .A2(net1175),
    .A1(\tdc_inst.stop_count_debug[65] ));
 sg13g2_nand2_1 _3853_ (.Y(_0406_),
    .A(net983),
    .B(net719));
 sg13g2_a22oi_1 _3854_ (.Y(_1131_),
    .B1(net1086),
    .B2(net1601),
    .A2(net1175),
    .A1(net718));
 sg13g2_nand2_1 _3855_ (.Y(_0407_),
    .A(net983),
    .B(_1131_));
 sg13g2_a22oi_1 _3856_ (.Y(_1132_),
    .B1(net1093),
    .B2(net728),
    .A2(net1182),
    .A1(\tdc_inst.stop_count_debug[67] ));
 sg13g2_nand2_1 _3857_ (.Y(_0408_),
    .A(net983),
    .B(net729));
 sg13g2_a22oi_1 _3858_ (.Y(_1133_),
    .B1(net1091),
    .B2(net853),
    .A2(net1182),
    .A1(net728));
 sg13g2_nand2_1 _3859_ (.Y(_0409_),
    .A(net982),
    .B(_1133_));
 sg13g2_a22oi_1 _3860_ (.Y(_1134_),
    .B1(net1091),
    .B2(net944),
    .A2(net1180),
    .A1(net853));
 sg13g2_nand2_1 _3861_ (.Y(_0410_),
    .A(net982),
    .B(_1134_));
 sg13g2_a22oi_1 _3862_ (.Y(_1135_),
    .B1(net1093),
    .B2(net1663),
    .A2(net1180),
    .A1(net944));
 sg13g2_nand2_1 _3863_ (.Y(_0411_),
    .A(net988),
    .B(_1135_));
 sg13g2_a22oi_1 _3864_ (.Y(_1136_),
    .B1(net1091),
    .B2(net618),
    .A2(net1180),
    .A1(\tdc_inst.stop_count_debug[71] ));
 sg13g2_nand2_1 _3865_ (.Y(_0412_),
    .A(net988),
    .B(net619));
 sg13g2_a22oi_1 _3866_ (.Y(_1137_),
    .B1(net1091),
    .B2(net891),
    .A2(net1180),
    .A1(net618));
 sg13g2_nand2_1 _3867_ (.Y(_0413_),
    .A(net987),
    .B(_1137_));
 sg13g2_a22oi_1 _3868_ (.Y(_1138_),
    .B1(net1091),
    .B2(net682),
    .A2(net1180),
    .A1(\tdc_inst.stop_count_debug[73] ));
 sg13g2_nand2_1 _3869_ (.Y(_0414_),
    .A(net988),
    .B(net683));
 sg13g2_a22oi_1 _3870_ (.Y(_1139_),
    .B1(net1091),
    .B2(net1620),
    .A2(net1180),
    .A1(net682));
 sg13g2_nand2_1 _3871_ (.Y(_0415_),
    .A(net987),
    .B(_1139_));
 sg13g2_a22oi_1 _3872_ (.Y(_1140_),
    .B1(net1088),
    .B2(net1463),
    .A2(net1177),
    .A1(\tdc_inst.stop_count_debug[75] ));
 sg13g2_nand2_1 _3873_ (.Y(_0416_),
    .A(net987),
    .B(net1464));
 sg13g2_a22oi_1 _3874_ (.Y(_1141_),
    .B1(net1090),
    .B2(net1378),
    .A2(net1178),
    .A1(\tdc_inst.stop_count_debug[76] ));
 sg13g2_nand2_1 _3875_ (.Y(_0417_),
    .A(net985),
    .B(net1379));
 sg13g2_a22oi_1 _3876_ (.Y(_1142_),
    .B1(net1089),
    .B2(net1510),
    .A2(net1178),
    .A1(net1378));
 sg13g2_nand2_1 _3877_ (.Y(_0418_),
    .A(net985),
    .B(_1142_));
 sg13g2_a22oi_1 _3878_ (.Y(_1143_),
    .B1(net1089),
    .B2(net1606),
    .A2(net1179),
    .A1(net1510));
 sg13g2_nand2_1 _3879_ (.Y(_0419_),
    .A(net986),
    .B(_1143_));
 sg13g2_a22oi_1 _3880_ (.Y(_1144_),
    .B1(net1090),
    .B2(net1480),
    .A2(net1179),
    .A1(\tdc_inst.stop_count_debug[79] ));
 sg13g2_nand2_1 _3881_ (.Y(_0420_),
    .A(net989),
    .B(net1481));
 sg13g2_a22oi_1 _3882_ (.Y(_1145_),
    .B1(net1092),
    .B2(net1669),
    .A2(net1181),
    .A1(net1480));
 sg13g2_nand2_1 _3883_ (.Y(_0421_),
    .A(net989),
    .B(_1145_));
 sg13g2_a22oi_1 _3884_ (.Y(_1146_),
    .B1(net1092),
    .B2(net684),
    .A2(net1181),
    .A1(\tdc_inst.stop_count_debug[81] ));
 sg13g2_nand2_1 _3885_ (.Y(_0422_),
    .A(net989),
    .B(net685));
 sg13g2_a22oi_1 _3886_ (.Y(_1147_),
    .B1(net1092),
    .B2(net1565),
    .A2(net1181),
    .A1(net684));
 sg13g2_nand2_1 _3887_ (.Y(_0423_),
    .A(net989),
    .B(_1147_));
 sg13g2_a22oi_1 _3888_ (.Y(_1148_),
    .B1(net1092),
    .B2(net1638),
    .A2(net1181),
    .A1(net1565));
 sg13g2_nand2_1 _3889_ (.Y(_0424_),
    .A(net989),
    .B(_1148_));
 sg13g2_a22oi_1 _3890_ (.Y(_1149_),
    .B1(net1092),
    .B2(net1310),
    .A2(net1181),
    .A1(\tdc_inst.stop_count_debug[84] ));
 sg13g2_nand2_1 _3891_ (.Y(_0425_),
    .A(net989),
    .B(net1311));
 sg13g2_a22oi_1 _3892_ (.Y(_1150_),
    .B1(net1092),
    .B2(net1720),
    .A2(net1181),
    .A1(net1310));
 sg13g2_nand2_1 _3893_ (.Y(_0426_),
    .A(net990),
    .B(_1150_));
 sg13g2_a22oi_1 _3894_ (.Y(_1151_),
    .B1(net1092),
    .B2(net1383),
    .A2(net1181),
    .A1(\tdc_inst.stop_count_debug[86] ));
 sg13g2_nand2_1 _3895_ (.Y(_0427_),
    .A(net990),
    .B(net1384));
 sg13g2_a22oi_1 _3896_ (.Y(_1152_),
    .B1(net1093),
    .B2(net1369),
    .A2(net1182),
    .A1(\tdc_inst.stop_count_debug[87] ));
 sg13g2_nand2_1 _3897_ (.Y(_0428_),
    .A(net987),
    .B(net1370));
 sg13g2_a22oi_1 _3898_ (.Y(_1153_),
    .B1(net1093),
    .B2(net698),
    .A2(net1182),
    .A1(\tdc_inst.stop_count_debug[88] ));
 sg13g2_nand2_1 _3899_ (.Y(_0429_),
    .A(net987),
    .B(net699));
 sg13g2_a22oi_1 _3900_ (.Y(_1154_),
    .B1(net1092),
    .B2(net1326),
    .A2(net1181),
    .A1(net698));
 sg13g2_nand2_1 _3901_ (.Y(_0430_),
    .A(net988),
    .B(_1154_));
 sg13g2_a22oi_1 _3902_ (.Y(_1155_),
    .B1(net1091),
    .B2(net1446),
    .A2(net1180),
    .A1(net1326));
 sg13g2_nand2_1 _3903_ (.Y(_0431_),
    .A(net987),
    .B(_1155_));
 sg13g2_a22oi_1 _3904_ (.Y(_1156_),
    .B1(net1091),
    .B2(net1717),
    .A2(net1180),
    .A1(net1446));
 sg13g2_nand2_1 _3905_ (.Y(_0432_),
    .A(net987),
    .B(_1156_));
 sg13g2_a22oi_1 _3906_ (.Y(_1157_),
    .B1(net1090),
    .B2(net1439),
    .A2(net1179),
    .A1(\tdc_inst.stop_count_debug[92] ));
 sg13g2_nand2_1 _3907_ (.Y(_0433_),
    .A(net987),
    .B(net1440));
 sg13g2_a22oi_1 _3908_ (.Y(_1158_),
    .B1(net1088),
    .B2(net781),
    .A2(net1177),
    .A1(\tdc_inst.stop_count_debug[93] ));
 sg13g2_nand2_1 _3909_ (.Y(_0434_),
    .A(net985),
    .B(net782));
 sg13g2_a22oi_1 _3910_ (.Y(_1159_),
    .B1(net1088),
    .B2(net1532),
    .A2(net1177),
    .A1(net781));
 sg13g2_nand2_1 _3911_ (.Y(_0435_),
    .A(net979),
    .B(_1159_));
 sg13g2_a22oi_1 _3912_ (.Y(_1160_),
    .B1(net1090),
    .B2(net1700),
    .A2(net1179),
    .A1(net1532));
 sg13g2_nand2_1 _3913_ (.Y(_0436_),
    .A(net982),
    .B(_1160_));
 sg13g2_a22oi_1 _3914_ (.Y(_1161_),
    .B1(net1086),
    .B2(net1406),
    .A2(net1175),
    .A1(\tdc_inst.stop_count_debug[96] ));
 sg13g2_nand2_1 _3915_ (.Y(_0437_),
    .A(net982),
    .B(net1407));
 sg13g2_a22oi_1 _3916_ (.Y(_1162_),
    .B1(net1086),
    .B2(net1438),
    .A2(net1175),
    .A1(net1406));
 sg13g2_nand2_1 _3917_ (.Y(_0438_),
    .A(net982),
    .B(_1162_));
 sg13g2_a22oi_1 _3918_ (.Y(_1163_),
    .B1(net1086),
    .B2(net1554),
    .A2(net1175),
    .A1(net1438));
 sg13g2_nand2_1 _3919_ (.Y(_0439_),
    .A(net982),
    .B(_1163_));
 sg13g2_a22oi_1 _3920_ (.Y(_1164_),
    .B1(net1083),
    .B2(net1441),
    .A2(net1172),
    .A1(\tdc_inst.stop_count_debug[99] ));
 sg13g2_nand2_1 _3921_ (.Y(_0440_),
    .A(net982),
    .B(net1442));
 sg13g2_a22oi_1 _3922_ (.Y(_1165_),
    .B1(net1084),
    .B2(net1575),
    .A2(net1172),
    .A1(net1441));
 sg13g2_nand2_1 _3923_ (.Y(_0441_),
    .A(net982),
    .B(_1165_));
 sg13g2_a22oi_1 _3924_ (.Y(_1166_),
    .B1(net1083),
    .B2(net1527),
    .A2(net1173),
    .A1(\tdc_inst.stop_count_debug[101] ));
 sg13g2_nand2_1 _3925_ (.Y(_0442_),
    .A(net978),
    .B(net1528));
 sg13g2_a22oi_1 _3926_ (.Y(_1167_),
    .B1(net1083),
    .B2(net1455),
    .A2(net1172),
    .A1(\tdc_inst.stop_count_debug[102] ));
 sg13g2_nand2_1 _3927_ (.Y(_0443_),
    .A(net978),
    .B(net1456));
 sg13g2_a22oi_1 _3928_ (.Y(_1168_),
    .B1(net1083),
    .B2(net1545),
    .A2(net1172),
    .A1(net1455));
 sg13g2_nand2_1 _3929_ (.Y(_0444_),
    .A(net978),
    .B(_1168_));
 sg13g2_a22oi_1 _3930_ (.Y(_1169_),
    .B1(net1083),
    .B2(net1574),
    .A2(net1172),
    .A1(net1545));
 sg13g2_nand2_1 _3931_ (.Y(_0445_),
    .A(net979),
    .B(_1169_));
 sg13g2_a22oi_1 _3932_ (.Y(_1170_),
    .B1(net1083),
    .B2(net1381),
    .A2(net1172),
    .A1(\tdc_inst.stop_count_debug[105] ));
 sg13g2_nand2_1 _3933_ (.Y(_0446_),
    .A(net979),
    .B(net1382));
 sg13g2_a22oi_1 _3934_ (.Y(_1171_),
    .B1(net1083),
    .B2(net1282),
    .A2(net1172),
    .A1(\tdc_inst.stop_count_debug[106] ));
 sg13g2_nand2_1 _3935_ (.Y(_0447_),
    .A(net979),
    .B(net1283));
 sg13g2_a22oi_1 _3936_ (.Y(_1172_),
    .B1(net1083),
    .B2(net1409),
    .A2(net1172),
    .A1(net1282));
 sg13g2_nand2_1 _3937_ (.Y(_0448_),
    .A(net979),
    .B(_1172_));
 sg13g2_a22oi_1 _3938_ (.Y(_1173_),
    .B1(net1088),
    .B2(net1465),
    .A2(net1177),
    .A1(net1409));
 sg13g2_nand2_1 _3939_ (.Y(_0449_),
    .A(net984),
    .B(_1173_));
 sg13g2_a22oi_1 _3940_ (.Y(_1174_),
    .B1(net1088),
    .B2(net1304),
    .A2(net1177),
    .A1(\tdc_inst.stop_count_debug[109] ));
 sg13g2_nand2_1 _3941_ (.Y(_0450_),
    .A(net984),
    .B(net1305));
 sg13g2_a22oi_1 _3942_ (.Y(_1175_),
    .B1(net1081),
    .B2(net1549),
    .A2(net1170),
    .A1(net1304));
 sg13g2_nand2_1 _3943_ (.Y(_0451_),
    .A(net979),
    .B(_1175_));
 sg13g2_a22oi_1 _3944_ (.Y(_1176_),
    .B1(net1074),
    .B2(net1732),
    .A2(net1163),
    .A1(net1549));
 sg13g2_nand2_1 _3945_ (.Y(_0452_),
    .A(net970),
    .B(_1176_));
 sg13g2_a22oi_1 _3946_ (.Y(_1177_),
    .B1(net1080),
    .B2(net558),
    .A2(net1169),
    .A1(\tdc_inst.stop_count_debug[112] ));
 sg13g2_nand2_1 _3947_ (.Y(_0453_),
    .A(net970),
    .B(net559));
 sg13g2_a22oi_1 _3948_ (.Y(_1178_),
    .B1(net1080),
    .B2(net1281),
    .A2(net1169),
    .A1(net558));
 sg13g2_nand2_1 _3949_ (.Y(_0454_),
    .A(net970),
    .B(_1178_));
 sg13g2_a22oi_1 _3950_ (.Y(_1179_),
    .B1(net1080),
    .B2(net1354),
    .A2(net1169),
    .A1(net1281));
 sg13g2_nand2_1 _3951_ (.Y(_0455_),
    .A(net970),
    .B(_1179_));
 sg13g2_a22oi_1 _3952_ (.Y(_1180_),
    .B1(net1080),
    .B2(net1426),
    .A2(net1169),
    .A1(net1354));
 sg13g2_nand2_1 _3953_ (.Y(_0456_),
    .A(net975),
    .B(_1180_));
 sg13g2_a22oi_1 _3954_ (.Y(_1181_),
    .B1(net1080),
    .B2(net1301),
    .A2(net1169),
    .A1(\tdc_inst.stop_count_debug[116] ));
 sg13g2_nand2_1 _3955_ (.Y(_0457_),
    .A(net975),
    .B(net1302));
 sg13g2_a22oi_1 _3956_ (.Y(_1182_),
    .B1(net1080),
    .B2(net1343),
    .A2(net1169),
    .A1(net1301));
 sg13g2_nand2_1 _3957_ (.Y(_0458_),
    .A(net974),
    .B(_1182_));
 sg13g2_a22oi_1 _3958_ (.Y(_1183_),
    .B1(net1080),
    .B2(net1694),
    .A2(net1169),
    .A1(net1343));
 sg13g2_nand2_1 _3959_ (.Y(_0459_),
    .A(net985),
    .B(_1183_));
 sg13g2_a22oi_1 _3960_ (.Y(_1184_),
    .B1(net1080),
    .B2(net1539),
    .A2(net1169),
    .A1(\tdc_inst.stop_count_debug[119] ));
 sg13g2_nand2_1 _3961_ (.Y(_0460_),
    .A(net985),
    .B(net1540));
 sg13g2_a22oi_1 _3962_ (.Y(_1185_),
    .B1(net1088),
    .B2(net861),
    .A2(net1177),
    .A1(\tdc_inst.stop_count_debug[120] ));
 sg13g2_nand2_1 _3963_ (.Y(_0461_),
    .A(net985),
    .B(net862));
 sg13g2_a22oi_1 _3964_ (.Y(_1186_),
    .B1(net1088),
    .B2(net574),
    .A2(net1177),
    .A1(\tdc_inst.stop_count_debug[121] ));
 sg13g2_nand2_1 _3965_ (.Y(_0462_),
    .A(net986),
    .B(net575));
 sg13g2_a22oi_1 _3966_ (.Y(_1187_),
    .B1(net1088),
    .B2(net1614),
    .A2(net1177),
    .A1(net574));
 sg13g2_nand2_1 _3967_ (.Y(_0463_),
    .A(net986),
    .B(_1187_));
 sg13g2_a22oi_1 _3968_ (.Y(_1188_),
    .B1(net1089),
    .B2(net931),
    .A2(net1178),
    .A1(\tdc_inst.stop_count_debug[123] ));
 sg13g2_nand2_1 _3969_ (.Y(_0464_),
    .A(net985),
    .B(net932));
 sg13g2_a22oi_1 _3970_ (.Y(_1189_),
    .B1(net1089),
    .B2(net1560),
    .A2(net1178),
    .A1(net931));
 sg13g2_nand2_1 _3971_ (.Y(_0465_),
    .A(net985),
    .B(_1189_));
 sg13g2_a22oi_1 _3972_ (.Y(_1190_),
    .B1(net1089),
    .B2(net1583),
    .A2(net1178),
    .A1(net1560));
 sg13g2_nand2_1 _3973_ (.Y(_0466_),
    .A(net986),
    .B(_1190_));
 sg13g2_a22oi_1 _3974_ (.Y(_1191_),
    .B1(net1081),
    .B2(net779),
    .A2(net1170),
    .A1(\tdc_inst.stop_count_debug[126] ));
 sg13g2_nand2_1 _3975_ (.Y(_0467_),
    .A(net986),
    .B(net780));
 sg13g2_a22oi_1 _3976_ (.Y(_1192_),
    .B1(net1081),
    .B2(net914),
    .A2(net1170),
    .A1(net779));
 sg13g2_nand2_1 _3977_ (.Y(_0468_),
    .A(net975),
    .B(_1192_));
 sg13g2_a22oi_1 _3978_ (.Y(_1193_),
    .B1(net1081),
    .B2(net1451),
    .A2(net1170),
    .A1(net914));
 sg13g2_nand2_1 _3979_ (.Y(_0469_),
    .A(net975),
    .B(_1193_));
 sg13g2_a22oi_1 _3980_ (.Y(_1194_),
    .B1(net1081),
    .B2(net841),
    .A2(net1170),
    .A1(\tdc_inst.stop_count_debug[129] ));
 sg13g2_nand2_1 _3981_ (.Y(_0470_),
    .A(net974),
    .B(net842));
 sg13g2_a22oi_1 _3982_ (.Y(_1195_),
    .B1(net1082),
    .B2(net1372),
    .A2(net1171),
    .A1(net841));
 sg13g2_nand2_1 _3983_ (.Y(_0471_),
    .A(net974),
    .B(_1195_));
 sg13g2_a22oi_1 _3984_ (.Y(_1196_),
    .B1(net1081),
    .B2(net1410),
    .A2(net1170),
    .A1(net1372));
 sg13g2_nand2_1 _3985_ (.Y(_0472_),
    .A(net976),
    .B(_1196_));
 sg13g2_a22oi_1 _3986_ (.Y(_1197_),
    .B1(net1081),
    .B2(net1639),
    .A2(net1170),
    .A1(net1410));
 sg13g2_nand2_1 _3987_ (.Y(_0473_),
    .A(net975),
    .B(_1197_));
 sg13g2_a22oi_1 _3988_ (.Y(_1198_),
    .B1(net1078),
    .B2(net874),
    .A2(net1167),
    .A1(\tdc_inst.stop_count_debug[133] ));
 sg13g2_nand2_1 _3989_ (.Y(_0474_),
    .A(net975),
    .B(net875));
 sg13g2_a22oi_1 _3990_ (.Y(_1199_),
    .B1(net1078),
    .B2(net1580),
    .A2(net1167),
    .A1(net874));
 sg13g2_nand2_1 _3991_ (.Y(_0475_),
    .A(net975),
    .B(_1199_));
 sg13g2_a22oi_1 _3992_ (.Y(_1200_),
    .B1(net1078),
    .B2(net800),
    .A2(net1167),
    .A1(\tdc_inst.stop_count_debug[135] ));
 sg13g2_nand2_1 _3993_ (.Y(_0476_),
    .A(net972),
    .B(net801));
 sg13g2_a22oi_1 _3994_ (.Y(_1201_),
    .B1(net1078),
    .B2(net1380),
    .A2(net1167),
    .A1(net800));
 sg13g2_nand2_1 _3995_ (.Y(_0477_),
    .A(net972),
    .B(_1201_));
 sg13g2_a22oi_1 _3996_ (.Y(_1202_),
    .B1(net1078),
    .B2(net1416),
    .A2(net1167),
    .A1(net1380));
 sg13g2_nand2_1 _3997_ (.Y(_0478_),
    .A(net976),
    .B(_1202_));
 sg13g2_a22oi_1 _3998_ (.Y(_1203_),
    .B1(net1095),
    .B2(net811),
    .A2(net1184),
    .A1(\tdc_inst.stop_count_debug[138] ));
 sg13g2_nand2_1 _3999_ (.Y(_0479_),
    .A(net976),
    .B(net812));
 sg13g2_a22oi_1 _4000_ (.Y(_1204_),
    .B1(net1095),
    .B2(net1596),
    .A2(net1184),
    .A1(net811));
 sg13g2_nand2_1 _4001_ (.Y(_0480_),
    .A(net972),
    .B(_1204_));
 sg13g2_a22oi_1 _4002_ (.Y(_1205_),
    .B1(net1071),
    .B2(net1612),
    .A2(net1158),
    .A1(net1596));
 sg13g2_nand2_1 _4003_ (.Y(_0481_),
    .A(net972),
    .B(_1205_));
 sg13g2_a221oi_1 _4004_ (.B2(net1318),
    .C1(_1063_),
    .B1(net1071),
    .A1(net1612),
    .Y(_1206_),
    .A2(net1158));
 sg13g2_inv_1 _4005_ (.Y(_0482_),
    .A(_1206_));
 sg13g2_xor2_1 _4006_ (.B(cpol_sync),
    .A(cpha_sync),
    .X(_1207_));
 sg13g2_nand3b_1 _4007_ (.B(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .C(_0007_),
    .Y(_1208_),
    .A_N(spi_clk_sync));
 sg13g2_nand3b_1 _4008_ (.B(_0007_),
    .C(spi_clk_sync),
    .Y(_1209_),
    .A_N(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_nand2b_1 _4009_ (.Y(_1210_),
    .B(_1209_),
    .A_N(_1207_));
 sg13g2_a21oi_1 _4010_ (.A1(_1207_),
    .A2(_1208_),
    .Y(_1211_),
    .B1(_0722_));
 sg13g2_nand2_1 _4011_ (.Y(_1212_),
    .A(_1210_),
    .B(_1211_));
 sg13g2_nor2_2 _4012_ (.A(_0725_),
    .B(net1043),
    .Y(_1213_));
 sg13g2_o21ai_1 _4013_ (.B1(_0725_),
    .Y(_1214_),
    .A1(_0742_),
    .A2(net1043));
 sg13g2_nor2b_1 _4014_ (.A(_1213_),
    .B_N(_1214_),
    .Y(_0483_));
 sg13g2_xor2_1 _4015_ (.B(_1213_),
    .A(net1760),
    .X(_0484_));
 sg13g2_nand3_1 _4016_ (.B(net1698),
    .C(_1213_),
    .A(net1760),
    .Y(_1215_));
 sg13g2_a21o_1 _4017_ (.A2(_1213_),
    .A1(net1760),
    .B1(net1698),
    .X(_1216_));
 sg13g2_and2_1 _4018_ (.A(_1215_),
    .B(_1216_),
    .X(_0485_));
 sg13g2_xnor2_1 _4019_ (.Y(_1217_),
    .A(_0726_),
    .B(_1215_));
 sg13g2_nor2_1 _4020_ (.A(_0749_),
    .B(_1217_),
    .Y(_0486_));
 sg13g2_nor2_1 _4021_ (.A(net1500),
    .B(net1041),
    .Y(_1218_));
 sg13g2_a21oi_1 _4022_ (.A1(_0721_),
    .A2(net1041),
    .Y(_0487_),
    .B1(_1218_));
 sg13g2_mux2_1 _4023_ (.A0(net1581),
    .A1(net1744),
    .S(net1041),
    .X(_0488_));
 sg13g2_mux2_1 _4024_ (.A0(net700),
    .A1(\spi_wrapper_i.reg_addr[1] ),
    .S(net1041),
    .X(_0489_));
 sg13g2_nor2_1 _4025_ (.A(net858),
    .B(net1041),
    .Y(_1219_));
 sg13g2_a21oi_1 _4026_ (.A1(_0730_),
    .A2(net1041),
    .Y(_0490_),
    .B1(_1219_));
 sg13g2_nor2_1 _4027_ (.A(net1666),
    .B(net1041),
    .Y(_1220_));
 sg13g2_a21oi_1 _4028_ (.A1(_0734_),
    .A2(net1041),
    .Y(_0491_),
    .B1(_1220_));
 sg13g2_nand2_1 _4029_ (.Y(_1221_),
    .A(_0722_),
    .B(net921));
 sg13g2_o21ai_1 _4030_ (.B1(_1221_),
    .Y(_0492_),
    .A1(_0721_),
    .A2(net1042));
 sg13g2_mux2_1 _4031_ (.A0(net1581),
    .A1(net1223),
    .S(net1042),
    .X(_0493_));
 sg13g2_mux2_1 _4032_ (.A0(net700),
    .A1(net1222),
    .S(net1042),
    .X(_0494_));
 sg13g2_mux2_1 _4033_ (.A0(net858),
    .A1(net1221),
    .S(_0750_),
    .X(_0495_));
 sg13g2_mux2_1 _4034_ (.A0(net1666),
    .A1(net1220),
    .S(net1042),
    .X(_0496_));
 sg13g2_mux2_1 _4035_ (.A0(net1524),
    .A1(net1219),
    .S(_0750_),
    .X(_0497_));
 sg13g2_mux2_1 _4036_ (.A0(net1270),
    .A1(net1218),
    .S(net1042),
    .X(_0498_));
 sg13g2_mux2_1 _4037_ (.A0(net1457),
    .A1(net1217),
    .S(net1042),
    .X(_0499_));
 sg13g2_mux2_1 _4038_ (.A0(net1500),
    .A1(net1216),
    .S(net1042),
    .X(_0500_));
 sg13g2_nor2_2 _4039_ (.A(_0724_),
    .B(net1043),
    .Y(_1222_));
 sg13g2_a21o_1 _4040_ (.A2(_0740_),
    .A1(net1809),
    .B1(net1043),
    .X(_1223_));
 sg13g2_a21oi_1 _4041_ (.A1(_0724_),
    .A2(_1223_),
    .Y(_0501_),
    .B1(_1222_));
 sg13g2_xor2_1 _4042_ (.B(_1222_),
    .A(net1695),
    .X(_0502_));
 sg13g2_a21oi_1 _4043_ (.A1(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .A2(_1222_),
    .Y(_1224_),
    .B1(net901));
 sg13g2_and2_1 _4044_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .B(net901),
    .X(_1225_));
 sg13g2_a21oi_1 _4045_ (.A1(_1222_),
    .A2(_1225_),
    .Y(_0503_),
    .B1(net902));
 sg13g2_nand3_1 _4046_ (.B(_0747_),
    .C(net1043),
    .A(net1781),
    .Y(_1226_));
 sg13g2_nand2_1 _4047_ (.Y(_1227_),
    .A(net1769),
    .B(_1225_));
 sg13g2_xor2_1 _4048_ (.B(_1227_),
    .A(net1781),
    .X(_1228_));
 sg13g2_o21ai_1 _4049_ (.B1(net1782),
    .Y(_0504_),
    .A1(_1223_),
    .A2(_1228_));
 sg13g2_nand2_2 _4050_ (.Y(_1229_),
    .A(\spi_wrapper_i.reg_addr[1] ),
    .B(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_nor2_2 _4051_ (.A(_0008_),
    .B(_1229_),
    .Y(_1230_));
 sg13g2_nand2_2 _4052_ (.Y(_1231_),
    .A(net1260),
    .B(\spi_wrapper_i.reg_data_o_vld ));
 sg13g2_nor3_2 _4053_ (.A(net1226),
    .B(_1229_),
    .C(_1231_),
    .Y(_1232_));
 sg13g2_mux2_1 _4054_ (.A0(net714),
    .A1(net1223),
    .S(_1232_),
    .X(_0505_));
 sg13g2_mux2_1 _4055_ (.A0(net855),
    .A1(net1222),
    .S(_1232_),
    .X(_0506_));
 sg13g2_mux2_1 _4056_ (.A0(net677),
    .A1(net1221),
    .S(_1232_),
    .X(_0507_));
 sg13g2_mux2_1 _4057_ (.A0(net754),
    .A1(net1220),
    .S(_1232_),
    .X(_0508_));
 sg13g2_mux2_1 _4058_ (.A0(net892),
    .A1(net1219),
    .S(_1232_),
    .X(_0509_));
 sg13g2_mux2_1 _4059_ (.A0(net813),
    .A1(net1218),
    .S(_1232_),
    .X(_0510_));
 sg13g2_mux2_1 _4060_ (.A0(net679),
    .A1(net1217),
    .S(_1232_),
    .X(_0511_));
 sg13g2_mux2_1 _4061_ (.A0(net666),
    .A1(net1216),
    .S(_1232_),
    .X(_0512_));
 sg13g2_mux2_1 _4062_ (.A0(_1208_),
    .A1(_1209_),
    .S(_1207_),
    .X(_1233_));
 sg13g2_nand2_1 _4063_ (.Y(_1234_),
    .A(net1133),
    .B(_1233_));
 sg13g2_o21ai_1 _4064_ (.B1(net1259),
    .Y(_1235_),
    .A1(_0751_),
    .A2(_1234_));
 sg13g2_nor2_1 _4065_ (.A(\spi_wrapper_i.reg_addr[1] ),
    .B(\spi_wrapper_i.reg_addr[0] ),
    .Y(_1236_));
 sg13g2_or2_1 _4066_ (.X(_1237_),
    .B(\spi_wrapper_i.reg_addr[0] ),
    .A(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_a21oi_1 _4067_ (.A1(_0730_),
    .A2(_1237_),
    .Y(_1238_),
    .B1(_0731_));
 sg13g2_o21ai_1 _4068_ (.B1(net1226),
    .Y(_1239_),
    .A1(net1227),
    .A2(_1236_));
 sg13g2_nand2b_2 _4069_ (.Y(_1240_),
    .B(\spi_wrapper_i.reg_addr[1] ),
    .A_N(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_nor2_1 _4070_ (.A(net1227),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_a22oi_1 _4071_ (.Y(_1242_),
    .B1(net1127),
    .B2(\config_regs[16] ),
    .A2(net1134),
    .A1(\config_regs[32] ));
 sg13g2_nor2_1 _4072_ (.A(net1227),
    .B(_1229_),
    .Y(_1243_));
 sg13g2_a22oi_1 _4073_ (.Y(_1244_),
    .B1(net1125),
    .B2(\config_regs[24] ),
    .A2(_1230_),
    .A1(\config_regs[56] ));
 sg13g2_nor2_2 _4074_ (.A(net1226),
    .B(_1240_),
    .Y(_1245_));
 sg13g2_nand2b_2 _4075_ (.Y(_1246_),
    .B(\spi_wrapper_i.reg_addr[0] ),
    .A_N(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_nor2_1 _4076_ (.A(net1227),
    .B(_1246_),
    .Y(_1247_));
 sg13g2_a22oi_1 _4077_ (.Y(_1248_),
    .B1(net1123),
    .B2(\config_regs[8] ),
    .A2(_1245_),
    .A1(\config_regs[48] ));
 sg13g2_nand3_1 _4078_ (.B(_1244_),
    .C(_1248_),
    .A(_1242_),
    .Y(_1249_));
 sg13g2_nor2_1 _4079_ (.A(net1226),
    .B(_1246_),
    .Y(_1250_));
 sg13g2_a21oi_1 _4080_ (.A1(\config_regs[40] ),
    .A2(net1121),
    .Y(_1251_),
    .B1(net1224));
 sg13g2_o21ai_1 _4081_ (.B1(_1251_),
    .Y(_1252_),
    .A1(_0009_),
    .A2(net1128));
 sg13g2_nor2_1 _4082_ (.A(net1226),
    .B(_1237_),
    .Y(_1253_));
 sg13g2_a21oi_1 _4083_ (.A1(_1239_),
    .A2(_1249_),
    .Y(_1254_),
    .B1(_1252_));
 sg13g2_a22oi_1 _4084_ (.Y(_1255_),
    .B1(net1122),
    .B2(\coarse_result[8] ),
    .A2(net1124),
    .A1(\coarse_result[24] ));
 sg13g2_a22oi_1 _4085_ (.Y(_1256_),
    .B1(net1120),
    .B2(\fine_result[0] ),
    .A2(net1126),
    .A1(net570));
 sg13g2_a221oi_1 _4086_ (.B2(\fine_result[8] ),
    .C1(_0734_),
    .B1(net1121),
    .A1(_0733_),
    .Y(_1257_),
    .A2(net1131));
 sg13g2_nand3_1 _4087_ (.B(_1256_),
    .C(_1257_),
    .A(_1255_),
    .Y(_1258_));
 sg13g2_nor4_1 _4088_ (.A(_0722_),
    .B(_0751_),
    .C(net1132),
    .D(_1254_),
    .Y(_1259_));
 sg13g2_a22oi_1 _4089_ (.Y(_1260_),
    .B1(_1258_),
    .B2(_1259_),
    .A2(net967),
    .A1(net602));
 sg13g2_inv_1 _4090_ (.Y(_0513_),
    .A(net603));
 sg13g2_a22oi_1 _4091_ (.Y(_1261_),
    .B1(net1120),
    .B2(\config_regs[33] ),
    .A2(net1121),
    .A1(\config_regs[41] ));
 sg13g2_a22oi_1 _4092_ (.Y(_1262_),
    .B1(net1125),
    .B2(\config_regs[25] ),
    .A2(_1230_),
    .A1(\config_regs[57] ));
 sg13g2_a22oi_1 _4093_ (.Y(_1263_),
    .B1(net1123),
    .B2(\config_regs[9] ),
    .A2(net1127),
    .A1(\config_regs[17] ));
 sg13g2_a21oi_1 _4094_ (.A1(\config_regs[49] ),
    .A2(_1245_),
    .Y(_1264_),
    .B1(net1225));
 sg13g2_nand4_1 _4095_ (.B(_1262_),
    .C(_1263_),
    .A(_1261_),
    .Y(_1265_),
    .D(_1264_));
 sg13g2_a22oi_1 _4096_ (.Y(_1266_),
    .B1(net1122),
    .B2(\coarse_result[9] ),
    .A2(net1134),
    .A1(\fine_result[1] ));
 sg13g2_a22oi_1 _4097_ (.Y(_1267_),
    .B1(net1124),
    .B2(\coarse_result[25] ),
    .A2(net1126),
    .A1(\coarse_result[17] ));
 sg13g2_nand3_1 _4098_ (.B(_1266_),
    .C(_1267_),
    .A(net1224),
    .Y(_1268_));
 sg13g2_nand3_1 _4099_ (.B(_1265_),
    .C(_1268_),
    .A(_1239_),
    .Y(_1269_));
 sg13g2_nand2_1 _4100_ (.Y(_1270_),
    .A(_0734_),
    .B(_0012_));
 sg13g2_a21oi_1 _4101_ (.A1(net1224),
    .A2(_0013_),
    .Y(_1271_),
    .B1(net1128));
 sg13g2_a21oi_1 _4102_ (.A1(_1270_),
    .A2(_1271_),
    .Y(_1272_),
    .B1(net1133));
 sg13g2_or2_2 _4103_ (.X(_1273_),
    .B(net967),
    .A(_0751_));
 sg13g2_a221oi_1 _4104_ (.B2(_1272_),
    .C1(_1273_),
    .B1(_1269_),
    .A1(_0011_),
    .Y(_1274_),
    .A2(net1132));
 sg13g2_a21o_1 _4105_ (.A2(net967),
    .A1(net706),
    .B1(_1274_),
    .X(_0514_));
 sg13g2_a22oi_1 _4106_ (.Y(_1275_),
    .B1(net1126),
    .B2(\coarse_result[18] ),
    .A2(net1134),
    .A1(\fine_result[2] ));
 sg13g2_a22oi_1 _4107_ (.Y(_1276_),
    .B1(net1122),
    .B2(\coarse_result[10] ),
    .A2(net1124),
    .A1(\coarse_result[26] ));
 sg13g2_a22oi_1 _4108_ (.Y(_1277_),
    .B1(net1125),
    .B2(\config_regs[26] ),
    .A2(net1127),
    .A1(\config_regs[18] ));
 sg13g2_a21oi_1 _4109_ (.A1(\config_regs[10] ),
    .A2(net1123),
    .Y(_1278_),
    .B1(net1129));
 sg13g2_a22oi_1 _4110_ (.Y(_1279_),
    .B1(_1253_),
    .B2(\config_regs[34] ),
    .A2(_1250_),
    .A1(\config_regs[42] ));
 sg13g2_a22oi_1 _4111_ (.Y(_1280_),
    .B1(_1245_),
    .B2(\config_regs[50] ),
    .A2(_1230_),
    .A1(\config_regs[58] ));
 sg13g2_nand4_1 _4112_ (.B(_1278_),
    .C(_1279_),
    .A(_1277_),
    .Y(_1281_),
    .D(_1280_));
 sg13g2_a21oi_1 _4113_ (.A1(_0015_),
    .A2(net1129),
    .Y(_1282_),
    .B1(net1225));
 sg13g2_nand2_1 _4114_ (.Y(_1283_),
    .A(_1281_),
    .B(_1282_));
 sg13g2_nand3_1 _4115_ (.B(_1275_),
    .C(_1276_),
    .A(net1128),
    .Y(_1284_));
 sg13g2_a21oi_1 _4116_ (.A1(_0016_),
    .A2(net1131),
    .Y(_1285_),
    .B1(_0734_));
 sg13g2_a21oi_1 _4117_ (.A1(_1284_),
    .A2(_1285_),
    .Y(_1286_),
    .B1(net1132));
 sg13g2_a221oi_1 _4118_ (.B2(_1286_),
    .C1(_1273_),
    .B1(_1283_),
    .A1(_0014_),
    .Y(_1287_),
    .A2(net1132));
 sg13g2_a21o_1 _4119_ (.A2(net967),
    .A1(net675),
    .B1(_1287_),
    .X(_0515_));
 sg13g2_a22oi_1 _4120_ (.Y(_1288_),
    .B1(net1124),
    .B2(\coarse_result[27] ),
    .A2(net1134),
    .A1(\fine_result[3] ));
 sg13g2_a22oi_1 _4121_ (.Y(_1289_),
    .B1(net1122),
    .B2(\coarse_result[11] ),
    .A2(net1126),
    .A1(\coarse_result[19] ));
 sg13g2_a21oi_1 _4122_ (.A1(_1288_),
    .A2(_1289_),
    .Y(_1290_),
    .B1(net1131));
 sg13g2_o21ai_1 _4123_ (.B1(net1224),
    .Y(_1291_),
    .A1(_0019_),
    .A2(net1128));
 sg13g2_nor2_1 _4124_ (.A(_1290_),
    .B(_1291_),
    .Y(_1292_));
 sg13g2_nand2_1 _4125_ (.Y(_1293_),
    .A(_0018_),
    .B(net1130));
 sg13g2_nand2_1 _4126_ (.Y(_1294_),
    .A(\config_regs[19] ),
    .B(net1127));
 sg13g2_a22oi_1 _4127_ (.Y(_1295_),
    .B1(net1125),
    .B2(\config_regs[27] ),
    .A2(_1230_),
    .A1(\config_regs[59] ));
 sg13g2_a22oi_1 _4128_ (.Y(_1296_),
    .B1(net1121),
    .B2(\config_regs[43] ),
    .A2(_1245_),
    .A1(\config_regs[51] ));
 sg13g2_a21oi_1 _4129_ (.A1(\config_regs[11] ),
    .A2(net1123),
    .Y(_1297_),
    .B1(net1130));
 sg13g2_nand4_1 _4130_ (.B(_1295_),
    .C(_1296_),
    .A(_1294_),
    .Y(_1298_),
    .D(_1297_));
 sg13g2_a221oi_1 _4131_ (.B2(_1298_),
    .C1(net1225),
    .B1(_1293_),
    .A1(\config_regs[35] ),
    .Y(_1299_),
    .A2(net1120));
 sg13g2_o21ai_1 _4132_ (.B1(_0755_),
    .Y(_1300_),
    .A1(_1292_),
    .A2(_1299_));
 sg13g2_a21oi_1 _4133_ (.A1(_0017_),
    .A2(net1132),
    .Y(_1301_),
    .B1(_1273_));
 sg13g2_a22oi_1 _4134_ (.Y(_1302_),
    .B1(_1300_),
    .B2(_1301_),
    .A2(net967),
    .A1(net582));
 sg13g2_inv_1 _4135_ (.Y(_0516_),
    .A(net583));
 sg13g2_and2_1 _4136_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ),
    .B(net967),
    .X(_1303_));
 sg13g2_nand2_1 _4137_ (.Y(_1304_),
    .A(_0021_),
    .B(net1129));
 sg13g2_nand2_1 _4138_ (.Y(_1305_),
    .A(\config_regs[44] ),
    .B(net1121));
 sg13g2_a22oi_1 _4139_ (.Y(_1306_),
    .B1(net1127),
    .B2(\config_regs[20] ),
    .A2(_1230_),
    .A1(\config_regs[60] ));
 sg13g2_a22oi_1 _4140_ (.Y(_1307_),
    .B1(net1123),
    .B2(\config_regs[12] ),
    .A2(net1125),
    .A1(\config_regs[28] ));
 sg13g2_a21oi_1 _4141_ (.A1(\config_regs[52] ),
    .A2(_1245_),
    .Y(_1308_),
    .B1(net1129));
 sg13g2_nand4_1 _4142_ (.B(_1306_),
    .C(_1307_),
    .A(_1305_),
    .Y(_1309_),
    .D(_1308_));
 sg13g2_a22oi_1 _4143_ (.Y(_1310_),
    .B1(net1124),
    .B2(\coarse_result[28] ),
    .A2(net1134),
    .A1(\fine_result[4] ));
 sg13g2_a22oi_1 _4144_ (.Y(_1311_),
    .B1(net1122),
    .B2(\coarse_result[12] ),
    .A2(net1126),
    .A1(\coarse_result[20] ));
 sg13g2_a21oi_1 _4145_ (.A1(_1310_),
    .A2(_1311_),
    .Y(_1312_),
    .B1(net1131));
 sg13g2_o21ai_1 _4146_ (.B1(net1224),
    .Y(_1313_),
    .A1(_0022_),
    .A2(net1128));
 sg13g2_nor2_1 _4147_ (.A(_1312_),
    .B(_1313_),
    .Y(_1314_));
 sg13g2_a221oi_1 _4148_ (.B2(_1309_),
    .C1(net1225),
    .B1(_1304_),
    .A1(\config_regs[36] ),
    .Y(_1315_),
    .A2(net1120));
 sg13g2_o21ai_1 _4149_ (.B1(_0755_),
    .Y(_1316_),
    .A1(_1314_),
    .A2(_1315_));
 sg13g2_a21oi_1 _4150_ (.A1(net1735),
    .A2(net1132),
    .Y(_1317_),
    .B1(_1273_));
 sg13g2_a21o_1 _4151_ (.A2(_1317_),
    .A1(_1316_),
    .B1(_1303_),
    .X(_0517_));
 sg13g2_a22oi_1 _4152_ (.Y(_1318_),
    .B1(net1122),
    .B2(\coarse_result[13] ),
    .A2(net1134),
    .A1(\fine_result[5] ));
 sg13g2_a22oi_1 _4153_ (.Y(_1319_),
    .B1(net1124),
    .B2(\coarse_result[29] ),
    .A2(net1126),
    .A1(\coarse_result[21] ));
 sg13g2_a21oi_1 _4154_ (.A1(_1318_),
    .A2(_1319_),
    .Y(_1320_),
    .B1(net1131));
 sg13g2_o21ai_1 _4155_ (.B1(net1224),
    .Y(_1321_),
    .A1(_0025_),
    .A2(net1128));
 sg13g2_nor2_1 _4156_ (.A(_1320_),
    .B(_1321_),
    .Y(_1322_));
 sg13g2_nand2_1 _4157_ (.Y(_1323_),
    .A(_0024_),
    .B(net1129));
 sg13g2_nand2_1 _4158_ (.Y(_1324_),
    .A(\config_regs[29] ),
    .B(net1125));
 sg13g2_a22oi_1 _4159_ (.Y(_1325_),
    .B1(net1127),
    .B2(\config_regs[21] ),
    .A2(_1230_),
    .A1(\config_regs[61] ));
 sg13g2_a22oi_1 _4160_ (.Y(_1326_),
    .B1(net1121),
    .B2(\config_regs[45] ),
    .A2(net1123),
    .A1(\config_regs[13] ));
 sg13g2_a21oi_1 _4161_ (.A1(\config_regs[53] ),
    .A2(_1245_),
    .Y(_1327_),
    .B1(net1130));
 sg13g2_nand4_1 _4162_ (.B(_1325_),
    .C(_1326_),
    .A(_1324_),
    .Y(_1328_),
    .D(_1327_));
 sg13g2_a221oi_1 _4163_ (.B2(_1328_),
    .C1(net1225),
    .B1(_1323_),
    .A1(\config_regs[37] ),
    .Y(_1329_),
    .A2(net1120));
 sg13g2_o21ai_1 _4164_ (.B1(_0755_),
    .Y(_1330_),
    .A1(_1322_),
    .A2(_1329_));
 sg13g2_a21oi_1 _4165_ (.A1(_0023_),
    .A2(net1132),
    .Y(_1331_),
    .B1(_1273_));
 sg13g2_a22oi_1 _4166_ (.Y(_1332_),
    .B1(_1330_),
    .B2(_1331_),
    .A2(_1235_),
    .A1(net576));
 sg13g2_inv_1 _4167_ (.Y(_0518_),
    .A(net577));
 sg13g2_nand2_1 _4168_ (.Y(_1333_),
    .A(_0027_),
    .B(net1129));
 sg13g2_a22oi_1 _4169_ (.Y(_1334_),
    .B1(net1120),
    .B2(\config_regs[38] ),
    .A2(net1121),
    .A1(\config_regs[46] ));
 sg13g2_a22oi_1 _4170_ (.Y(_1335_),
    .B1(net1123),
    .B2(\config_regs[14] ),
    .A2(net1125),
    .A1(\config_regs[30] ));
 sg13g2_a22oi_1 _4171_ (.Y(_1336_),
    .B1(net1127),
    .B2(\config_regs[22] ),
    .A2(_1230_),
    .A1(\config_regs[62] ));
 sg13g2_a21oi_1 _4172_ (.A1(\config_regs[54] ),
    .A2(_1245_),
    .Y(_1337_),
    .B1(net1129));
 sg13g2_nand4_1 _4173_ (.B(_1335_),
    .C(_1336_),
    .A(_1334_),
    .Y(_1338_),
    .D(_1337_));
 sg13g2_a21oi_2 _4174_ (.B1(net1225),
    .Y(_1339_),
    .A2(_1338_),
    .A1(_1333_));
 sg13g2_a22oi_1 _4175_ (.Y(_1340_),
    .B1(net1124),
    .B2(\coarse_result[30] ),
    .A2(net1134),
    .A1(\fine_result[6] ));
 sg13g2_a22oi_1 _4176_ (.Y(_1341_),
    .B1(net1122),
    .B2(\coarse_result[14] ),
    .A2(net1126),
    .A1(\coarse_result[22] ));
 sg13g2_a21oi_1 _4177_ (.A1(_1340_),
    .A2(_1341_),
    .Y(_1342_),
    .B1(net1131));
 sg13g2_o21ai_1 _4178_ (.B1(net1224),
    .Y(_1343_),
    .A1(_0028_),
    .A2(net1128));
 sg13g2_nor2_1 _4179_ (.A(_1342_),
    .B(_1343_),
    .Y(_1344_));
 sg13g2_o21ai_1 _4180_ (.B1(_0755_),
    .Y(_1345_),
    .A1(_1339_),
    .A2(_1344_));
 sg13g2_a21oi_1 _4181_ (.A1(_0026_),
    .A2(net1133),
    .Y(_1346_),
    .B1(_1273_));
 sg13g2_a22oi_1 _4182_ (.Y(_1347_),
    .B1(_1345_),
    .B2(_1346_),
    .A2(net967),
    .A1(net584));
 sg13g2_inv_1 _4183_ (.Y(_0519_),
    .A(net585));
 sg13g2_nand2_1 _4184_ (.Y(_1348_),
    .A(net590),
    .B(net967));
 sg13g2_and2_1 _4185_ (.A(_0030_),
    .B(net1130),
    .X(_1349_));
 sg13g2_a22oi_1 _4186_ (.Y(_1350_),
    .B1(_1245_),
    .B2(\config_regs[55] ),
    .A2(_1230_),
    .A1(\config_regs[63] ));
 sg13g2_a22oi_1 _4187_ (.Y(_1351_),
    .B1(net1123),
    .B2(\config_regs[15] ),
    .A2(net1125),
    .A1(\config_regs[31] ));
 sg13g2_a21oi_1 _4188_ (.A1(\config_regs[47] ),
    .A2(net1121),
    .Y(_1352_),
    .B1(net1129));
 sg13g2_nand3_1 _4189_ (.B(_1351_),
    .C(_1352_),
    .A(_1350_),
    .Y(_1353_));
 sg13g2_a21oi_1 _4190_ (.A1(\config_regs[23] ),
    .A2(net1127),
    .Y(_1354_),
    .B1(_1353_));
 sg13g2_a22oi_1 _4191_ (.Y(_1355_),
    .B1(net1124),
    .B2(\coarse_result[31] ),
    .A2(net1126),
    .A1(\coarse_result[23] ));
 sg13g2_a22oi_1 _4192_ (.Y(_1356_),
    .B1(net1122),
    .B2(\coarse_result[15] ),
    .A2(net1134),
    .A1(\fine_result[7] ));
 sg13g2_a21oi_1 _4193_ (.A1(_1355_),
    .A2(_1356_),
    .Y(_1357_),
    .B1(net1131));
 sg13g2_nor2_1 _4194_ (.A(_0734_),
    .B(_1357_),
    .Y(_1358_));
 sg13g2_o21ai_1 _4195_ (.B1(_1358_),
    .Y(_1359_),
    .A1(_0031_),
    .A2(net1128));
 sg13g2_a21oi_1 _4196_ (.A1(\config_regs[39] ),
    .A2(net1120),
    .Y(_1360_),
    .B1(net1225));
 sg13g2_o21ai_1 _4197_ (.B1(_1360_),
    .Y(_1361_),
    .A1(_1349_),
    .A2(_1354_));
 sg13g2_a21oi_1 _4198_ (.A1(_1359_),
    .A2(_1361_),
    .Y(_1362_),
    .B1(net1132));
 sg13g2_a21o_1 _4199_ (.A2(net1133),
    .A1(_0029_),
    .B1(_1273_),
    .X(_1363_));
 sg13g2_o21ai_1 _4200_ (.B1(_1348_),
    .Y(_0520_),
    .A1(_1362_),
    .A2(_1363_));
 sg13g2_nor2b_1 _4201_ (.A(\tdc_inst.fine_procedure_counter[1] ),
    .B_N(\tdc_inst.fine_procedure_counter[4] ),
    .Y(_1364_));
 sg13g2_a221oi_1 _4202_ (.B2(_1364_),
    .C1(_0713_),
    .B1(_0766_),
    .A1(_0005_),
    .Y(_1365_),
    .A2(_0765_));
 sg13g2_nor2_1 _4203_ (.A(\tdc_inst.fine_procedure_counter[8] ),
    .B(_1365_),
    .Y(_1366_));
 sg13g2_nand4_1 _4204_ (.B(\tdc_inst.fine_procedure_counter[0] ),
    .C(_0766_),
    .A(\tdc_inst.fine_procedure_counter[7] ),
    .Y(_1367_),
    .D(_1364_));
 sg13g2_nand3_1 _4205_ (.B(\tdc_inst.fine_procedure_counter[4] ),
    .C(_0766_),
    .A(\tdc_inst.fine_procedure_counter[7] ),
    .Y(_1368_));
 sg13g2_and2_1 _4206_ (.A(_1366_),
    .B(_1367_),
    .X(_1369_));
 sg13g2_nand2b_1 _4207_ (.Y(_1370_),
    .B(net1210),
    .A_N(_1369_));
 sg13g2_nor2_1 _4208_ (.A(net1160),
    .B(_1369_),
    .Y(_1371_));
 sg13g2_mux2_1 _4209_ (.A0(net1686),
    .A1(\tdc_inst.fine_another_counter[0] ),
    .S(net964),
    .X(_0521_));
 sg13g2_mux2_1 _4210_ (.A0(net1650),
    .A1(\tdc_inst.fine_another_counter[1] ),
    .S(net964),
    .X(_0522_));
 sg13g2_mux2_1 _4211_ (.A0(net1330),
    .A1(\tdc_inst.fine_another_counter[2] ),
    .S(net964),
    .X(_0523_));
 sg13g2_mux2_1 _4212_ (.A0(net912),
    .A1(\tdc_inst.fine_another_counter[3] ),
    .S(net964),
    .X(_0524_));
 sg13g2_mux2_1 _4213_ (.A0(net766),
    .A1(\tdc_inst.fine_another_counter[4] ),
    .S(net961),
    .X(_0525_));
 sg13g2_mux2_1 _4214_ (.A0(net1722),
    .A1(\tdc_inst.fine_another_counter[5] ),
    .S(net964),
    .X(_0526_));
 sg13g2_mux2_1 _4215_ (.A0(net1356),
    .A1(\tdc_inst.fine_another_counter[6] ),
    .S(net964),
    .X(_0527_));
 sg13g2_mux2_1 _4216_ (.A0(net1673),
    .A1(\tdc_inst.fine_another_counter[7] ),
    .S(net964),
    .X(_0528_));
 sg13g2_mux2_1 _4217_ (.A0(net859),
    .A1(\tdc_inst.fine_another_counter[8] ),
    .S(net965),
    .X(_0529_));
 sg13g2_mux2_1 _4218_ (.A0(net604),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .S(net1043),
    .X(_0530_));
 sg13g2_mux2_1 _4219_ (.A0(net1581),
    .A1(net700),
    .S(net1043),
    .X(_0531_));
 sg13g2_mux2_1 _4220_ (.A0(net700),
    .A1(net858),
    .S(net1044),
    .X(_0532_));
 sg13g2_mux2_1 _4221_ (.A0(net858),
    .A1(net1666),
    .S(net1043),
    .X(_0533_));
 sg13g2_mux2_1 _4222_ (.A0(net1666),
    .A1(net1524),
    .S(net1044),
    .X(_0534_));
 sg13g2_mux2_1 _4223_ (.A0(net1524),
    .A1(net1270),
    .S(net1044),
    .X(_0535_));
 sg13g2_mux2_1 _4224_ (.A0(net1270),
    .A1(net1457),
    .S(net1044),
    .X(_0536_));
 sg13g2_mux2_1 _4225_ (.A0(net1457),
    .A1(net1500),
    .S(net1044),
    .X(_0537_));
 sg13g2_mux2_1 _4226_ (.A0(net1640),
    .A1(net1487),
    .S(net1261),
    .X(_0538_));
 sg13g2_nand2b_2 _4227_ (.Y(_1372_),
    .B(net1120),
    .A_N(_1231_));
 sg13g2_mux2_1 _4228_ (.A0(net1223),
    .A1(net1629),
    .S(_1372_),
    .X(_0539_));
 sg13g2_mux2_1 _4229_ (.A0(net1222),
    .A1(net1660),
    .S(_1372_),
    .X(_0540_));
 sg13g2_mux2_1 _4230_ (.A0(net1221),
    .A1(net1664),
    .S(_1372_),
    .X(_0541_));
 sg13g2_mux2_1 _4231_ (.A0(net1360),
    .A1(\config_regs[35] ),
    .S(_1372_),
    .X(_0542_));
 sg13g2_mux2_1 _4232_ (.A0(net833),
    .A1(\config_regs[36] ),
    .S(_1372_),
    .X(_0543_));
 sg13g2_mux2_1 _4233_ (.A0(net1503),
    .A1(\config_regs[37] ),
    .S(_1372_),
    .X(_0544_));
 sg13g2_mux2_1 _4234_ (.A0(net669),
    .A1(\config_regs[38] ),
    .S(_1372_),
    .X(_0545_));
 sg13g2_mux2_1 _4235_ (.A0(net659),
    .A1(\config_regs[39] ),
    .S(_1372_),
    .X(_0546_));
 sg13g2_nor3_2 _4236_ (.A(net1226),
    .B(_1231_),
    .C(_1246_),
    .Y(_1373_));
 sg13g2_mux2_1 _4237_ (.A0(net794),
    .A1(\spi_wrapper_i.reg_data_o[0] ),
    .S(_1373_),
    .X(_0547_));
 sg13g2_mux2_1 _4238_ (.A0(net710),
    .A1(net1222),
    .S(_1373_),
    .X(_0548_));
 sg13g2_mux2_1 _4239_ (.A0(net722),
    .A1(net1221),
    .S(_1373_),
    .X(_0549_));
 sg13g2_mux2_1 _4240_ (.A0(net739),
    .A1(net1220),
    .S(_1373_),
    .X(_0550_));
 sg13g2_mux2_1 _4241_ (.A0(net815),
    .A1(net1219),
    .S(_1373_),
    .X(_0551_));
 sg13g2_mux2_1 _4242_ (.A0(net825),
    .A1(net1218),
    .S(_1373_),
    .X(_0552_));
 sg13g2_mux2_1 _4243_ (.A0(net747),
    .A1(net1217),
    .S(_1373_),
    .X(_0553_));
 sg13g2_mux2_1 _4244_ (.A0(net838),
    .A1(net1216),
    .S(_1373_),
    .X(_0554_));
 sg13g2_nor3_2 _4245_ (.A(net1227),
    .B(_1229_),
    .C(_1231_),
    .Y(_1374_));
 sg13g2_mux2_1 _4246_ (.A0(net752),
    .A1(net1223),
    .S(_1374_),
    .X(_0555_));
 sg13g2_mux2_1 _4247_ (.A0(net724),
    .A1(net1222),
    .S(_1374_),
    .X(_0556_));
 sg13g2_mux2_1 _4248_ (.A0(net758),
    .A1(net1221),
    .S(_1374_),
    .X(_0557_));
 sg13g2_mux2_1 _4249_ (.A0(net1334),
    .A1(net1220),
    .S(_1374_),
    .X(_0558_));
 sg13g2_mux2_1 _4250_ (.A0(net726),
    .A1(net1219),
    .S(_1374_),
    .X(_0559_));
 sg13g2_mux2_1 _4251_ (.A0(net1287),
    .A1(net1218),
    .S(_1374_),
    .X(_0560_));
 sg13g2_mux2_1 _4252_ (.A0(net693),
    .A1(net1217),
    .S(_1374_),
    .X(_0561_));
 sg13g2_mux2_1 _4253_ (.A0(net817),
    .A1(net1216),
    .S(_1374_),
    .X(_0562_));
 sg13g2_nor3_2 _4254_ (.A(net1226),
    .B(_1231_),
    .C(_1240_),
    .Y(_1375_));
 sg13g2_mux2_1 _4255_ (.A0(net777),
    .A1(net1223),
    .S(_1375_),
    .X(_0563_));
 sg13g2_mux2_1 _4256_ (.A0(net884),
    .A1(net1222),
    .S(_1375_),
    .X(_0564_));
 sg13g2_mux2_1 _4257_ (.A0(net1347),
    .A1(net1221),
    .S(_1375_),
    .X(_0565_));
 sg13g2_mux2_1 _4258_ (.A0(net737),
    .A1(net1220),
    .S(_1375_),
    .X(_0566_));
 sg13g2_mux2_1 _4259_ (.A0(net865),
    .A1(net1219),
    .S(_1375_),
    .X(_0567_));
 sg13g2_mux2_1 _4260_ (.A0(net788),
    .A1(net1218),
    .S(_1375_),
    .X(_0568_));
 sg13g2_mux2_1 _4261_ (.A0(net849),
    .A1(net1217),
    .S(_1375_),
    .X(_0569_));
 sg13g2_mux2_1 _4262_ (.A0(net818),
    .A1(net1216),
    .S(_1375_),
    .X(_0570_));
 sg13g2_nor3_2 _4263_ (.A(net1227),
    .B(_1231_),
    .C(_1240_),
    .Y(_1376_));
 sg13g2_mux2_1 _4264_ (.A0(net929),
    .A1(net1223),
    .S(_1376_),
    .X(_0571_));
 sg13g2_mux2_1 _4265_ (.A0(net743),
    .A1(net1222),
    .S(_1376_),
    .X(_0572_));
 sg13g2_mux2_1 _4266_ (.A0(net720),
    .A1(net1221),
    .S(_1376_),
    .X(_0573_));
 sg13g2_mux2_1 _4267_ (.A0(net937),
    .A1(net1220),
    .S(_1376_),
    .X(_0574_));
 sg13g2_mux2_1 _4268_ (.A0(net773),
    .A1(net1219),
    .S(_1376_),
    .X(_0575_));
 sg13g2_mux2_1 _4269_ (.A0(net819),
    .A1(net1218),
    .S(_1376_),
    .X(_0576_));
 sg13g2_mux2_1 _4270_ (.A0(net837),
    .A1(net1217),
    .S(_1376_),
    .X(_0577_));
 sg13g2_mux2_1 _4271_ (.A0(net850),
    .A1(net1216),
    .S(_1376_),
    .X(_0578_));
 sg13g2_nor3_2 _4272_ (.A(net1227),
    .B(_1231_),
    .C(_1246_),
    .Y(_1377_));
 sg13g2_mux2_1 _4273_ (.A0(net879),
    .A1(net1223),
    .S(_1377_),
    .X(_0579_));
 sg13g2_mux2_1 _4274_ (.A0(net750),
    .A1(net1222),
    .S(_1377_),
    .X(_0580_));
 sg13g2_mux2_1 _4275_ (.A0(net796),
    .A1(net1221),
    .S(_1377_),
    .X(_0581_));
 sg13g2_mux2_1 _4276_ (.A0(net863),
    .A1(net1220),
    .S(_1377_),
    .X(_0582_));
 sg13g2_mux2_1 _4277_ (.A0(net696),
    .A1(net1219),
    .S(_1377_),
    .X(_0583_));
 sg13g2_mux2_1 _4278_ (.A0(net654),
    .A1(net1218),
    .S(_1377_),
    .X(_0584_));
 sg13g2_mux2_1 _4279_ (.A0(net1483),
    .A1(net1217),
    .S(_1377_),
    .X(_0585_));
 sg13g2_mux2_1 _4280_ (.A0(net1355),
    .A1(net1216),
    .S(_1377_),
    .X(_0586_));
 sg13g2_nor3_2 _4281_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(_1231_),
    .C(_1237_),
    .Y(_1378_));
 sg13g2_mux2_1 _4282_ (.A0(net626),
    .A1(net1223),
    .S(_1378_),
    .X(_0587_));
 sg13g2_mux2_1 _4283_ (.A0(net614),
    .A1(\spi_wrapper_i.reg_data_o[1] ),
    .S(_1378_),
    .X(_0588_));
 sg13g2_mux2_1 _4284_ (.A0(net606),
    .A1(\spi_wrapper_i.reg_data_o[2] ),
    .S(_1378_),
    .X(_0589_));
 sg13g2_mux2_1 _4285_ (.A0(net608),
    .A1(net1220),
    .S(_1378_),
    .X(_0590_));
 sg13g2_mux2_1 _4286_ (.A0(net620),
    .A1(net1219),
    .S(_1378_),
    .X(_0591_));
 sg13g2_mux2_1 _4287_ (.A0(net610),
    .A1(net1218),
    .S(_1378_),
    .X(_0592_));
 sg13g2_mux2_1 _4288_ (.A0(net587),
    .A1(net1217),
    .S(_1378_),
    .X(_0593_));
 sg13g2_mux2_1 _4289_ (.A0(net616),
    .A1(net1216),
    .S(_1378_),
    .X(_0594_));
 sg13g2_and2_1 _4290_ (.A(net1238),
    .B(_1370_),
    .X(_1379_));
 sg13g2_nand2_2 _4291_ (.Y(_1380_),
    .A(net1238),
    .B(_1370_));
 sg13g2_nor4_1 _4292_ (.A(\tdc_inst.coarse_count[29] ),
    .B(\tdc_inst.coarse_count[28] ),
    .C(\tdc_inst.coarse_count[30] ),
    .D(\tdc_inst.coarse_count[31] ),
    .Y(_1381_));
 sg13g2_nor4_1 _4293_ (.A(\tdc_inst.coarse_count[25] ),
    .B(\tdc_inst.coarse_count[24] ),
    .C(\tdc_inst.coarse_count[27] ),
    .D(\tdc_inst.coarse_count[26] ),
    .Y(_1382_));
 sg13g2_nor4_1 _4294_ (.A(\tdc_inst.coarse_count[21] ),
    .B(\tdc_inst.coarse_count[20] ),
    .C(\tdc_inst.coarse_count[23] ),
    .D(\tdc_inst.coarse_count[22] ),
    .Y(_1383_));
 sg13g2_nand3_1 _4295_ (.B(_1382_),
    .C(_1383_),
    .A(_1381_),
    .Y(_1384_));
 sg13g2_nor4_2 _4296_ (.A(_0720_),
    .B(\tdc_inst.coarse_count[1] ),
    .C(\tdc_inst.coarse_count[3] ),
    .Y(_1385_),
    .D(\tdc_inst.coarse_count[2] ));
 sg13g2_nand3b_1 _4297_ (.B(_1385_),
    .C(\tdc_inst.stop_signal_sampling_clock_level ),
    .Y(_1386_),
    .A_N(\tdc_inst.start_signal_sampling_clock_level ));
 sg13g2_nor4_1 _4298_ (.A(\tdc_inst.coarse_count[9] ),
    .B(\tdc_inst.coarse_count[8] ),
    .C(\tdc_inst.coarse_count[11] ),
    .D(\tdc_inst.coarse_count[10] ),
    .Y(_1387_));
 sg13g2_nor4_1 _4299_ (.A(\tdc_inst.coarse_count[5] ),
    .B(\tdc_inst.coarse_count[4] ),
    .C(\tdc_inst.coarse_count[7] ),
    .D(\tdc_inst.coarse_count[6] ),
    .Y(_1388_));
 sg13g2_nor4_1 _4300_ (.A(\tdc_inst.coarse_count[16] ),
    .B(\tdc_inst.coarse_count[17] ),
    .C(\tdc_inst.coarse_count[19] ),
    .D(\tdc_inst.coarse_count[18] ),
    .Y(_1389_));
 sg13g2_nor4_1 _4301_ (.A(\tdc_inst.coarse_count[13] ),
    .B(\tdc_inst.coarse_count[12] ),
    .C(\tdc_inst.coarse_count[15] ),
    .D(\tdc_inst.coarse_count[14] ),
    .Y(_1390_));
 sg13g2_nand4_1 _4302_ (.B(_1388_),
    .C(_1389_),
    .A(_1387_),
    .Y(_1391_),
    .D(_1390_));
 sg13g2_nor3_2 _4303_ (.A(_1384_),
    .B(_1386_),
    .C(_1391_),
    .Y(_1392_));
 sg13g2_xnor2_1 _4304_ (.Y(_1393_),
    .A(_0044_),
    .B(_1392_));
 sg13g2_a22oi_1 _4305_ (.Y(_1394_),
    .B1(_1393_),
    .B2(net965),
    .A2(net959),
    .A1(net571));
 sg13g2_inv_1 _4306_ (.Y(_0595_),
    .A(_1394_));
 sg13g2_a22oi_1 _4307_ (.Y(_1395_),
    .B1(net959),
    .B2(net547),
    .A2(net965),
    .A1(\tdc_inst.coarse_count[1] ));
 sg13g2_inv_1 _4308_ (.Y(_0596_),
    .A(_1395_));
 sg13g2_a22oi_1 _4309_ (.Y(_1396_),
    .B1(net957),
    .B2(net551),
    .A2(net965),
    .A1(\tdc_inst.coarse_count[2] ));
 sg13g2_inv_1 _4310_ (.Y(_0597_),
    .A(_1396_));
 sg13g2_a22oi_1 _4311_ (.Y(_1397_),
    .B1(net957),
    .B2(net546),
    .A2(net965),
    .A1(\tdc_inst.coarse_count[3] ));
 sg13g2_inv_1 _4312_ (.Y(_0598_),
    .A(_1397_));
 sg13g2_a22oi_1 _4313_ (.Y(_1398_),
    .B1(net957),
    .B2(net550),
    .A2(net963),
    .A1(\tdc_inst.coarse_count[4] ));
 sg13g2_inv_1 _4314_ (.Y(_0599_),
    .A(_1398_));
 sg13g2_a22oi_1 _4315_ (.Y(_1399_),
    .B1(net956),
    .B2(net549),
    .A2(net963),
    .A1(\tdc_inst.coarse_count[5] ));
 sg13g2_inv_1 _4316_ (.Y(_0600_),
    .A(_1399_));
 sg13g2_a22oi_1 _4317_ (.Y(_1400_),
    .B1(net956),
    .B2(net548),
    .A2(net963),
    .A1(\tdc_inst.coarse_count[6] ));
 sg13g2_inv_1 _4318_ (.Y(_0601_),
    .A(_1400_));
 sg13g2_a22oi_1 _4319_ (.Y(_1401_),
    .B1(net957),
    .B2(net554),
    .A2(net963),
    .A1(\tdc_inst.coarse_count[7] ));
 sg13g2_inv_1 _4320_ (.Y(_0602_),
    .A(_1401_));
 sg13g2_a22oi_1 _4321_ (.Y(_1402_),
    .B1(net957),
    .B2(net641),
    .A2(net962),
    .A1(\tdc_inst.coarse_count[8] ));
 sg13g2_inv_1 _4322_ (.Y(_0603_),
    .A(_1402_));
 sg13g2_a22oi_1 _4323_ (.Y(_1403_),
    .B1(net959),
    .B2(net562),
    .A2(net965),
    .A1(\tdc_inst.coarse_count[9] ));
 sg13g2_inv_1 _4324_ (.Y(_0604_),
    .A(_1403_));
 sg13g2_a22oi_1 _4325_ (.Y(_1404_),
    .B1(net956),
    .B2(net656),
    .A2(net963),
    .A1(\tdc_inst.coarse_count[10] ));
 sg13g2_inv_1 _4326_ (.Y(_0605_),
    .A(_1404_));
 sg13g2_a22oi_1 _4327_ (.Y(_1405_),
    .B1(net957),
    .B2(net593),
    .A2(net962),
    .A1(\tdc_inst.coarse_count[11] ));
 sg13g2_inv_1 _4328_ (.Y(_0606_),
    .A(_1405_));
 sg13g2_a22oi_1 _4329_ (.Y(_1406_),
    .B1(net956),
    .B2(net592),
    .A2(net962),
    .A1(\tdc_inst.coarse_count[12] ));
 sg13g2_inv_1 _4330_ (.Y(_0607_),
    .A(_1406_));
 sg13g2_a22oi_1 _4331_ (.Y(_1407_),
    .B1(net956),
    .B2(net561),
    .A2(net963),
    .A1(\tdc_inst.coarse_count[13] ));
 sg13g2_inv_1 _4332_ (.Y(_0608_),
    .A(_1407_));
 sg13g2_nor2b_1 _4333_ (.A(_0039_),
    .B_N(_1392_),
    .Y(_1408_));
 sg13g2_o21ai_1 _4334_ (.B1(net962),
    .Y(_1409_),
    .A1(\tdc_inst.coarse_count[14] ),
    .A2(_1408_));
 sg13g2_o21ai_1 _4335_ (.B1(_1409_),
    .Y(_0609_),
    .A1(_0719_),
    .A2(_1380_));
 sg13g2_a22oi_1 _4336_ (.Y(_1410_),
    .B1(net957),
    .B2(net566),
    .A2(net966),
    .A1(\tdc_inst.coarse_count[15] ));
 sg13g2_inv_1 _4337_ (.Y(_0610_),
    .A(_1410_));
 sg13g2_a22oi_1 _4338_ (.Y(_1411_),
    .B1(net959),
    .B2(net570),
    .A2(net965),
    .A1(\tdc_inst.coarse_count[16] ));
 sg13g2_inv_1 _4339_ (.Y(_0611_),
    .A(_1411_));
 sg13g2_a22oi_1 _4340_ (.Y(_1412_),
    .B1(net956),
    .B2(net557),
    .A2(net962),
    .A1(\tdc_inst.coarse_count[17] ));
 sg13g2_inv_1 _4341_ (.Y(_0612_),
    .A(_1412_));
 sg13g2_nor2b_1 _4342_ (.A(_0040_),
    .B_N(_1392_),
    .Y(_1413_));
 sg13g2_o21ai_1 _4343_ (.B1(net962),
    .Y(_1414_),
    .A1(\tdc_inst.coarse_count[18] ),
    .A2(_1413_));
 sg13g2_o21ai_1 _4344_ (.B1(_1414_),
    .Y(_0613_),
    .A1(_0718_),
    .A2(_1380_));
 sg13g2_a22oi_1 _4345_ (.Y(_1415_),
    .B1(net956),
    .B2(net589),
    .A2(net962),
    .A1(\tdc_inst.coarse_count[19] ));
 sg13g2_inv_1 _4346_ (.Y(_0614_),
    .A(_1415_));
 sg13g2_a22oi_1 _4347_ (.Y(_1416_),
    .B1(net956),
    .B2(net572),
    .A2(net962),
    .A1(\tdc_inst.coarse_count[20] ));
 sg13g2_inv_1 _4348_ (.Y(_0615_),
    .A(_1416_));
 sg13g2_a22oi_1 _4349_ (.Y(_1417_),
    .B1(net958),
    .B2(net560),
    .A2(net960),
    .A1(\tdc_inst.coarse_count[21] ));
 sg13g2_inv_1 _4350_ (.Y(_0616_),
    .A(_1417_));
 sg13g2_nor2b_1 _4351_ (.A(_0041_),
    .B_N(_1392_),
    .Y(_1418_));
 sg13g2_o21ai_1 _4352_ (.B1(net960),
    .Y(_1419_),
    .A1(\tdc_inst.coarse_count[22] ),
    .A2(_1418_));
 sg13g2_o21ai_1 _4353_ (.B1(_1419_),
    .Y(_0617_),
    .A1(_0717_),
    .A2(_1380_));
 sg13g2_a22oi_1 _4354_ (.Y(_1420_),
    .B1(net958),
    .B2(net565),
    .A2(net960),
    .A1(\tdc_inst.coarse_count[23] ));
 sg13g2_inv_1 _4355_ (.Y(_0618_),
    .A(_1420_));
 sg13g2_a22oi_1 _4356_ (.Y(_1421_),
    .B1(net958),
    .B2(net647),
    .A2(net960),
    .A1(\tdc_inst.coarse_count[24] ));
 sg13g2_inv_1 _4357_ (.Y(_0619_),
    .A(_1421_));
 sg13g2_dfrbp_1 _4358_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net316),
    .D(_0047_),
    .Q_N(_2248_),
    .Q(\tdc_inst.start_count_debug[0] ));
 sg13g2_dfrbp_1 _4359_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net73),
    .D(_0048_),
    .Q_N(_2247_),
    .Q(\tdc_inst.start_count_debug[1] ));
 sg13g2_dfrbp_1 _4360_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net72),
    .D(_0049_),
    .Q_N(_2246_),
    .Q(\tdc_inst.start_count_debug[2] ));
 sg13g2_dfrbp_1 _4361_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net71),
    .D(_0050_),
    .Q_N(_2245_),
    .Q(\tdc_inst.start_count_debug[3] ));
 sg13g2_dfrbp_1 _4362_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net70),
    .D(_0051_),
    .Q_N(_2244_),
    .Q(\tdc_inst.start_count_debug[4] ));
 sg13g2_dfrbp_1 _4363_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net69),
    .D(_0052_),
    .Q_N(_2243_),
    .Q(\tdc_inst.start_count_debug[5] ));
 sg13g2_dfrbp_1 _4364_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net68),
    .D(_0053_),
    .Q_N(_2242_),
    .Q(\tdc_inst.start_count_debug[6] ));
 sg13g2_dfrbp_1 _4365_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net67),
    .D(_0054_),
    .Q_N(_2241_),
    .Q(\tdc_inst.start_count_debug[7] ));
 sg13g2_dfrbp_1 _4366_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net66),
    .D(_0055_),
    .Q_N(_2240_),
    .Q(\tdc_inst.start_count_debug[8] ));
 sg13g2_dfrbp_1 _4367_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net65),
    .D(_0056_),
    .Q_N(_2239_),
    .Q(\tdc_inst.start_count_debug[9] ));
 sg13g2_dfrbp_1 _4368_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net64),
    .D(_0057_),
    .Q_N(_2238_),
    .Q(\tdc_inst.start_count_debug[10] ));
 sg13g2_dfrbp_1 _4369_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net63),
    .D(_0058_),
    .Q_N(_2237_),
    .Q(\tdc_inst.start_count_debug[11] ));
 sg13g2_dfrbp_1 _4370_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net62),
    .D(_0059_),
    .Q_N(_2236_),
    .Q(\tdc_inst.start_count_debug[12] ));
 sg13g2_dfrbp_1 _4371_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net61),
    .D(_0060_),
    .Q_N(_2235_),
    .Q(\tdc_inst.start_count_debug[13] ));
 sg13g2_dfrbp_1 _4372_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net60),
    .D(_0061_),
    .Q_N(_2234_),
    .Q(\tdc_inst.start_count_debug[14] ));
 sg13g2_dfrbp_1 _4373_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net59),
    .D(_0062_),
    .Q_N(_2233_),
    .Q(\tdc_inst.start_count_debug[15] ));
 sg13g2_dfrbp_1 _4374_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net58),
    .D(_0063_),
    .Q_N(_2232_),
    .Q(\tdc_inst.start_count_debug[16] ));
 sg13g2_dfrbp_1 _4375_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net57),
    .D(_0064_),
    .Q_N(_2231_),
    .Q(\tdc_inst.start_count_debug[17] ));
 sg13g2_dfrbp_1 _4376_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net56),
    .D(_0065_),
    .Q_N(_2230_),
    .Q(\tdc_inst.start_count_debug[18] ));
 sg13g2_dfrbp_1 _4377_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net55),
    .D(_0066_),
    .Q_N(_2229_),
    .Q(\tdc_inst.start_count_debug[19] ));
 sg13g2_dfrbp_1 _4378_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net54),
    .D(_0067_),
    .Q_N(_2228_),
    .Q(\tdc_inst.start_count_debug[20] ));
 sg13g2_dfrbp_1 _4379_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net53),
    .D(_0068_),
    .Q_N(_2227_),
    .Q(\tdc_inst.start_count_debug[21] ));
 sg13g2_dfrbp_1 _4380_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net52),
    .D(_0069_),
    .Q_N(_2226_),
    .Q(\tdc_inst.start_count_debug[22] ));
 sg13g2_dfrbp_1 _4381_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net51),
    .D(_0070_),
    .Q_N(_2225_),
    .Q(\tdc_inst.start_count_debug[23] ));
 sg13g2_dfrbp_1 _4382_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net50),
    .D(_0071_),
    .Q_N(_2224_),
    .Q(\tdc_inst.start_count_debug[24] ));
 sg13g2_dfrbp_1 _4383_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net49),
    .D(_0072_),
    .Q_N(_2223_),
    .Q(\tdc_inst.start_count_debug[25] ));
 sg13g2_dfrbp_1 _4384_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net48),
    .D(_0073_),
    .Q_N(_2222_),
    .Q(\tdc_inst.start_count_debug[26] ));
 sg13g2_dfrbp_1 _4385_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net47),
    .D(_0074_),
    .Q_N(_2221_),
    .Q(\tdc_inst.start_count_debug[27] ));
 sg13g2_dfrbp_1 _4386_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net46),
    .D(_0075_),
    .Q_N(_2220_),
    .Q(\tdc_inst.start_count_debug[28] ));
 sg13g2_dfrbp_1 _4387_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net45),
    .D(_0076_),
    .Q_N(_2219_),
    .Q(\tdc_inst.start_count_debug[29] ));
 sg13g2_dfrbp_1 _4388_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net44),
    .D(_0077_),
    .Q_N(_2218_),
    .Q(\tdc_inst.start_count_debug[30] ));
 sg13g2_dfrbp_1 _4389_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net43),
    .D(_0078_),
    .Q_N(_2217_),
    .Q(\tdc_inst.start_count_debug[31] ));
 sg13g2_dfrbp_1 _4390_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net42),
    .D(_0079_),
    .Q_N(_2216_),
    .Q(\tdc_inst.start_count_debug[32] ));
 sg13g2_dfrbp_1 _4391_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net41),
    .D(_0080_),
    .Q_N(_2215_),
    .Q(\tdc_inst.start_count_debug[33] ));
 sg13g2_dfrbp_1 _4392_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net40),
    .D(_0081_),
    .Q_N(_2214_),
    .Q(\tdc_inst.start_count_debug[34] ));
 sg13g2_dfrbp_1 _4393_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net39),
    .D(_0082_),
    .Q_N(_2213_),
    .Q(\tdc_inst.start_count_debug[35] ));
 sg13g2_dfrbp_1 _4394_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net38),
    .D(_0083_),
    .Q_N(_2212_),
    .Q(\tdc_inst.start_count_debug[36] ));
 sg13g2_dfrbp_1 _4395_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net37),
    .D(_0084_),
    .Q_N(_2211_),
    .Q(\tdc_inst.start_count_debug[37] ));
 sg13g2_dfrbp_1 _4396_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net36),
    .D(_0085_),
    .Q_N(_2210_),
    .Q(\tdc_inst.start_count_debug[38] ));
 sg13g2_dfrbp_1 _4397_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net35),
    .D(_0086_),
    .Q_N(_2209_),
    .Q(\tdc_inst.start_count_debug[39] ));
 sg13g2_dfrbp_1 _4398_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net34),
    .D(_0087_),
    .Q_N(_2208_),
    .Q(\tdc_inst.start_count_debug[40] ));
 sg13g2_dfrbp_1 _4399_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net33),
    .D(_0088_),
    .Q_N(_2207_),
    .Q(\tdc_inst.start_count_debug[41] ));
 sg13g2_dfrbp_1 _4400_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net32),
    .D(_0089_),
    .Q_N(_2206_),
    .Q(\tdc_inst.start_count_debug[42] ));
 sg13g2_dfrbp_1 _4401_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net31),
    .D(_0090_),
    .Q_N(_2205_),
    .Q(\tdc_inst.start_count_debug[43] ));
 sg13g2_dfrbp_1 _4402_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net30),
    .D(_0091_),
    .Q_N(_2204_),
    .Q(\tdc_inst.start_count_debug[44] ));
 sg13g2_dfrbp_1 _4403_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net29),
    .D(_0092_),
    .Q_N(_2203_),
    .Q(\tdc_inst.start_count_debug[45] ));
 sg13g2_dfrbp_1 _4404_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net28),
    .D(_0093_),
    .Q_N(_2202_),
    .Q(\tdc_inst.start_count_debug[46] ));
 sg13g2_dfrbp_1 _4405_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net27),
    .D(_0094_),
    .Q_N(_2201_),
    .Q(\tdc_inst.start_count_debug[47] ));
 sg13g2_dfrbp_1 _4406_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net26),
    .D(_0095_),
    .Q_N(_2200_),
    .Q(\tdc_inst.start_count_debug[48] ));
 sg13g2_dfrbp_1 _4407_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net25),
    .D(_0096_),
    .Q_N(_2199_),
    .Q(\tdc_inst.start_count_debug[49] ));
 sg13g2_dfrbp_1 _4408_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net540),
    .D(_0097_),
    .Q_N(_2198_),
    .Q(\tdc_inst.start_count_debug[50] ));
 sg13g2_dfrbp_1 _4409_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net539),
    .D(_0098_),
    .Q_N(_2197_),
    .Q(\tdc_inst.start_count_debug[51] ));
 sg13g2_dfrbp_1 _4410_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net538),
    .D(_0099_),
    .Q_N(_2196_),
    .Q(\tdc_inst.start_count_debug[52] ));
 sg13g2_dfrbp_1 _4411_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net537),
    .D(_0100_),
    .Q_N(_2195_),
    .Q(\tdc_inst.start_count_debug[53] ));
 sg13g2_dfrbp_1 _4412_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net536),
    .D(_0101_),
    .Q_N(_2194_),
    .Q(\tdc_inst.start_count_debug[54] ));
 sg13g2_dfrbp_1 _4413_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net535),
    .D(_0102_),
    .Q_N(_2193_),
    .Q(\tdc_inst.start_count_debug[55] ));
 sg13g2_dfrbp_1 _4414_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net534),
    .D(_0103_),
    .Q_N(_2192_),
    .Q(\tdc_inst.start_count_debug[56] ));
 sg13g2_dfrbp_1 _4415_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net533),
    .D(_0104_),
    .Q_N(_2191_),
    .Q(\tdc_inst.start_count_debug[57] ));
 sg13g2_dfrbp_1 _4416_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net532),
    .D(_0105_),
    .Q_N(_2190_),
    .Q(\tdc_inst.start_count_debug[58] ));
 sg13g2_dfrbp_1 _4417_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net531),
    .D(_0106_),
    .Q_N(_2189_),
    .Q(\tdc_inst.start_count_debug[59] ));
 sg13g2_dfrbp_1 _4418_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net530),
    .D(_0107_),
    .Q_N(_2188_),
    .Q(\tdc_inst.start_count_debug[60] ));
 sg13g2_dfrbp_1 _4419_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net529),
    .D(_0108_),
    .Q_N(_2187_),
    .Q(\tdc_inst.start_count_debug[61] ));
 sg13g2_dfrbp_1 _4420_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net528),
    .D(_0109_),
    .Q_N(_2186_),
    .Q(\tdc_inst.start_count_debug[62] ));
 sg13g2_dfrbp_1 _4421_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net527),
    .D(_0110_),
    .Q_N(_2185_),
    .Q(\tdc_inst.start_count_debug[63] ));
 sg13g2_dfrbp_1 _4422_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net526),
    .D(_0111_),
    .Q_N(_2184_),
    .Q(\tdc_inst.start_count_debug[64] ));
 sg13g2_dfrbp_1 _4423_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net525),
    .D(_0112_),
    .Q_N(_2183_),
    .Q(\tdc_inst.start_count_debug[65] ));
 sg13g2_dfrbp_1 _4424_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net524),
    .D(_0113_),
    .Q_N(_2182_),
    .Q(\tdc_inst.start_count_debug[66] ));
 sg13g2_dfrbp_1 _4425_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net523),
    .D(_0114_),
    .Q_N(_2181_),
    .Q(\tdc_inst.start_count_debug[67] ));
 sg13g2_dfrbp_1 _4426_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net522),
    .D(_0115_),
    .Q_N(_2180_),
    .Q(\tdc_inst.start_count_debug[68] ));
 sg13g2_dfrbp_1 _4427_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net521),
    .D(_0116_),
    .Q_N(_2179_),
    .Q(\tdc_inst.start_count_debug[69] ));
 sg13g2_dfrbp_1 _4428_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net520),
    .D(_0117_),
    .Q_N(_2178_),
    .Q(\tdc_inst.start_count_debug[70] ));
 sg13g2_dfrbp_1 _4429_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net519),
    .D(_0118_),
    .Q_N(_2177_),
    .Q(\tdc_inst.start_count_debug[71] ));
 sg13g2_dfrbp_1 _4430_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net518),
    .D(_0119_),
    .Q_N(_2176_),
    .Q(\tdc_inst.start_count_debug[72] ));
 sg13g2_dfrbp_1 _4431_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net517),
    .D(_0120_),
    .Q_N(_2175_),
    .Q(\tdc_inst.start_count_debug[73] ));
 sg13g2_dfrbp_1 _4432_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net516),
    .D(_0121_),
    .Q_N(_2174_),
    .Q(\tdc_inst.start_count_debug[74] ));
 sg13g2_dfrbp_1 _4433_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net515),
    .D(_0122_),
    .Q_N(_2173_),
    .Q(\tdc_inst.start_count_debug[75] ));
 sg13g2_dfrbp_1 _4434_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net514),
    .D(_0123_),
    .Q_N(_2172_),
    .Q(\tdc_inst.start_count_debug[76] ));
 sg13g2_dfrbp_1 _4435_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net513),
    .D(_0124_),
    .Q_N(_2171_),
    .Q(\tdc_inst.start_count_debug[77] ));
 sg13g2_dfrbp_1 _4436_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net512),
    .D(_0125_),
    .Q_N(_2170_),
    .Q(\tdc_inst.start_count_debug[78] ));
 sg13g2_dfrbp_1 _4437_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net511),
    .D(_0126_),
    .Q_N(_2169_),
    .Q(\tdc_inst.start_count_debug[79] ));
 sg13g2_dfrbp_1 _4438_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net510),
    .D(_0127_),
    .Q_N(_2168_),
    .Q(\tdc_inst.start_count_debug[80] ));
 sg13g2_dfrbp_1 _4439_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net509),
    .D(_0128_),
    .Q_N(_2167_),
    .Q(\tdc_inst.start_count_debug[81] ));
 sg13g2_dfrbp_1 _4440_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net508),
    .D(_0129_),
    .Q_N(_2166_),
    .Q(\tdc_inst.start_count_debug[82] ));
 sg13g2_dfrbp_1 _4441_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net507),
    .D(_0130_),
    .Q_N(_2165_),
    .Q(\tdc_inst.start_count_debug[83] ));
 sg13g2_dfrbp_1 _4442_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net506),
    .D(_0131_),
    .Q_N(_2164_),
    .Q(\tdc_inst.start_count_debug[84] ));
 sg13g2_dfrbp_1 _4443_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net505),
    .D(_0132_),
    .Q_N(_2163_),
    .Q(\tdc_inst.start_count_debug[85] ));
 sg13g2_dfrbp_1 _4444_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net504),
    .D(_0133_),
    .Q_N(_2162_),
    .Q(\tdc_inst.start_count_debug[86] ));
 sg13g2_dfrbp_1 _4445_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net503),
    .D(_0134_),
    .Q_N(_2161_),
    .Q(\tdc_inst.start_count_debug[87] ));
 sg13g2_dfrbp_1 _4446_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net502),
    .D(_0135_),
    .Q_N(_2160_),
    .Q(\tdc_inst.start_count_debug[88] ));
 sg13g2_dfrbp_1 _4447_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net501),
    .D(_0136_),
    .Q_N(_2159_),
    .Q(\tdc_inst.start_count_debug[89] ));
 sg13g2_dfrbp_1 _4448_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net500),
    .D(_0137_),
    .Q_N(_2158_),
    .Q(\tdc_inst.start_count_debug[90] ));
 sg13g2_dfrbp_1 _4449_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net499),
    .D(_0138_),
    .Q_N(_2157_),
    .Q(\tdc_inst.start_count_debug[91] ));
 sg13g2_dfrbp_1 _4450_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net498),
    .D(_0139_),
    .Q_N(_2156_),
    .Q(\tdc_inst.start_count_debug[92] ));
 sg13g2_dfrbp_1 _4451_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net497),
    .D(_0140_),
    .Q_N(_2155_),
    .Q(\tdc_inst.start_count_debug[93] ));
 sg13g2_dfrbp_1 _4452_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net496),
    .D(_0141_),
    .Q_N(_2154_),
    .Q(\tdc_inst.start_count_debug[94] ));
 sg13g2_dfrbp_1 _4453_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net495),
    .D(_0142_),
    .Q_N(_2153_),
    .Q(\tdc_inst.start_count_debug[95] ));
 sg13g2_dfrbp_1 _4454_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net494),
    .D(_0143_),
    .Q_N(_2152_),
    .Q(\tdc_inst.start_count_debug[96] ));
 sg13g2_dfrbp_1 _4455_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net493),
    .D(_0144_),
    .Q_N(_2151_),
    .Q(\tdc_inst.start_count_debug[97] ));
 sg13g2_dfrbp_1 _4456_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net492),
    .D(_0145_),
    .Q_N(_2150_),
    .Q(\tdc_inst.start_count_debug[98] ));
 sg13g2_dfrbp_1 _4457_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net491),
    .D(_0146_),
    .Q_N(_2149_),
    .Q(\tdc_inst.start_count_debug[99] ));
 sg13g2_dfrbp_1 _4458_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net490),
    .D(_0147_),
    .Q_N(_2148_),
    .Q(\tdc_inst.start_count_debug[100] ));
 sg13g2_dfrbp_1 _4459_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net489),
    .D(_0148_),
    .Q_N(_2147_),
    .Q(\tdc_inst.start_count_debug[101] ));
 sg13g2_dfrbp_1 _4460_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net488),
    .D(_0149_),
    .Q_N(_2146_),
    .Q(\tdc_inst.start_count_debug[102] ));
 sg13g2_dfrbp_1 _4461_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net487),
    .D(_0150_),
    .Q_N(_2145_),
    .Q(\tdc_inst.start_count_debug[103] ));
 sg13g2_dfrbp_1 _4462_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net486),
    .D(_0151_),
    .Q_N(_2144_),
    .Q(\tdc_inst.start_count_debug[104] ));
 sg13g2_dfrbp_1 _4463_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net485),
    .D(_0152_),
    .Q_N(_2143_),
    .Q(\tdc_inst.start_count_debug[105] ));
 sg13g2_dfrbp_1 _4464_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net484),
    .D(_0153_),
    .Q_N(_2142_),
    .Q(\tdc_inst.start_count_debug[106] ));
 sg13g2_dfrbp_1 _4465_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net483),
    .D(_0154_),
    .Q_N(_2141_),
    .Q(\tdc_inst.start_count_debug[107] ));
 sg13g2_dfrbp_1 _4466_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net482),
    .D(_0155_),
    .Q_N(_2140_),
    .Q(\tdc_inst.start_count_debug[108] ));
 sg13g2_dfrbp_1 _4467_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net481),
    .D(_0156_),
    .Q_N(_2139_),
    .Q(\tdc_inst.start_count_debug[109] ));
 sg13g2_dfrbp_1 _4468_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net480),
    .D(_0157_),
    .Q_N(_2138_),
    .Q(\tdc_inst.start_count_debug[110] ));
 sg13g2_dfrbp_1 _4469_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net479),
    .D(_0158_),
    .Q_N(_2137_),
    .Q(\tdc_inst.start_count_debug[111] ));
 sg13g2_dfrbp_1 _4470_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net478),
    .D(_0159_),
    .Q_N(_2136_),
    .Q(\tdc_inst.start_count_debug[112] ));
 sg13g2_dfrbp_1 _4471_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net477),
    .D(_0160_),
    .Q_N(_2135_),
    .Q(\tdc_inst.start_count_debug[113] ));
 sg13g2_dfrbp_1 _4472_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net476),
    .D(_0161_),
    .Q_N(_2134_),
    .Q(\tdc_inst.start_count_debug[114] ));
 sg13g2_dfrbp_1 _4473_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net475),
    .D(_0162_),
    .Q_N(_2133_),
    .Q(\tdc_inst.start_count_debug[115] ));
 sg13g2_dfrbp_1 _4474_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net474),
    .D(_0163_),
    .Q_N(_2132_),
    .Q(\tdc_inst.start_count_debug[116] ));
 sg13g2_dfrbp_1 _4475_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net473),
    .D(_0164_),
    .Q_N(_2131_),
    .Q(\tdc_inst.start_count_debug[117] ));
 sg13g2_dfrbp_1 _4476_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net472),
    .D(_0165_),
    .Q_N(_2130_),
    .Q(\tdc_inst.start_count_debug[118] ));
 sg13g2_dfrbp_1 _4477_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net471),
    .D(_0166_),
    .Q_N(_2129_),
    .Q(\tdc_inst.start_count_debug[119] ));
 sg13g2_dfrbp_1 _4478_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net470),
    .D(_0167_),
    .Q_N(_2128_),
    .Q(\tdc_inst.start_count_debug[120] ));
 sg13g2_dfrbp_1 _4479_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net469),
    .D(_0168_),
    .Q_N(_2127_),
    .Q(\tdc_inst.start_count_debug[121] ));
 sg13g2_dfrbp_1 _4480_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net468),
    .D(_0169_),
    .Q_N(_2126_),
    .Q(\tdc_inst.start_count_debug[122] ));
 sg13g2_dfrbp_1 _4481_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net467),
    .D(_0170_),
    .Q_N(_2125_),
    .Q(\tdc_inst.start_count_debug[123] ));
 sg13g2_dfrbp_1 _4482_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net466),
    .D(_0171_),
    .Q_N(_2124_),
    .Q(\tdc_inst.start_count_debug[124] ));
 sg13g2_dfrbp_1 _4483_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net465),
    .D(_0172_),
    .Q_N(_2123_),
    .Q(\tdc_inst.start_count_debug[125] ));
 sg13g2_dfrbp_1 _4484_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net464),
    .D(_0173_),
    .Q_N(_2122_),
    .Q(\tdc_inst.start_count_debug[126] ));
 sg13g2_dfrbp_1 _4485_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net463),
    .D(_0174_),
    .Q_N(_2121_),
    .Q(\tdc_inst.start_count_debug[127] ));
 sg13g2_dfrbp_1 _4486_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net462),
    .D(_0175_),
    .Q_N(_2120_),
    .Q(\tdc_inst.start_count_debug[128] ));
 sg13g2_dfrbp_1 _4487_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net461),
    .D(_0176_),
    .Q_N(_2119_),
    .Q(\tdc_inst.start_count_debug[129] ));
 sg13g2_dfrbp_1 _4488_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net460),
    .D(_0177_),
    .Q_N(_2118_),
    .Q(\tdc_inst.start_count_debug[130] ));
 sg13g2_dfrbp_1 _4489_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net459),
    .D(_0178_),
    .Q_N(_2117_),
    .Q(\tdc_inst.start_count_debug[131] ));
 sg13g2_dfrbp_1 _4490_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net458),
    .D(_0179_),
    .Q_N(_2116_),
    .Q(\tdc_inst.start_count_debug[132] ));
 sg13g2_dfrbp_1 _4491_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net457),
    .D(_0180_),
    .Q_N(_2115_),
    .Q(\tdc_inst.start_count_debug[133] ));
 sg13g2_dfrbp_1 _4492_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net456),
    .D(_0181_),
    .Q_N(_2114_),
    .Q(\tdc_inst.start_count_debug[134] ));
 sg13g2_dfrbp_1 _4493_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net455),
    .D(_0182_),
    .Q_N(_2113_),
    .Q(\tdc_inst.start_count_debug[135] ));
 sg13g2_dfrbp_1 _4494_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net454),
    .D(_0183_),
    .Q_N(_2112_),
    .Q(\tdc_inst.start_count_debug[136] ));
 sg13g2_dfrbp_1 _4495_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net453),
    .D(_0184_),
    .Q_N(_2111_),
    .Q(\tdc_inst.start_count_debug[137] ));
 sg13g2_dfrbp_1 _4496_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net452),
    .D(_0185_),
    .Q_N(_2110_),
    .Q(\tdc_inst.start_count_debug[138] ));
 sg13g2_dfrbp_1 _4497_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net451),
    .D(_0186_),
    .Q_N(_2109_),
    .Q(\tdc_inst.start_count_debug[139] ));
 sg13g2_dfrbp_1 _4498_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net450),
    .D(_0187_),
    .Q_N(_2108_),
    .Q(\tdc_inst.start_count_debug[140] ));
 sg13g2_dfrbp_1 _4499_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net449),
    .D(_0188_),
    .Q_N(_2107_),
    .Q(\tdc_inst.start_count_debug[141] ));
 sg13g2_dfrbp_1 _4500_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net448),
    .D(_0189_),
    .Q_N(_2106_),
    .Q(\tdc_inst.tdc_xor_result[0] ));
 sg13g2_dfrbp_1 _4501_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net447),
    .D(_0190_),
    .Q_N(_2105_),
    .Q(\tdc_inst.tdc_xor_result[1] ));
 sg13g2_dfrbp_1 _4502_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net446),
    .D(_0191_),
    .Q_N(_2104_),
    .Q(\tdc_inst.tdc_xor_result[2] ));
 sg13g2_dfrbp_1 _4503_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net445),
    .D(_0192_),
    .Q_N(_2103_),
    .Q(\tdc_inst.tdc_xor_result[3] ));
 sg13g2_dfrbp_1 _4504_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net444),
    .D(_0193_),
    .Q_N(_2102_),
    .Q(\tdc_inst.tdc_xor_result[4] ));
 sg13g2_dfrbp_1 _4505_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net443),
    .D(_0194_),
    .Q_N(_2101_),
    .Q(\tdc_inst.tdc_xor_result[5] ));
 sg13g2_dfrbp_1 _4506_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net442),
    .D(_0195_),
    .Q_N(_2100_),
    .Q(\tdc_inst.tdc_xor_result[6] ));
 sg13g2_dfrbp_1 _4507_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net441),
    .D(_0196_),
    .Q_N(_2099_),
    .Q(\tdc_inst.tdc_xor_result[7] ));
 sg13g2_dfrbp_1 _4508_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net440),
    .D(_0197_),
    .Q_N(_2098_),
    .Q(\tdc_inst.tdc_xor_result[8] ));
 sg13g2_dfrbp_1 _4509_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net439),
    .D(_0198_),
    .Q_N(_2097_),
    .Q(\tdc_inst.tdc_xor_result[9] ));
 sg13g2_dfrbp_1 _4510_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net438),
    .D(_0199_),
    .Q_N(_2096_),
    .Q(\tdc_inst.tdc_xor_result[10] ));
 sg13g2_dfrbp_1 _4511_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net437),
    .D(_0200_),
    .Q_N(_2095_),
    .Q(\tdc_inst.tdc_xor_result[11] ));
 sg13g2_dfrbp_1 _4512_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net436),
    .D(_0201_),
    .Q_N(_2094_),
    .Q(\tdc_inst.tdc_xor_result[12] ));
 sg13g2_dfrbp_1 _4513_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net435),
    .D(_0202_),
    .Q_N(_2093_),
    .Q(\tdc_inst.tdc_xor_result[13] ));
 sg13g2_dfrbp_1 _4514_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net434),
    .D(_0203_),
    .Q_N(_2092_),
    .Q(\tdc_inst.tdc_xor_result[14] ));
 sg13g2_dfrbp_1 _4515_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net433),
    .D(_0204_),
    .Q_N(_2091_),
    .Q(\tdc_inst.tdc_xor_result[15] ));
 sg13g2_dfrbp_1 _4516_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net432),
    .D(_0205_),
    .Q_N(_2090_),
    .Q(\tdc_inst.tdc_xor_result[16] ));
 sg13g2_dfrbp_1 _4517_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net431),
    .D(_0206_),
    .Q_N(_2089_),
    .Q(\tdc_inst.tdc_xor_result[17] ));
 sg13g2_dfrbp_1 _4518_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net430),
    .D(_0207_),
    .Q_N(_2088_),
    .Q(\tdc_inst.tdc_xor_result[18] ));
 sg13g2_dfrbp_1 _4519_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net429),
    .D(_0208_),
    .Q_N(_2087_),
    .Q(\tdc_inst.tdc_xor_result[19] ));
 sg13g2_dfrbp_1 _4520_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net428),
    .D(_0209_),
    .Q_N(_2086_),
    .Q(\tdc_inst.tdc_xor_result[20] ));
 sg13g2_dfrbp_1 _4521_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net427),
    .D(_0210_),
    .Q_N(_2085_),
    .Q(\tdc_inst.tdc_xor_result[21] ));
 sg13g2_dfrbp_1 _4522_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net426),
    .D(_0211_),
    .Q_N(_2084_),
    .Q(\tdc_inst.tdc_xor_result[22] ));
 sg13g2_dfrbp_1 _4523_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net425),
    .D(_0212_),
    .Q_N(_2083_),
    .Q(\tdc_inst.tdc_xor_result[23] ));
 sg13g2_dfrbp_1 _4524_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net424),
    .D(_0213_),
    .Q_N(_2082_),
    .Q(\tdc_inst.tdc_xor_result[24] ));
 sg13g2_dfrbp_1 _4525_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net423),
    .D(_0214_),
    .Q_N(_2081_),
    .Q(\tdc_inst.tdc_xor_result[25] ));
 sg13g2_dfrbp_1 _4526_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net422),
    .D(_0215_),
    .Q_N(_2080_),
    .Q(\tdc_inst.tdc_xor_result[26] ));
 sg13g2_dfrbp_1 _4527_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net421),
    .D(_0216_),
    .Q_N(_2079_),
    .Q(\tdc_inst.tdc_xor_result[27] ));
 sg13g2_dfrbp_1 _4528_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net420),
    .D(_0217_),
    .Q_N(_2078_),
    .Q(\tdc_inst.tdc_xor_result[28] ));
 sg13g2_dfrbp_1 _4529_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net419),
    .D(_0218_),
    .Q_N(_2077_),
    .Q(\tdc_inst.tdc_xor_result[29] ));
 sg13g2_dfrbp_1 _4530_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net418),
    .D(_0219_),
    .Q_N(_2076_),
    .Q(\tdc_inst.tdc_xor_result[30] ));
 sg13g2_dfrbp_1 _4531_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net417),
    .D(_0220_),
    .Q_N(_2075_),
    .Q(\tdc_inst.tdc_xor_result[31] ));
 sg13g2_dfrbp_1 _4532_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net416),
    .D(_0221_),
    .Q_N(_2074_),
    .Q(\tdc_inst.tdc_xor_result[32] ));
 sg13g2_dfrbp_1 _4533_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net415),
    .D(_0222_),
    .Q_N(_2073_),
    .Q(\tdc_inst.tdc_xor_result[33] ));
 sg13g2_dfrbp_1 _4534_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net414),
    .D(_0223_),
    .Q_N(_2072_),
    .Q(\tdc_inst.tdc_xor_result[34] ));
 sg13g2_dfrbp_1 _4535_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net413),
    .D(_0224_),
    .Q_N(_2071_),
    .Q(\tdc_inst.tdc_xor_result[35] ));
 sg13g2_dfrbp_1 _4536_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net412),
    .D(_0225_),
    .Q_N(_2070_),
    .Q(\tdc_inst.tdc_xor_result[36] ));
 sg13g2_dfrbp_1 _4537_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net411),
    .D(_0226_),
    .Q_N(_2069_),
    .Q(\tdc_inst.tdc_xor_result[37] ));
 sg13g2_dfrbp_1 _4538_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net410),
    .D(_0227_),
    .Q_N(_2068_),
    .Q(\tdc_inst.tdc_xor_result[38] ));
 sg13g2_dfrbp_1 _4539_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net409),
    .D(_0228_),
    .Q_N(_2067_),
    .Q(\tdc_inst.tdc_xor_result[39] ));
 sg13g2_dfrbp_1 _4540_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net408),
    .D(_0229_),
    .Q_N(_2066_),
    .Q(\tdc_inst.tdc_xor_result[40] ));
 sg13g2_dfrbp_1 _4541_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net407),
    .D(_0230_),
    .Q_N(_2065_),
    .Q(\tdc_inst.tdc_xor_result[41] ));
 sg13g2_dfrbp_1 _4542_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net406),
    .D(_0231_),
    .Q_N(_2064_),
    .Q(\tdc_inst.tdc_xor_result[42] ));
 sg13g2_dfrbp_1 _4543_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net405),
    .D(_0232_),
    .Q_N(_2063_),
    .Q(\tdc_inst.tdc_xor_result[43] ));
 sg13g2_dfrbp_1 _4544_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net404),
    .D(_0233_),
    .Q_N(_2062_),
    .Q(\tdc_inst.tdc_xor_result[44] ));
 sg13g2_dfrbp_1 _4545_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net403),
    .D(_0234_),
    .Q_N(_2061_),
    .Q(\tdc_inst.tdc_xor_result[45] ));
 sg13g2_dfrbp_1 _4546_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net402),
    .D(_0235_),
    .Q_N(_2060_),
    .Q(\tdc_inst.tdc_xor_result[46] ));
 sg13g2_dfrbp_1 _4547_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net401),
    .D(_0236_),
    .Q_N(_2059_),
    .Q(\tdc_inst.tdc_xor_result[47] ));
 sg13g2_dfrbp_1 _4548_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net400),
    .D(_0237_),
    .Q_N(_2058_),
    .Q(\tdc_inst.tdc_xor_result[48] ));
 sg13g2_dfrbp_1 _4549_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net399),
    .D(_0238_),
    .Q_N(_2057_),
    .Q(\tdc_inst.tdc_xor_result[49] ));
 sg13g2_dfrbp_1 _4550_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net398),
    .D(_0239_),
    .Q_N(_2056_),
    .Q(\tdc_inst.tdc_xor_result[50] ));
 sg13g2_dfrbp_1 _4551_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net397),
    .D(_0240_),
    .Q_N(_2055_),
    .Q(\tdc_inst.tdc_xor_result[51] ));
 sg13g2_dfrbp_1 _4552_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net396),
    .D(_0241_),
    .Q_N(_2054_),
    .Q(\tdc_inst.tdc_xor_result[52] ));
 sg13g2_dfrbp_1 _4553_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net395),
    .D(_0242_),
    .Q_N(_2053_),
    .Q(\tdc_inst.tdc_xor_result[53] ));
 sg13g2_dfrbp_1 _4554_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net394),
    .D(_0243_),
    .Q_N(_2052_),
    .Q(\tdc_inst.tdc_xor_result[54] ));
 sg13g2_dfrbp_1 _4555_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net393),
    .D(_0244_),
    .Q_N(_2051_),
    .Q(\tdc_inst.tdc_xor_result[55] ));
 sg13g2_dfrbp_1 _4556_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net392),
    .D(_0245_),
    .Q_N(_2050_),
    .Q(\tdc_inst.tdc_xor_result[56] ));
 sg13g2_dfrbp_1 _4557_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net391),
    .D(_0246_),
    .Q_N(_2049_),
    .Q(\tdc_inst.tdc_xor_result[57] ));
 sg13g2_dfrbp_1 _4558_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net390),
    .D(_0247_),
    .Q_N(_2048_),
    .Q(\tdc_inst.tdc_xor_result[58] ));
 sg13g2_dfrbp_1 _4559_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net389),
    .D(_0248_),
    .Q_N(_2047_),
    .Q(\tdc_inst.tdc_xor_result[59] ));
 sg13g2_dfrbp_1 _4560_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net388),
    .D(_0249_),
    .Q_N(_2046_),
    .Q(\tdc_inst.tdc_xor_result[60] ));
 sg13g2_dfrbp_1 _4561_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net387),
    .D(_0250_),
    .Q_N(_2045_),
    .Q(\tdc_inst.tdc_xor_result[61] ));
 sg13g2_dfrbp_1 _4562_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net386),
    .D(_0251_),
    .Q_N(_2044_),
    .Q(\tdc_inst.tdc_xor_result[62] ));
 sg13g2_dfrbp_1 _4563_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net385),
    .D(_0252_),
    .Q_N(_2043_),
    .Q(\tdc_inst.tdc_xor_result[63] ));
 sg13g2_dfrbp_1 _4564_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net384),
    .D(_0253_),
    .Q_N(_2042_),
    .Q(\tdc_inst.tdc_xor_result[64] ));
 sg13g2_dfrbp_1 _4565_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net383),
    .D(_0254_),
    .Q_N(_2041_),
    .Q(\tdc_inst.tdc_xor_result[65] ));
 sg13g2_dfrbp_1 _4566_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net382),
    .D(_0255_),
    .Q_N(_2040_),
    .Q(\tdc_inst.tdc_xor_result[66] ));
 sg13g2_dfrbp_1 _4567_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net381),
    .D(_0256_),
    .Q_N(_2039_),
    .Q(\tdc_inst.tdc_xor_result[67] ));
 sg13g2_dfrbp_1 _4568_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net380),
    .D(_0257_),
    .Q_N(_2038_),
    .Q(\tdc_inst.tdc_xor_result[68] ));
 sg13g2_dfrbp_1 _4569_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net379),
    .D(_0258_),
    .Q_N(_2037_),
    .Q(\tdc_inst.tdc_xor_result[69] ));
 sg13g2_dfrbp_1 _4570_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net378),
    .D(_0259_),
    .Q_N(_2036_),
    .Q(\tdc_inst.tdc_xor_result[70] ));
 sg13g2_dfrbp_1 _4571_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net377),
    .D(_0260_),
    .Q_N(_2035_),
    .Q(\tdc_inst.tdc_xor_result[71] ));
 sg13g2_dfrbp_1 _4572_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net376),
    .D(_0261_),
    .Q_N(_2034_),
    .Q(\tdc_inst.tdc_xor_result[72] ));
 sg13g2_dfrbp_1 _4573_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net375),
    .D(_0262_),
    .Q_N(_2033_),
    .Q(\tdc_inst.tdc_xor_result[73] ));
 sg13g2_dfrbp_1 _4574_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net374),
    .D(_0263_),
    .Q_N(_2032_),
    .Q(\tdc_inst.tdc_xor_result[74] ));
 sg13g2_dfrbp_1 _4575_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net373),
    .D(_0264_),
    .Q_N(_2031_),
    .Q(\tdc_inst.tdc_xor_result[75] ));
 sg13g2_dfrbp_1 _4576_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net372),
    .D(_0265_),
    .Q_N(_2030_),
    .Q(\tdc_inst.tdc_xor_result[76] ));
 sg13g2_dfrbp_1 _4577_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net371),
    .D(_0266_),
    .Q_N(_2029_),
    .Q(\tdc_inst.tdc_xor_result[77] ));
 sg13g2_dfrbp_1 _4578_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net370),
    .D(_0267_),
    .Q_N(_2028_),
    .Q(\tdc_inst.tdc_xor_result[78] ));
 sg13g2_dfrbp_1 _4579_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net369),
    .D(_0268_),
    .Q_N(_2027_),
    .Q(\tdc_inst.tdc_xor_result[79] ));
 sg13g2_dfrbp_1 _4580_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net368),
    .D(_0269_),
    .Q_N(_2026_),
    .Q(\tdc_inst.tdc_xor_result[80] ));
 sg13g2_dfrbp_1 _4581_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net367),
    .D(_0270_),
    .Q_N(_2025_),
    .Q(\tdc_inst.tdc_xor_result[81] ));
 sg13g2_dfrbp_1 _4582_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net366),
    .D(_0271_),
    .Q_N(_2024_),
    .Q(\tdc_inst.tdc_xor_result[82] ));
 sg13g2_dfrbp_1 _4583_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net365),
    .D(_0272_),
    .Q_N(_2023_),
    .Q(\tdc_inst.tdc_xor_result[83] ));
 sg13g2_dfrbp_1 _4584_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net364),
    .D(_0273_),
    .Q_N(_2022_),
    .Q(\tdc_inst.tdc_xor_result[84] ));
 sg13g2_dfrbp_1 _4585_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net363),
    .D(_0274_),
    .Q_N(_2021_),
    .Q(\tdc_inst.tdc_xor_result[85] ));
 sg13g2_dfrbp_1 _4586_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net362),
    .D(_0275_),
    .Q_N(_2020_),
    .Q(\tdc_inst.tdc_xor_result[86] ));
 sg13g2_dfrbp_1 _4587_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net361),
    .D(_0276_),
    .Q_N(_2019_),
    .Q(\tdc_inst.tdc_xor_result[87] ));
 sg13g2_dfrbp_1 _4588_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net360),
    .D(_0277_),
    .Q_N(_2018_),
    .Q(\tdc_inst.tdc_xor_result[88] ));
 sg13g2_dfrbp_1 _4589_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net359),
    .D(_0278_),
    .Q_N(_2017_),
    .Q(\tdc_inst.tdc_xor_result[89] ));
 sg13g2_dfrbp_1 _4590_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net358),
    .D(_0279_),
    .Q_N(_2016_),
    .Q(\tdc_inst.tdc_xor_result[90] ));
 sg13g2_dfrbp_1 _4591_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net357),
    .D(_0280_),
    .Q_N(_2015_),
    .Q(\tdc_inst.tdc_xor_result[91] ));
 sg13g2_dfrbp_1 _4592_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net356),
    .D(_0281_),
    .Q_N(_2014_),
    .Q(\tdc_inst.tdc_xor_result[92] ));
 sg13g2_dfrbp_1 _4593_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net355),
    .D(_0282_),
    .Q_N(_2013_),
    .Q(\tdc_inst.tdc_xor_result[93] ));
 sg13g2_dfrbp_1 _4594_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net354),
    .D(_0283_),
    .Q_N(_2012_),
    .Q(\tdc_inst.tdc_xor_result[94] ));
 sg13g2_dfrbp_1 _4595_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net353),
    .D(_0284_),
    .Q_N(_2011_),
    .Q(\tdc_inst.tdc_xor_result[95] ));
 sg13g2_dfrbp_1 _4596_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net352),
    .D(_0285_),
    .Q_N(_2010_),
    .Q(\tdc_inst.tdc_xor_result[96] ));
 sg13g2_dfrbp_1 _4597_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net351),
    .D(_0286_),
    .Q_N(_2009_),
    .Q(\tdc_inst.tdc_xor_result[97] ));
 sg13g2_dfrbp_1 _4598_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net350),
    .D(_0287_),
    .Q_N(_2008_),
    .Q(\tdc_inst.tdc_xor_result[98] ));
 sg13g2_dfrbp_1 _4599_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net349),
    .D(_0288_),
    .Q_N(_2007_),
    .Q(\tdc_inst.tdc_xor_result[99] ));
 sg13g2_dfrbp_1 _4600_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net348),
    .D(_0289_),
    .Q_N(_2006_),
    .Q(\tdc_inst.tdc_xor_result[100] ));
 sg13g2_dfrbp_1 _4601_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net347),
    .D(_0290_),
    .Q_N(_2005_),
    .Q(\tdc_inst.tdc_xor_result[101] ));
 sg13g2_dfrbp_1 _4602_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net346),
    .D(_0291_),
    .Q_N(_2004_),
    .Q(\tdc_inst.tdc_xor_result[102] ));
 sg13g2_dfrbp_1 _4603_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net345),
    .D(_0292_),
    .Q_N(_2003_),
    .Q(\tdc_inst.tdc_xor_result[103] ));
 sg13g2_dfrbp_1 _4604_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net344),
    .D(_0293_),
    .Q_N(_2002_),
    .Q(\tdc_inst.tdc_xor_result[104] ));
 sg13g2_dfrbp_1 _4605_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net343),
    .D(_0294_),
    .Q_N(_2001_),
    .Q(\tdc_inst.tdc_xor_result[105] ));
 sg13g2_dfrbp_1 _4606_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net342),
    .D(_0295_),
    .Q_N(_2000_),
    .Q(\tdc_inst.tdc_xor_result[106] ));
 sg13g2_dfrbp_1 _4607_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net341),
    .D(_0296_),
    .Q_N(_1999_),
    .Q(\tdc_inst.tdc_xor_result[107] ));
 sg13g2_dfrbp_1 _4608_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net340),
    .D(_0297_),
    .Q_N(_1998_),
    .Q(\tdc_inst.tdc_xor_result[108] ));
 sg13g2_dfrbp_1 _4609_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net339),
    .D(_0298_),
    .Q_N(_1997_),
    .Q(\tdc_inst.tdc_xor_result[109] ));
 sg13g2_dfrbp_1 _4610_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net338),
    .D(_0299_),
    .Q_N(_1996_),
    .Q(\tdc_inst.tdc_xor_result[110] ));
 sg13g2_dfrbp_1 _4611_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net337),
    .D(_0300_),
    .Q_N(_1995_),
    .Q(\tdc_inst.tdc_xor_result[111] ));
 sg13g2_dfrbp_1 _4612_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net336),
    .D(_0301_),
    .Q_N(_1994_),
    .Q(\tdc_inst.tdc_xor_result[112] ));
 sg13g2_dfrbp_1 _4613_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net335),
    .D(_0302_),
    .Q_N(_1993_),
    .Q(\tdc_inst.tdc_xor_result[113] ));
 sg13g2_dfrbp_1 _4614_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net334),
    .D(_0303_),
    .Q_N(_1992_),
    .Q(\tdc_inst.tdc_xor_result[114] ));
 sg13g2_dfrbp_1 _4615_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net333),
    .D(_0304_),
    .Q_N(_1991_),
    .Q(\tdc_inst.tdc_xor_result[115] ));
 sg13g2_dfrbp_1 _4616_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net332),
    .D(_0305_),
    .Q_N(_1990_),
    .Q(\tdc_inst.tdc_xor_result[116] ));
 sg13g2_dfrbp_1 _4617_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net331),
    .D(_0306_),
    .Q_N(_1989_),
    .Q(\tdc_inst.tdc_xor_result[117] ));
 sg13g2_dfrbp_1 _4618_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net330),
    .D(_0307_),
    .Q_N(_1988_),
    .Q(\tdc_inst.tdc_xor_result[118] ));
 sg13g2_dfrbp_1 _4619_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net329),
    .D(_0308_),
    .Q_N(_1987_),
    .Q(\tdc_inst.tdc_xor_result[119] ));
 sg13g2_dfrbp_1 _4620_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net328),
    .D(_0309_),
    .Q_N(_1986_),
    .Q(\tdc_inst.tdc_xor_result[120] ));
 sg13g2_dfrbp_1 _4621_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net327),
    .D(_0310_),
    .Q_N(_1985_),
    .Q(\tdc_inst.tdc_xor_result[121] ));
 sg13g2_dfrbp_1 _4622_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net326),
    .D(_0311_),
    .Q_N(_1984_),
    .Q(\tdc_inst.tdc_xor_result[122] ));
 sg13g2_dfrbp_1 _4623_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net325),
    .D(_0312_),
    .Q_N(_1983_),
    .Q(\tdc_inst.tdc_xor_result[123] ));
 sg13g2_dfrbp_1 _4624_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net324),
    .D(_0313_),
    .Q_N(_1982_),
    .Q(\tdc_inst.tdc_xor_result[124] ));
 sg13g2_dfrbp_1 _4625_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net323),
    .D(_0314_),
    .Q_N(_1981_),
    .Q(\tdc_inst.tdc_xor_result[125] ));
 sg13g2_dfrbp_1 _4626_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net322),
    .D(_0315_),
    .Q_N(_1980_),
    .Q(\tdc_inst.tdc_xor_result[126] ));
 sg13g2_dfrbp_1 _4627_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net321),
    .D(_0316_),
    .Q_N(_1979_),
    .Q(\tdc_inst.tdc_xor_result[127] ));
 sg13g2_dfrbp_1 _4628_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net320),
    .D(_0317_),
    .Q_N(_1978_),
    .Q(\tdc_inst.tdc_xor_result[128] ));
 sg13g2_dfrbp_1 _4629_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net319),
    .D(_0318_),
    .Q_N(_1977_),
    .Q(\tdc_inst.tdc_xor_result[129] ));
 sg13g2_dfrbp_1 _4630_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net318),
    .D(_0319_),
    .Q_N(_1976_),
    .Q(\tdc_inst.tdc_xor_result[130] ));
 sg13g2_dfrbp_1 _4631_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net317),
    .D(_0320_),
    .Q_N(_1975_),
    .Q(\tdc_inst.tdc_xor_result[131] ));
 sg13g2_dfrbp_1 _4632_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net315),
    .D(_0321_),
    .Q_N(_1974_),
    .Q(\tdc_inst.tdc_xor_result[132] ));
 sg13g2_dfrbp_1 _4633_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net314),
    .D(_0322_),
    .Q_N(_1973_),
    .Q(\tdc_inst.tdc_xor_result[133] ));
 sg13g2_dfrbp_1 _4634_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net313),
    .D(_0323_),
    .Q_N(_1972_),
    .Q(\tdc_inst.tdc_xor_result[134] ));
 sg13g2_dfrbp_1 _4635_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net312),
    .D(_0324_),
    .Q_N(_1971_),
    .Q(\tdc_inst.tdc_xor_result[135] ));
 sg13g2_dfrbp_1 _4636_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net311),
    .D(_0325_),
    .Q_N(_1970_),
    .Q(\tdc_inst.tdc_xor_result[136] ));
 sg13g2_dfrbp_1 _4637_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net310),
    .D(_0326_),
    .Q_N(_1969_),
    .Q(\tdc_inst.tdc_xor_result[137] ));
 sg13g2_dfrbp_1 _4638_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net309),
    .D(_0327_),
    .Q_N(_1968_),
    .Q(\tdc_inst.tdc_xor_result[138] ));
 sg13g2_dfrbp_1 _4639_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net308),
    .D(_0328_),
    .Q_N(_1967_),
    .Q(\tdc_inst.tdc_xor_result[139] ));
 sg13g2_dfrbp_1 _4640_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net307),
    .D(_0329_),
    .Q_N(_1966_),
    .Q(\tdc_inst.tdc_xor_result[140] ));
 sg13g2_dfrbp_1 _4641_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net306),
    .D(_0330_),
    .Q_N(_1965_),
    .Q(\tdc_inst.tdc_xor_result[141] ));
 sg13g2_dfrbp_1 _4642_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1245),
    .D(_0331_),
    .Q_N(_1964_),
    .Q(\synchronizer_spi_cs_n_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _4643_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1246),
    .D(_0332_),
    .Q_N(_1963_),
    .Q(spi_clk_sync));
 sg13g2_dfrbp_1 _4644_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1245),
    .D(_0333_),
    .Q_N(_1962_),
    .Q(\synchronizer_spi_clk_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _4645_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1249),
    .D(_0334_),
    .Q_N(_1961_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_dfrbp_1 _4646_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1245),
    .D(_0335_),
    .Q_N(_1960_),
    .Q(\synchronizer_spi_mosi_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _4647_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1248),
    .D(_0336_),
    .Q_N(_1959_),
    .Q(cpol_sync));
 sg13g2_dfrbp_1 _4648_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1248),
    .D(_0337_),
    .Q_N(_1958_),
    .Q(\synchronizer_spi_mode_cpol.data_sync[1] ));
 sg13g2_dfrbp_1 _4649_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1248),
    .D(_0338_),
    .Q_N(_1957_),
    .Q(cpha_sync));
 sg13g2_dfrbp_1 _4650_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1248),
    .D(_0339_),
    .Q_N(_1956_),
    .Q(\synchronizer_spi_mode_cpha.data_sync[1] ));
 sg13g2_dfrbp_1 _4651_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1246),
    .D(_0340_),
    .Q_N(_0007_),
    .Q(spi_cs_n_sync));
 sg13g2_dfrbp_1 _4652_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net305),
    .D(_0341_),
    .Q_N(_1955_),
    .Q(\tdc_inst.stop_count_debug[0] ));
 sg13g2_dfrbp_1 _4653_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net304),
    .D(_0342_),
    .Q_N(_1954_),
    .Q(\tdc_inst.stop_count_debug[1] ));
 sg13g2_dfrbp_1 _4654_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net303),
    .D(_0343_),
    .Q_N(_1953_),
    .Q(\tdc_inst.stop_count_debug[2] ));
 sg13g2_dfrbp_1 _4655_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net302),
    .D(_0344_),
    .Q_N(_1952_),
    .Q(\tdc_inst.stop_count_debug[3] ));
 sg13g2_dfrbp_1 _4656_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net301),
    .D(_0345_),
    .Q_N(_1951_),
    .Q(\tdc_inst.stop_count_debug[4] ));
 sg13g2_dfrbp_1 _4657_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net300),
    .D(_0346_),
    .Q_N(_1950_),
    .Q(\tdc_inst.stop_count_debug[5] ));
 sg13g2_dfrbp_1 _4658_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net299),
    .D(_0347_),
    .Q_N(_1949_),
    .Q(\tdc_inst.stop_count_debug[6] ));
 sg13g2_dfrbp_1 _4659_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net298),
    .D(_0348_),
    .Q_N(_1948_),
    .Q(\tdc_inst.stop_count_debug[7] ));
 sg13g2_dfrbp_1 _4660_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net297),
    .D(_0349_),
    .Q_N(_1947_),
    .Q(\tdc_inst.stop_count_debug[8] ));
 sg13g2_dfrbp_1 _4661_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net296),
    .D(_0350_),
    .Q_N(_1946_),
    .Q(\tdc_inst.stop_count_debug[9] ));
 sg13g2_dfrbp_1 _4662_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net295),
    .D(_0351_),
    .Q_N(_1945_),
    .Q(\tdc_inst.stop_count_debug[10] ));
 sg13g2_dfrbp_1 _4663_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net294),
    .D(_0352_),
    .Q_N(_1944_),
    .Q(\tdc_inst.stop_count_debug[11] ));
 sg13g2_dfrbp_1 _4664_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net293),
    .D(_0353_),
    .Q_N(_1943_),
    .Q(\tdc_inst.stop_count_debug[12] ));
 sg13g2_dfrbp_1 _4665_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net292),
    .D(_0354_),
    .Q_N(_1942_),
    .Q(\tdc_inst.stop_count_debug[13] ));
 sg13g2_dfrbp_1 _4666_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net291),
    .D(_0355_),
    .Q_N(_1941_),
    .Q(\tdc_inst.stop_count_debug[14] ));
 sg13g2_dfrbp_1 _4667_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net290),
    .D(_0356_),
    .Q_N(_1940_),
    .Q(\tdc_inst.stop_count_debug[15] ));
 sg13g2_dfrbp_1 _4668_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net289),
    .D(_0357_),
    .Q_N(_1939_),
    .Q(\tdc_inst.stop_count_debug[16] ));
 sg13g2_dfrbp_1 _4669_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net288),
    .D(_0358_),
    .Q_N(_1938_),
    .Q(\tdc_inst.stop_count_debug[17] ));
 sg13g2_dfrbp_1 _4670_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net287),
    .D(_0359_),
    .Q_N(_1937_),
    .Q(\tdc_inst.stop_count_debug[18] ));
 sg13g2_dfrbp_1 _4671_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net286),
    .D(_0360_),
    .Q_N(_1936_),
    .Q(\tdc_inst.stop_count_debug[19] ));
 sg13g2_dfrbp_1 _4672_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net285),
    .D(_0361_),
    .Q_N(_1935_),
    .Q(\tdc_inst.stop_count_debug[20] ));
 sg13g2_dfrbp_1 _4673_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net284),
    .D(_0362_),
    .Q_N(_1934_),
    .Q(\tdc_inst.stop_count_debug[21] ));
 sg13g2_dfrbp_1 _4674_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net283),
    .D(_0363_),
    .Q_N(_1933_),
    .Q(\tdc_inst.stop_count_debug[22] ));
 sg13g2_dfrbp_1 _4675_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net282),
    .D(_0364_),
    .Q_N(_1932_),
    .Q(\tdc_inst.stop_count_debug[23] ));
 sg13g2_dfrbp_1 _4676_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net281),
    .D(_0365_),
    .Q_N(_1931_),
    .Q(\tdc_inst.stop_count_debug[24] ));
 sg13g2_dfrbp_1 _4677_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net280),
    .D(_0366_),
    .Q_N(_1930_),
    .Q(\tdc_inst.stop_count_debug[25] ));
 sg13g2_dfrbp_1 _4678_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net279),
    .D(_0367_),
    .Q_N(_1929_),
    .Q(\tdc_inst.stop_count_debug[26] ));
 sg13g2_dfrbp_1 _4679_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net278),
    .D(_0368_),
    .Q_N(_1928_),
    .Q(\tdc_inst.stop_count_debug[27] ));
 sg13g2_dfrbp_1 _4680_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net277),
    .D(_0369_),
    .Q_N(_1927_),
    .Q(\tdc_inst.stop_count_debug[28] ));
 sg13g2_dfrbp_1 _4681_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net276),
    .D(_0370_),
    .Q_N(_1926_),
    .Q(\tdc_inst.stop_count_debug[29] ));
 sg13g2_dfrbp_1 _4682_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net275),
    .D(_0371_),
    .Q_N(_1925_),
    .Q(\tdc_inst.stop_count_debug[30] ));
 sg13g2_dfrbp_1 _4683_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net274),
    .D(_0372_),
    .Q_N(_1924_),
    .Q(\tdc_inst.stop_count_debug[31] ));
 sg13g2_dfrbp_1 _4684_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net273),
    .D(_0373_),
    .Q_N(_1923_),
    .Q(\tdc_inst.stop_count_debug[32] ));
 sg13g2_dfrbp_1 _4685_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net272),
    .D(_0374_),
    .Q_N(_1922_),
    .Q(\tdc_inst.stop_count_debug[33] ));
 sg13g2_dfrbp_1 _4686_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net271),
    .D(_0375_),
    .Q_N(_1921_),
    .Q(\tdc_inst.stop_count_debug[34] ));
 sg13g2_dfrbp_1 _4687_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net270),
    .D(_0376_),
    .Q_N(_1920_),
    .Q(\tdc_inst.stop_count_debug[35] ));
 sg13g2_dfrbp_1 _4688_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net269),
    .D(_0377_),
    .Q_N(_1919_),
    .Q(\tdc_inst.stop_count_debug[36] ));
 sg13g2_dfrbp_1 _4689_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net268),
    .D(_0378_),
    .Q_N(_1918_),
    .Q(\tdc_inst.stop_count_debug[37] ));
 sg13g2_dfrbp_1 _4690_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net267),
    .D(_0379_),
    .Q_N(_1917_),
    .Q(\tdc_inst.stop_count_debug[38] ));
 sg13g2_dfrbp_1 _4691_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net266),
    .D(_0380_),
    .Q_N(_1916_),
    .Q(\tdc_inst.stop_count_debug[39] ));
 sg13g2_dfrbp_1 _4692_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net265),
    .D(_0381_),
    .Q_N(_1915_),
    .Q(\tdc_inst.stop_count_debug[40] ));
 sg13g2_dfrbp_1 _4693_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net264),
    .D(_0382_),
    .Q_N(_1914_),
    .Q(\tdc_inst.stop_count_debug[41] ));
 sg13g2_dfrbp_1 _4694_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net263),
    .D(_0383_),
    .Q_N(_1913_),
    .Q(\tdc_inst.stop_count_debug[42] ));
 sg13g2_dfrbp_1 _4695_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net262),
    .D(_0384_),
    .Q_N(_1912_),
    .Q(\tdc_inst.stop_count_debug[43] ));
 sg13g2_dfrbp_1 _4696_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net261),
    .D(_0385_),
    .Q_N(_1911_),
    .Q(\tdc_inst.stop_count_debug[44] ));
 sg13g2_dfrbp_1 _4697_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net260),
    .D(_0386_),
    .Q_N(_1910_),
    .Q(\tdc_inst.stop_count_debug[45] ));
 sg13g2_dfrbp_1 _4698_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net259),
    .D(_0387_),
    .Q_N(_1909_),
    .Q(\tdc_inst.stop_count_debug[46] ));
 sg13g2_dfrbp_1 _4699_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net258),
    .D(_0388_),
    .Q_N(_1908_),
    .Q(\tdc_inst.stop_count_debug[47] ));
 sg13g2_dfrbp_1 _4700_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net257),
    .D(_0389_),
    .Q_N(_1907_),
    .Q(\tdc_inst.stop_count_debug[48] ));
 sg13g2_dfrbp_1 _4701_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net256),
    .D(_0390_),
    .Q_N(_1906_),
    .Q(\tdc_inst.stop_count_debug[49] ));
 sg13g2_dfrbp_1 _4702_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net255),
    .D(_0391_),
    .Q_N(_1905_),
    .Q(\tdc_inst.stop_count_debug[50] ));
 sg13g2_dfrbp_1 _4703_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net254),
    .D(_0392_),
    .Q_N(_1904_),
    .Q(\tdc_inst.stop_count_debug[51] ));
 sg13g2_dfrbp_1 _4704_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net253),
    .D(_0393_),
    .Q_N(_1903_),
    .Q(\tdc_inst.stop_count_debug[52] ));
 sg13g2_dfrbp_1 _4705_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net252),
    .D(_0394_),
    .Q_N(_1902_),
    .Q(\tdc_inst.stop_count_debug[53] ));
 sg13g2_dfrbp_1 _4706_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net251),
    .D(_0395_),
    .Q_N(_1901_),
    .Q(\tdc_inst.stop_count_debug[54] ));
 sg13g2_dfrbp_1 _4707_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net250),
    .D(_0396_),
    .Q_N(_1900_),
    .Q(\tdc_inst.stop_count_debug[55] ));
 sg13g2_dfrbp_1 _4708_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net249),
    .D(_0397_),
    .Q_N(_1899_),
    .Q(\tdc_inst.stop_count_debug[56] ));
 sg13g2_dfrbp_1 _4709_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net248),
    .D(_0398_),
    .Q_N(_1898_),
    .Q(\tdc_inst.stop_count_debug[57] ));
 sg13g2_dfrbp_1 _4710_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net247),
    .D(_0399_),
    .Q_N(_1897_),
    .Q(\tdc_inst.stop_count_debug[58] ));
 sg13g2_dfrbp_1 _4711_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net246),
    .D(_0400_),
    .Q_N(_1896_),
    .Q(\tdc_inst.stop_count_debug[59] ));
 sg13g2_dfrbp_1 _4712_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net245),
    .D(_0401_),
    .Q_N(_1895_),
    .Q(\tdc_inst.stop_count_debug[60] ));
 sg13g2_dfrbp_1 _4713_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net244),
    .D(_0402_),
    .Q_N(_1894_),
    .Q(\tdc_inst.stop_count_debug[61] ));
 sg13g2_dfrbp_1 _4714_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net243),
    .D(_0403_),
    .Q_N(_1893_),
    .Q(\tdc_inst.stop_count_debug[62] ));
 sg13g2_dfrbp_1 _4715_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net242),
    .D(_0404_),
    .Q_N(_1892_),
    .Q(\tdc_inst.stop_count_debug[63] ));
 sg13g2_dfrbp_1 _4716_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net241),
    .D(_0405_),
    .Q_N(_1891_),
    .Q(\tdc_inst.stop_count_debug[64] ));
 sg13g2_dfrbp_1 _4717_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net240),
    .D(_0406_),
    .Q_N(_1890_),
    .Q(\tdc_inst.stop_count_debug[65] ));
 sg13g2_dfrbp_1 _4718_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net239),
    .D(_0407_),
    .Q_N(_1889_),
    .Q(\tdc_inst.stop_count_debug[66] ));
 sg13g2_dfrbp_1 _4719_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net238),
    .D(_0408_),
    .Q_N(_1888_),
    .Q(\tdc_inst.stop_count_debug[67] ));
 sg13g2_dfrbp_1 _4720_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net237),
    .D(_0409_),
    .Q_N(_1887_),
    .Q(\tdc_inst.stop_count_debug[68] ));
 sg13g2_dfrbp_1 _4721_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net236),
    .D(_0410_),
    .Q_N(_1886_),
    .Q(\tdc_inst.stop_count_debug[69] ));
 sg13g2_dfrbp_1 _4722_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net235),
    .D(_0411_),
    .Q_N(_1885_),
    .Q(\tdc_inst.stop_count_debug[70] ));
 sg13g2_dfrbp_1 _4723_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net234),
    .D(_0412_),
    .Q_N(_1884_),
    .Q(\tdc_inst.stop_count_debug[71] ));
 sg13g2_dfrbp_1 _4724_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net233),
    .D(_0413_),
    .Q_N(_1883_),
    .Q(\tdc_inst.stop_count_debug[72] ));
 sg13g2_dfrbp_1 _4725_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net232),
    .D(_0414_),
    .Q_N(_1882_),
    .Q(\tdc_inst.stop_count_debug[73] ));
 sg13g2_dfrbp_1 _4726_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net231),
    .D(_0415_),
    .Q_N(_1881_),
    .Q(\tdc_inst.stop_count_debug[74] ));
 sg13g2_dfrbp_1 _4727_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net230),
    .D(_0416_),
    .Q_N(_1880_),
    .Q(\tdc_inst.stop_count_debug[75] ));
 sg13g2_dfrbp_1 _4728_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net229),
    .D(_0417_),
    .Q_N(_1879_),
    .Q(\tdc_inst.stop_count_debug[76] ));
 sg13g2_dfrbp_1 _4729_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net228),
    .D(_0418_),
    .Q_N(_1878_),
    .Q(\tdc_inst.stop_count_debug[77] ));
 sg13g2_dfrbp_1 _4730_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net227),
    .D(_0419_),
    .Q_N(_1877_),
    .Q(\tdc_inst.stop_count_debug[78] ));
 sg13g2_dfrbp_1 _4731_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net226),
    .D(_0420_),
    .Q_N(_1876_),
    .Q(\tdc_inst.stop_count_debug[79] ));
 sg13g2_dfrbp_1 _4732_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net225),
    .D(_0421_),
    .Q_N(_1875_),
    .Q(\tdc_inst.stop_count_debug[80] ));
 sg13g2_dfrbp_1 _4733_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net224),
    .D(_0422_),
    .Q_N(_1874_),
    .Q(\tdc_inst.stop_count_debug[81] ));
 sg13g2_dfrbp_1 _4734_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net223),
    .D(_0423_),
    .Q_N(_1873_),
    .Q(\tdc_inst.stop_count_debug[82] ));
 sg13g2_dfrbp_1 _4735_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net222),
    .D(_0424_),
    .Q_N(_1872_),
    .Q(\tdc_inst.stop_count_debug[83] ));
 sg13g2_dfrbp_1 _4736_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net221),
    .D(_0425_),
    .Q_N(_1871_),
    .Q(\tdc_inst.stop_count_debug[84] ));
 sg13g2_dfrbp_1 _4737_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net220),
    .D(_0426_),
    .Q_N(_1870_),
    .Q(\tdc_inst.stop_count_debug[85] ));
 sg13g2_dfrbp_1 _4738_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net219),
    .D(_0427_),
    .Q_N(_1869_),
    .Q(\tdc_inst.stop_count_debug[86] ));
 sg13g2_dfrbp_1 _4739_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net218),
    .D(_0428_),
    .Q_N(_1868_),
    .Q(\tdc_inst.stop_count_debug[87] ));
 sg13g2_dfrbp_1 _4740_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net217),
    .D(_0429_),
    .Q_N(_1867_),
    .Q(\tdc_inst.stop_count_debug[88] ));
 sg13g2_dfrbp_1 _4741_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net216),
    .D(_0430_),
    .Q_N(_1866_),
    .Q(\tdc_inst.stop_count_debug[89] ));
 sg13g2_dfrbp_1 _4742_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net215),
    .D(_0431_),
    .Q_N(_1865_),
    .Q(\tdc_inst.stop_count_debug[90] ));
 sg13g2_dfrbp_1 _4743_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net214),
    .D(_0432_),
    .Q_N(_1864_),
    .Q(\tdc_inst.stop_count_debug[91] ));
 sg13g2_dfrbp_1 _4744_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net213),
    .D(_0433_),
    .Q_N(_1863_),
    .Q(\tdc_inst.stop_count_debug[92] ));
 sg13g2_dfrbp_1 _4745_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net212),
    .D(_0434_),
    .Q_N(_1862_),
    .Q(\tdc_inst.stop_count_debug[93] ));
 sg13g2_dfrbp_1 _4746_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net211),
    .D(_0435_),
    .Q_N(_1861_),
    .Q(\tdc_inst.stop_count_debug[94] ));
 sg13g2_dfrbp_1 _4747_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net210),
    .D(_0436_),
    .Q_N(_1860_),
    .Q(\tdc_inst.stop_count_debug[95] ));
 sg13g2_dfrbp_1 _4748_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net209),
    .D(_0437_),
    .Q_N(_1859_),
    .Q(\tdc_inst.stop_count_debug[96] ));
 sg13g2_dfrbp_1 _4749_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net208),
    .D(_0438_),
    .Q_N(_1858_),
    .Q(\tdc_inst.stop_count_debug[97] ));
 sg13g2_dfrbp_1 _4750_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net207),
    .D(_0439_),
    .Q_N(_1857_),
    .Q(\tdc_inst.stop_count_debug[98] ));
 sg13g2_dfrbp_1 _4751_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net206),
    .D(_0440_),
    .Q_N(_1856_),
    .Q(\tdc_inst.stop_count_debug[99] ));
 sg13g2_dfrbp_1 _4752_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net205),
    .D(_0441_),
    .Q_N(_1855_),
    .Q(\tdc_inst.stop_count_debug[100] ));
 sg13g2_dfrbp_1 _4753_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net204),
    .D(_0442_),
    .Q_N(_1854_),
    .Q(\tdc_inst.stop_count_debug[101] ));
 sg13g2_dfrbp_1 _4754_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net203),
    .D(_0443_),
    .Q_N(_1853_),
    .Q(\tdc_inst.stop_count_debug[102] ));
 sg13g2_dfrbp_1 _4755_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net202),
    .D(_0444_),
    .Q_N(_1852_),
    .Q(\tdc_inst.stop_count_debug[103] ));
 sg13g2_dfrbp_1 _4756_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net201),
    .D(_0445_),
    .Q_N(_1851_),
    .Q(\tdc_inst.stop_count_debug[104] ));
 sg13g2_dfrbp_1 _4757_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net200),
    .D(_0446_),
    .Q_N(_1850_),
    .Q(\tdc_inst.stop_count_debug[105] ));
 sg13g2_dfrbp_1 _4758_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net199),
    .D(_0447_),
    .Q_N(_1849_),
    .Q(\tdc_inst.stop_count_debug[106] ));
 sg13g2_dfrbp_1 _4759_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net198),
    .D(_0448_),
    .Q_N(_1848_),
    .Q(\tdc_inst.stop_count_debug[107] ));
 sg13g2_dfrbp_1 _4760_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net197),
    .D(_0449_),
    .Q_N(_1847_),
    .Q(\tdc_inst.stop_count_debug[108] ));
 sg13g2_dfrbp_1 _4761_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net196),
    .D(_0450_),
    .Q_N(_1846_),
    .Q(\tdc_inst.stop_count_debug[109] ));
 sg13g2_dfrbp_1 _4762_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net195),
    .D(_0451_),
    .Q_N(_1845_),
    .Q(\tdc_inst.stop_count_debug[110] ));
 sg13g2_dfrbp_1 _4763_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net194),
    .D(_0452_),
    .Q_N(_1844_),
    .Q(\tdc_inst.stop_count_debug[111] ));
 sg13g2_dfrbp_1 _4764_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net193),
    .D(_0453_),
    .Q_N(_1843_),
    .Q(\tdc_inst.stop_count_debug[112] ));
 sg13g2_dfrbp_1 _4765_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net192),
    .D(_0454_),
    .Q_N(_1842_),
    .Q(\tdc_inst.stop_count_debug[113] ));
 sg13g2_dfrbp_1 _4766_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net191),
    .D(_0455_),
    .Q_N(_1841_),
    .Q(\tdc_inst.stop_count_debug[114] ));
 sg13g2_dfrbp_1 _4767_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net190),
    .D(_0456_),
    .Q_N(_1840_),
    .Q(\tdc_inst.stop_count_debug[115] ));
 sg13g2_dfrbp_1 _4768_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net189),
    .D(_0457_),
    .Q_N(_1839_),
    .Q(\tdc_inst.stop_count_debug[116] ));
 sg13g2_dfrbp_1 _4769_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net188),
    .D(_0458_),
    .Q_N(_1838_),
    .Q(\tdc_inst.stop_count_debug[117] ));
 sg13g2_dfrbp_1 _4770_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net187),
    .D(_0459_),
    .Q_N(_1837_),
    .Q(\tdc_inst.stop_count_debug[118] ));
 sg13g2_dfrbp_1 _4771_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net186),
    .D(_0460_),
    .Q_N(_1836_),
    .Q(\tdc_inst.stop_count_debug[119] ));
 sg13g2_dfrbp_1 _4772_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net185),
    .D(_0461_),
    .Q_N(_1835_),
    .Q(\tdc_inst.stop_count_debug[120] ));
 sg13g2_dfrbp_1 _4773_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net184),
    .D(_0462_),
    .Q_N(_1834_),
    .Q(\tdc_inst.stop_count_debug[121] ));
 sg13g2_dfrbp_1 _4774_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net183),
    .D(_0463_),
    .Q_N(_1833_),
    .Q(\tdc_inst.stop_count_debug[122] ));
 sg13g2_dfrbp_1 _4775_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net182),
    .D(_0464_),
    .Q_N(_1832_),
    .Q(\tdc_inst.stop_count_debug[123] ));
 sg13g2_dfrbp_1 _4776_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net181),
    .D(_0465_),
    .Q_N(_1831_),
    .Q(\tdc_inst.stop_count_debug[124] ));
 sg13g2_dfrbp_1 _4777_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net180),
    .D(_0466_),
    .Q_N(_1830_),
    .Q(\tdc_inst.stop_count_debug[125] ));
 sg13g2_dfrbp_1 _4778_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net179),
    .D(_0467_),
    .Q_N(_1829_),
    .Q(\tdc_inst.stop_count_debug[126] ));
 sg13g2_dfrbp_1 _4779_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net178),
    .D(_0468_),
    .Q_N(_1828_),
    .Q(\tdc_inst.stop_count_debug[127] ));
 sg13g2_dfrbp_1 _4780_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net177),
    .D(_0469_),
    .Q_N(_1827_),
    .Q(\tdc_inst.stop_count_debug[128] ));
 sg13g2_dfrbp_1 _4781_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net176),
    .D(_0470_),
    .Q_N(_1826_),
    .Q(\tdc_inst.stop_count_debug[129] ));
 sg13g2_dfrbp_1 _4782_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net175),
    .D(_0471_),
    .Q_N(_1825_),
    .Q(\tdc_inst.stop_count_debug[130] ));
 sg13g2_dfrbp_1 _4783_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net174),
    .D(_0472_),
    .Q_N(_1824_),
    .Q(\tdc_inst.stop_count_debug[131] ));
 sg13g2_dfrbp_1 _4784_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net173),
    .D(_0473_),
    .Q_N(_1823_),
    .Q(\tdc_inst.stop_count_debug[132] ));
 sg13g2_dfrbp_1 _4785_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net172),
    .D(_0474_),
    .Q_N(_1822_),
    .Q(\tdc_inst.stop_count_debug[133] ));
 sg13g2_dfrbp_1 _4786_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net171),
    .D(_0475_),
    .Q_N(_1821_),
    .Q(\tdc_inst.stop_count_debug[134] ));
 sg13g2_dfrbp_1 _4787_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net170),
    .D(_0476_),
    .Q_N(_1820_),
    .Q(\tdc_inst.stop_count_debug[135] ));
 sg13g2_dfrbp_1 _4788_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net169),
    .D(_0477_),
    .Q_N(_1819_),
    .Q(\tdc_inst.stop_count_debug[136] ));
 sg13g2_dfrbp_1 _4789_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net168),
    .D(_0478_),
    .Q_N(_1818_),
    .Q(\tdc_inst.stop_count_debug[137] ));
 sg13g2_dfrbp_1 _4790_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net167),
    .D(_0479_),
    .Q_N(_1817_),
    .Q(\tdc_inst.stop_count_debug[138] ));
 sg13g2_dfrbp_1 _4791_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net166),
    .D(_0480_),
    .Q_N(_1816_),
    .Q(\tdc_inst.stop_count_debug[139] ));
 sg13g2_dfrbp_1 _4792_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net165),
    .D(_0481_),
    .Q_N(_1815_),
    .Q(\tdc_inst.stop_count_debug[140] ));
 sg13g2_dfrbp_1 _4793_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net164),
    .D(_0482_),
    .Q_N(_1814_),
    .Q(\tdc_inst.stop_count_debug[141] ));
 sg13g2_dfrbp_1 _4794_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1248),
    .D(_0046_),
    .Q_N(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .Q(_0045_));
 sg13g2_dfrbp_1 _4795_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1247),
    .D(_0000_),
    .Q_N(_2249_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[1] ));
 sg13g2_dfrbp_1 _4796_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1247),
    .D(_0001_),
    .Q_N(_2250_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_dfrbp_1 _4797_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1248),
    .D(net556),
    .Q_N(_2251_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_dfrbp_1 _4798_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1248),
    .D(net663),
    .Q_N(_1813_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_dfrbp_1 _4799_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1255),
    .D(_0483_),
    .Q_N(_1812_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ));
 sg13g2_dfrbp_1 _4800_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1256),
    .D(net1761),
    .Q_N(_1811_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ));
 sg13g2_dfrbp_1 _4801_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1256),
    .D(_0485_),
    .Q_N(_1810_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ));
 sg13g2_dfrbp_1 _4802_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1256),
    .D(_0486_),
    .Q_N(_1809_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_dfrbp_1 _4803_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1247),
    .D(_0487_),
    .Q_N(_1808_),
    .Q(\spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_dfrbp_1 _4804_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1243),
    .D(_0488_),
    .Q_N(_1807_),
    .Q(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_dfrbp_1 _4805_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1247),
    .D(net701),
    .Q_N(_1806_),
    .Q(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_dfrbp_1 _4806_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1243),
    .D(_0490_),
    .Q_N(_0008_),
    .Q(\spi_wrapper_i.reg_addr[2] ));
 sg13g2_dfrbp_1 _4807_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1251),
    .D(_0491_),
    .Q_N(_1805_),
    .Q(\spi_wrapper_i.reg_addr[3] ));
 sg13g2_dfrbp_1 _4808_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1247),
    .D(net922),
    .Q_N(_1804_),
    .Q(\spi_wrapper_i.reg_data_o_vld ));
 sg13g2_dfrbp_1 _4809_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1247),
    .D(_0493_),
    .Q_N(_1803_),
    .Q(\spi_wrapper_i.reg_data_o[0] ));
 sg13g2_dfrbp_1 _4810_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1247),
    .D(_0494_),
    .Q_N(_1802_),
    .Q(\spi_wrapper_i.reg_data_o[1] ));
 sg13g2_dfrbp_1 _4811_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1255),
    .D(_0495_),
    .Q_N(_1801_),
    .Q(\spi_wrapper_i.reg_data_o[2] ));
 sg13g2_dfrbp_1 _4812_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1255),
    .D(_0496_),
    .Q_N(_1800_),
    .Q(\spi_wrapper_i.reg_data_o[3] ));
 sg13g2_dfrbp_1 _4813_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1255),
    .D(_0497_),
    .Q_N(_1799_),
    .Q(\spi_wrapper_i.reg_data_o[4] ));
 sg13g2_dfrbp_1 _4814_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1256),
    .D(net1271),
    .Q_N(_1798_),
    .Q(\spi_wrapper_i.reg_data_o[5] ));
 sg13g2_dfrbp_1 _4815_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1256),
    .D(_0499_),
    .Q_N(_1797_),
    .Q(\spi_wrapper_i.reg_data_o[6] ));
 sg13g2_dfrbp_1 _4816_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1256),
    .D(_0500_),
    .Q_N(_1796_),
    .Q(\spi_wrapper_i.reg_data_o[7] ));
 sg13g2_dfrbp_1 _4817_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1245),
    .D(_0501_),
    .Q_N(_1795_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ));
 sg13g2_dfrbp_1 _4818_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1245),
    .D(net1696),
    .Q_N(_1794_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ));
 sg13g2_dfrbp_1 _4819_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1245),
    .D(net903),
    .Q_N(_1793_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ));
 sg13g2_dfrbp_1 _4820_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1246),
    .D(net1783),
    .Q_N(_1792_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ));
 sg13g2_dfrbp_1 _4821_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1237),
    .D(net715),
    .Q_N(_1791_),
    .Q(\config_regs[56] ));
 sg13g2_dfrbp_1 _4822_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1237),
    .D(_0506_),
    .Q_N(_1790_),
    .Q(\config_regs[57] ));
 sg13g2_dfrbp_1 _4823_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1250),
    .D(net678),
    .Q_N(_1789_),
    .Q(\config_regs[58] ));
 sg13g2_dfrbp_1 _4824_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1239),
    .D(net755),
    .Q_N(_1788_),
    .Q(\config_regs[59] ));
 sg13g2_dfrbp_1 _4825_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1240),
    .D(_0509_),
    .Q_N(_1787_),
    .Q(\config_regs[60] ));
 sg13g2_dfrbp_1 _4826_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1241),
    .D(net814),
    .Q_N(_1786_),
    .Q(\config_regs[61] ));
 sg13g2_dfrbp_1 _4827_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1252),
    .D(_0511_),
    .Q_N(_1785_),
    .Q(\config_regs[62] ));
 sg13g2_dfrbp_1 _4828_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1252),
    .D(_0512_),
    .Q_N(_1784_),
    .Q(\config_regs[63] ));
 sg13g2_dfrbp_1 _4829_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1244),
    .D(_0513_),
    .Q_N(_0011_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ));
 sg13g2_dfrbp_1 _4830_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1244),
    .D(net707),
    .Q_N(_0014_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ));
 sg13g2_dfrbp_1 _4831_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1244),
    .D(net676),
    .Q_N(_0017_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ));
 sg13g2_dfrbp_1 _4832_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1244),
    .D(_0516_),
    .Q_N(_0020_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ));
 sg13g2_dfrbp_1 _4833_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1244),
    .D(net1736),
    .Q_N(_0023_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ));
 sg13g2_dfrbp_1 _4834_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1246),
    .D(_0518_),
    .Q_N(_0026_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ));
 sg13g2_dfrbp_1 _4835_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1246),
    .D(_0519_),
    .Q_N(_0029_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ));
 sg13g2_dfrbp_1 _4836_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1246),
    .D(net591),
    .Q_N(_1783_),
    .Q(spi_miso));
 sg13g2_dfrbp_1 _4837_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net163),
    .D(net1687),
    .Q_N(_1782_),
    .Q(\fine_result[0] ));
 sg13g2_dfrbp_1 _4838_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net162),
    .D(net1651),
    .Q_N(_1781_),
    .Q(\fine_result[1] ));
 sg13g2_dfrbp_1 _4839_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net161),
    .D(net1331),
    .Q_N(_1780_),
    .Q(\fine_result[2] ));
 sg13g2_dfrbp_1 _4840_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net160),
    .D(net913),
    .Q_N(_1779_),
    .Q(\fine_result[3] ));
 sg13g2_dfrbp_1 _4841_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net159),
    .D(net767),
    .Q_N(_1778_),
    .Q(\fine_result[4] ));
 sg13g2_dfrbp_1 _4842_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net158),
    .D(net1723),
    .Q_N(_1777_),
    .Q(\fine_result[5] ));
 sg13g2_dfrbp_1 _4843_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net157),
    .D(net1357),
    .Q_N(_1776_),
    .Q(\fine_result[6] ));
 sg13g2_dfrbp_1 _4844_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net156),
    .D(net1674),
    .Q_N(_1775_),
    .Q(\fine_result[7] ));
 sg13g2_dfrbp_1 _4845_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net155),
    .D(net860),
    .Q_N(_1774_),
    .Q(\fine_result[8] ));
 sg13g2_dfrbp_1 _4846_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1246),
    .D(net605),
    .Q_N(_1773_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ));
 sg13g2_dfrbp_1 _4847_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1247),
    .D(_0531_),
    .Q_N(_1772_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ));
 sg13g2_dfrbp_1 _4848_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1255),
    .D(_0532_),
    .Q_N(_1771_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ));
 sg13g2_dfrbp_1 _4849_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1255),
    .D(_0533_),
    .Q_N(_1770_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ));
 sg13g2_dfrbp_1 _4850_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1255),
    .D(_0534_),
    .Q_N(_1769_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ));
 sg13g2_dfrbp_1 _4851_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1255),
    .D(_0535_),
    .Q_N(_1768_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ));
 sg13g2_dfrbp_1 _4852_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1256),
    .D(_0536_),
    .Q_N(_1767_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ));
 sg13g2_dfrbp_1 _4853_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1257),
    .D(_0537_),
    .Q_N(_1766_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ));
 sg13g2_dfrbp_1 _4854_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1245),
    .D(_0538_),
    .Q_N(_1765_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ));
 sg13g2_dfrbp_1 _4855_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1242),
    .D(net1630),
    .Q_N(_1764_),
    .Q(\config_regs[32] ));
 sg13g2_dfrbp_1 _4856_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1242),
    .D(_0540_),
    .Q_N(_1763_),
    .Q(\config_regs[33] ));
 sg13g2_dfrbp_1 _4857_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1250),
    .D(net1665),
    .Q_N(_1762_),
    .Q(\config_regs[34] ));
 sg13g2_dfrbp_1 _4858_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1251),
    .D(net1361),
    .Q_N(_1761_),
    .Q(\config_regs[35] ));
 sg13g2_dfrbp_1 _4859_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1251),
    .D(net834),
    .Q_N(_1760_),
    .Q(\config_regs[36] ));
 sg13g2_dfrbp_1 _4860_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1254),
    .D(net1504),
    .Q_N(_1759_),
    .Q(\config_regs[37] ));
 sg13g2_dfrbp_1 _4861_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1253),
    .D(net670),
    .Q_N(_1758_),
    .Q(\config_regs[38] ));
 sg13g2_dfrbp_1 _4862_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1253),
    .D(net660),
    .Q_N(_1757_),
    .Q(\config_regs[39] ));
 sg13g2_dfrbp_1 _4863_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1243),
    .D(net795),
    .Q_N(_1756_),
    .Q(\config_regs[40] ));
 sg13g2_dfrbp_1 _4864_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1242),
    .D(net711),
    .Q_N(_1755_),
    .Q(\config_regs[41] ));
 sg13g2_dfrbp_1 _4865_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1250),
    .D(net723),
    .Q_N(_1754_),
    .Q(\config_regs[42] ));
 sg13g2_dfrbp_1 _4866_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1239),
    .D(net740),
    .Q_N(_1753_),
    .Q(\config_regs[43] ));
 sg13g2_dfrbp_1 _4867_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1239),
    .D(net816),
    .Q_N(_1752_),
    .Q(\config_regs[44] ));
 sg13g2_dfrbp_1 _4868_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1241),
    .D(net826),
    .Q_N(_1751_),
    .Q(\config_regs[45] ));
 sg13g2_dfrbp_1 _4869_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1253),
    .D(_0553_),
    .Q_N(_1750_),
    .Q(\config_regs[46] ));
 sg13g2_dfrbp_1 _4870_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1253),
    .D(_0554_),
    .Q_N(_1749_),
    .Q(\config_regs[47] ));
 sg13g2_dfrbp_1 _4871_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1242),
    .D(net753),
    .Q_N(_1748_),
    .Q(\config_regs[24] ));
 sg13g2_dfrbp_1 _4872_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1237),
    .D(net725),
    .Q_N(_1747_),
    .Q(\config_regs[25] ));
 sg13g2_dfrbp_1 _4873_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1250),
    .D(net759),
    .Q_N(_1746_),
    .Q(\config_regs[26] ));
 sg13g2_dfrbp_1 _4874_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1239),
    .D(net1335),
    .Q_N(_1745_),
    .Q(\config_regs[27] ));
 sg13g2_dfrbp_1 _4875_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1240),
    .D(net727),
    .Q_N(_1744_),
    .Q(\config_regs[28] ));
 sg13g2_dfrbp_1 _4876_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1241),
    .D(net1288),
    .Q_N(_1743_),
    .Q(\config_regs[29] ));
 sg13g2_dfrbp_1 _4877_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1252),
    .D(_0561_),
    .Q_N(_1742_),
    .Q(\config_regs[30] ));
 sg13g2_dfrbp_1 _4878_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1252),
    .D(_0562_),
    .Q_N(_1741_),
    .Q(\config_regs[31] ));
 sg13g2_dfrbp_1 _4879_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1242),
    .D(net778),
    .Q_N(_1740_),
    .Q(\config_regs[48] ));
 sg13g2_dfrbp_1 _4880_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1242),
    .D(_0564_),
    .Q_N(_1739_),
    .Q(\config_regs[49] ));
 sg13g2_dfrbp_1 _4881_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1250),
    .D(net1348),
    .Q_N(_1738_),
    .Q(\config_regs[50] ));
 sg13g2_dfrbp_1 _4882_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1239),
    .D(net738),
    .Q_N(_1737_),
    .Q(\config_regs[51] ));
 sg13g2_dfrbp_1 _4883_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1239),
    .D(_0567_),
    .Q_N(_1736_),
    .Q(\config_regs[52] ));
 sg13g2_dfrbp_1 _4884_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1241),
    .D(net789),
    .Q_N(_1735_),
    .Q(\config_regs[53] ));
 sg13g2_dfrbp_1 _4885_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1252),
    .D(_0569_),
    .Q_N(_1734_),
    .Q(\config_regs[54] ));
 sg13g2_dfrbp_1 _4886_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1252),
    .D(_0570_),
    .Q_N(_1733_),
    .Q(\config_regs[55] ));
 sg13g2_dfrbp_1 _4887_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1242),
    .D(net930),
    .Q_N(_1732_),
    .Q(\config_regs[16] ));
 sg13g2_dfrbp_1 _4888_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1237),
    .D(net744),
    .Q_N(_1731_),
    .Q(\config_regs[17] ));
 sg13g2_dfrbp_1 _4889_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1250),
    .D(net721),
    .Q_N(_1730_),
    .Q(\config_regs[18] ));
 sg13g2_dfrbp_1 _4890_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1239),
    .D(net938),
    .Q_N(_1729_),
    .Q(\config_regs[19] ));
 sg13g2_dfrbp_1 _4891_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1241),
    .D(net774),
    .Q_N(_1728_),
    .Q(\config_regs[20] ));
 sg13g2_dfrbp_1 _4892_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1241),
    .D(net820),
    .Q_N(_1727_),
    .Q(\config_regs[21] ));
 sg13g2_dfrbp_1 _4893_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1252),
    .D(_0577_),
    .Q_N(_1726_),
    .Q(\config_regs[22] ));
 sg13g2_dfrbp_1 _4894_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1253),
    .D(_0578_),
    .Q_N(_1725_),
    .Q(\config_regs[23] ));
 sg13g2_dfrbp_1 _4895_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1242),
    .D(net880),
    .Q_N(_1724_),
    .Q(\config_regs[8] ));
 sg13g2_dfrbp_1 _4896_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1237),
    .D(net751),
    .Q_N(_1723_),
    .Q(\config_regs[9] ));
 sg13g2_dfrbp_1 _4897_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1250),
    .D(net797),
    .Q_N(_1722_),
    .Q(\config_regs[10] ));
 sg13g2_dfrbp_1 _4898_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1239),
    .D(net864),
    .Q_N(_1721_),
    .Q(\config_regs[11] ));
 sg13g2_dfrbp_1 _4899_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1240),
    .D(net697),
    .Q_N(_1720_),
    .Q(\config_regs[12] ));
 sg13g2_dfrbp_1 _4900_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1241),
    .D(net655),
    .Q_N(_1719_),
    .Q(\config_regs[13] ));
 sg13g2_dfrbp_1 _4901_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1252),
    .D(_0585_),
    .Q_N(_1718_),
    .Q(\config_regs[14] ));
 sg13g2_dfrbp_1 _4902_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1254),
    .D(_0586_),
    .Q_N(_1717_),
    .Q(\config_regs[15] ));
 sg13g2_dfrbp_1 _4903_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1243),
    .D(net627),
    .Q_N(_0009_),
    .Q(\config_regs[0] ));
 sg13g2_dfrbp_1 _4904_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1243),
    .D(net615),
    .Q_N(_0012_),
    .Q(\config_regs[1] ));
 sg13g2_dfrbp_1 _4905_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1251),
    .D(net607),
    .Q_N(_0015_),
    .Q(\config_regs[2] ));
 sg13g2_dfrbp_1 _4906_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1251),
    .D(net609),
    .Q_N(_0018_),
    .Q(\config_regs[3] ));
 sg13g2_dfrbp_1 _4907_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1250),
    .D(net621),
    .Q_N(_0021_),
    .Q(\config_regs[4] ));
 sg13g2_dfrbp_1 _4908_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1253),
    .D(net611),
    .Q_N(_0024_),
    .Q(\config_regs[5] ));
 sg13g2_dfrbp_1 _4909_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1253),
    .D(net588),
    .Q_N(_0027_),
    .Q(\config_regs[6] ));
 sg13g2_dfrbp_1 _4910_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1253),
    .D(net617),
    .Q_N(_0030_),
    .Q(\config_regs[7] ));
 sg13g2_dfrbp_1 _4911_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net154),
    .D(_0595_),
    .Q_N(_0010_),
    .Q(\coarse_result[0] ));
 sg13g2_dfrbp_1 _4912_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net152),
    .D(_0596_),
    .Q_N(_0013_),
    .Q(\coarse_result[1] ));
 sg13g2_dfrbp_1 _4913_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net151),
    .D(_0597_),
    .Q_N(_0016_),
    .Q(\coarse_result[2] ));
 sg13g2_dfrbp_1 _4914_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net149),
    .D(_0598_),
    .Q_N(_0019_),
    .Q(\coarse_result[3] ));
 sg13g2_dfrbp_1 _4915_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net148),
    .D(_0599_),
    .Q_N(_0022_),
    .Q(\coarse_result[4] ));
 sg13g2_dfrbp_1 _4916_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0600_),
    .Q_N(_0025_),
    .Q(\coarse_result[5] ));
 sg13g2_dfrbp_1 _4917_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net145),
    .D(_0601_),
    .Q_N(_0028_),
    .Q(\coarse_result[6] ));
 sg13g2_dfrbp_1 _4918_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net143),
    .D(_0602_),
    .Q_N(_0031_),
    .Q(\coarse_result[7] ));
 sg13g2_dfrbp_1 _4919_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net142),
    .D(_0603_),
    .Q_N(_1716_),
    .Q(\coarse_result[8] ));
 sg13g2_dfrbp_1 _4920_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net140),
    .D(_0604_),
    .Q_N(_1715_),
    .Q(\coarse_result[9] ));
 sg13g2_dfrbp_1 _4921_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net139),
    .D(_0605_),
    .Q_N(_1714_),
    .Q(\coarse_result[10] ));
 sg13g2_dfrbp_1 _4922_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net137),
    .D(_0606_),
    .Q_N(_1713_),
    .Q(\coarse_result[11] ));
 sg13g2_dfrbp_1 _4923_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net136),
    .D(_0607_),
    .Q_N(_1712_),
    .Q(\coarse_result[12] ));
 sg13g2_dfrbp_1 _4924_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net134),
    .D(_0608_),
    .Q_N(_1711_),
    .Q(\coarse_result[13] ));
 sg13g2_dfrbp_1 _4925_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net133),
    .D(_0609_),
    .Q_N(_1710_),
    .Q(\coarse_result[14] ));
 sg13g2_dfrbp_1 _4926_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net131),
    .D(_0610_),
    .Q_N(_1709_),
    .Q(\coarse_result[15] ));
 sg13g2_dfrbp_1 _4927_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net130),
    .D(_0611_),
    .Q_N(_1708_),
    .Q(\coarse_result[16] ));
 sg13g2_dfrbp_1 _4928_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net128),
    .D(_0612_),
    .Q_N(_1707_),
    .Q(\coarse_result[17] ));
 sg13g2_dfrbp_1 _4929_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net127),
    .D(_0613_),
    .Q_N(_1706_),
    .Q(\coarse_result[18] ));
 sg13g2_dfrbp_1 _4930_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net125),
    .D(_0614_),
    .Q_N(_1705_),
    .Q(\coarse_result[19] ));
 sg13g2_dfrbp_1 _4931_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net124),
    .D(_0615_),
    .Q_N(_1704_),
    .Q(\coarse_result[20] ));
 sg13g2_dfrbp_1 _4932_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net122),
    .D(_0616_),
    .Q_N(_1703_),
    .Q(\coarse_result[21] ));
 sg13g2_dfrbp_1 _4933_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net121),
    .D(_0617_),
    .Q_N(_1702_),
    .Q(\coarse_result[22] ));
 sg13g2_dfrbp_1 _4934_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net119),
    .D(_0618_),
    .Q_N(_1701_),
    .Q(\coarse_result[23] ));
 sg13g2_dfrbp_1 _4935_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net117),
    .D(_0619_),
    .Q_N(_1700_),
    .Q(\coarse_result[24] ));
 sg13g2_dfrbp_1 _4936_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net115),
    .D(_0620_),
    .Q_N(_1699_),
    .Q(\coarse_result[25] ));
 sg13g2_dfrbp_1 _4937_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net113),
    .D(_0621_),
    .Q_N(_1698_),
    .Q(\coarse_result[26] ));
 sg13g2_dfrbp_1 _4938_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net111),
    .D(_0622_),
    .Q_N(_1697_),
    .Q(\coarse_result[27] ));
 sg13g2_dfrbp_1 _4939_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net109),
    .D(_0623_),
    .Q_N(_1696_),
    .Q(\coarse_result[28] ));
 sg13g2_dfrbp_1 _4940_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net108),
    .D(_0624_),
    .Q_N(_1695_),
    .Q(\coarse_result[29] ));
 sg13g2_dfrbp_1 _4941_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net106),
    .D(_0625_),
    .Q_N(_1694_),
    .Q(\coarse_result[30] ));
 sg13g2_dfrbp_1 _4942_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net104),
    .D(_0626_),
    .Q_N(_1693_),
    .Q(\coarse_result[31] ));
 sg13g2_dfrbp_1 _4943_ (.CLK(net3),
    .RESET_B(net102),
    .D(_0627_),
    .Q_N(_1692_),
    .Q(\tdc_inst.start_signal_sampling_clock_level ));
 sg13g2_dfrbp_1 _4944_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net101),
    .D(_0628_),
    .Q_N(_1691_),
    .Q(\tdc_inst.tdc_xor_result[142] ));
 sg13g2_dfrbp_1 _4945_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net99),
    .D(_0629_),
    .Q_N(_1690_),
    .Q(\tdc_inst.start_count_debug[142] ));
 sg13g2_dfrbp_1 _4946_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net97),
    .D(_0630_),
    .Q_N(_1689_),
    .Q(\tdc_inst.stop_count_debug[142] ));
 sg13g2_dfrbp_1 _4947_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net95),
    .D(_0631_),
    .Q_N(_1688_),
    .Q(\tdc_inst.fine_procedure_counter[0] ));
 sg13g2_dfrbp_1 _4948_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net93),
    .D(_0632_),
    .Q_N(_1687_),
    .Q(\tdc_inst.fine_procedure_counter[1] ));
 sg13g2_dfrbp_1 _4949_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net92),
    .D(_0633_),
    .Q_N(_1686_),
    .Q(\tdc_inst.fine_procedure_counter[2] ));
 sg13g2_dfrbp_1 _4950_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net91),
    .D(_0634_),
    .Q_N(_1685_),
    .Q(\tdc_inst.fine_procedure_counter[3] ));
 sg13g2_dfrbp_1 _4951_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net90),
    .D(_0635_),
    .Q_N(_0005_),
    .Q(\tdc_inst.fine_procedure_counter[4] ));
 sg13g2_dfrbp_1 _4952_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net89),
    .D(_0636_),
    .Q_N(_1684_),
    .Q(\tdc_inst.fine_procedure_counter[5] ));
 sg13g2_dfrbp_1 _4953_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net88),
    .D(net1775),
    .Q_N(_1683_),
    .Q(\tdc_inst.fine_procedure_counter[6] ));
 sg13g2_dfrbp_1 _4954_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net87),
    .D(_0638_),
    .Q_N(_1682_),
    .Q(\tdc_inst.fine_procedure_counter[7] ));
 sg13g2_dfrbp_1 _4955_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net86),
    .D(_0639_),
    .Q_N(_0006_),
    .Q(\tdc_inst.fine_procedure_counter[8] ));
 sg13g2_dfrbp_1 _4956_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net85),
    .D(_0640_),
    .Q_N(_0032_),
    .Q(\tdc_inst.fine_another_counter[1] ));
 sg13g2_dfrbp_1 _4957_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net84),
    .D(_0641_),
    .Q_N(_0033_),
    .Q(\tdc_inst.fine_another_counter[2] ));
 sg13g2_dfrbp_1 _4958_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net83),
    .D(_0642_),
    .Q_N(_0034_),
    .Q(\tdc_inst.fine_another_counter[3] ));
 sg13g2_dfrbp_1 _4959_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net82),
    .D(_0643_),
    .Q_N(_0035_),
    .Q(\tdc_inst.fine_another_counter[4] ));
 sg13g2_dfrbp_1 _4960_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net81),
    .D(_0644_),
    .Q_N(_1681_),
    .Q(\tdc_inst.fine_another_counter[5] ));
 sg13g2_dfrbp_1 _4961_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net80),
    .D(_0645_),
    .Q_N(_0036_),
    .Q(\tdc_inst.fine_another_counter[6] ));
 sg13g2_dfrbp_1 _4962_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net79),
    .D(_0646_),
    .Q_N(_0037_),
    .Q(\tdc_inst.fine_another_counter[7] ));
 sg13g2_dfrbp_1 _4963_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net78),
    .D(net1777),
    .Q_N(_0038_),
    .Q(\tdc_inst.fine_another_counter[8] ));
 sg13g2_dfrbp_1 _4964_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net77),
    .D(net1636),
    .Q_N(_1680_),
    .Q(\tdc_inst.fine_start_counter[0] ));
 sg13g2_dfrbp_1 _4965_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net76),
    .D(net1748),
    .Q_N(_1679_),
    .Q(\tdc_inst.fine_start_counter[1] ));
 sg13g2_dfrbp_1 _4966_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net75),
    .D(_0650_),
    .Q_N(_1678_),
    .Q(\tdc_inst.fine_start_counter[2] ));
 sg13g2_dfrbp_1 _4967_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net74),
    .D(net1708),
    .Q_N(_1677_),
    .Q(\tdc_inst.fine_start_counter[3] ));
 sg13g2_dfrbp_1 _4968_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net153),
    .D(net1753),
    .Q_N(_1676_),
    .Q(\tdc_inst.fine_start_counter[4] ));
 sg13g2_dfrbp_1 _4969_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net150),
    .D(_0653_),
    .Q_N(_1675_),
    .Q(\tdc_inst.fine_start_counter[5] ));
 sg13g2_dfrbp_1 _4970_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net147),
    .D(net1739),
    .Q_N(_1674_),
    .Q(\tdc_inst.fine_start_counter[6] ));
 sg13g2_dfrbp_1 _4971_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net144),
    .D(_0655_),
    .Q_N(_1673_),
    .Q(\tdc_inst.fine_start_counter[7] ));
 sg13g2_dfrbp_1 _4972_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net141),
    .D(net1538),
    .Q_N(_1672_),
    .Q(\tdc_inst.fine_start_counter[8] ));
 sg13g2_dfrbp_1 _4973_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net138),
    .D(net1429),
    .Q_N(_1671_),
    .Q(\tdc_inst.fine_stop_counter[0] ));
 sg13g2_dfrbp_1 _4974_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net135),
    .D(net1711),
    .Q_N(_1670_),
    .Q(\tdc_inst.fine_stop_counter[1] ));
 sg13g2_dfrbp_1 _4975_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net132),
    .D(_0659_),
    .Q_N(_1669_),
    .Q(\tdc_inst.fine_stop_counter[2] ));
 sg13g2_dfrbp_1 _4976_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net129),
    .D(_0660_),
    .Q_N(_1668_),
    .Q(\tdc_inst.fine_stop_counter[3] ));
 sg13g2_dfrbp_1 _4977_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net126),
    .D(_0661_),
    .Q_N(_1667_),
    .Q(\tdc_inst.fine_stop_counter[4] ));
 sg13g2_dfrbp_1 _4978_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net123),
    .D(_0662_),
    .Q_N(_1666_),
    .Q(\tdc_inst.fine_stop_counter[5] ));
 sg13g2_dfrbp_1 _4979_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net120),
    .D(_0663_),
    .Q_N(_1665_),
    .Q(\tdc_inst.fine_stop_counter[6] ));
 sg13g2_dfrbp_1 _4980_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net116),
    .D(net1797),
    .Q_N(_1664_),
    .Q(\tdc_inst.fine_stop_counter[7] ));
 sg13g2_dfrbp_1 _4981_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net112),
    .D(net1713),
    .Q_N(_1663_),
    .Q(\tdc_inst.fine_stop_counter[8] ));
 sg13g2_dfrbp_1 _4982_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1245),
    .D(_0666_),
    .Q_N(_1662_),
    .Q(spi_mosi_sync));
 sg13g2_dfrbp_1 _4983_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net107),
    .D(_0667_),
    .Q_N(_1661_),
    .Q(\tdc_inst.reset_internal_logic ));
 sg13g2_dfrbp_1 _4984_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net103),
    .D(_0668_),
    .Q_N(_1660_),
    .Q(\tdc_inst.positions_sum[4] ));
 sg13g2_dfrbp_1 _4985_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net100),
    .D(_0669_),
    .Q_N(_1659_),
    .Q(\tdc_inst.positions_sum[5] ));
 sg13g2_dfrbp_1 _4986_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net98),
    .D(_0670_),
    .Q_N(_1658_),
    .Q(\tdc_inst.positions_sum[6] ));
 sg13g2_dfrbp_1 _4987_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net96),
    .D(_0671_),
    .Q_N(_1657_),
    .Q(\tdc_inst.positions_sum[7] ));
 sg13g2_dfrbp_1 _4988_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net94),
    .D(net1625),
    .Q_N(_1656_),
    .Q(\tdc_inst.positions_sum[8] ));
 sg13g2_dfrbp_1 _4989_ (.CLK(net1235),
    .RESET_B(\tdc_inst.reset_internal_logic ),
    .D(_0673_),
    .Q_N(_0044_),
    .Q(\tdc_inst.coarse_count[0] ));
 sg13g2_dfrbp_1 _4990_ (.CLK(net1235),
    .RESET_B(net1215),
    .D(_0674_),
    .Q_N(_1655_),
    .Q(\tdc_inst.coarse_count[1] ));
 sg13g2_dfrbp_1 _4991_ (.CLK(net1235),
    .RESET_B(\tdc_inst.reset_internal_logic ),
    .D(_0675_),
    .Q_N(_1654_),
    .Q(\tdc_inst.coarse_count[2] ));
 sg13g2_dfrbp_1 _4992_ (.CLK(net1235),
    .RESET_B(net1214),
    .D(_0676_),
    .Q_N(_1653_),
    .Q(\tdc_inst.coarse_count[3] ));
 sg13g2_dfrbp_1 _4993_ (.CLK(net1233),
    .RESET_B(net1214),
    .D(_0677_),
    .Q_N(_1652_),
    .Q(\tdc_inst.coarse_count[4] ));
 sg13g2_dfrbp_1 _4994_ (.CLK(net1233),
    .RESET_B(net1214),
    .D(_0678_),
    .Q_N(_1651_),
    .Q(\tdc_inst.coarse_count[5] ));
 sg13g2_dfrbp_1 _4995_ (.CLK(net1233),
    .RESET_B(net1214),
    .D(_0679_),
    .Q_N(_1650_),
    .Q(\tdc_inst.coarse_count[6] ));
 sg13g2_dfrbp_1 _4996_ (.CLK(net1233),
    .RESET_B(net1214),
    .D(_0680_),
    .Q_N(_1649_),
    .Q(\tdc_inst.coarse_count[7] ));
 sg13g2_dfrbp_1 _4997_ (.CLK(net1233),
    .RESET_B(net1213),
    .D(_0681_),
    .Q_N(_1648_),
    .Q(\tdc_inst.coarse_count[8] ));
 sg13g2_dfrbp_1 _4998_ (.CLK(net1232),
    .RESET_B(net1214),
    .D(_0682_),
    .Q_N(_1647_),
    .Q(\tdc_inst.coarse_count[9] ));
 sg13g2_dfrbp_1 _4999_ (.CLK(net1232),
    .RESET_B(net1213),
    .D(_0683_),
    .Q_N(_1646_),
    .Q(\tdc_inst.coarse_count[10] ));
 sg13g2_dfrbp_1 _5000_ (.CLK(net1232),
    .RESET_B(net1213),
    .D(_0684_),
    .Q_N(_1645_),
    .Q(\tdc_inst.coarse_count[11] ));
 sg13g2_dfrbp_1 _5001_ (.CLK(net1232),
    .RESET_B(net1213),
    .D(_0685_),
    .Q_N(_1644_),
    .Q(\tdc_inst.coarse_count[12] ));
 sg13g2_dfrbp_1 _5002_ (.CLK(net1232),
    .RESET_B(net1213),
    .D(_0686_),
    .Q_N(_1643_),
    .Q(\tdc_inst.coarse_count[13] ));
 sg13g2_dfrbp_1 _5003_ (.CLK(net1232),
    .RESET_B(net1213),
    .D(_0687_),
    .Q_N(_0039_),
    .Q(\tdc_inst.coarse_count[14] ));
 sg13g2_dfrbp_1 _5004_ (.CLK(net1232),
    .RESET_B(net1213),
    .D(_0688_),
    .Q_N(_1642_),
    .Q(\tdc_inst.coarse_count[15] ));
 sg13g2_dfrbp_1 _5005_ (.CLK(net1232),
    .RESET_B(net1213),
    .D(_0689_),
    .Q_N(_1641_),
    .Q(\tdc_inst.coarse_count[16] ));
 sg13g2_dfrbp_1 _5006_ (.CLK(net1231),
    .RESET_B(net1212),
    .D(_0690_),
    .Q_N(_1640_),
    .Q(\tdc_inst.coarse_count[17] ));
 sg13g2_dfrbp_1 _5007_ (.CLK(net1231),
    .RESET_B(net1212),
    .D(_0691_),
    .Q_N(_0040_),
    .Q(\tdc_inst.coarse_count[18] ));
 sg13g2_dfrbp_1 _5008_ (.CLK(net1230),
    .RESET_B(net1212),
    .D(_0692_),
    .Q_N(_1639_),
    .Q(\tdc_inst.coarse_count[19] ));
 sg13g2_dfrbp_1 _5009_ (.CLK(net1231),
    .RESET_B(net1212),
    .D(_0693_),
    .Q_N(_1638_),
    .Q(\tdc_inst.coarse_count[20] ));
 sg13g2_dfrbp_1 _5010_ (.CLK(net1231),
    .RESET_B(net1211),
    .D(_0694_),
    .Q_N(_1637_),
    .Q(\tdc_inst.coarse_count[21] ));
 sg13g2_dfrbp_1 _5011_ (.CLK(net1231),
    .RESET_B(net1212),
    .D(_0695_),
    .Q_N(_0041_),
    .Q(\tdc_inst.coarse_count[22] ));
 sg13g2_dfrbp_1 _5012_ (.CLK(net1231),
    .RESET_B(net1211),
    .D(_0696_),
    .Q_N(_1636_),
    .Q(\tdc_inst.coarse_count[23] ));
 sg13g2_dfrbp_1 _5013_ (.CLK(net1230),
    .RESET_B(net1211),
    .D(_0697_),
    .Q_N(_1635_),
    .Q(\tdc_inst.coarse_count[24] ));
 sg13g2_dfrbp_1 _5014_ (.CLK(net1230),
    .RESET_B(net1211),
    .D(_0698_),
    .Q_N(_1634_),
    .Q(\tdc_inst.coarse_count[25] ));
 sg13g2_dfrbp_1 _5015_ (.CLK(net1230),
    .RESET_B(net1211),
    .D(_0699_),
    .Q_N(_0042_),
    .Q(\tdc_inst.coarse_count[26] ));
 sg13g2_dfrbp_1 _5016_ (.CLK(net1230),
    .RESET_B(net1211),
    .D(_0700_),
    .Q_N(_1633_),
    .Q(\tdc_inst.coarse_count[27] ));
 sg13g2_dfrbp_1 _5017_ (.CLK(net1230),
    .RESET_B(net1211),
    .D(_0701_),
    .Q_N(_1632_),
    .Q(\tdc_inst.coarse_count[28] ));
 sg13g2_dfrbp_1 _5018_ (.CLK(net1230),
    .RESET_B(net1212),
    .D(_0702_),
    .Q_N(_1631_),
    .Q(\tdc_inst.coarse_count[29] ));
 sg13g2_dfrbp_1 _5019_ (.CLK(net1230),
    .RESET_B(net1211),
    .D(_0703_),
    .Q_N(_0043_),
    .Q(\tdc_inst.coarse_count[30] ));
 sg13g2_dfrbp_1 _5020_ (.CLK(net1234),
    .RESET_B(net1215),
    .D(_0704_),
    .Q_N(_2252_),
    .Q(\tdc_inst.coarse_count[31] ));
 sg13g2_dfrbp_1 _5021_ (.CLK(net4),
    .RESET_B(net1215),
    .D(net118),
    .Q_N(_0004_),
    .Q(\tdc_inst.stop_signal_activated ));
 sg13g2_dfrbp_1 _5022_ (.CLK(net4),
    .RESET_B(net105),
    .D(_0705_),
    .Q_N(_2253_),
    .Q(\tdc_inst.stop_signal_sampling_clock_level ));
 sg13g2_dfrbp_1 _5023_ (.CLK(net3),
    .RESET_B(\tdc_inst.reset_internal_logic ),
    .D(net114),
    .Q_N(_1630_),
    .Q(\tdc_inst.start_signal_activated ));
 sg13g2_dfrbp_1 _5024_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net110),
    .D(net1768),
    .Q_N(_1629_),
    .Q(\tdc_inst.fine_another_counter[0] ));
 sg13g2_tiehi _4406__26 (.L_HI(net26));
 sg13g2_tiehi _4405__27 (.L_HI(net27));
 sg13g2_tiehi _4404__28 (.L_HI(net28));
 sg13g2_tiehi _4403__29 (.L_HI(net29));
 sg13g2_tiehi _4402__30 (.L_HI(net30));
 sg13g2_tiehi _4401__31 (.L_HI(net31));
 sg13g2_tiehi _4400__32 (.L_HI(net32));
 sg13g2_tiehi _4399__33 (.L_HI(net33));
 sg13g2_tiehi _4398__34 (.L_HI(net34));
 sg13g2_tiehi _4397__35 (.L_HI(net35));
 sg13g2_tiehi _4396__36 (.L_HI(net36));
 sg13g2_tiehi _4395__37 (.L_HI(net37));
 sg13g2_tiehi _4394__38 (.L_HI(net38));
 sg13g2_tiehi _4393__39 (.L_HI(net39));
 sg13g2_tiehi _4392__40 (.L_HI(net40));
 sg13g2_tiehi _4391__41 (.L_HI(net41));
 sg13g2_tiehi _4390__42 (.L_HI(net42));
 sg13g2_tiehi _4389__43 (.L_HI(net43));
 sg13g2_tiehi _4388__44 (.L_HI(net44));
 sg13g2_tiehi _4387__45 (.L_HI(net45));
 sg13g2_tiehi _4386__46 (.L_HI(net46));
 sg13g2_tiehi _4385__47 (.L_HI(net47));
 sg13g2_tiehi _4384__48 (.L_HI(net48));
 sg13g2_tiehi _4383__49 (.L_HI(net49));
 sg13g2_tiehi _4382__50 (.L_HI(net50));
 sg13g2_tiehi _4381__51 (.L_HI(net51));
 sg13g2_tiehi _4380__52 (.L_HI(net52));
 sg13g2_tiehi _4379__53 (.L_HI(net53));
 sg13g2_tiehi _4378__54 (.L_HI(net54));
 sg13g2_tiehi _4377__55 (.L_HI(net55));
 sg13g2_tiehi _4376__56 (.L_HI(net56));
 sg13g2_tiehi _4375__57 (.L_HI(net57));
 sg13g2_tiehi _4374__58 (.L_HI(net58));
 sg13g2_tiehi _4373__59 (.L_HI(net59));
 sg13g2_tiehi _4372__60 (.L_HI(net60));
 sg13g2_tiehi _4371__61 (.L_HI(net61));
 sg13g2_tiehi _4370__62 (.L_HI(net62));
 sg13g2_tiehi _4369__63 (.L_HI(net63));
 sg13g2_tiehi _4368__64 (.L_HI(net64));
 sg13g2_tiehi _4367__65 (.L_HI(net65));
 sg13g2_tiehi _4366__66 (.L_HI(net66));
 sg13g2_tiehi _4365__67 (.L_HI(net67));
 sg13g2_tiehi _4364__68 (.L_HI(net68));
 sg13g2_tiehi _4363__69 (.L_HI(net69));
 sg13g2_tiehi _4362__70 (.L_HI(net70));
 sg13g2_tiehi _4361__71 (.L_HI(net71));
 sg13g2_tiehi _4360__72 (.L_HI(net72));
 sg13g2_tiehi _4359__73 (.L_HI(net73));
 sg13g2_tiehi _4967__74 (.L_HI(net74));
 sg13g2_tiehi _4966__75 (.L_HI(net75));
 sg13g2_tiehi _4965__76 (.L_HI(net76));
 sg13g2_tiehi _4964__77 (.L_HI(net77));
 sg13g2_tiehi _4963__78 (.L_HI(net78));
 sg13g2_tiehi _4962__79 (.L_HI(net79));
 sg13g2_tiehi _4961__80 (.L_HI(net80));
 sg13g2_tiehi _4960__81 (.L_HI(net81));
 sg13g2_tiehi _4959__82 (.L_HI(net82));
 sg13g2_tiehi _4958__83 (.L_HI(net83));
 sg13g2_tiehi _4957__84 (.L_HI(net84));
 sg13g2_tiehi _4956__85 (.L_HI(net85));
 sg13g2_tiehi _4955__86 (.L_HI(net86));
 sg13g2_tiehi _4954__87 (.L_HI(net87));
 sg13g2_tiehi _4953__88 (.L_HI(net88));
 sg13g2_tiehi _4952__89 (.L_HI(net89));
 sg13g2_tiehi _4951__90 (.L_HI(net90));
 sg13g2_tiehi _4950__91 (.L_HI(net91));
 sg13g2_tiehi _4949__92 (.L_HI(net92));
 sg13g2_tiehi _4948__93 (.L_HI(net93));
 sg13g2_tiehi _4988__94 (.L_HI(net94));
 sg13g2_tiehi _4947__95 (.L_HI(net95));
 sg13g2_tiehi _4987__96 (.L_HI(net96));
 sg13g2_tiehi _4946__97 (.L_HI(net97));
 sg13g2_tiehi _4986__98 (.L_HI(net98));
 sg13g2_tiehi _4945__99 (.L_HI(net99));
 sg13g2_tiehi _4985__100 (.L_HI(net100));
 sg13g2_tiehi _4944__101 (.L_HI(net101));
 sg13g2_tiehi _4943__102 (.L_HI(net102));
 sg13g2_tiehi _4984__103 (.L_HI(net103));
 sg13g2_tiehi _4942__104 (.L_HI(net104));
 sg13g2_tiehi _5022__105 (.L_HI(net105));
 sg13g2_tiehi _4941__106 (.L_HI(net106));
 sg13g2_tiehi _4983__107 (.L_HI(net107));
 sg13g2_tiehi _4940__108 (.L_HI(net108));
 sg13g2_tiehi _4939__109 (.L_HI(net109));
 sg13g2_tiehi _5024__110 (.L_HI(net110));
 sg13g2_tiehi _4938__111 (.L_HI(net111));
 sg13g2_tiehi _4981__112 (.L_HI(net112));
 sg13g2_tiehi _4937__113 (.L_HI(net113));
 sg13g2_tiehi _5023__114 (.L_HI(net114));
 sg13g2_tiehi _4936__115 (.L_HI(net115));
 sg13g2_tiehi _4980__116 (.L_HI(net116));
 sg13g2_tiehi _4935__117 (.L_HI(net117));
 sg13g2_tiehi _5021__118 (.L_HI(net118));
 sg13g2_tiehi _4934__119 (.L_HI(net119));
 sg13g2_tiehi _4979__120 (.L_HI(net120));
 sg13g2_tiehi _4933__121 (.L_HI(net121));
 sg13g2_tiehi _4932__122 (.L_HI(net122));
 sg13g2_tiehi _4978__123 (.L_HI(net123));
 sg13g2_tiehi _4931__124 (.L_HI(net124));
 sg13g2_tiehi _4930__125 (.L_HI(net125));
 sg13g2_tiehi _4977__126 (.L_HI(net126));
 sg13g2_tiehi _4929__127 (.L_HI(net127));
 sg13g2_tiehi _4928__128 (.L_HI(net128));
 sg13g2_tiehi _4976__129 (.L_HI(net129));
 sg13g2_tiehi _4927__130 (.L_HI(net130));
 sg13g2_tiehi _4926__131 (.L_HI(net131));
 sg13g2_tiehi _4975__132 (.L_HI(net132));
 sg13g2_tiehi _4925__133 (.L_HI(net133));
 sg13g2_tiehi _4924__134 (.L_HI(net134));
 sg13g2_tiehi _4974__135 (.L_HI(net135));
 sg13g2_tiehi _4923__136 (.L_HI(net136));
 sg13g2_tiehi _4922__137 (.L_HI(net137));
 sg13g2_tiehi _4973__138 (.L_HI(net138));
 sg13g2_tiehi _4921__139 (.L_HI(net139));
 sg13g2_tiehi _4920__140 (.L_HI(net140));
 sg13g2_tiehi _4972__141 (.L_HI(net141));
 sg13g2_tiehi _4919__142 (.L_HI(net142));
 sg13g2_tiehi _4918__143 (.L_HI(net143));
 sg13g2_tiehi _4971__144 (.L_HI(net144));
 sg13g2_tiehi _4917__145 (.L_HI(net145));
 sg13g2_tiehi _4916__146 (.L_HI(net146));
 sg13g2_tiehi _4970__147 (.L_HI(net147));
 sg13g2_tiehi _4915__148 (.L_HI(net148));
 sg13g2_tiehi _4914__149 (.L_HI(net149));
 sg13g2_tiehi _4969__150 (.L_HI(net150));
 sg13g2_tiehi _4913__151 (.L_HI(net151));
 sg13g2_tiehi _4912__152 (.L_HI(net152));
 sg13g2_tiehi _4968__153 (.L_HI(net153));
 sg13g2_tiehi _4911__154 (.L_HI(net154));
 sg13g2_tiehi _4845__155 (.L_HI(net155));
 sg13g2_tiehi _4844__156 (.L_HI(net156));
 sg13g2_tiehi _4843__157 (.L_HI(net157));
 sg13g2_tiehi _4842__158 (.L_HI(net158));
 sg13g2_tiehi _4841__159 (.L_HI(net159));
 sg13g2_tiehi _4840__160 (.L_HI(net160));
 sg13g2_tiehi _4839__161 (.L_HI(net161));
 sg13g2_tiehi _4838__162 (.L_HI(net162));
 sg13g2_tiehi _4837__163 (.L_HI(net163));
 sg13g2_tiehi _4793__164 (.L_HI(net164));
 sg13g2_tiehi _4792__165 (.L_HI(net165));
 sg13g2_tiehi _4791__166 (.L_HI(net166));
 sg13g2_tiehi _4790__167 (.L_HI(net167));
 sg13g2_tiehi _4789__168 (.L_HI(net168));
 sg13g2_tiehi _4788__169 (.L_HI(net169));
 sg13g2_tiehi _4787__170 (.L_HI(net170));
 sg13g2_tiehi _4786__171 (.L_HI(net171));
 sg13g2_tiehi _4785__172 (.L_HI(net172));
 sg13g2_tiehi _4784__173 (.L_HI(net173));
 sg13g2_tiehi _4783__174 (.L_HI(net174));
 sg13g2_tiehi _4782__175 (.L_HI(net175));
 sg13g2_tiehi _4781__176 (.L_HI(net176));
 sg13g2_tiehi _4780__177 (.L_HI(net177));
 sg13g2_tiehi _4779__178 (.L_HI(net178));
 sg13g2_tiehi _4778__179 (.L_HI(net179));
 sg13g2_tiehi _4777__180 (.L_HI(net180));
 sg13g2_tiehi _4776__181 (.L_HI(net181));
 sg13g2_tiehi _4775__182 (.L_HI(net182));
 sg13g2_tiehi _4774__183 (.L_HI(net183));
 sg13g2_tiehi _4773__184 (.L_HI(net184));
 sg13g2_tiehi _4772__185 (.L_HI(net185));
 sg13g2_tiehi _4771__186 (.L_HI(net186));
 sg13g2_tiehi _4770__187 (.L_HI(net187));
 sg13g2_tiehi _4769__188 (.L_HI(net188));
 sg13g2_tiehi _4768__189 (.L_HI(net189));
 sg13g2_tiehi _4767__190 (.L_HI(net190));
 sg13g2_tiehi _4766__191 (.L_HI(net191));
 sg13g2_tiehi _4765__192 (.L_HI(net192));
 sg13g2_tiehi _4764__193 (.L_HI(net193));
 sg13g2_tiehi _4763__194 (.L_HI(net194));
 sg13g2_tiehi _4762__195 (.L_HI(net195));
 sg13g2_tiehi _4761__196 (.L_HI(net196));
 sg13g2_tiehi _4760__197 (.L_HI(net197));
 sg13g2_tiehi _4759__198 (.L_HI(net198));
 sg13g2_tiehi _4758__199 (.L_HI(net199));
 sg13g2_tiehi _4757__200 (.L_HI(net200));
 sg13g2_tiehi _4756__201 (.L_HI(net201));
 sg13g2_tiehi _4755__202 (.L_HI(net202));
 sg13g2_tiehi _4754__203 (.L_HI(net203));
 sg13g2_tiehi _4753__204 (.L_HI(net204));
 sg13g2_tiehi _4752__205 (.L_HI(net205));
 sg13g2_tiehi _4751__206 (.L_HI(net206));
 sg13g2_tiehi _4750__207 (.L_HI(net207));
 sg13g2_tiehi _4749__208 (.L_HI(net208));
 sg13g2_tiehi _4748__209 (.L_HI(net209));
 sg13g2_tiehi _4747__210 (.L_HI(net210));
 sg13g2_tiehi _4746__211 (.L_HI(net211));
 sg13g2_tiehi _4745__212 (.L_HI(net212));
 sg13g2_tiehi _4744__213 (.L_HI(net213));
 sg13g2_tiehi _4743__214 (.L_HI(net214));
 sg13g2_tiehi _4742__215 (.L_HI(net215));
 sg13g2_tiehi _4741__216 (.L_HI(net216));
 sg13g2_tiehi _4740__217 (.L_HI(net217));
 sg13g2_tiehi _4739__218 (.L_HI(net218));
 sg13g2_tiehi _4738__219 (.L_HI(net219));
 sg13g2_tiehi _4737__220 (.L_HI(net220));
 sg13g2_tiehi _4736__221 (.L_HI(net221));
 sg13g2_tiehi _4735__222 (.L_HI(net222));
 sg13g2_tiehi _4734__223 (.L_HI(net223));
 sg13g2_tiehi _4733__224 (.L_HI(net224));
 sg13g2_tiehi _4732__225 (.L_HI(net225));
 sg13g2_tiehi _4731__226 (.L_HI(net226));
 sg13g2_tiehi _4730__227 (.L_HI(net227));
 sg13g2_tiehi _4729__228 (.L_HI(net228));
 sg13g2_tiehi _4728__229 (.L_HI(net229));
 sg13g2_tiehi _4727__230 (.L_HI(net230));
 sg13g2_tiehi _4726__231 (.L_HI(net231));
 sg13g2_tiehi _4725__232 (.L_HI(net232));
 sg13g2_tiehi _4724__233 (.L_HI(net233));
 sg13g2_tiehi _4723__234 (.L_HI(net234));
 sg13g2_tiehi _4722__235 (.L_HI(net235));
 sg13g2_tiehi _4721__236 (.L_HI(net236));
 sg13g2_tiehi _4720__237 (.L_HI(net237));
 sg13g2_tiehi _4719__238 (.L_HI(net238));
 sg13g2_tiehi _4718__239 (.L_HI(net239));
 sg13g2_tiehi _4717__240 (.L_HI(net240));
 sg13g2_tiehi _4716__241 (.L_HI(net241));
 sg13g2_tiehi _4715__242 (.L_HI(net242));
 sg13g2_tiehi _4714__243 (.L_HI(net243));
 sg13g2_tiehi _4713__244 (.L_HI(net244));
 sg13g2_tiehi _4712__245 (.L_HI(net245));
 sg13g2_tiehi _4711__246 (.L_HI(net246));
 sg13g2_tiehi _4710__247 (.L_HI(net247));
 sg13g2_tiehi _4709__248 (.L_HI(net248));
 sg13g2_tiehi _4708__249 (.L_HI(net249));
 sg13g2_tiehi _4707__250 (.L_HI(net250));
 sg13g2_tiehi _4706__251 (.L_HI(net251));
 sg13g2_tiehi _4705__252 (.L_HI(net252));
 sg13g2_tiehi _4704__253 (.L_HI(net253));
 sg13g2_tiehi _4703__254 (.L_HI(net254));
 sg13g2_tiehi _4702__255 (.L_HI(net255));
 sg13g2_tiehi _4701__256 (.L_HI(net256));
 sg13g2_tiehi _4700__257 (.L_HI(net257));
 sg13g2_tiehi _4699__258 (.L_HI(net258));
 sg13g2_tiehi _4698__259 (.L_HI(net259));
 sg13g2_tiehi _4697__260 (.L_HI(net260));
 sg13g2_tiehi _4696__261 (.L_HI(net261));
 sg13g2_tiehi _4695__262 (.L_HI(net262));
 sg13g2_tiehi _4694__263 (.L_HI(net263));
 sg13g2_tiehi _4693__264 (.L_HI(net264));
 sg13g2_tiehi _4692__265 (.L_HI(net265));
 sg13g2_tiehi _4691__266 (.L_HI(net266));
 sg13g2_tiehi _4690__267 (.L_HI(net267));
 sg13g2_tiehi _4689__268 (.L_HI(net268));
 sg13g2_tiehi _4688__269 (.L_HI(net269));
 sg13g2_tiehi _4687__270 (.L_HI(net270));
 sg13g2_tiehi _4686__271 (.L_HI(net271));
 sg13g2_tiehi _4685__272 (.L_HI(net272));
 sg13g2_tiehi _4684__273 (.L_HI(net273));
 sg13g2_tiehi _4683__274 (.L_HI(net274));
 sg13g2_tiehi _4682__275 (.L_HI(net275));
 sg13g2_tiehi _4681__276 (.L_HI(net276));
 sg13g2_tiehi _4680__277 (.L_HI(net277));
 sg13g2_tiehi _4679__278 (.L_HI(net278));
 sg13g2_tiehi _4678__279 (.L_HI(net279));
 sg13g2_tiehi _4677__280 (.L_HI(net280));
 sg13g2_tiehi _4676__281 (.L_HI(net281));
 sg13g2_tiehi _4675__282 (.L_HI(net282));
 sg13g2_tiehi _4674__283 (.L_HI(net283));
 sg13g2_tiehi _4673__284 (.L_HI(net284));
 sg13g2_tiehi _4672__285 (.L_HI(net285));
 sg13g2_tiehi _4671__286 (.L_HI(net286));
 sg13g2_tiehi _4670__287 (.L_HI(net287));
 sg13g2_tiehi _4669__288 (.L_HI(net288));
 sg13g2_tiehi _4668__289 (.L_HI(net289));
 sg13g2_tiehi _4667__290 (.L_HI(net290));
 sg13g2_tiehi _4666__291 (.L_HI(net291));
 sg13g2_tiehi _4665__292 (.L_HI(net292));
 sg13g2_tiehi _4664__293 (.L_HI(net293));
 sg13g2_tiehi _4663__294 (.L_HI(net294));
 sg13g2_tiehi _4662__295 (.L_HI(net295));
 sg13g2_tiehi _4661__296 (.L_HI(net296));
 sg13g2_tiehi _4660__297 (.L_HI(net297));
 sg13g2_tiehi _4659__298 (.L_HI(net298));
 sg13g2_tiehi _4658__299 (.L_HI(net299));
 sg13g2_tiehi _4657__300 (.L_HI(net300));
 sg13g2_tiehi _4656__301 (.L_HI(net301));
 sg13g2_tiehi _4655__302 (.L_HI(net302));
 sg13g2_tiehi _4654__303 (.L_HI(net303));
 sg13g2_tiehi _4653__304 (.L_HI(net304));
 sg13g2_tiehi _4652__305 (.L_HI(net305));
 sg13g2_tiehi _4641__306 (.L_HI(net306));
 sg13g2_tiehi _4640__307 (.L_HI(net307));
 sg13g2_tiehi _4639__308 (.L_HI(net308));
 sg13g2_tiehi _4638__309 (.L_HI(net309));
 sg13g2_tiehi _4637__310 (.L_HI(net310));
 sg13g2_tiehi _4636__311 (.L_HI(net311));
 sg13g2_tiehi _4635__312 (.L_HI(net312));
 sg13g2_tiehi _4634__313 (.L_HI(net313));
 sg13g2_tiehi _4633__314 (.L_HI(net314));
 sg13g2_tiehi _4632__315 (.L_HI(net315));
 sg13g2_tiehi _4358__316 (.L_HI(net316));
 sg13g2_tiehi _4631__317 (.L_HI(net317));
 sg13g2_tiehi _4630__318 (.L_HI(net318));
 sg13g2_tiehi _4629__319 (.L_HI(net319));
 sg13g2_tiehi _4628__320 (.L_HI(net320));
 sg13g2_tiehi _4627__321 (.L_HI(net321));
 sg13g2_tiehi _4626__322 (.L_HI(net322));
 sg13g2_tiehi _4625__323 (.L_HI(net323));
 sg13g2_tiehi _4624__324 (.L_HI(net324));
 sg13g2_tiehi _4623__325 (.L_HI(net325));
 sg13g2_tiehi _4622__326 (.L_HI(net326));
 sg13g2_tiehi _4621__327 (.L_HI(net327));
 sg13g2_tiehi _4620__328 (.L_HI(net328));
 sg13g2_tiehi _4619__329 (.L_HI(net329));
 sg13g2_tiehi _4618__330 (.L_HI(net330));
 sg13g2_tiehi _4617__331 (.L_HI(net331));
 sg13g2_tiehi _4616__332 (.L_HI(net332));
 sg13g2_tiehi _4615__333 (.L_HI(net333));
 sg13g2_tiehi _4614__334 (.L_HI(net334));
 sg13g2_tiehi _4613__335 (.L_HI(net335));
 sg13g2_tiehi _4612__336 (.L_HI(net336));
 sg13g2_tiehi _4611__337 (.L_HI(net337));
 sg13g2_tiehi _4610__338 (.L_HI(net338));
 sg13g2_tiehi _4609__339 (.L_HI(net339));
 sg13g2_tiehi _4608__340 (.L_HI(net340));
 sg13g2_tiehi _4607__341 (.L_HI(net341));
 sg13g2_tiehi _4606__342 (.L_HI(net342));
 sg13g2_tiehi _4605__343 (.L_HI(net343));
 sg13g2_tiehi _4604__344 (.L_HI(net344));
 sg13g2_tiehi _4603__345 (.L_HI(net345));
 sg13g2_tiehi _4602__346 (.L_HI(net346));
 sg13g2_tiehi _4601__347 (.L_HI(net347));
 sg13g2_tiehi _4600__348 (.L_HI(net348));
 sg13g2_tiehi _4599__349 (.L_HI(net349));
 sg13g2_tiehi _4598__350 (.L_HI(net350));
 sg13g2_tiehi _4597__351 (.L_HI(net351));
 sg13g2_tiehi _4596__352 (.L_HI(net352));
 sg13g2_tiehi _4595__353 (.L_HI(net353));
 sg13g2_tiehi _4594__354 (.L_HI(net354));
 sg13g2_tiehi _4593__355 (.L_HI(net355));
 sg13g2_tiehi _4592__356 (.L_HI(net356));
 sg13g2_tiehi _4591__357 (.L_HI(net357));
 sg13g2_tiehi _4590__358 (.L_HI(net358));
 sg13g2_tiehi _4589__359 (.L_HI(net359));
 sg13g2_tiehi _4588__360 (.L_HI(net360));
 sg13g2_tiehi _4587__361 (.L_HI(net361));
 sg13g2_tiehi _4586__362 (.L_HI(net362));
 sg13g2_tiehi _4585__363 (.L_HI(net363));
 sg13g2_tiehi _4584__364 (.L_HI(net364));
 sg13g2_tiehi _4583__365 (.L_HI(net365));
 sg13g2_tiehi _4582__366 (.L_HI(net366));
 sg13g2_tiehi _4581__367 (.L_HI(net367));
 sg13g2_tiehi _4580__368 (.L_HI(net368));
 sg13g2_tiehi _4579__369 (.L_HI(net369));
 sg13g2_tiehi _4578__370 (.L_HI(net370));
 sg13g2_tiehi _4577__371 (.L_HI(net371));
 sg13g2_tiehi _4576__372 (.L_HI(net372));
 sg13g2_tiehi _4575__373 (.L_HI(net373));
 sg13g2_tiehi _4574__374 (.L_HI(net374));
 sg13g2_tiehi _4573__375 (.L_HI(net375));
 sg13g2_tiehi _4572__376 (.L_HI(net376));
 sg13g2_tiehi _4571__377 (.L_HI(net377));
 sg13g2_tiehi _4570__378 (.L_HI(net378));
 sg13g2_tiehi _4569__379 (.L_HI(net379));
 sg13g2_tiehi _4568__380 (.L_HI(net380));
 sg13g2_tiehi _4567__381 (.L_HI(net381));
 sg13g2_tiehi _4566__382 (.L_HI(net382));
 sg13g2_tiehi _4565__383 (.L_HI(net383));
 sg13g2_tiehi _4564__384 (.L_HI(net384));
 sg13g2_tiehi _4563__385 (.L_HI(net385));
 sg13g2_tiehi _4562__386 (.L_HI(net386));
 sg13g2_tiehi _4561__387 (.L_HI(net387));
 sg13g2_tiehi _4560__388 (.L_HI(net388));
 sg13g2_tiehi _4559__389 (.L_HI(net389));
 sg13g2_tiehi _4558__390 (.L_HI(net390));
 sg13g2_tiehi _4557__391 (.L_HI(net391));
 sg13g2_tiehi _4556__392 (.L_HI(net392));
 sg13g2_tiehi _4555__393 (.L_HI(net393));
 sg13g2_tiehi _4554__394 (.L_HI(net394));
 sg13g2_tiehi _4553__395 (.L_HI(net395));
 sg13g2_tiehi _4552__396 (.L_HI(net396));
 sg13g2_tiehi _4551__397 (.L_HI(net397));
 sg13g2_tiehi _4550__398 (.L_HI(net398));
 sg13g2_tiehi _4549__399 (.L_HI(net399));
 sg13g2_tiehi _4548__400 (.L_HI(net400));
 sg13g2_tiehi _4547__401 (.L_HI(net401));
 sg13g2_tiehi _4546__402 (.L_HI(net402));
 sg13g2_tiehi _4545__403 (.L_HI(net403));
 sg13g2_tiehi _4544__404 (.L_HI(net404));
 sg13g2_tiehi _4543__405 (.L_HI(net405));
 sg13g2_tiehi _4542__406 (.L_HI(net406));
 sg13g2_tiehi _4541__407 (.L_HI(net407));
 sg13g2_tiehi _4540__408 (.L_HI(net408));
 sg13g2_tiehi _4539__409 (.L_HI(net409));
 sg13g2_tiehi _4538__410 (.L_HI(net410));
 sg13g2_tiehi _4537__411 (.L_HI(net411));
 sg13g2_tiehi _4536__412 (.L_HI(net412));
 sg13g2_tiehi _4535__413 (.L_HI(net413));
 sg13g2_tiehi _4534__414 (.L_HI(net414));
 sg13g2_tiehi _4533__415 (.L_HI(net415));
 sg13g2_tiehi _4532__416 (.L_HI(net416));
 sg13g2_tiehi _4531__417 (.L_HI(net417));
 sg13g2_tiehi _4530__418 (.L_HI(net418));
 sg13g2_tiehi _4529__419 (.L_HI(net419));
 sg13g2_tiehi _4528__420 (.L_HI(net420));
 sg13g2_tiehi _4527__421 (.L_HI(net421));
 sg13g2_tiehi _4526__422 (.L_HI(net422));
 sg13g2_tiehi _4525__423 (.L_HI(net423));
 sg13g2_tiehi _4524__424 (.L_HI(net424));
 sg13g2_tiehi _4523__425 (.L_HI(net425));
 sg13g2_tiehi _4522__426 (.L_HI(net426));
 sg13g2_tiehi _4521__427 (.L_HI(net427));
 sg13g2_tiehi _4520__428 (.L_HI(net428));
 sg13g2_tiehi _4519__429 (.L_HI(net429));
 sg13g2_tiehi _4518__430 (.L_HI(net430));
 sg13g2_tiehi _4517__431 (.L_HI(net431));
 sg13g2_tiehi _4516__432 (.L_HI(net432));
 sg13g2_tiehi _4515__433 (.L_HI(net433));
 sg13g2_tiehi _4514__434 (.L_HI(net434));
 sg13g2_tiehi _4513__435 (.L_HI(net435));
 sg13g2_tiehi _4512__436 (.L_HI(net436));
 sg13g2_tiehi _4511__437 (.L_HI(net437));
 sg13g2_tiehi _4510__438 (.L_HI(net438));
 sg13g2_tiehi _4509__439 (.L_HI(net439));
 sg13g2_tiehi _4508__440 (.L_HI(net440));
 sg13g2_tiehi _4507__441 (.L_HI(net441));
 sg13g2_tiehi _4506__442 (.L_HI(net442));
 sg13g2_tiehi _4505__443 (.L_HI(net443));
 sg13g2_tiehi _4504__444 (.L_HI(net444));
 sg13g2_tiehi _4503__445 (.L_HI(net445));
 sg13g2_tiehi _4502__446 (.L_HI(net446));
 sg13g2_tiehi _4501__447 (.L_HI(net447));
 sg13g2_tiehi _4500__448 (.L_HI(net448));
 sg13g2_tiehi _4499__449 (.L_HI(net449));
 sg13g2_tiehi _4498__450 (.L_HI(net450));
 sg13g2_tiehi _4497__451 (.L_HI(net451));
 sg13g2_tiehi _4496__452 (.L_HI(net452));
 sg13g2_tiehi _4495__453 (.L_HI(net453));
 sg13g2_tiehi _4494__454 (.L_HI(net454));
 sg13g2_tiehi _4493__455 (.L_HI(net455));
 sg13g2_tiehi _4492__456 (.L_HI(net456));
 sg13g2_tiehi _4491__457 (.L_HI(net457));
 sg13g2_tiehi _4490__458 (.L_HI(net458));
 sg13g2_tiehi _4489__459 (.L_HI(net459));
 sg13g2_tiehi _4488__460 (.L_HI(net460));
 sg13g2_tiehi _4487__461 (.L_HI(net461));
 sg13g2_tiehi _4486__462 (.L_HI(net462));
 sg13g2_tiehi _4485__463 (.L_HI(net463));
 sg13g2_tiehi _4484__464 (.L_HI(net464));
 sg13g2_tiehi _4483__465 (.L_HI(net465));
 sg13g2_tiehi _4482__466 (.L_HI(net466));
 sg13g2_tiehi _4481__467 (.L_HI(net467));
 sg13g2_tiehi _4480__468 (.L_HI(net468));
 sg13g2_tiehi _4479__469 (.L_HI(net469));
 sg13g2_tiehi _4478__470 (.L_HI(net470));
 sg13g2_tiehi _4477__471 (.L_HI(net471));
 sg13g2_tiehi _4476__472 (.L_HI(net472));
 sg13g2_tiehi _4475__473 (.L_HI(net473));
 sg13g2_tiehi _4474__474 (.L_HI(net474));
 sg13g2_tiehi _4473__475 (.L_HI(net475));
 sg13g2_tiehi _4472__476 (.L_HI(net476));
 sg13g2_tiehi _4471__477 (.L_HI(net477));
 sg13g2_tiehi _4470__478 (.L_HI(net478));
 sg13g2_tiehi _4469__479 (.L_HI(net479));
 sg13g2_tiehi _4468__480 (.L_HI(net480));
 sg13g2_tiehi _4467__481 (.L_HI(net481));
 sg13g2_tiehi _4466__482 (.L_HI(net482));
 sg13g2_tiehi _4465__483 (.L_HI(net483));
 sg13g2_tiehi _4464__484 (.L_HI(net484));
 sg13g2_tiehi _4463__485 (.L_HI(net485));
 sg13g2_tiehi _4462__486 (.L_HI(net486));
 sg13g2_tiehi _4461__487 (.L_HI(net487));
 sg13g2_tiehi _4460__488 (.L_HI(net488));
 sg13g2_tiehi _4459__489 (.L_HI(net489));
 sg13g2_tiehi _4458__490 (.L_HI(net490));
 sg13g2_tiehi _4457__491 (.L_HI(net491));
 sg13g2_tiehi _4456__492 (.L_HI(net492));
 sg13g2_tiehi _4455__493 (.L_HI(net493));
 sg13g2_tiehi _4454__494 (.L_HI(net494));
 sg13g2_tiehi _4453__495 (.L_HI(net495));
 sg13g2_tiehi _4452__496 (.L_HI(net496));
 sg13g2_tiehi _4451__497 (.L_HI(net497));
 sg13g2_tiehi _4450__498 (.L_HI(net498));
 sg13g2_tiehi _4449__499 (.L_HI(net499));
 sg13g2_tiehi _4448__500 (.L_HI(net500));
 sg13g2_tiehi _4447__501 (.L_HI(net501));
 sg13g2_tiehi _4446__502 (.L_HI(net502));
 sg13g2_tiehi _4445__503 (.L_HI(net503));
 sg13g2_tiehi _4444__504 (.L_HI(net504));
 sg13g2_tiehi _4443__505 (.L_HI(net505));
 sg13g2_tiehi _4442__506 (.L_HI(net506));
 sg13g2_tiehi _4441__507 (.L_HI(net507));
 sg13g2_tiehi _4440__508 (.L_HI(net508));
 sg13g2_tiehi _4439__509 (.L_HI(net509));
 sg13g2_tiehi _4438__510 (.L_HI(net510));
 sg13g2_tiehi _4437__511 (.L_HI(net511));
 sg13g2_tiehi _4436__512 (.L_HI(net512));
 sg13g2_tiehi _4435__513 (.L_HI(net513));
 sg13g2_tiehi _4434__514 (.L_HI(net514));
 sg13g2_tiehi _4433__515 (.L_HI(net515));
 sg13g2_tiehi _4432__516 (.L_HI(net516));
 sg13g2_tiehi _4431__517 (.L_HI(net517));
 sg13g2_tiehi _4430__518 (.L_HI(net518));
 sg13g2_tiehi _4429__519 (.L_HI(net519));
 sg13g2_tiehi _4428__520 (.L_HI(net520));
 sg13g2_tiehi _4427__521 (.L_HI(net521));
 sg13g2_tiehi _4426__522 (.L_HI(net522));
 sg13g2_tiehi _4425__523 (.L_HI(net523));
 sg13g2_tiehi _4424__524 (.L_HI(net524));
 sg13g2_tiehi _4423__525 (.L_HI(net525));
 sg13g2_tiehi _4422__526 (.L_HI(net526));
 sg13g2_tiehi _4421__527 (.L_HI(net527));
 sg13g2_tiehi _4420__528 (.L_HI(net528));
 sg13g2_tiehi _4419__529 (.L_HI(net529));
 sg13g2_tiehi _4418__530 (.L_HI(net530));
 sg13g2_tiehi _4417__531 (.L_HI(net531));
 sg13g2_tiehi _4416__532 (.L_HI(net532));
 sg13g2_tiehi _4415__533 (.L_HI(net533));
 sg13g2_tiehi _4414__534 (.L_HI(net534));
 sg13g2_tiehi _4413__535 (.L_HI(net535));
 sg13g2_tiehi _4412__536 (.L_HI(net536));
 sg13g2_tiehi _4411__537 (.L_HI(net537));
 sg13g2_tiehi _4410__538 (.L_HI(net538));
 sg13g2_tiehi _4409__539 (.L_HI(net539));
 sg13g2_tiehi _4408__540 (.L_HI(net540));
 sg13g2_tiehi tt_um_brukstus_tdc_with_spi_541 (.L_HI(net541));
 sg13g2_tiehi tt_um_brukstus_tdc_with_spi_542 (.L_HI(net542));
 sg13g2_tiehi tt_um_brukstus_tdc_with_spi_543 (.L_HI(net543));
 sg13g2_tiehi tt_um_brukstus_tdc_with_spi_544 (.L_HI(net544));
 sg13g2_tiehi tt_um_brukstus_tdc_with_spi_545 (.L_HI(net545));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_9 (.L_LO(net9));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_10 (.L_LO(net10));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_11 (.L_LO(net11));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_12 (.L_LO(net12));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_13 (.L_LO(net13));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_14 (.L_LO(net14));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_15 (.L_LO(net15));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_16 (.L_LO(net16));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_17 (.L_LO(net17));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_18 (.L_LO(net18));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_19 (.L_LO(net19));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_20 (.L_LO(net20));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_21 (.L_LO(net21));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_22 (.L_LO(net22));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_23 (.L_LO(net23));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_24 (.L_LO(net24));
 sg13g2_tiehi _4407__25 (.L_HI(net25));
 sg13g2_buf_2 _5563_ (.A(spi_miso),
    .X(uio_out[3]));
 sg13g2_buf_2 _5564_ (.A(\tdc_inst.busy ),
    .X(uo_out[0]));
 sg13g2_buf_4 fanout956 (.X(net956),
    .A(net957));
 sg13g2_buf_4 fanout957 (.X(net957),
    .A(net959));
 sg13g2_buf_4 fanout958 (.X(net958),
    .A(net959));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(_1379_));
 sg13g2_buf_2 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(net966),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(net963),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(net966),
    .X(net963));
 sg13g2_buf_4 fanout964 (.X(net964),
    .A(net965));
 sg13g2_buf_4 fanout965 (.X(net965),
    .A(net966));
 sg13g2_buf_2 fanout966 (.A(_1371_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_1235_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(net969),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(net977),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(net971),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(net977),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(net976),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(net976),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(net975),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(net976),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_1064_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(net979),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(net984),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(net981),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(net984),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(net984),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(net984),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_1064_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(net986),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(net990),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(net989),
    .X(net987));
 sg13g2_buf_1 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(net990),
    .X(net989));
 sg13g2_buf_1 fanout990 (.A(_1064_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(net994),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(net994),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(net994),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(net1015),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(net997),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(net997),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(net1015),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(net1002),
    .X(net998));
 sg13g2_buf_1 fanout999 (.A(net1002),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(net1002),
    .X(net1000));
 sg13g2_buf_1 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_1 fanout1002 (.A(net1003),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(net1015),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(net1006),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(net1006),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(net1015),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(net1011),
    .X(net1007));
 sg13g2_buf_1 fanout1008 (.A(net1011),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(net1011),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(net1011),
    .X(net1010));
 sg13g2_buf_1 fanout1011 (.A(net1015),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(net1013),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(net1015),
    .X(net1014));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(_0920_));
 sg13g2_buf_2 fanout1016 (.A(net1021),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(net1020),
    .X(net1017));
 sg13g2_buf_1 fanout1018 (.A(net1020),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(net1020),
    .X(net1019));
 sg13g2_buf_1 fanout1020 (.A(net1021),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(net1040),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(net1026),
    .X(net1023));
 sg13g2_buf_1 fanout1024 (.A(net1026),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(net1040),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(net1030),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(net1030),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(net1040),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(net1034),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net1033),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(net1039),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(net1039),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(net1039),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(net1038),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(net1040),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_0775_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_0760_),
    .X(net1041));
 sg13g2_buf_4 fanout1042 (.X(net1042),
    .A(_0750_));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(_1212_));
 sg13g2_buf_2 fanout1044 (.A(_1212_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(net1049),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(net1049),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(net1049),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(net1049),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(net1069),
    .X(net1049));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(net1052));
 sg13g2_buf_1 fanout1051 (.A(net1052),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(net1069),
    .X(net1052));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(net1055));
 sg13g2_buf_2 fanout1054 (.A(net1055),
    .X(net1054));
 sg13g2_buf_4 fanout1055 (.X(net1055),
    .A(net1058));
 sg13g2_buf_2 fanout1056 (.A(net1057),
    .X(net1056));
 sg13g2_buf_4 fanout1057 (.X(net1057),
    .A(net1058));
 sg13g2_buf_2 fanout1058 (.A(net1069),
    .X(net1058));
 sg13g2_buf_4 fanout1059 (.X(net1059),
    .A(net1061));
 sg13g2_buf_4 fanout1060 (.X(net1060),
    .A(net1061));
 sg13g2_buf_2 fanout1061 (.A(net1064),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(net1064),
    .X(net1062));
 sg13g2_buf_4 fanout1063 (.X(net1063),
    .A(net1064));
 sg13g2_buf_2 fanout1064 (.A(net1068),
    .X(net1064));
 sg13g2_buf_4 fanout1065 (.X(net1065),
    .A(net1068));
 sg13g2_buf_2 fanout1066 (.A(net1067),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(net1069),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(net1118),
    .X(net1069));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(net1118));
 sg13g2_buf_2 fanout1071 (.A(net1118),
    .X(net1071));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(net1075));
 sg13g2_buf_2 fanout1073 (.A(net1075),
    .X(net1073));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(net1075));
 sg13g2_buf_2 fanout1075 (.A(net1082),
    .X(net1075));
 sg13g2_buf_4 fanout1076 (.X(net1076),
    .A(net1079));
 sg13g2_buf_1 fanout1077 (.A(net1079),
    .X(net1077));
 sg13g2_buf_4 fanout1078 (.X(net1078),
    .A(net1079));
 sg13g2_buf_2 fanout1079 (.A(net1082),
    .X(net1079));
 sg13g2_buf_4 fanout1080 (.X(net1080),
    .A(net1081));
 sg13g2_buf_4 fanout1081 (.X(net1081),
    .A(net1082));
 sg13g2_buf_2 fanout1082 (.A(net1118),
    .X(net1082));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(net1084));
 sg13g2_buf_4 fanout1084 (.X(net1084),
    .A(net1094));
 sg13g2_buf_2 fanout1085 (.A(net1087),
    .X(net1085));
 sg13g2_buf_4 fanout1086 (.X(net1086),
    .A(net1087));
 sg13g2_buf_2 fanout1087 (.A(net1094),
    .X(net1087));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(net1090));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(net1090));
 sg13g2_buf_2 fanout1090 (.A(net1094),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(net1093),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(net1093),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(net1118),
    .X(net1094));
 sg13g2_buf_4 fanout1095 (.X(net1095),
    .A(net1097));
 sg13g2_buf_1 fanout1096 (.A(net1097),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(net1100),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(net1099),
    .X(net1098));
 sg13g2_buf_4 fanout1099 (.X(net1099),
    .A(net1100));
 sg13g2_buf_2 fanout1100 (.A(net1117),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(net1117),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(net1117),
    .X(net1102));
 sg13g2_buf_4 fanout1103 (.X(net1103),
    .A(net1105));
 sg13g2_buf_4 fanout1104 (.X(net1104),
    .A(net1105));
 sg13g2_buf_2 fanout1105 (.A(net1117),
    .X(net1105));
 sg13g2_buf_4 fanout1106 (.X(net1106),
    .A(net1108));
 sg13g2_buf_4 fanout1107 (.X(net1107),
    .A(net1108));
 sg13g2_buf_2 fanout1108 (.A(net1117),
    .X(net1108));
 sg13g2_buf_4 fanout1109 (.X(net1109),
    .A(net1110));
 sg13g2_buf_2 fanout1110 (.A(net1116),
    .X(net1110));
 sg13g2_buf_4 fanout1111 (.X(net1111),
    .A(net1115));
 sg13g2_buf_2 fanout1112 (.A(net1115),
    .X(net1112));
 sg13g2_buf_4 fanout1113 (.X(net1113),
    .A(net1115));
 sg13g2_buf_2 fanout1114 (.A(net1115),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(net1117),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(net1118),
    .X(net1117));
 sg13g2_buf_4 fanout1118 (.X(net1118),
    .A(_0772_));
 sg13g2_buf_2 fanout1119 (.A(_0770_),
    .X(net1119));
 sg13g2_buf_4 fanout1120 (.X(net1120),
    .A(_1253_));
 sg13g2_buf_4 fanout1121 (.X(net1121),
    .A(_1250_));
 sg13g2_buf_4 fanout1122 (.X(net1122),
    .A(_1247_));
 sg13g2_buf_4 fanout1123 (.X(net1123),
    .A(_1247_));
 sg13g2_buf_4 fanout1124 (.X(net1124),
    .A(_1243_));
 sg13g2_buf_4 fanout1125 (.X(net1125),
    .A(_1243_));
 sg13g2_buf_2 fanout1126 (.A(_1241_),
    .X(net1126));
 sg13g2_buf_4 fanout1127 (.X(net1127),
    .A(_1241_));
 sg13g2_buf_4 fanout1128 (.X(net1128),
    .A(_1239_));
 sg13g2_buf_2 fanout1129 (.A(net1130),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(net1131),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_1238_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(net1133),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_0756_),
    .X(net1133));
 sg13g2_buf_4 fanout1134 (.X(net1134),
    .A(_1236_));
 sg13g2_buf_2 fanout1135 (.A(net1139),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(net1139),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(net1139),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(net1139),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(net1157),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(net1142),
    .X(net1140));
 sg13g2_buf_1 fanout1141 (.A(net1142),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(net1157),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(net1145),
    .X(net1143));
 sg13g2_buf_1 fanout1144 (.A(net1145),
    .X(net1144));
 sg13g2_buf_2 fanout1145 (.A(net1147),
    .X(net1145));
 sg13g2_buf_2 fanout1146 (.A(net1147),
    .X(net1146));
 sg13g2_buf_2 fanout1147 (.A(net1157),
    .X(net1147));
 sg13g2_buf_2 fanout1148 (.A(net1150),
    .X(net1148));
 sg13g2_buf_2 fanout1149 (.A(net1150),
    .X(net1149));
 sg13g2_buf_2 fanout1150 (.A(net1153),
    .X(net1150));
 sg13g2_buf_2 fanout1151 (.A(net1153),
    .X(net1151));
 sg13g2_buf_2 fanout1152 (.A(net1153),
    .X(net1152));
 sg13g2_buf_2 fanout1153 (.A(net1157),
    .X(net1153));
 sg13g2_buf_2 fanout1154 (.A(net1157),
    .X(net1154));
 sg13g2_buf_2 fanout1155 (.A(net1156),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(net1207),
    .X(net1157));
 sg13g2_buf_2 fanout1158 (.A(net1159),
    .X(net1158));
 sg13g2_buf_2 fanout1159 (.A(net1207),
    .X(net1159));
 sg13g2_buf_2 fanout1160 (.A(net1207),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(net1164),
    .X(net1161));
 sg13g2_buf_1 fanout1162 (.A(net1164),
    .X(net1162));
 sg13g2_buf_2 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(net1171),
    .X(net1164));
 sg13g2_buf_2 fanout1165 (.A(net1168),
    .X(net1165));
 sg13g2_buf_1 fanout1166 (.A(net1168),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(net1168),
    .X(net1167));
 sg13g2_buf_1 fanout1168 (.A(net1171),
    .X(net1168));
 sg13g2_buf_2 fanout1169 (.A(net1170),
    .X(net1169));
 sg13g2_buf_2 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_buf_2 fanout1171 (.A(net1207),
    .X(net1171));
 sg13g2_buf_2 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_2 fanout1173 (.A(net1183),
    .X(net1173));
 sg13g2_buf_2 fanout1174 (.A(net1176),
    .X(net1174));
 sg13g2_buf_2 fanout1175 (.A(net1176),
    .X(net1175));
 sg13g2_buf_2 fanout1176 (.A(net1183),
    .X(net1176));
 sg13g2_buf_2 fanout1177 (.A(net1179),
    .X(net1177));
 sg13g2_buf_2 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_buf_2 fanout1179 (.A(net1183),
    .X(net1179));
 sg13g2_buf_2 fanout1180 (.A(net1182),
    .X(net1180));
 sg13g2_buf_2 fanout1181 (.A(net1182),
    .X(net1181));
 sg13g2_buf_2 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_2 fanout1183 (.A(net1207),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(net1186),
    .X(net1184));
 sg13g2_buf_1 fanout1185 (.A(net1186),
    .X(net1185));
 sg13g2_buf_2 fanout1186 (.A(net1189),
    .X(net1186));
 sg13g2_buf_2 fanout1187 (.A(net1188),
    .X(net1187));
 sg13g2_buf_2 fanout1188 (.A(net1189),
    .X(net1188));
 sg13g2_buf_2 fanout1189 (.A(net1206),
    .X(net1189));
 sg13g2_buf_2 fanout1190 (.A(net1206),
    .X(net1190));
 sg13g2_buf_2 fanout1191 (.A(net1206),
    .X(net1191));
 sg13g2_buf_2 fanout1192 (.A(net1194),
    .X(net1192));
 sg13g2_buf_2 fanout1193 (.A(net1194),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(net1206),
    .X(net1194));
 sg13g2_buf_2 fanout1195 (.A(net1197),
    .X(net1195));
 sg13g2_buf_2 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_buf_2 fanout1197 (.A(net1206),
    .X(net1197));
 sg13g2_buf_2 fanout1198 (.A(net1199),
    .X(net1198));
 sg13g2_buf_2 fanout1199 (.A(net1205),
    .X(net1199));
 sg13g2_buf_2 fanout1200 (.A(net1204),
    .X(net1200));
 sg13g2_buf_1 fanout1201 (.A(net1204),
    .X(net1201));
 sg13g2_buf_2 fanout1202 (.A(net1204),
    .X(net1202));
 sg13g2_buf_2 fanout1203 (.A(net1204),
    .X(net1203));
 sg13g2_buf_1 fanout1204 (.A(net1205),
    .X(net1204));
 sg13g2_buf_2 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_buf_2 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_4 fanout1207 (.X(net1207),
    .A(_0771_));
 sg13g2_buf_2 fanout1208 (.A(_0712_),
    .X(net1208));
 sg13g2_buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_2 fanout1210 (.A(\tdc_inst.stop_signal_activated ),
    .X(net1210));
 sg13g2_buf_4 fanout1211 (.X(net1211),
    .A(net1212));
 sg13g2_buf_4 fanout1212 (.X(net1212),
    .A(net1215));
 sg13g2_buf_4 fanout1213 (.X(net1213),
    .A(net1214));
 sg13g2_buf_4 fanout1214 (.X(net1214),
    .A(net1215));
 sg13g2_buf_4 fanout1215 (.X(net1215),
    .A(\tdc_inst.reset_internal_logic ));
 sg13g2_buf_4 fanout1216 (.X(net1216),
    .A(net659));
 sg13g2_buf_4 fanout1217 (.X(net1217),
    .A(net669));
 sg13g2_buf_4 fanout1218 (.X(net1218),
    .A(\spi_wrapper_i.reg_data_o[5] ));
 sg13g2_buf_4 fanout1219 (.X(net1219),
    .A(net833));
 sg13g2_buf_4 fanout1220 (.X(net1220),
    .A(net1360));
 sg13g2_buf_2 fanout1221 (.A(net1728),
    .X(net1221));
 sg13g2_buf_4 fanout1222 (.X(net1222),
    .A(net854));
 sg13g2_buf_2 fanout1223 (.A(net1718),
    .X(net1223));
 sg13g2_buf_4 fanout1224 (.X(net1224),
    .A(net1678));
 sg13g2_buf_2 fanout1225 (.A(\spi_wrapper_i.reg_addr[3] ),
    .X(net1225));
 sg13g2_buf_2 fanout1226 (.A(_0008_),
    .X(net1226));
 sg13g2_buf_2 fanout1227 (.A(net1727),
    .X(net1227));
 sg13g2_buf_4 fanout1228 (.X(net1228),
    .A(_0729_));
 sg13g2_buf_4 fanout1229 (.X(net1229),
    .A(_0729_));
 sg13g2_buf_2 fanout1230 (.A(net1234),
    .X(net1230));
 sg13g2_buf_2 fanout1231 (.A(net1234),
    .X(net1231));
 sg13g2_buf_2 fanout1232 (.A(net1233),
    .X(net1232));
 sg13g2_buf_2 fanout1233 (.A(net1234),
    .X(net1233));
 sg13g2_buf_1 fanout1234 (.A(net1235),
    .X(net1234));
 sg13g2_buf_2 fanout1235 (.A(ui_in[2]),
    .X(net1235));
 sg13g2_buf_4 fanout1236 (.X(net1236),
    .A(net1238));
 sg13g2_buf_4 fanout1237 (.X(net1237),
    .A(net1238));
 sg13g2_buf_2 fanout1238 (.A(net1258),
    .X(net1238));
 sg13g2_buf_4 fanout1239 (.X(net1239),
    .A(net1240));
 sg13g2_buf_2 fanout1240 (.A(net1241),
    .X(net1240));
 sg13g2_buf_4 fanout1241 (.X(net1241),
    .A(net1258));
 sg13g2_buf_4 fanout1242 (.X(net1242),
    .A(net1244));
 sg13g2_buf_2 fanout1243 (.A(net1244),
    .X(net1243));
 sg13g2_buf_4 fanout1244 (.X(net1244),
    .A(net1258));
 sg13g2_buf_4 fanout1245 (.X(net1245),
    .A(net1246));
 sg13g2_buf_4 fanout1246 (.X(net1246),
    .A(net1249));
 sg13g2_buf_4 fanout1247 (.X(net1247),
    .A(net1249));
 sg13g2_buf_4 fanout1248 (.X(net1248),
    .A(net1249));
 sg13g2_buf_2 fanout1249 (.A(net1258),
    .X(net1249));
 sg13g2_buf_4 fanout1250 (.X(net1250),
    .A(net1257));
 sg13g2_buf_2 fanout1251 (.A(net1257),
    .X(net1251));
 sg13g2_buf_4 fanout1252 (.X(net1252),
    .A(net1254));
 sg13g2_buf_4 fanout1253 (.X(net1253),
    .A(net1254));
 sg13g2_buf_2 fanout1254 (.A(net1257),
    .X(net1254));
 sg13g2_buf_4 fanout1255 (.X(net1255),
    .A(net1256));
 sg13g2_buf_4 fanout1256 (.X(net1256),
    .A(net1257));
 sg13g2_buf_2 fanout1257 (.A(net1258),
    .X(net1257));
 sg13g2_buf_4 fanout1258 (.X(net1258),
    .A(rst_n));
 sg13g2_buf_2 fanout1259 (.A(net1261),
    .X(net1259));
 sg13g2_buf_1 fanout1260 (.A(net1261),
    .X(net1260));
 sg13g2_buf_4 fanout1261 (.X(net1261),
    .A(ena));
 sg13g2_buf_4 fanout1262 (.X(net1262),
    .A(ena));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[6]),
    .X(net7));
 sg13g2_tielo tt_um_brukstus_tdc_with_spi_8 (.L_LO(net8));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_4_9_0_clk));
 sg13g2_buf_2 clkload7 (.A(clknet_4_10_0_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_4_13_0_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_4_14_0_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_3_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_76_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_77_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_13_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_14_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_22_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_68_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_71_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_54_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_33_clk));
 sg13g2_inv_8 clkload26 (.A(clknet_leaf_36_clk));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_43_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_39_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_41_clk));
 sg13g2_inv_2 clkload30 (.A(clknet_leaf_46_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\coarse_result[3] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold2 (.A(\coarse_result[1] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold3 (.A(\coarse_result[6] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold4 (.A(\coarse_result[5] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold5 (.A(\coarse_result[4] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold6 (.A(\coarse_result[2] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold7 (.A(\tdc_inst.stop_count_debug[35] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold8 (.A(_1099_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold9 (.A(\coarse_result[7] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold10 (.A(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0002_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold12 (.A(\coarse_result[17] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold13 (.A(\tdc_inst.stop_count_debug[113] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold14 (.A(_1177_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold15 (.A(\coarse_result[21] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold16 (.A(\coarse_result[13] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold17 (.A(\coarse_result[9] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold18 (.A(\tdc_inst.start_count_debug[82] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0857_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold20 (.A(\coarse_result[23] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold21 (.A(\coarse_result[15] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold22 (.A(\coarse_result[27] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold23 (.A(\tdc_inst.start_count_debug[120] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0895_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold25 (.A(\coarse_result[16] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold26 (.A(\coarse_result[0] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold27 (.A(\coarse_result[20] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold28 (.A(\coarse_result[31] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold29 (.A(\tdc_inst.stop_count_debug[122] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold30 (.A(_1186_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold31 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold32 (.A(_1332_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold33 (.A(\tdc_inst.start_count_debug[101] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0876_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold35 (.A(\tdc_inst.start_count_debug[4] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0779_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold37 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold38 (.A(_1302_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold39 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold40 (.A(_1347_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold41 (.A(\coarse_result[28] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold42 (.A(\config_regs[6] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0593_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold44 (.A(\coarse_result[19] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold45 (.A(spi_miso),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0520_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold47 (.A(\coarse_result[12] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold48 (.A(\coarse_result[11] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold49 (.A(\tdc_inst.start_count_debug[57] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0832_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0006_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold52 (.A(_1447_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold53 (.A(\tdc_inst.tdc_xor_result[122] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold54 (.A(_1042_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold55 (.A(\tdc_inst.start_count_debug[115] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0890_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold57 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold58 (.A(_1260_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold59 (.A(spi_mosi_sync),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0530_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold61 (.A(\config_regs[2] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0589_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold63 (.A(\config_regs[3] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0590_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold65 (.A(\config_regs[5] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0592_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold67 (.A(\tdc_inst.start_count_debug[26] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0801_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold69 (.A(\config_regs[1] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0588_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold71 (.A(\config_regs[7] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0594_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold73 (.A(\tdc_inst.stop_count_debug[72] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold74 (.A(_1136_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold75 (.A(\config_regs[4] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0591_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold77 (.A(\tdc_inst.tdc_xor_result[17] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0937_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold79 (.A(\tdc_inst.start_count_debug[9] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0784_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold81 (.A(\config_regs[0] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0587_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold83 (.A(\tdc_inst.start_count_debug[38] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0813_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold85 (.A(\tdc_inst.stop_count_debug[22] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold86 (.A(_1086_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold87 (.A(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold88 (.A(\tdc_inst.start_count_debug[118] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0893_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold90 (.A(\tdc_inst.tdc_xor_result[82] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold91 (.A(_1002_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold92 (.A(\tdc_inst.tdc_xor_result[50] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0970_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold94 (.A(\tdc_inst.start_count_debug[48] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0823_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold96 (.A(\coarse_result[8] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold97 (.A(\tdc_inst.tdc_xor_result[72] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0992_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold99 (.A(\coarse_result[25] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold100 (.A(\tdc_inst.tdc_xor_result[88] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold101 (.A(_1008_),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold102 (.A(\coarse_result[24] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold103 (.A(\tdc_inst.tdc_xor_result[108] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold104 (.A(_1028_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold105 (.A(\tdc_inst.tdc_xor_result[92] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold106 (.A(_1012_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold107 (.A(\tdc_inst.start_count_debug[75] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0850_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold109 (.A(\config_regs[13] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0584_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold111 (.A(\coarse_result[10] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold112 (.A(\tdc_inst.stop_count_debug[64] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold113 (.A(_1128_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold114 (.A(\spi_wrapper_i.reg_data_o[7] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0546_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold116 (.A(\spi_wrapper_i.spi_reg_inst.reg_rw ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0764_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0003_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold119 (.A(\tdc_inst.tdc_xor_result[78] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0998_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold121 (.A(\config_regs[63] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold122 (.A(\tdc_inst.tdc_xor_result[23] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0943_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold124 (.A(\spi_wrapper_i.reg_data_o[6] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0545_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold126 (.A(\tdc_inst.tdc_xor_result[61] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0981_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold128 (.A(\tdc_inst.tdc_xor_result[28] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0948_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold130 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0515_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold132 (.A(\config_regs[58] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0507_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold134 (.A(\config_regs[62] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold135 (.A(\tdc_inst.start_count_debug[92] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0867_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold137 (.A(\tdc_inst.stop_count_debug[74] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold138 (.A(_1138_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold139 (.A(\tdc_inst.stop_count_debug[82] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold140 (.A(_1146_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold141 (.A(\tdc_inst.tdc_xor_result[106] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold142 (.A(_1026_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold143 (.A(\tdc_inst.tdc_xor_result[52] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0972_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold145 (.A(\tdc_inst.tdc_xor_result[138] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold146 (.A(_1058_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold147 (.A(\tdc_inst.start_count_debug[27] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold148 (.A(\config_regs[30] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold149 (.A(\tdc_inst.start_count_debug[98] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0873_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold151 (.A(\config_regs[12] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0583_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold153 (.A(\tdc_inst.stop_count_debug[89] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold154 (.A(_1153_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold155 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0489_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold157 (.A(\tdc_inst.tdc_xor_result[20] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0940_),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold159 (.A(\tdc_inst.tdc_xor_result[85] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold160 (.A(_1005_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold161 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0514_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold163 (.A(\tdc_inst.stop_count_debug[46] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold164 (.A(_1110_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold165 (.A(\config_regs[41] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0548_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold167 (.A(\tdc_inst.stop_count_debug[59] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold168 (.A(_1123_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold169 (.A(\config_regs[56] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0505_),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold171 (.A(\tdc_inst.tdc_xor_result[74] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0994_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold173 (.A(\tdc_inst.stop_count_debug[66] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold174 (.A(_1130_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold175 (.A(\config_regs[18] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0573_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold177 (.A(\config_regs[42] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0549_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold179 (.A(\config_regs[25] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0556_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold181 (.A(\config_regs[28] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0559_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold183 (.A(\tdc_inst.stop_count_debug[68] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold184 (.A(_1132_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold185 (.A(\tdc_inst.positions_sum[6] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold186 (.A(\tdc_inst.stop_count_debug[62] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold187 (.A(_1126_),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold188 (.A(\tdc_inst.stop_count_debug[40] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1104_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold190 (.A(\tdc_inst.start_count_debug[81] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0856_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold192 (.A(\config_regs[51] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0566_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold194 (.A(\config_regs[43] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0550_),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold196 (.A(\tdc_inst.start_count_debug[95] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0870_),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold198 (.A(\config_regs[17] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0572_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold200 (.A(\tdc_inst.start_count_debug[31] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0806_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold202 (.A(\config_regs[46] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold203 (.A(\tdc_inst.tdc_xor_result[66] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0986_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold205 (.A(\config_regs[9] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0580_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold207 (.A(\config_regs[24] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0555_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold209 (.A(\config_regs[59] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0508_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold211 (.A(\tdc_inst.tdc_xor_result[131] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold212 (.A(_1051_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold213 (.A(\config_regs[26] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0557_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold215 (.A(\tdc_inst.start_count_debug[124] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0899_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold217 (.A(\tdc_inst.stop_count_debug[25] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1089_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold219 (.A(\tdc_inst.start_count_debug[40] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0815_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold221 (.A(\fine_result[4] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0525_),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold223 (.A(\tdc_inst.start_count_debug[63] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0838_),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold225 (.A(\coarse_result[30] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold226 (.A(\tdc_inst.start_count_debug[97] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0872_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold228 (.A(\config_regs[20] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0575_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold230 (.A(\tdc_inst.tdc_xor_result[49] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0969_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold232 (.A(\config_regs[48] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0563_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold234 (.A(\tdc_inst.stop_count_debug[127] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold235 (.A(_1191_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold236 (.A(\tdc_inst.stop_count_debug[94] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold237 (.A(_1158_),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold238 (.A(\tdc_inst.start_count_debug[58] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold239 (.A(\tdc_inst.start_count_debug[70] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0845_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold241 (.A(\tdc_inst.start_count_debug[15] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0790_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold243 (.A(\config_regs[53] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0568_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold245 (.A(\tdc_inst.start_count_debug[127] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0902_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold247 (.A(\tdc_inst.tdc_xor_result[128] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold248 (.A(_1048_),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold249 (.A(\config_regs[40] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0547_),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold251 (.A(\config_regs[10] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0581_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold253 (.A(\tdc_inst.start_count_debug[29] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0804_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold255 (.A(\tdc_inst.stop_count_debug[136] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold256 (.A(_1200_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold257 (.A(\tdc_inst.start_count_debug[69] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0844_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold259 (.A(\tdc_inst.stop_count_debug[14] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold260 (.A(_1078_),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold261 (.A(\tdc_inst.tdc_xor_result[70] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0990_),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold263 (.A(\tdc_inst.start_count_debug[11] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0786_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold265 (.A(\coarse_result[18] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold266 (.A(\tdc_inst.stop_count_debug[139] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold267 (.A(_1203_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold268 (.A(\config_regs[61] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0510_),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold270 (.A(\config_regs[44] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0551_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold272 (.A(\config_regs[31] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold273 (.A(\config_regs[55] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold274 (.A(\config_regs[21] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0576_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold276 (.A(\tdc_inst.tdc_xor_result[15] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0935_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold278 (.A(\tdc_inst.start_count_debug[62] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0837_),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold280 (.A(\config_regs[45] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0552_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold282 (.A(\tdc_inst.start_count_debug[137] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0912_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold284 (.A(\tdc_inst.tdc_xor_result[32] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0952_),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold286 (.A(\tdc_inst.stop_count_debug[63] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold287 (.A(\tdc_inst.start_count_debug[125] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold288 (.A(\spi_wrapper_i.reg_data_o[4] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0543_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold290 (.A(\tdc_inst.tdc_xor_result[90] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold291 (.A(_1010_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold292 (.A(\config_regs[22] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold293 (.A(\config_regs[47] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold294 (.A(\tdc_inst.start_count_debug[60] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0835_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold296 (.A(\tdc_inst.stop_count_debug[130] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold297 (.A(_1194_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold298 (.A(\tdc_inst.positions_sum[4] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold299 (.A(\tdc_inst.stop_count_debug[16] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold300 (.A(_1080_),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold301 (.A(\tdc_inst.tdc_xor_result[120] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold302 (.A(_1040_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold303 (.A(\tdc_inst.start_count_debug[102] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold304 (.A(\config_regs[54] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold305 (.A(\config_regs[23] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold306 (.A(\tdc_inst.stop_count_debug[56] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold307 (.A(_1120_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold308 (.A(\tdc_inst.stop_count_debug[69] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold309 (.A(\spi_wrapper_i.reg_data_o[1] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold310 (.A(\config_regs[57] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold311 (.A(\tdc_inst.start_count_debug[134] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0909_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold313 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold314 (.A(\fine_result[8] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0529_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold316 (.A(\tdc_inst.stop_count_debug[121] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold317 (.A(_1185_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold318 (.A(\config_regs[11] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0582_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold320 (.A(\config_regs[52] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold321 (.A(\tdc_inst.tdc_xor_result[27] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0947_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold323 (.A(\tdc_inst.tdc_xor_result[58] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0978_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold325 (.A(\tdc_inst.tdc_xor_result[116] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold326 (.A(_1036_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold327 (.A(\tdc_inst.tdc_xor_result[113] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold328 (.A(_1033_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold329 (.A(\tdc_inst.stop_count_debug[134] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold330 (.A(_1198_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold331 (.A(\tdc_inst.stop_count_debug[48] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold332 (.A(_1112_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold333 (.A(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold334 (.A(\config_regs[8] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0579_),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold336 (.A(\coarse_result[29] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold337 (.A(\tdc_inst.tdc_xor_result[96] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold338 (.A(_1016_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold339 (.A(\config_regs[49] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold340 (.A(\tdc_inst.tdc_xor_result[36] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0956_),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold342 (.A(\tdc_inst.start_count_debug[56] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0831_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold344 (.A(\tdc_inst.tdc_xor_result[115] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold345 (.A(_1035_),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold346 (.A(\tdc_inst.stop_count_debug[73] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold347 (.A(\config_regs[60] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold348 (.A(\tdc_inst.stop_count_debug[4] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold349 (.A(_1068_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold350 (.A(\tdc_inst.tdc_xor_result[134] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold351 (.A(_1054_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold352 (.A(\tdc_inst.start_count_debug[2] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0777_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold354 (.A(\tdc_inst.tdc_xor_result[39] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0959_),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold356 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold357 (.A(_1224_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0503_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold359 (.A(\tdc_inst.tdc_xor_result[29] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold360 (.A(\tdc_inst.start_count_debug[105] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0880_),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold362 (.A(\tdc_inst.tdc_xor_result[57] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0977_),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold364 (.A(\tdc_inst.tdc_xor_result[126] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold365 (.A(_1046_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold366 (.A(\tdc_inst.tdc_xor_result[33] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold367 (.A(\fine_result[3] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0524_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold369 (.A(\tdc_inst.stop_count_debug[128] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold370 (.A(\tdc_inst.start_count_debug[85] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0860_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold372 (.A(\tdc_inst.start_count_debug[73] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0848_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold374 (.A(\tdc_inst.start_count_debug[99] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold375 (.A(\tdc_inst.stop_count_debug[41] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold376 (.A(\spi_wrapper_i.reg_data_o_vld ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0492_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold378 (.A(\tdc_inst.stop_count_debug[32] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold379 (.A(_1096_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold380 (.A(\tdc_inst.start_count_debug[136] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0911_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold382 (.A(\tdc_inst.tdc_xor_result[119] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold383 (.A(_1039_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold384 (.A(\config_regs[16] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0571_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold386 (.A(\tdc_inst.stop_count_debug[124] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold387 (.A(_1188_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold388 (.A(\tdc_inst.tdc_xor_result[103] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold389 (.A(_1023_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold390 (.A(\coarse_result[22] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold391 (.A(\tdc_inst.positions_sum[5] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold392 (.A(\config_regs[19] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0574_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold394 (.A(\tdc_inst.start_count_debug[133] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0908_),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold396 (.A(\tdc_inst.start_count_debug[33] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0808_),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold398 (.A(\synchronizer_spi_clk_inst.data_sync[1] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold399 (.A(\tdc_inst.stop_count_debug[70] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold400 (.A(\tdc_inst.start_count_debug[17] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0792_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold402 (.A(\tdc_inst.start_count_debug[52] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0827_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold404 (.A(\tdc_inst.start_count_debug[13] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0788_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold406 (.A(\tdc_inst.start_count_debug[45] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0820_),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold408 (.A(\tdc_inst.start_count_debug[90] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0865_),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold410 (.A(\tdc_inst.stop_count_debug[13] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold411 (.A(_1077_),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold412 (.A(\tdc_inst.start_count_debug[54] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0829_),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold414 (.A(\tdc_inst.stop_count_debug[28] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold415 (.A(_1092_),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold416 (.A(\tdc_inst.tdc_xor_result[7] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0927_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold418 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0498_),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold420 (.A(\tdc_inst.tdc_xor_result[26] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0946_),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold422 (.A(\coarse_result[14] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold423 (.A(\tdc_inst.start_count_debug[141] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold424 (.A(_0916_),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold425 (.A(\tdc_inst.tdc_xor_result[93] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold426 (.A(\tdc_inst.start_count_debug[74] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold427 (.A(\tdc_inst.start_count_debug[65] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0840_),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold429 (.A(\tdc_inst.stop_count_debug[114] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold430 (.A(\tdc_inst.stop_count_debug[107] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold431 (.A(_1171_),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold432 (.A(\tdc_inst.stop_count_debug[17] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold433 (.A(\tdc_inst.tdc_xor_result[13] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0933_),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold435 (.A(\config_regs[29] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0560_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold437 (.A(\tdc_inst.stop_count_debug[30] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold438 (.A(_1094_),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold439 (.A(\tdc_inst.tdc_xor_result[84] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold440 (.A(_1004_),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold441 (.A(\tdc_inst.start_count_debug[72] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0847_),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold443 (.A(\coarse_result[26] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold444 (.A(\tdc_inst.stop_count_debug[55] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold445 (.A(_1119_),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold446 (.A(\tdc_inst.tdc_xor_result[11] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0931_),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold448 (.A(\tdc_inst.start_count_debug[14] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold449 (.A(\tdc_inst.stop_count_debug[117] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold450 (.A(_1181_),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold451 (.A(\tdc_inst.stop_count_debug[33] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold452 (.A(\tdc_inst.stop_count_debug[110] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold453 (.A(_1174_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold454 (.A(spi_clk_sync),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold455 (.A(\tdc_inst.tdc_xor_result[94] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold456 (.A(\tdc_inst.tdc_xor_result[9] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0929_),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold458 (.A(\tdc_inst.stop_count_debug[85] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold459 (.A(_1149_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold460 (.A(\tdc_inst.tdc_xor_result[46] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0966_),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold462 (.A(\tdc_inst.tdc_xor_result[4] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0924_),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold464 (.A(\tdc_inst.tdc_xor_result[53] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold465 (.A(\synchronizer_spi_mode_cpha.data_sync[1] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold466 (.A(\tdc_inst.stop_count_debug[142] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold467 (.A(\tdc_inst.tdc_xor_result[124] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold468 (.A(_1044_),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold469 (.A(\tdc_inst.start_count_debug[114] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0889_),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold471 (.A(\tdc_inst.start_count_debug[138] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold472 (.A(\tdc_inst.tdc_xor_result[55] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0975_),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold474 (.A(\tdc_inst.stop_count_debug[90] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold475 (.A(\tdc_inst.tdc_xor_result[43] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0963_),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold477 (.A(\tdc_inst.tdc_xor_result[104] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold478 (.A(\fine_result[2] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0523_),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold480 (.A(\tdc_inst.stop_count_debug[29] ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold481 (.A(\tdc_inst.stop_count_debug[5] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold482 (.A(\config_regs[27] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0558_),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold484 (.A(\tdc_inst.start_count_debug[93] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold485 (.A(\tdc_inst.tdc_xor_result[112] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold486 (.A(_1032_),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold487 (.A(\tdc_inst.tdc_xor_result[142] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold488 (.A(\tdc_inst.start_count_debug[61] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold489 (.A(\tdc_inst.stop_count_debug[19] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold490 (.A(_1083_),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold491 (.A(\tdc_inst.stop_count_debug[118] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold492 (.A(\tdc_inst.tdc_xor_result[123] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold493 (.A(\tdc_inst.start_count_debug[77] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold494 (.A(_0852_),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold495 (.A(\config_regs[50] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0565_),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold497 (.A(\tdc_inst.start_count_debug[87] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0862_),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold499 (.A(\tdc_inst.stop_count_debug[2] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold500 (.A(_1066_),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold501 (.A(\tdc_inst.tdc_xor_result[91] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold502 (.A(\tdc_inst.stop_count_debug[115] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold503 (.A(\config_regs[15] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold504 (.A(\fine_result[6] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0527_),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold506 (.A(\tdc_inst.start_count_debug[68] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold507 (.A(_0843_),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold508 (.A(\spi_wrapper_i.reg_data_o[3] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0542_),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold510 (.A(\tdc_inst.tdc_xor_result[136] ),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold511 (.A(_1056_),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold512 (.A(\tdc_inst.tdc_xor_result[1] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0921_),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold514 (.A(\tdc_inst.stop_count_debug[26] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold515 (.A(\tdc_inst.tdc_xor_result[111] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold516 (.A(_1031_),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold517 (.A(\tdc_inst.stop_count_debug[88] ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold518 (.A(_1152_),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold519 (.A(\tdc_inst.tdc_xor_result[105] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold520 (.A(\tdc_inst.stop_count_debug[131] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold521 (.A(\tdc_inst.start_count_debug[7] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0782_),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold523 (.A(\tdc_inst.start_count_debug[20] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0795_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold525 (.A(\tdc_inst.start_count_debug[142] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold526 (.A(\tdc_inst.stop_count_debug[77] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold527 (.A(_1141_),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold528 (.A(\tdc_inst.stop_count_debug[137] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold529 (.A(\tdc_inst.stop_count_debug[106] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold530 (.A(_1170_),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold531 (.A(\tdc_inst.stop_count_debug[87] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold532 (.A(_1151_),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold533 (.A(\tdc_inst.start_count_debug[109] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold534 (.A(_0884_),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold535 (.A(\tdc_inst.stop_count_debug[58] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold536 (.A(_1122_),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold537 (.A(\tdc_inst.start_count_debug[59] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold538 (.A(\tdc_inst.start_count_debug[41] ),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold539 (.A(\tdc_inst.tdc_xor_result[109] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold540 (.A(\tdc_inst.start_count_debug[126] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold541 (.A(\tdc_inst.tdc_xor_result[139] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold542 (.A(\tdc_inst.tdc_xor_result[69] ),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0989_),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold544 (.A(\tdc_inst.start_count_debug[78] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold545 (.A(\tdc_inst.start_count_debug[46] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold546 (.A(\tdc_inst.tdc_xor_result[12] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold547 (.A(\tdc_inst.start_count_debug[35] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0810_),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold549 (.A(\tdc_inst.tdc_xor_result[110] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold550 (.A(\tdc_inst.stop_count_debug[20] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold551 (.A(\tdc_inst.start_count_debug[130] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold552 (.A(_0905_),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold553 (.A(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold554 (.A(\tdc_inst.stop_count_debug[97] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold555 (.A(_1161_),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold556 (.A(\tdc_inst.start_count_debug[66] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold557 (.A(\tdc_inst.stop_count_debug[108] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold558 (.A(\tdc_inst.stop_count_debug[132] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold559 (.A(\tdc_inst.start_count_debug[42] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold560 (.A(\tdc_inst.start_count_debug[111] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0886_),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold562 (.A(\synchronizer_spi_mode_cpol.data_sync[1] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold563 (.A(\tdc_inst.tdc_xor_result[127] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold564 (.A(\tdc_inst.stop_count_debug[138] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold565 (.A(\tdc_inst.start_count_debug[112] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold566 (.A(\tdc_inst.stop_count_debug[60] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold567 (.A(\tdc_inst.start_count_debug[23] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold568 (.A(_0798_),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold569 (.A(\tdc_inst.stop_count_debug[51] ),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold570 (.A(_1115_),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold571 (.A(\tdc_inst.stop_count_debug[39] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold572 (.A(_1103_),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold573 (.A(\tdc_inst.tdc_xor_result[125] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold574 (.A(\tdc_inst.stop_count_debug[116] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold575 (.A(\tdc_inst.fine_stop_counter[0] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold576 (.A(_1532_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold577 (.A(_0657_),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold578 (.A(\tdc_inst.tdc_xor_result[47] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold579 (.A(\tdc_inst.start_count_debug[139] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold580 (.A(\tdc_inst.stop_count_debug[18] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold581 (.A(\tdc_inst.start_count_debug[129] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold582 (.A(_0904_),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold583 (.A(\tdc_inst.stop_count_debug[38] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold584 (.A(_1102_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold585 (.A(\tdc_inst.stop_count_debug[21] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold586 (.A(\tdc_inst.stop_count_debug[98] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold587 (.A(\tdc_inst.stop_count_debug[93] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold588 (.A(_1157_),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold589 (.A(\tdc_inst.stop_count_debug[100] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold590 (.A(_1164_),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold591 (.A(\tdc_inst.start_count_debug[51] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold592 (.A(_0826_),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold593 (.A(cpha_sync),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold594 (.A(\tdc_inst.stop_count_debug[91] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold595 (.A(\tdc_inst.tdc_xor_result[100] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold596 (.A(_1020_),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold597 (.A(\tdc_inst.tdc_xor_result[54] ),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold598 (.A(\tdc_inst.stop_count_debug[49] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold599 (.A(\tdc_inst.stop_count_debug[129] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold600 (.A(\tdc_inst.start_count_debug[43] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold601 (.A(\tdc_inst.start_count_debug[117] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0892_),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold603 (.A(\tdc_inst.stop_count_debug[103] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold604 (.A(_1167_),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold605 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold606 (.A(\tdc_inst.stop_count_debug[6] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold607 (.A(\tdc_inst.start_count_debug[108] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold608 (.A(_0883_),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold609 (.A(\tdc_inst.start_count_debug[91] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold610 (.A(\tdc_inst.tdc_xor_result[79] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold611 (.A(\tdc_inst.stop_count_debug[76] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold612 (.A(_1140_),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold613 (.A(\tdc_inst.stop_count_debug[109] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold614 (.A(\tdc_inst.start_count_debug[83] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold615 (.A(\tdc_inst.tdc_xor_result[81] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold616 (.A(_1001_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold617 (.A(\tdc_inst.tdc_xor_result[130] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold618 (.A(_1050_),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold619 (.A(\tdc_inst.tdc_xor_result[22] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold620 (.A(_0942_),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold621 (.A(\tdc_inst.start_count_debug[22] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold622 (.A(_0797_),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold623 (.A(\spi_wrapper_i.spi_reg_inst.state[4] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold624 (.A(\tdc_inst.start_count_debug[64] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold625 (.A(\tdc_inst.stop_count_debug[8] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold626 (.A(_1072_),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold627 (.A(\tdc_inst.start_count_debug[128] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold628 (.A(\tdc_inst.stop_count_debug[80] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold629 (.A(_1144_),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold630 (.A(\tdc_inst.tdc_xor_result[56] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold631 (.A(\config_regs[14] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold632 (.A(\tdc_inst.start_count_debug[88] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold633 (.A(\tdc_inst.tdc_xor_result[99] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold634 (.A(_1019_),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold635 (.A(spi_cs_n_sync),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold636 (.A(\tdc_inst.start_count_debug[49] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold637 (.A(\tdc_inst.stop_count_debug[24] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold638 (.A(_1088_),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold639 (.A(\tdc_inst.start_count_debug[32] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold640 (.A(\tdc_inst.tdc_xor_result[3] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold641 (.A(_0923_),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold642 (.A(\tdc_inst.tdc_xor_result[10] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold643 (.A(\tdc_inst.start_count_debug[103] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold644 (.A(\tdc_inst.start_count_debug[79] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold645 (.A(\tdc_inst.tdc_xor_result[76] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold646 (.A(_0996_),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold647 (.A(\tdc_inst.start_count_debug[104] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold648 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold649 (.A(\tdc_inst.tdc_xor_result[40] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold650 (.A(\tdc_inst.start_count_debug[34] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold651 (.A(\spi_wrapper_i.reg_data_o[5] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold652 (.A(_0544_),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold653 (.A(\tdc_inst.tdc_xor_result[38] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold654 (.A(_0958_),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold655 (.A(\tdc_inst.tdc_xor_result[77] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold656 (.A(\tdc_inst.tdc_xor_result[133] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold657 (.A(_1053_),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold658 (.A(\tdc_inst.stop_count_debug[78] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold659 (.A(\tdc_inst.tdc_xor_result[63] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold660 (.A(_0983_),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold661 (.A(\tdc_inst.start_count_debug[24] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold662 (.A(\tdc_inst.start_count_debug[135] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold663 (.A(\tdc_inst.start_count_debug[21] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold664 (.A(\tdc_inst.stop_count_debug[27] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold665 (.A(\tdc_inst.tdc_xor_result[68] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold666 (.A(_0988_),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold667 (.A(\tdc_inst.start_count_debug[107] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold668 (.A(_0882_),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold669 (.A(\tdc_inst.tdc_xor_result[97] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold670 (.A(\tdc_inst.stop_count_debug[10] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold671 (.A(_1074_),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold672 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold673 (.A(\tdc_inst.stop_count_debug[54] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold674 (.A(_1118_),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold675 (.A(\tdc_inst.stop_count_debug[102] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold676 (.A(_1166_),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold677 (.A(\tdc_inst.tdc_xor_result[25] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold678 (.A(_0945_),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold679 (.A(\tdc_inst.start_count_debug[113] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold680 (.A(\tdc_inst.stop_count_debug[95] ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold681 (.A(\tdc_inst.start_count_debug[19] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold682 (.A(_0794_),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold683 (.A(\tdc_inst.start_count_debug[28] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold684 (.A(\tdc_inst.tdc_xor_result[2] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold685 (.A(\tdc_inst.fine_start_counter[8] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold686 (.A(_0656_),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold687 (.A(\tdc_inst.stop_count_debug[120] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold688 (.A(_1184_),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold689 (.A(cpol_sync),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold690 (.A(\tdc_inst.stop_count_debug[43] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold691 (.A(_1107_),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold692 (.A(\tdc_inst.stop_count_debug[57] ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold693 (.A(\tdc_inst.stop_count_debug[104] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold694 (.A(_0036_),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold695 (.A(_1499_),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold696 (.A(_1500_),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold697 (.A(\tdc_inst.stop_count_debug[111] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold698 (.A(\tdc_inst.tdc_xor_result[102] ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold699 (.A(_1022_),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold700 (.A(\tdc_inst.tdc_xor_result[65] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold701 (.A(_0985_),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold702 (.A(\tdc_inst.stop_count_debug[99] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold703 (.A(\tdc_inst.start_count_debug[10] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold704 (.A(\tdc_inst.start_count_debug[122] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold705 (.A(_0897_),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold706 (.A(\tdc_inst.stop_count_debug[37] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold707 (.A(_1101_),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold708 (.A(\tdc_inst.stop_count_debug[125] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold709 (.A(\tdc_inst.stop_count_debug[12] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold710 (.A(_1076_),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold711 (.A(\tdc_inst.tdc_xor_result[117] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold712 (.A(\tdc_inst.stop_count_debug[11] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold713 (.A(\tdc_inst.stop_count_debug[83] ),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold714 (.A(\tdc_inst.tdc_xor_result[48] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold715 (.A(\tdc_inst.stop_count_debug[53] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold716 (.A(_1117_),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold717 (.A(\tdc_inst.tdc_xor_result[16] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold718 (.A(\tdc_inst.stop_count_debug[7] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold719 (.A(\tdc_inst.tdc_xor_result[6] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold720 (.A(_0926_),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold721 (.A(\tdc_inst.tdc_xor_result[59] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold722 (.A(\tdc_inst.stop_count_debug[105] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold723 (.A(\tdc_inst.stop_count_debug[101] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold724 (.A(\tdc_inst.stop_count_debug[52] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold725 (.A(\tdc_inst.tdc_xor_result[14] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold726 (.A(\tdc_inst.stop_count_debug[9] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold727 (.A(\tdc_inst.start_count_debug[76] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold728 (.A(\tdc_inst.stop_count_debug[135] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold729 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold730 (.A(\tdc_inst.start_count_debug[3] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold731 (.A(\tdc_inst.stop_count_debug[126] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold732 (.A(\tdc_inst.start_count_debug[25] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold733 (.A(\tdc_inst.tdc_xor_result[98] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold734 (.A(\tdc_inst.tdc_xor_result[67] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold735 (.A(\tdc_inst.start_count_debug[8] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold736 (.A(\tdc_inst.tdc_xor_result[80] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold737 (.A(\tdc_inst.tdc_xor_result[107] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold738 (.A(\tdc_inst.stop_count_debug[50] ),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold739 (.A(\tdc_inst.tdc_xor_result[19] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold740 (.A(_0939_),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold741 (.A(\tdc_inst.tdc_xor_result[129] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold742 (.A(\tdc_inst.tdc_xor_result[41] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold743 (.A(\tdc_inst.tdc_xor_result[135] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold744 (.A(\tdc_inst.stop_count_debug[140] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold745 (.A(\tdc_inst.start_count_debug[36] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold746 (.A(\tdc_inst.tdc_xor_result[8] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold747 (.A(\tdc_inst.tdc_xor_result[87] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold748 (.A(_1007_),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold749 (.A(\tdc_inst.stop_count_debug[67] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold750 (.A(\tdc_inst.stop_count_debug[65] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold751 (.A(\tdc_inst.tdc_xor_result[101] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold752 (.A(\tdc_inst.start_count_debug[50] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold753 (.A(\tdc_inst.start_count_debug[18] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold754 (.A(\tdc_inst.stop_count_debug[79] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold755 (.A(\tdc_inst.stop_count_debug[47] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold756 (.A(\tdc_inst.tdc_xor_result[24] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold757 (.A(\tdc_inst.tdc_xor_result[30] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold758 (.A(\tdc_inst.tdc_xor_result[60] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold759 (.A(\tdc_inst.stop_count_debug[31] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold760 (.A(\tdc_inst.stop_count_debug[141] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold761 (.A(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold762 (.A(\tdc_inst.stop_count_debug[123] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold763 (.A(\tdc_inst.stop_count_debug[1] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold764 (.A(_1065_),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold765 (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold766 (.A(\tdc_inst.tdc_xor_result[35] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold767 (.A(_0955_),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold768 (.A(\tdc_inst.stop_count_debug[75] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold769 (.A(\tdc_inst.stop_count_debug[45] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold770 (.A(_1109_),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold771 (.A(\tdc_inst.start_count_debug[94] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold772 (.A(\tdc_inst.positions_sum[8] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold773 (.A(_0672_),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold774 (.A(\tdc_inst.tdc_xor_result[137] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold775 (.A(\spi_wrapper_i.spi_reg_inst.state[2] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold776 (.A(\tdc_inst.tdc_xor_result[5] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold777 (.A(\config_regs[32] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold778 (.A(_0539_),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold779 (.A(\tdc_inst.start_count_debug[6] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold780 (.A(_0781_),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold781 (.A(\tdc_inst.tdc_xor_result[34] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold782 (.A(\tdc_inst.fine_start_counter[0] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold783 (.A(_1514_),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold784 (.A(_0648_),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold785 (.A(\tdc_inst.tdc_xor_result[37] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold786 (.A(\tdc_inst.stop_count_debug[84] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold787 (.A(\tdc_inst.stop_count_debug[133] ),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold788 (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold789 (.A(\tdc_inst.stop_count_debug[42] ),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold790 (.A(\tdc_inst.start_count_debug[47] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold791 (.A(\tdc_inst.start_count_debug[140] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold792 (.A(\tdc_inst.tdc_xor_result[31] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold793 (.A(\tdc_inst.tdc_xor_result[132] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold794 (.A(\tdc_inst.tdc_xor_result[44] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold795 (.A(\tdc_inst.start_count_debug[131] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold796 (.A(\tdc_inst.start_count_debug[89] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold797 (.A(\tdc_inst.tdc_xor_result[121] ),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold798 (.A(\fine_result[1] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold799 (.A(_0522_),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold800 (.A(\tdc_inst.tdc_xor_result[141] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold801 (.A(_1061_),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold802 (.A(\tdc_inst.stop_count_debug[3] ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold803 (.A(\tdc_inst.tdc_xor_result[51] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold804 (.A(\tdc_inst.tdc_xor_result[83] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold805 (.A(\tdc_inst.positions_sum[7] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold806 (.A(\tdc_inst.stop_count_debug[61] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold807 (.A(\tdc_inst.tdc_xor_result[64] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold808 (.A(\config_regs[33] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold809 (.A(\tdc_inst.stop_count_debug[36] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold810 (.A(\tdc_inst.tdc_xor_result[95] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold811 (.A(\tdc_inst.stop_count_debug[71] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold812 (.A(\config_regs[34] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold813 (.A(_0541_),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold814 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold815 (.A(\tdc_inst.tdc_xor_result[86] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold816 (.A(\tdc_inst.tdc_xor_result[42] ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold817 (.A(\tdc_inst.stop_count_debug[81] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold818 (.A(\tdc_inst.start_count_debug[30] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold819 (.A(\tdc_inst.start_count_debug[123] ),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold820 (.A(\tdc_inst.tdc_xor_result[73] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold821 (.A(\fine_result[7] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold822 (.A(_0528_),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold823 (.A(\tdc_inst.tdc_xor_result[89] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold824 (.A(\tdc_inst.tdc_xor_result[114] ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold825 (.A(\tdc_inst.start_count_debug[53] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold826 (.A(\spi_wrapper_i.reg_addr[3] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold827 (.A(\tdc_inst.start_count_debug[71] ),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold828 (.A(\tdc_inst.tdc_xor_result[18] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold829 (.A(\tdc_inst.start_count_debug[44] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold830 (.A(\tdc_inst.start_count_debug[132] ),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold831 (.A(\tdc_inst.tdc_xor_result[118] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold832 (.A(\tdc_inst.stop_count_debug[44] ),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold833 (.A(\tdc_inst.start_count_debug[106] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold834 (.A(\fine_result[0] ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold835 (.A(_0521_),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold836 (.A(\tdc_inst.fine_stop_counter[3] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold837 (.A(_1538_),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold838 (.A(\tdc_inst.start_count_debug[80] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold839 (.A(\tdc_inst.start_count_debug[100] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold840 (.A(\tdc_inst.stop_count_debug[34] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold841 (.A(\tdc_inst.start_count_debug[16] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold842 (.A(\tdc_inst.stop_count_debug[119] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold843 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold844 (.A(_0502_),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold845 (.A(\tdc_inst.tdc_xor_result[75] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold846 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold847 (.A(_0742_),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold848 (.A(\tdc_inst.stop_count_debug[96] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold849 (.A(\tdc_inst.start_count_debug[37] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold850 (.A(\tdc_inst.tdc_xor_result[140] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold851 (.A(\tdc_inst.start_count_debug[12] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold852 (.A(\tdc_inst.start_count_debug[5] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold853 (.A(\tdc_inst.tdc_xor_result[21] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold854 (.A(\tdc_inst.fine_start_counter[3] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold855 (.A(_1520_),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold856 (.A(_0651_),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold857 (.A(\tdc_inst.fine_stop_counter[1] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold858 (.A(_1535_),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold859 (.A(_0658_),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold860 (.A(\tdc_inst.fine_stop_counter[8] ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold861 (.A(_0665_),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold862 (.A(\tdc_inst.start_count_debug[96] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold863 (.A(\tdc_inst.tdc_xor_result[71] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold864 (.A(\tdc_inst.start_count_debug[67] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold865 (.A(\tdc_inst.stop_count_debug[92] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold866 (.A(\spi_wrapper_i.reg_data_o[0] ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold867 (.A(\tdc_inst.start_count_debug[86] ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold868 (.A(\tdc_inst.stop_count_debug[86] ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold869 (.A(\tdc_inst.start_count_debug[39] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold870 (.A(\fine_result[5] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold871 (.A(_0526_),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold872 (.A(\tdc_inst.stop_count_debug[15] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold873 (.A(_0034_),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold874 (.A(_1480_),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold875 (.A(\spi_wrapper_i.reg_addr[2] ),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold876 (.A(\spi_wrapper_i.reg_data_o[2] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold877 (.A(\tdc_inst.tdc_xor_result[45] ),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold878 (.A(\tdc_inst.start_count_debug[55] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold879 (.A(\tdc_inst.tdc_xor_result[62] ),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold880 (.A(\tdc_inst.stop_count_debug[112] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold881 (.A(\tdc_inst.start_count_debug[116] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold882 (.A(\tdc_inst.start_count_debug[121] ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold883 (.A(_0020_),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold884 (.A(_0517_),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold885 (.A(\tdc_inst.fine_start_counter[6] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold886 (.A(_1526_),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold887 (.A(_0654_),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold888 (.A(\tdc_inst.start_count_debug[110] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold889 (.A(\tdc_inst.start_count_debug[1] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold890 (.A(_0776_),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold891 (.A(\tdc_inst.start_count_debug[119] ),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold892 (.A(\spi_wrapper_i.reg_addr[0] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold893 (.A(\tdc_inst.start_count_debug[84] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold894 (.A(\tdc_inst.fine_start_counter[1] ),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold895 (.A(_1517_),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold896 (.A(_0649_),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold897 (.A(\tdc_inst.fine_procedure_counter[0] ),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold898 (.A(_1431_),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold899 (.A(\tdc_inst.fine_start_counter[4] ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold900 (.A(_1523_),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold901 (.A(_0652_),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold902 (.A(\tdc_inst.stop_count_debug[23] ),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold903 (.A(_0005_),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold904 (.A(_1441_),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold905 (.A(_1442_),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold906 (.A(\tdc_inst.fine_stop_counter[6] ),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold907 (.A(_1544_),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold908 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold909 (.A(_0484_),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold910 (.A(\tdc_inst.fine_stop_counter[4] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold911 (.A(_1541_),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold912 (.A(\tdc_inst.fine_another_counter[2] ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold913 (.A(_1471_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold914 (.A(\tdc_inst.tdc_xor_result[0] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold915 (.A(_1627_),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold916 (.A(_0706_),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold917 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold918 (.A(\tdc_inst.fine_procedure_counter[3] ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold919 (.A(_1437_),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold920 (.A(\tdc_inst.fine_procedure_counter[2] ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold921 (.A(_1436_),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold922 (.A(\tdc_inst.fine_procedure_counter[6] ),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold923 (.A(_0637_),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold924 (.A(\tdc_inst.fine_another_counter[8] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold925 (.A(_0647_),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold926 (.A(\tdc_inst.fine_another_counter[1] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold927 (.A(_1463_),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold928 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold929 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold930 (.A(_1226_),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold931 (.A(_0504_),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold932 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold933 (.A(\tdc_inst.fine_stop_counter[2] ),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold934 (.A(_1537_),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold935 (.A(\tdc_inst.fine_procedure_counter[1] ),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold936 (.A(\tdc_inst.fine_start_counter[2] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold937 (.A(_1519_),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold938 (.A(\tdc_inst.fine_start_counter[5] ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold939 (.A(_1525_),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold940 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold941 (.A(\tdc_inst.fine_start_counter[7] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold942 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold943 (.A(\tdc_inst.fine_stop_counter[7] ),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold944 (.A(_1547_),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold945 (.A(_0664_),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold946 (.A(\tdc_inst.fine_stop_counter[5] ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold947 (.A(\tdc_inst.fine_procedure_counter[7] ),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold948 (.A(_1446_),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold949 (.A(\tdc_inst.fine_procedure_counter[5] ),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold950 (.A(_1444_),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold951 (.A(\tdc_inst.fine_another_counter[7] ),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold952 (.A(_1505_),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold953 (.A(\tdc_inst.fine_another_counter[5] ),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold954 (.A(_1492_),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold955 (.A(\tdc_inst.fine_another_counter[4] ),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold956 (.A(_1487_),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold957 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold958 (.A(\tdc_inst.fine_stop_counter[2] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold959 (.A(\tdc_inst.fine_stop_counter[5] ),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold960 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .X(net1812));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_830 ();
 sg13g2_decap_8 FILLER_14_837 ();
 sg13g2_decap_8 FILLER_14_844 ();
 sg13g2_decap_8 FILLER_14_851 ();
 sg13g2_decap_4 FILLER_14_858 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_4 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_473 ();
 sg13g2_decap_8 FILLER_15_480 ();
 sg13g2_decap_8 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_494 ();
 sg13g2_decap_8 FILLER_15_501 ();
 sg13g2_decap_8 FILLER_15_508 ();
 sg13g2_decap_8 FILLER_15_515 ();
 sg13g2_decap_8 FILLER_15_522 ();
 sg13g2_decap_8 FILLER_15_529 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_decap_8 FILLER_15_564 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_decap_8 FILLER_15_578 ();
 sg13g2_decap_8 FILLER_15_585 ();
 sg13g2_decap_8 FILLER_15_592 ();
 sg13g2_decap_8 FILLER_15_599 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_decap_8 FILLER_15_613 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_8 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_decap_8 FILLER_15_669 ();
 sg13g2_decap_8 FILLER_15_676 ();
 sg13g2_decap_8 FILLER_15_683 ();
 sg13g2_decap_8 FILLER_15_690 ();
 sg13g2_decap_8 FILLER_15_697 ();
 sg13g2_decap_8 FILLER_15_704 ();
 sg13g2_decap_8 FILLER_15_711 ();
 sg13g2_decap_8 FILLER_15_718 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_8 FILLER_15_732 ();
 sg13g2_decap_8 FILLER_15_739 ();
 sg13g2_decap_8 FILLER_15_746 ();
 sg13g2_decap_8 FILLER_15_753 ();
 sg13g2_decap_8 FILLER_15_760 ();
 sg13g2_decap_8 FILLER_15_767 ();
 sg13g2_decap_8 FILLER_15_774 ();
 sg13g2_decap_8 FILLER_15_781 ();
 sg13g2_decap_8 FILLER_15_788 ();
 sg13g2_decap_8 FILLER_15_795 ();
 sg13g2_fill_1 FILLER_15_802 ();
 sg13g2_decap_4 FILLER_15_807 ();
 sg13g2_fill_1 FILLER_15_811 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_fill_2 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_281 ();
 sg13g2_decap_4 FILLER_16_291 ();
 sg13g2_fill_2 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_fill_1 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_414 ();
 sg13g2_decap_8 FILLER_16_421 ();
 sg13g2_decap_8 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_16_435 ();
 sg13g2_decap_8 FILLER_16_442 ();
 sg13g2_decap_8 FILLER_16_449 ();
 sg13g2_decap_8 FILLER_16_456 ();
 sg13g2_decap_8 FILLER_16_463 ();
 sg13g2_decap_8 FILLER_16_470 ();
 sg13g2_decap_8 FILLER_16_477 ();
 sg13g2_fill_1 FILLER_16_484 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_decap_8 FILLER_16_506 ();
 sg13g2_decap_8 FILLER_16_513 ();
 sg13g2_decap_8 FILLER_16_520 ();
 sg13g2_decap_8 FILLER_16_527 ();
 sg13g2_decap_8 FILLER_16_534 ();
 sg13g2_decap_8 FILLER_16_541 ();
 sg13g2_decap_8 FILLER_16_548 ();
 sg13g2_decap_8 FILLER_16_555 ();
 sg13g2_decap_8 FILLER_16_562 ();
 sg13g2_decap_8 FILLER_16_569 ();
 sg13g2_decap_8 FILLER_16_576 ();
 sg13g2_decap_8 FILLER_16_583 ();
 sg13g2_decap_8 FILLER_16_590 ();
 sg13g2_decap_8 FILLER_16_597 ();
 sg13g2_decap_8 FILLER_16_604 ();
 sg13g2_decap_8 FILLER_16_611 ();
 sg13g2_decap_8 FILLER_16_618 ();
 sg13g2_decap_8 FILLER_16_625 ();
 sg13g2_decap_8 FILLER_16_632 ();
 sg13g2_decap_8 FILLER_16_639 ();
 sg13g2_decap_8 FILLER_16_646 ();
 sg13g2_decap_8 FILLER_16_653 ();
 sg13g2_decap_8 FILLER_16_660 ();
 sg13g2_decap_8 FILLER_16_667 ();
 sg13g2_decap_8 FILLER_16_674 ();
 sg13g2_decap_8 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_688 ();
 sg13g2_decap_8 FILLER_16_695 ();
 sg13g2_decap_8 FILLER_16_702 ();
 sg13g2_decap_8 FILLER_16_709 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_730 ();
 sg13g2_decap_8 FILLER_16_737 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_fill_2 FILLER_16_772 ();
 sg13g2_fill_1 FILLER_16_774 ();
 sg13g2_fill_2 FILLER_16_779 ();
 sg13g2_fill_1 FILLER_16_781 ();
 sg13g2_decap_4 FILLER_16_786 ();
 sg13g2_fill_1 FILLER_16_790 ();
 sg13g2_fill_2 FILLER_16_823 ();
 sg13g2_decap_8 FILLER_16_855 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_261 ();
 sg13g2_fill_2 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_285 ();
 sg13g2_fill_2 FILLER_17_295 ();
 sg13g2_fill_1 FILLER_17_297 ();
 sg13g2_fill_1 FILLER_17_313 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_decap_4 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_349 ();
 sg13g2_fill_1 FILLER_17_362 ();
 sg13g2_fill_2 FILLER_17_393 ();
 sg13g2_fill_1 FILLER_17_395 ();
 sg13g2_fill_1 FILLER_17_431 ();
 sg13g2_decap_4 FILLER_17_436 ();
 sg13g2_fill_2 FILLER_17_440 ();
 sg13g2_decap_8 FILLER_17_446 ();
 sg13g2_fill_2 FILLER_17_453 ();
 sg13g2_fill_2 FILLER_17_459 ();
 sg13g2_fill_2 FILLER_17_473 ();
 sg13g2_fill_1 FILLER_17_475 ();
 sg13g2_fill_2 FILLER_17_480 ();
 sg13g2_fill_1 FILLER_17_482 ();
 sg13g2_decap_8 FILLER_17_505 ();
 sg13g2_decap_8 FILLER_17_512 ();
 sg13g2_decap_8 FILLER_17_519 ();
 sg13g2_decap_8 FILLER_17_526 ();
 sg13g2_decap_8 FILLER_17_533 ();
 sg13g2_decap_8 FILLER_17_540 ();
 sg13g2_decap_8 FILLER_17_547 ();
 sg13g2_decap_8 FILLER_17_554 ();
 sg13g2_decap_8 FILLER_17_561 ();
 sg13g2_decap_8 FILLER_17_568 ();
 sg13g2_decap_8 FILLER_17_575 ();
 sg13g2_decap_8 FILLER_17_582 ();
 sg13g2_decap_4 FILLER_17_589 ();
 sg13g2_decap_8 FILLER_17_597 ();
 sg13g2_decap_8 FILLER_17_604 ();
 sg13g2_decap_8 FILLER_17_611 ();
 sg13g2_decap_8 FILLER_17_618 ();
 sg13g2_decap_8 FILLER_17_625 ();
 sg13g2_decap_8 FILLER_17_632 ();
 sg13g2_decap_8 FILLER_17_639 ();
 sg13g2_decap_8 FILLER_17_646 ();
 sg13g2_decap_8 FILLER_17_653 ();
 sg13g2_fill_2 FILLER_17_660 ();
 sg13g2_fill_1 FILLER_17_662 ();
 sg13g2_decap_8 FILLER_17_669 ();
 sg13g2_decap_8 FILLER_17_676 ();
 sg13g2_decap_8 FILLER_17_683 ();
 sg13g2_decap_8 FILLER_17_690 ();
 sg13g2_decap_8 FILLER_17_697 ();
 sg13g2_decap_8 FILLER_17_704 ();
 sg13g2_decap_8 FILLER_17_711 ();
 sg13g2_decap_8 FILLER_17_718 ();
 sg13g2_decap_4 FILLER_17_725 ();
 sg13g2_fill_2 FILLER_17_729 ();
 sg13g2_decap_4 FILLER_17_747 ();
 sg13g2_fill_1 FILLER_17_751 ();
 sg13g2_fill_2 FILLER_17_757 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_fill_1 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_423 ();
 sg13g2_fill_1 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_514 ();
 sg13g2_decap_8 FILLER_18_521 ();
 sg13g2_decap_8 FILLER_18_528 ();
 sg13g2_decap_8 FILLER_18_535 ();
 sg13g2_decap_8 FILLER_18_542 ();
 sg13g2_decap_8 FILLER_18_549 ();
 sg13g2_decap_4 FILLER_18_556 ();
 sg13g2_fill_1 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_565 ();
 sg13g2_fill_1 FILLER_18_572 ();
 sg13g2_fill_1 FILLER_18_577 ();
 sg13g2_fill_1 FILLER_18_582 ();
 sg13g2_fill_2 FILLER_18_587 ();
 sg13g2_decap_8 FILLER_18_603 ();
 sg13g2_decap_8 FILLER_18_610 ();
 sg13g2_decap_8 FILLER_18_617 ();
 sg13g2_fill_2 FILLER_18_624 ();
 sg13g2_fill_1 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_639 ();
 sg13g2_decap_8 FILLER_18_646 ();
 sg13g2_fill_2 FILLER_18_653 ();
 sg13g2_fill_1 FILLER_18_655 ();
 sg13g2_decap_4 FILLER_18_662 ();
 sg13g2_decap_8 FILLER_18_675 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_fill_2 FILLER_18_693 ();
 sg13g2_fill_1 FILLER_18_695 ();
 sg13g2_fill_2 FILLER_18_736 ();
 sg13g2_fill_1 FILLER_18_738 ();
 sg13g2_fill_2 FILLER_18_751 ();
 sg13g2_fill_1 FILLER_18_762 ();
 sg13g2_fill_1 FILLER_18_798 ();
 sg13g2_fill_1 FILLER_18_808 ();
 sg13g2_fill_2 FILLER_18_840 ();
 sg13g2_fill_1 FILLER_18_842 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_4 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_235 ();
 sg13g2_fill_2 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_270 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_304 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_fill_2 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_422 ();
 sg13g2_fill_2 FILLER_19_479 ();
 sg13g2_fill_2 FILLER_19_490 ();
 sg13g2_fill_1 FILLER_19_492 ();
 sg13g2_decap_8 FILLER_19_523 ();
 sg13g2_decap_8 FILLER_19_530 ();
 sg13g2_decap_8 FILLER_19_537 ();
 sg13g2_decap_4 FILLER_19_544 ();
 sg13g2_fill_1 FILLER_19_560 ();
 sg13g2_fill_2 FILLER_19_593 ();
 sg13g2_fill_1 FILLER_19_595 ();
 sg13g2_fill_2 FILLER_19_622 ();
 sg13g2_fill_1 FILLER_19_624 ();
 sg13g2_decap_4 FILLER_19_763 ();
 sg13g2_fill_2 FILLER_19_860 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_fill_2 FILLER_20_168 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_decap_8 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_215 ();
 sg13g2_fill_1 FILLER_20_217 ();
 sg13g2_fill_2 FILLER_20_222 ();
 sg13g2_decap_4 FILLER_20_228 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_fill_2 FILLER_20_341 ();
 sg13g2_fill_1 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_20_379 ();
 sg13g2_fill_1 FILLER_20_381 ();
 sg13g2_fill_2 FILLER_20_448 ();
 sg13g2_fill_1 FILLER_20_480 ();
 sg13g2_fill_1 FILLER_20_535 ();
 sg13g2_fill_1 FILLER_20_540 ();
 sg13g2_fill_1 FILLER_20_600 ();
 sg13g2_fill_2 FILLER_20_629 ();
 sg13g2_fill_1 FILLER_20_631 ();
 sg13g2_fill_2 FILLER_20_666 ();
 sg13g2_fill_1 FILLER_20_668 ();
 sg13g2_fill_2 FILLER_20_699 ();
 sg13g2_fill_1 FILLER_20_705 ();
 sg13g2_fill_2 FILLER_20_730 ();
 sg13g2_fill_2 FILLER_20_750 ();
 sg13g2_fill_1 FILLER_20_752 ();
 sg13g2_fill_2 FILLER_20_792 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_239 ();
 sg13g2_fill_1 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_291 ();
 sg13g2_fill_2 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_392 ();
 sg13g2_fill_1 FILLER_21_437 ();
 sg13g2_fill_1 FILLER_21_465 ();
 sg13g2_fill_1 FILLER_21_533 ();
 sg13g2_fill_2 FILLER_21_590 ();
 sg13g2_fill_1 FILLER_21_592 ();
 sg13g2_fill_2 FILLER_21_619 ();
 sg13g2_fill_1 FILLER_21_621 ();
 sg13g2_fill_1 FILLER_21_648 ();
 sg13g2_fill_1 FILLER_21_658 ();
 sg13g2_fill_2 FILLER_21_694 ();
 sg13g2_fill_1 FILLER_21_696 ();
 sg13g2_fill_1 FILLER_21_729 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_fill_1 FILLER_22_156 ();
 sg13g2_fill_2 FILLER_22_219 ();
 sg13g2_fill_1 FILLER_22_282 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_fill_2 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_364 ();
 sg13g2_fill_1 FILLER_22_366 ();
 sg13g2_fill_1 FILLER_22_412 ();
 sg13g2_fill_1 FILLER_22_439 ();
 sg13g2_fill_2 FILLER_22_466 ();
 sg13g2_fill_1 FILLER_22_468 ();
 sg13g2_fill_2 FILLER_22_540 ();
 sg13g2_fill_1 FILLER_22_542 ();
 sg13g2_fill_2 FILLER_22_552 ();
 sg13g2_fill_1 FILLER_22_554 ();
 sg13g2_fill_2 FILLER_22_608 ();
 sg13g2_fill_1 FILLER_22_610 ();
 sg13g2_fill_2 FILLER_22_641 ();
 sg13g2_fill_1 FILLER_22_700 ();
 sg13g2_decap_4 FILLER_22_799 ();
 sg13g2_fill_2 FILLER_22_832 ();
 sg13g2_fill_1 FILLER_22_856 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_4 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_186 ();
 sg13g2_fill_2 FILLER_23_196 ();
 sg13g2_fill_1 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_fill_1 FILLER_23_290 ();
 sg13g2_fill_2 FILLER_23_304 ();
 sg13g2_fill_1 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_435 ();
 sg13g2_fill_1 FILLER_23_437 ();
 sg13g2_fill_2 FILLER_23_447 ();
 sg13g2_fill_1 FILLER_23_449 ();
 sg13g2_fill_1 FILLER_23_455 ();
 sg13g2_fill_2 FILLER_23_497 ();
 sg13g2_fill_2 FILLER_23_534 ();
 sg13g2_fill_2 FILLER_23_577 ();
 sg13g2_fill_1 FILLER_23_641 ();
 sg13g2_fill_1 FILLER_23_648 ();
 sg13g2_fill_1 FILLER_23_677 ();
 sg13g2_fill_2 FILLER_23_704 ();
 sg13g2_fill_1 FILLER_23_706 ();
 sg13g2_fill_2 FILLER_23_733 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_4 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_fill_1 FILLER_24_298 ();
 sg13g2_fill_2 FILLER_24_375 ();
 sg13g2_fill_1 FILLER_24_377 ();
 sg13g2_fill_2 FILLER_24_417 ();
 sg13g2_fill_1 FILLER_24_419 ();
 sg13g2_fill_1 FILLER_24_451 ();
 sg13g2_fill_2 FILLER_24_467 ();
 sg13g2_fill_1 FILLER_24_469 ();
 sg13g2_fill_1 FILLER_24_535 ();
 sg13g2_fill_2 FILLER_24_545 ();
 sg13g2_fill_1 FILLER_24_559 ();
 sg13g2_fill_1 FILLER_24_610 ();
 sg13g2_fill_1 FILLER_24_680 ();
 sg13g2_fill_2 FILLER_24_751 ();
 sg13g2_fill_1 FILLER_24_753 ();
 sg13g2_fill_1 FILLER_24_767 ();
 sg13g2_fill_2 FILLER_24_785 ();
 sg13g2_fill_1 FILLER_24_787 ();
 sg13g2_fill_1 FILLER_24_823 ();
 sg13g2_fill_1 FILLER_24_830 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_140 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_173 ();
 sg13g2_fill_2 FILLER_25_208 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_fill_2 FILLER_25_350 ();
 sg13g2_fill_2 FILLER_25_402 ();
 sg13g2_fill_2 FILLER_25_441 ();
 sg13g2_fill_1 FILLER_25_443 ();
 sg13g2_fill_2 FILLER_25_483 ();
 sg13g2_fill_2 FILLER_25_523 ();
 sg13g2_fill_1 FILLER_25_525 ();
 sg13g2_fill_2 FILLER_25_561 ();
 sg13g2_fill_1 FILLER_25_563 ();
 sg13g2_fill_2 FILLER_25_590 ();
 sg13g2_fill_1 FILLER_25_592 ();
 sg13g2_fill_1 FILLER_25_632 ();
 sg13g2_fill_1 FILLER_25_650 ();
 sg13g2_fill_2 FILLER_25_660 ();
 sg13g2_fill_1 FILLER_25_689 ();
 sg13g2_fill_1 FILLER_25_751 ();
 sg13g2_fill_2 FILLER_25_804 ();
 sg13g2_fill_1 FILLER_25_806 ();
 sg13g2_fill_1 FILLER_25_820 ();
 sg13g2_fill_2 FILLER_25_833 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_fill_2 FILLER_26_204 ();
 sg13g2_fill_2 FILLER_26_225 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_232 ();
 sg13g2_fill_2 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_291 ();
 sg13g2_fill_1 FILLER_26_293 ();
 sg13g2_fill_2 FILLER_26_353 ();
 sg13g2_fill_2 FILLER_26_456 ();
 sg13g2_fill_1 FILLER_26_458 ();
 sg13g2_fill_1 FILLER_26_538 ();
 sg13g2_fill_2 FILLER_26_606 ();
 sg13g2_fill_1 FILLER_26_608 ();
 sg13g2_fill_2 FILLER_26_624 ();
 sg13g2_fill_1 FILLER_26_626 ();
 sg13g2_fill_2 FILLER_26_636 ();
 sg13g2_fill_1 FILLER_26_638 ();
 sg13g2_fill_1 FILLER_26_758 ();
 sg13g2_fill_1 FILLER_26_800 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_1 FILLER_27_157 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_fill_2 FILLER_27_364 ();
 sg13g2_fill_2 FILLER_27_375 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_27_416 ();
 sg13g2_fill_1 FILLER_27_418 ();
 sg13g2_fill_2 FILLER_27_441 ();
 sg13g2_fill_1 FILLER_27_443 ();
 sg13g2_fill_1 FILLER_27_453 ();
 sg13g2_fill_2 FILLER_27_460 ();
 sg13g2_fill_2 FILLER_27_518 ();
 sg13g2_fill_2 FILLER_27_546 ();
 sg13g2_fill_1 FILLER_27_548 ();
 sg13g2_fill_1 FILLER_27_568 ();
 sg13g2_fill_1 FILLER_27_663 ();
 sg13g2_fill_2 FILLER_27_675 ();
 sg13g2_fill_2 FILLER_27_706 ();
 sg13g2_fill_1 FILLER_27_708 ();
 sg13g2_fill_1 FILLER_27_739 ();
 sg13g2_fill_1 FILLER_27_753 ();
 sg13g2_fill_1 FILLER_27_814 ();
 sg13g2_fill_1 FILLER_27_827 ();
 sg13g2_decap_4 FILLER_27_858 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_fill_1 FILLER_28_332 ();
 sg13g2_fill_2 FILLER_28_348 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_fill_2 FILLER_28_390 ();
 sg13g2_fill_2 FILLER_28_416 ();
 sg13g2_fill_1 FILLER_28_479 ();
 sg13g2_fill_2 FILLER_28_536 ();
 sg13g2_fill_2 FILLER_28_599 ();
 sg13g2_fill_1 FILLER_28_601 ();
 sg13g2_fill_1 FILLER_28_637 ();
 sg13g2_fill_2 FILLER_28_659 ();
 sg13g2_fill_1 FILLER_28_661 ();
 sg13g2_fill_1 FILLER_28_692 ();
 sg13g2_fill_2 FILLER_28_697 ();
 sg13g2_fill_2 FILLER_28_708 ();
 sg13g2_fill_1 FILLER_28_740 ();
 sg13g2_fill_2 FILLER_28_793 ();
 sg13g2_fill_2 FILLER_28_839 ();
 sg13g2_fill_2 FILLER_28_859 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_294 ();
 sg13g2_fill_1 FILLER_29_296 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_361 ();
 sg13g2_fill_1 FILLER_29_363 ();
 sg13g2_fill_2 FILLER_29_442 ();
 sg13g2_fill_1 FILLER_29_444 ();
 sg13g2_fill_1 FILLER_29_466 ();
 sg13g2_fill_2 FILLER_29_479 ();
 sg13g2_fill_1 FILLER_29_533 ();
 sg13g2_fill_1 FILLER_29_616 ();
 sg13g2_fill_1 FILLER_29_691 ();
 sg13g2_fill_1 FILLER_29_758 ();
 sg13g2_fill_2 FILLER_29_776 ();
 sg13g2_fill_2 FILLER_29_809 ();
 sg13g2_fill_1 FILLER_29_811 ();
 sg13g2_fill_1 FILLER_29_818 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_4 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_130 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_fill_2 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_333 ();
 sg13g2_fill_2 FILLER_30_347 ();
 sg13g2_fill_1 FILLER_30_349 ();
 sg13g2_fill_1 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_fill_2 FILLER_30_383 ();
 sg13g2_fill_2 FILLER_30_415 ();
 sg13g2_fill_1 FILLER_30_417 ();
 sg13g2_fill_1 FILLER_30_433 ();
 sg13g2_fill_1 FILLER_30_491 ();
 sg13g2_fill_2 FILLER_30_544 ();
 sg13g2_fill_2 FILLER_30_570 ();
 sg13g2_fill_1 FILLER_30_572 ();
 sg13g2_fill_2 FILLER_30_736 ();
 sg13g2_fill_1 FILLER_30_743 ();
 sg13g2_fill_1 FILLER_30_795 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_4 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_130 ();
 sg13g2_fill_1 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_300 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_379 ();
 sg13g2_fill_2 FILLER_31_385 ();
 sg13g2_fill_1 FILLER_31_387 ();
 sg13g2_fill_2 FILLER_31_393 ();
 sg13g2_fill_1 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_452 ();
 sg13g2_fill_2 FILLER_31_471 ();
 sg13g2_fill_1 FILLER_31_473 ();
 sg13g2_decap_8 FILLER_31_520 ();
 sg13g2_decap_4 FILLER_31_527 ();
 sg13g2_fill_1 FILLER_31_531 ();
 sg13g2_fill_1 FILLER_31_687 ();
 sg13g2_fill_2 FILLER_31_698 ();
 sg13g2_fill_1 FILLER_31_741 ();
 sg13g2_fill_2 FILLER_31_771 ();
 sg13g2_fill_1 FILLER_31_773 ();
 sg13g2_fill_1 FILLER_31_800 ();
 sg13g2_fill_1 FILLER_31_810 ();
 sg13g2_fill_2 FILLER_31_859 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_4 FILLER_32_126 ();
 sg13g2_fill_1 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_253 ();
 sg13g2_fill_2 FILLER_32_309 ();
 sg13g2_fill_1 FILLER_32_311 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_390 ();
 sg13g2_fill_1 FILLER_32_392 ();
 sg13g2_fill_2 FILLER_32_403 ();
 sg13g2_fill_1 FILLER_32_405 ();
 sg13g2_fill_2 FILLER_32_415 ();
 sg13g2_fill_1 FILLER_32_417 ();
 sg13g2_decap_4 FILLER_32_430 ();
 sg13g2_fill_1 FILLER_32_434 ();
 sg13g2_fill_1 FILLER_32_483 ();
 sg13g2_fill_2 FILLER_32_511 ();
 sg13g2_fill_1 FILLER_32_513 ();
 sg13g2_fill_2 FILLER_32_518 ();
 sg13g2_fill_1 FILLER_32_520 ();
 sg13g2_fill_1 FILLER_32_564 ();
 sg13g2_fill_2 FILLER_32_579 ();
 sg13g2_fill_1 FILLER_32_581 ();
 sg13g2_fill_2 FILLER_32_639 ();
 sg13g2_fill_2 FILLER_32_656 ();
 sg13g2_fill_1 FILLER_32_658 ();
 sg13g2_fill_2 FILLER_32_696 ();
 sg13g2_fill_2 FILLER_32_722 ();
 sg13g2_fill_2 FILLER_32_782 ();
 sg13g2_fill_1 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_153 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_fill_2 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_432 ();
 sg13g2_fill_2 FILLER_33_465 ();
 sg13g2_fill_2 FILLER_33_501 ();
 sg13g2_fill_2 FILLER_33_529 ();
 sg13g2_fill_2 FILLER_33_555 ();
 sg13g2_fill_1 FILLER_33_589 ();
 sg13g2_fill_2 FILLER_33_599 ();
 sg13g2_fill_1 FILLER_33_601 ();
 sg13g2_fill_1 FILLER_33_621 ();
 sg13g2_fill_2 FILLER_33_695 ();
 sg13g2_fill_2 FILLER_33_823 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_fill_1 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_2 FILLER_34_264 ();
 sg13g2_fill_1 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_34_399 ();
 sg13g2_fill_1 FILLER_34_435 ();
 sg13g2_fill_1 FILLER_34_463 ();
 sg13g2_fill_1 FILLER_34_487 ();
 sg13g2_fill_2 FILLER_34_567 ();
 sg13g2_fill_2 FILLER_34_605 ();
 sg13g2_fill_2 FILLER_34_646 ();
 sg13g2_fill_1 FILLER_34_648 ();
 sg13g2_fill_2 FILLER_34_729 ();
 sg13g2_fill_1 FILLER_34_731 ();
 sg13g2_fill_2 FILLER_34_745 ();
 sg13g2_fill_1 FILLER_34_747 ();
 sg13g2_fill_2 FILLER_34_770 ();
 sg13g2_fill_2 FILLER_34_798 ();
 sg13g2_fill_1 FILLER_34_800 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_4 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_159 ();
 sg13g2_fill_2 FILLER_35_186 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_258 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_fill_2 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_fill_2 FILLER_35_387 ();
 sg13g2_fill_1 FILLER_35_424 ();
 sg13g2_fill_2 FILLER_35_503 ();
 sg13g2_fill_1 FILLER_35_555 ();
 sg13g2_fill_1 FILLER_35_562 ();
 sg13g2_fill_1 FILLER_35_576 ();
 sg13g2_fill_2 FILLER_35_629 ();
 sg13g2_fill_1 FILLER_35_724 ();
 sg13g2_fill_2 FILLER_35_782 ();
 sg13g2_fill_1 FILLER_35_784 ();
 sg13g2_fill_2 FILLER_35_837 ();
 sg13g2_fill_2 FILLER_35_860 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_173 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_370 ();
 sg13g2_fill_1 FILLER_36_372 ();
 sg13g2_fill_2 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_36_410 ();
 sg13g2_fill_2 FILLER_36_437 ();
 sg13g2_fill_1 FILLER_36_480 ();
 sg13g2_fill_2 FILLER_36_507 ();
 sg13g2_fill_1 FILLER_36_509 ();
 sg13g2_fill_1 FILLER_36_571 ();
 sg13g2_fill_2 FILLER_36_602 ();
 sg13g2_fill_1 FILLER_36_604 ();
 sg13g2_fill_1 FILLER_36_631 ();
 sg13g2_fill_1 FILLER_36_651 ();
 sg13g2_fill_1 FILLER_36_754 ();
 sg13g2_fill_2 FILLER_36_769 ();
 sg13g2_fill_1 FILLER_36_775 ();
 sg13g2_fill_2 FILLER_36_789 ();
 sg13g2_fill_2 FILLER_36_832 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_221 ();
 sg13g2_fill_2 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_233 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_fill_1 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_356 ();
 sg13g2_fill_2 FILLER_37_374 ();
 sg13g2_fill_1 FILLER_37_376 ();
 sg13g2_fill_2 FILLER_37_432 ();
 sg13g2_fill_1 FILLER_37_434 ();
 sg13g2_fill_2 FILLER_37_439 ();
 sg13g2_fill_2 FILLER_37_445 ();
 sg13g2_fill_2 FILLER_37_519 ();
 sg13g2_fill_1 FILLER_37_521 ();
 sg13g2_fill_1 FILLER_37_531 ();
 sg13g2_fill_1 FILLER_37_547 ();
 sg13g2_fill_2 FILLER_37_552 ();
 sg13g2_fill_2 FILLER_37_571 ();
 sg13g2_fill_1 FILLER_37_573 ();
 sg13g2_fill_1 FILLER_37_585 ();
 sg13g2_fill_2 FILLER_37_616 ();
 sg13g2_fill_1 FILLER_37_618 ();
 sg13g2_fill_2 FILLER_37_658 ();
 sg13g2_fill_2 FILLER_37_758 ();
 sg13g2_fill_2 FILLER_37_792 ();
 sg13g2_fill_2 FILLER_37_859 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_259 ();
 sg13g2_fill_1 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_362 ();
 sg13g2_fill_1 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_399 ();
 sg13g2_fill_1 FILLER_38_401 ();
 sg13g2_fill_2 FILLER_38_428 ();
 sg13g2_fill_1 FILLER_38_480 ();
 sg13g2_fill_2 FILLER_38_513 ();
 sg13g2_fill_2 FILLER_38_519 ();
 sg13g2_fill_1 FILLER_38_560 ();
 sg13g2_fill_1 FILLER_38_604 ();
 sg13g2_fill_2 FILLER_38_630 ();
 sg13g2_fill_1 FILLER_38_640 ();
 sg13g2_fill_1 FILLER_38_679 ();
 sg13g2_fill_2 FILLER_38_718 ();
 sg13g2_fill_1 FILLER_38_720 ();
 sg13g2_fill_2 FILLER_38_752 ();
 sg13g2_fill_1 FILLER_38_754 ();
 sg13g2_fill_2 FILLER_38_802 ();
 sg13g2_fill_1 FILLER_38_804 ();
 sg13g2_fill_2 FILLER_38_820 ();
 sg13g2_fill_1 FILLER_38_822 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_4 FILLER_39_133 ();
 sg13g2_fill_1 FILLER_39_137 ();
 sg13g2_fill_2 FILLER_39_142 ();
 sg13g2_fill_1 FILLER_39_144 ();
 sg13g2_fill_2 FILLER_39_158 ();
 sg13g2_fill_2 FILLER_39_194 ();
 sg13g2_fill_1 FILLER_39_211 ();
 sg13g2_fill_2 FILLER_39_226 ();
 sg13g2_fill_2 FILLER_39_283 ();
 sg13g2_fill_2 FILLER_39_294 ();
 sg13g2_fill_2 FILLER_39_311 ();
 sg13g2_fill_1 FILLER_39_313 ();
 sg13g2_fill_2 FILLER_39_323 ();
 sg13g2_fill_2 FILLER_39_367 ();
 sg13g2_fill_1 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_fill_2 FILLER_39_405 ();
 sg13g2_fill_1 FILLER_39_407 ();
 sg13g2_fill_2 FILLER_39_417 ();
 sg13g2_fill_1 FILLER_39_419 ();
 sg13g2_fill_2 FILLER_39_434 ();
 sg13g2_fill_1 FILLER_39_444 ();
 sg13g2_fill_2 FILLER_39_474 ();
 sg13g2_fill_1 FILLER_39_476 ();
 sg13g2_fill_2 FILLER_39_499 ();
 sg13g2_fill_1 FILLER_39_542 ();
 sg13g2_fill_1 FILLER_39_574 ();
 sg13g2_fill_1 FILLER_39_779 ();
 sg13g2_fill_2 FILLER_39_789 ();
 sg13g2_fill_1 FILLER_39_791 ();
 sg13g2_fill_1 FILLER_39_801 ();
 sg13g2_decap_8 FILLER_39_845 ();
 sg13g2_decap_8 FILLER_39_852 ();
 sg13g2_fill_2 FILLER_39_859 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_fill_2 FILLER_40_147 ();
 sg13g2_fill_1 FILLER_40_149 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_fill_2 FILLER_40_228 ();
 sg13g2_fill_1 FILLER_40_230 ();
 sg13g2_fill_1 FILLER_40_261 ();
 sg13g2_fill_2 FILLER_40_302 ();
 sg13g2_fill_1 FILLER_40_304 ();
 sg13g2_fill_2 FILLER_40_314 ();
 sg13g2_fill_1 FILLER_40_316 ();
 sg13g2_fill_1 FILLER_40_325 ();
 sg13g2_fill_1 FILLER_40_358 ();
 sg13g2_fill_1 FILLER_40_368 ();
 sg13g2_fill_2 FILLER_40_383 ();
 sg13g2_fill_1 FILLER_40_395 ();
 sg13g2_fill_2 FILLER_40_487 ();
 sg13g2_decap_4 FILLER_40_515 ();
 sg13g2_fill_2 FILLER_40_519 ();
 sg13g2_fill_2 FILLER_40_526 ();
 sg13g2_fill_2 FILLER_40_576 ();
 sg13g2_fill_1 FILLER_40_578 ();
 sg13g2_fill_2 FILLER_40_592 ();
 sg13g2_fill_1 FILLER_40_598 ();
 sg13g2_decap_8 FILLER_40_605 ();
 sg13g2_fill_2 FILLER_40_612 ();
 sg13g2_fill_1 FILLER_40_614 ();
 sg13g2_decap_4 FILLER_40_628 ();
 sg13g2_fill_2 FILLER_40_632 ();
 sg13g2_fill_2 FILLER_40_642 ();
 sg13g2_fill_1 FILLER_40_678 ();
 sg13g2_fill_2 FILLER_40_688 ();
 sg13g2_fill_2 FILLER_40_718 ();
 sg13g2_fill_1 FILLER_40_720 ();
 sg13g2_decap_4 FILLER_40_741 ();
 sg13g2_fill_2 FILLER_40_745 ();
 sg13g2_fill_1 FILLER_40_751 ();
 sg13g2_fill_2 FILLER_40_796 ();
 sg13g2_fill_1 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_845 ();
 sg13g2_decap_8 FILLER_40_852 ();
 sg13g2_fill_2 FILLER_40_859 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_fill_2 FILLER_41_208 ();
 sg13g2_fill_1 FILLER_41_240 ();
 sg13g2_fill_2 FILLER_41_279 ();
 sg13g2_fill_1 FILLER_41_409 ();
 sg13g2_fill_1 FILLER_41_419 ();
 sg13g2_fill_1 FILLER_41_441 ();
 sg13g2_decap_4 FILLER_41_446 ();
 sg13g2_decap_8 FILLER_41_508 ();
 sg13g2_fill_2 FILLER_41_567 ();
 sg13g2_fill_2 FILLER_41_573 ();
 sg13g2_fill_2 FILLER_41_579 ();
 sg13g2_fill_1 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_664 ();
 sg13g2_decap_4 FILLER_41_671 ();
 sg13g2_fill_2 FILLER_41_675 ();
 sg13g2_fill_1 FILLER_41_755 ();
 sg13g2_fill_1 FILLER_41_790 ();
 sg13g2_decap_8 FILLER_41_835 ();
 sg13g2_decap_8 FILLER_41_842 ();
 sg13g2_decap_8 FILLER_41_849 ();
 sg13g2_decap_4 FILLER_41_856 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_4 FILLER_42_161 ();
 sg13g2_fill_2 FILLER_42_165 ();
 sg13g2_fill_2 FILLER_42_187 ();
 sg13g2_fill_1 FILLER_42_204 ();
 sg13g2_fill_2 FILLER_42_223 ();
 sg13g2_fill_1 FILLER_42_225 ();
 sg13g2_fill_1 FILLER_42_235 ();
 sg13g2_fill_1 FILLER_42_251 ();
 sg13g2_fill_1 FILLER_42_278 ();
 sg13g2_fill_2 FILLER_42_337 ();
 sg13g2_fill_1 FILLER_42_339 ();
 sg13g2_decap_4 FILLER_42_491 ();
 sg13g2_fill_1 FILLER_42_495 ();
 sg13g2_fill_2 FILLER_42_537 ();
 sg13g2_fill_2 FILLER_42_544 ();
 sg13g2_fill_2 FILLER_42_590 ();
 sg13g2_fill_1 FILLER_42_620 ();
 sg13g2_fill_1 FILLER_42_637 ();
 sg13g2_fill_1 FILLER_42_644 ();
 sg13g2_decap_8 FILLER_42_671 ();
 sg13g2_decap_4 FILLER_42_678 ();
 sg13g2_fill_1 FILLER_42_682 ();
 sg13g2_decap_4 FILLER_42_701 ();
 sg13g2_fill_2 FILLER_42_709 ();
 sg13g2_fill_1 FILLER_42_711 ();
 sg13g2_fill_1 FILLER_42_720 ();
 sg13g2_fill_2 FILLER_42_742 ();
 sg13g2_fill_1 FILLER_42_744 ();
 sg13g2_decap_4 FILLER_42_762 ();
 sg13g2_fill_1 FILLER_42_766 ();
 sg13g2_fill_2 FILLER_42_775 ();
 sg13g2_fill_1 FILLER_42_777 ();
 sg13g2_decap_4 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_827 ();
 sg13g2_decap_8 FILLER_42_834 ();
 sg13g2_decap_8 FILLER_42_841 ();
 sg13g2_decap_8 FILLER_42_848 ();
 sg13g2_decap_8 FILLER_42_855 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_4 FILLER_43_161 ();
 sg13g2_fill_2 FILLER_43_165 ();
 sg13g2_fill_1 FILLER_43_209 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_fill_1 FILLER_43_309 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_fill_1 FILLER_43_366 ();
 sg13g2_fill_2 FILLER_43_390 ();
 sg13g2_fill_1 FILLER_43_418 ();
 sg13g2_decap_8 FILLER_43_436 ();
 sg13g2_fill_2 FILLER_43_443 ();
 sg13g2_fill_1 FILLER_43_453 ();
 sg13g2_fill_2 FILLER_43_472 ();
 sg13g2_fill_2 FILLER_43_505 ();
 sg13g2_fill_2 FILLER_43_520 ();
 sg13g2_fill_2 FILLER_43_582 ();
 sg13g2_fill_1 FILLER_43_584 ();
 sg13g2_fill_2 FILLER_43_600 ();
 sg13g2_fill_2 FILLER_43_634 ();
 sg13g2_fill_1 FILLER_43_735 ();
 sg13g2_fill_1 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_779 ();
 sg13g2_decap_8 FILLER_43_786 ();
 sg13g2_decap_8 FILLER_43_793 ();
 sg13g2_decap_8 FILLER_43_800 ();
 sg13g2_decap_8 FILLER_43_807 ();
 sg13g2_decap_8 FILLER_43_814 ();
 sg13g2_decap_8 FILLER_43_821 ();
 sg13g2_decap_8 FILLER_43_828 ();
 sg13g2_decap_8 FILLER_43_835 ();
 sg13g2_decap_8 FILLER_43_842 ();
 sg13g2_decap_8 FILLER_43_849 ();
 sg13g2_decap_4 FILLER_43_856 ();
 sg13g2_fill_2 FILLER_43_860 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_fill_1 FILLER_44_168 ();
 sg13g2_fill_2 FILLER_44_204 ();
 sg13g2_fill_2 FILLER_44_283 ();
 sg13g2_fill_2 FILLER_44_315 ();
 sg13g2_fill_1 FILLER_44_317 ();
 sg13g2_fill_1 FILLER_44_344 ();
 sg13g2_fill_2 FILLER_44_399 ();
 sg13g2_fill_1 FILLER_44_443 ();
 sg13g2_decap_4 FILLER_44_448 ();
 sg13g2_fill_1 FILLER_44_461 ();
 sg13g2_decap_4 FILLER_44_496 ();
 sg13g2_fill_1 FILLER_44_504 ();
 sg13g2_decap_8 FILLER_44_511 ();
 sg13g2_fill_1 FILLER_44_518 ();
 sg13g2_fill_1 FILLER_44_549 ();
 sg13g2_fill_2 FILLER_44_627 ();
 sg13g2_fill_1 FILLER_44_635 ();
 sg13g2_fill_2 FILLER_44_674 ();
 sg13g2_fill_2 FILLER_44_702 ();
 sg13g2_fill_2 FILLER_44_730 ();
 sg13g2_fill_2 FILLER_44_758 ();
 sg13g2_fill_1 FILLER_44_760 ();
 sg13g2_decap_8 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_decap_8 FILLER_44_831 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_fill_2 FILLER_44_859 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_4 FILLER_45_175 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_fill_2 FILLER_45_184 ();
 sg13g2_fill_1 FILLER_45_186 ();
 sg13g2_fill_2 FILLER_45_293 ();
 sg13g2_fill_2 FILLER_45_299 ();
 sg13g2_fill_1 FILLER_45_331 ();
 sg13g2_fill_1 FILLER_45_340 ();
 sg13g2_fill_2 FILLER_45_362 ();
 sg13g2_fill_1 FILLER_45_364 ();
 sg13g2_fill_2 FILLER_45_374 ();
 sg13g2_fill_2 FILLER_45_419 ();
 sg13g2_fill_2 FILLER_45_430 ();
 sg13g2_fill_1 FILLER_45_432 ();
 sg13g2_fill_2 FILLER_45_475 ();
 sg13g2_fill_2 FILLER_45_574 ();
 sg13g2_fill_2 FILLER_45_580 ();
 sg13g2_fill_2 FILLER_45_619 ();
 sg13g2_fill_1 FILLER_45_655 ();
 sg13g2_fill_1 FILLER_45_696 ();
 sg13g2_fill_1 FILLER_45_720 ();
 sg13g2_fill_1 FILLER_45_727 ();
 sg13g2_fill_2 FILLER_45_741 ();
 sg13g2_fill_1 FILLER_45_743 ();
 sg13g2_fill_2 FILLER_45_783 ();
 sg13g2_fill_2 FILLER_45_813 ();
 sg13g2_fill_1 FILLER_45_815 ();
 sg13g2_fill_1 FILLER_45_846 ();
 sg13g2_decap_8 FILLER_45_851 ();
 sg13g2_decap_4 FILLER_45_858 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_fill_1 FILLER_46_182 ();
 sg13g2_fill_2 FILLER_46_206 ();
 sg13g2_fill_2 FILLER_46_347 ();
 sg13g2_fill_1 FILLER_46_442 ();
 sg13g2_fill_1 FILLER_46_458 ();
 sg13g2_fill_2 FILLER_46_466 ();
 sg13g2_decap_4 FILLER_46_498 ();
 sg13g2_fill_1 FILLER_46_502 ();
 sg13g2_fill_2 FILLER_46_511 ();
 sg13g2_fill_1 FILLER_46_627 ();
 sg13g2_fill_2 FILLER_46_741 ();
 sg13g2_fill_1 FILLER_46_743 ();
 sg13g2_fill_2 FILLER_46_818 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_fill_2 FILLER_47_189 ();
 sg13g2_fill_1 FILLER_47_191 ();
 sg13g2_fill_1 FILLER_47_268 ();
 sg13g2_fill_1 FILLER_47_302 ();
 sg13g2_fill_2 FILLER_47_326 ();
 sg13g2_fill_1 FILLER_47_351 ();
 sg13g2_fill_1 FILLER_47_410 ();
 sg13g2_fill_1 FILLER_47_425 ();
 sg13g2_fill_2 FILLER_47_431 ();
 sg13g2_fill_1 FILLER_47_441 ();
 sg13g2_fill_2 FILLER_47_468 ();
 sg13g2_fill_1 FILLER_47_550 ();
 sg13g2_fill_2 FILLER_47_560 ();
 sg13g2_fill_2 FILLER_47_617 ();
 sg13g2_fill_1 FILLER_47_657 ();
 sg13g2_decap_8 FILLER_47_662 ();
 sg13g2_fill_1 FILLER_47_669 ();
 sg13g2_fill_2 FILLER_47_687 ();
 sg13g2_fill_2 FILLER_47_744 ();
 sg13g2_fill_2 FILLER_47_770 ();
 sg13g2_fill_1 FILLER_47_772 ();
 sg13g2_fill_1 FILLER_47_797 ();
 sg13g2_fill_1 FILLER_47_830 ();
 sg13g2_fill_2 FILLER_47_844 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_fill_2 FILLER_48_189 ();
 sg13g2_fill_1 FILLER_48_191 ();
 sg13g2_fill_2 FILLER_48_273 ();
 sg13g2_fill_1 FILLER_48_275 ();
 sg13g2_fill_2 FILLER_48_295 ();
 sg13g2_fill_1 FILLER_48_297 ();
 sg13g2_fill_2 FILLER_48_327 ();
 sg13g2_fill_1 FILLER_48_329 ();
 sg13g2_fill_2 FILLER_48_365 ();
 sg13g2_fill_2 FILLER_48_417 ();
 sg13g2_fill_2 FILLER_48_483 ();
 sg13g2_fill_2 FILLER_48_526 ();
 sg13g2_fill_1 FILLER_48_536 ();
 sg13g2_fill_1 FILLER_48_687 ();
 sg13g2_fill_1 FILLER_48_760 ();
 sg13g2_fill_1 FILLER_48_804 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_4 FILLER_49_182 ();
 sg13g2_fill_2 FILLER_49_186 ();
 sg13g2_fill_2 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_262 ();
 sg13g2_fill_2 FILLER_49_276 ();
 sg13g2_fill_2 FILLER_49_313 ();
 sg13g2_fill_2 FILLER_49_343 ();
 sg13g2_fill_1 FILLER_49_432 ();
 sg13g2_fill_2 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_461 ();
 sg13g2_fill_1 FILLER_49_543 ();
 sg13g2_fill_1 FILLER_49_554 ();
 sg13g2_fill_1 FILLER_49_586 ();
 sg13g2_fill_2 FILLER_49_625 ();
 sg13g2_fill_1 FILLER_49_627 ();
 sg13g2_fill_2 FILLER_49_649 ();
 sg13g2_fill_1 FILLER_49_651 ();
 sg13g2_fill_2 FILLER_49_681 ();
 sg13g2_fill_1 FILLER_49_683 ();
 sg13g2_fill_2 FILLER_49_723 ();
 sg13g2_fill_1 FILLER_49_733 ();
 sg13g2_fill_1 FILLER_49_765 ();
 sg13g2_fill_1 FILLER_49_775 ();
 sg13g2_fill_2 FILLER_49_796 ();
 sg13g2_fill_1 FILLER_49_828 ();
 sg13g2_fill_2 FILLER_49_844 ();
 sg13g2_fill_2 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_fill_1 FILLER_50_182 ();
 sg13g2_fill_1 FILLER_50_253 ();
 sg13g2_fill_2 FILLER_50_280 ();
 sg13g2_fill_2 FILLER_50_296 ();
 sg13g2_fill_2 FILLER_50_303 ();
 sg13g2_fill_1 FILLER_50_305 ();
 sg13g2_fill_1 FILLER_50_317 ();
 sg13g2_fill_2 FILLER_50_347 ();
 sg13g2_fill_2 FILLER_50_366 ();
 sg13g2_decap_4 FILLER_50_440 ();
 sg13g2_fill_1 FILLER_50_448 ();
 sg13g2_fill_2 FILLER_50_499 ();
 sg13g2_fill_1 FILLER_50_510 ();
 sg13g2_fill_2 FILLER_50_525 ();
 sg13g2_fill_1 FILLER_50_527 ();
 sg13g2_fill_1 FILLER_50_564 ();
 sg13g2_fill_2 FILLER_50_591 ();
 sg13g2_fill_2 FILLER_50_608 ();
 sg13g2_fill_1 FILLER_50_625 ();
 sg13g2_fill_2 FILLER_50_631 ();
 sg13g2_fill_2 FILLER_50_646 ();
 sg13g2_fill_1 FILLER_50_648 ();
 sg13g2_fill_1 FILLER_50_688 ();
 sg13g2_fill_2 FILLER_50_721 ();
 sg13g2_fill_1 FILLER_50_723 ();
 sg13g2_fill_2 FILLER_50_761 ();
 sg13g2_fill_1 FILLER_50_763 ();
 sg13g2_fill_2 FILLER_50_824 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_decap_8 FILLER_51_182 ();
 sg13g2_fill_2 FILLER_51_189 ();
 sg13g2_fill_1 FILLER_51_191 ();
 sg13g2_fill_2 FILLER_51_264 ();
 sg13g2_fill_1 FILLER_51_266 ();
 sg13g2_fill_2 FILLER_51_281 ();
 sg13g2_fill_2 FILLER_51_297 ();
 sg13g2_fill_1 FILLER_51_436 ();
 sg13g2_decap_4 FILLER_51_442 ();
 sg13g2_fill_1 FILLER_51_446 ();
 sg13g2_fill_1 FILLER_51_458 ();
 sg13g2_fill_2 FILLER_51_498 ();
 sg13g2_fill_1 FILLER_51_504 ();
 sg13g2_fill_2 FILLER_51_531 ();
 sg13g2_fill_1 FILLER_51_533 ();
 sg13g2_fill_2 FILLER_51_556 ();
 sg13g2_fill_2 FILLER_51_576 ();
 sg13g2_fill_2 FILLER_51_729 ();
 sg13g2_fill_1 FILLER_51_745 ();
 sg13g2_fill_2 FILLER_51_802 ();
 sg13g2_fill_1 FILLER_51_804 ();
 sg13g2_fill_1 FILLER_51_831 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_4 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_95 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_fill_2 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_129 ();
 sg13g2_decap_8 FILLER_52_136 ();
 sg13g2_decap_8 FILLER_52_143 ();
 sg13g2_decap_8 FILLER_52_150 ();
 sg13g2_decap_8 FILLER_52_186 ();
 sg13g2_decap_8 FILLER_52_193 ();
 sg13g2_fill_2 FILLER_52_281 ();
 sg13g2_fill_1 FILLER_52_327 ();
 sg13g2_fill_1 FILLER_52_398 ();
 sg13g2_decap_8 FILLER_52_429 ();
 sg13g2_fill_1 FILLER_52_436 ();
 sg13g2_fill_2 FILLER_52_523 ();
 sg13g2_fill_2 FILLER_52_616 ();
 sg13g2_fill_1 FILLER_52_618 ();
 sg13g2_fill_2 FILLER_52_625 ();
 sg13g2_fill_1 FILLER_52_636 ();
 sg13g2_fill_2 FILLER_52_696 ();
 sg13g2_fill_1 FILLER_52_722 ();
 sg13g2_fill_2 FILLER_52_775 ();
 sg13g2_fill_1 FILLER_52_777 ();
 sg13g2_fill_1 FILLER_52_796 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_78 ();
 sg13g2_decap_8 FILLER_53_85 ();
 sg13g2_fill_2 FILLER_53_92 ();
 sg13g2_fill_1 FILLER_53_94 ();
 sg13g2_fill_2 FILLER_53_121 ();
 sg13g2_decap_8 FILLER_53_152 ();
 sg13g2_fill_1 FILLER_53_159 ();
 sg13g2_fill_2 FILLER_53_163 ();
 sg13g2_fill_1 FILLER_53_165 ();
 sg13g2_fill_2 FILLER_53_207 ();
 sg13g2_fill_1 FILLER_53_209 ();
 sg13g2_fill_2 FILLER_53_233 ();
 sg13g2_fill_1 FILLER_53_235 ();
 sg13g2_fill_2 FILLER_53_298 ();
 sg13g2_fill_1 FILLER_53_324 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_fill_2 FILLER_53_379 ();
 sg13g2_fill_1 FILLER_53_388 ();
 sg13g2_fill_1 FILLER_53_399 ();
 sg13g2_decap_4 FILLER_53_427 ();
 sg13g2_fill_1 FILLER_53_431 ();
 sg13g2_fill_1 FILLER_53_514 ();
 sg13g2_fill_1 FILLER_53_553 ();
 sg13g2_fill_2 FILLER_53_577 ();
 sg13g2_fill_1 FILLER_53_579 ();
 sg13g2_fill_2 FILLER_53_590 ();
 sg13g2_fill_1 FILLER_53_592 ();
 sg13g2_fill_2 FILLER_53_703 ();
 sg13g2_fill_1 FILLER_53_787 ();
 sg13g2_fill_1 FILLER_53_792 ();
 sg13g2_fill_1 FILLER_53_832 ();
 sg13g2_fill_1 FILLER_53_846 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_4 FILLER_54_63 ();
 sg13g2_decap_4 FILLER_54_96 ();
 sg13g2_fill_1 FILLER_54_100 ();
 sg13g2_decap_8 FILLER_54_106 ();
 sg13g2_fill_1 FILLER_54_113 ();
 sg13g2_decap_4 FILLER_54_157 ();
 sg13g2_fill_1 FILLER_54_161 ();
 sg13g2_decap_4 FILLER_54_168 ();
 sg13g2_fill_2 FILLER_54_239 ();
 sg13g2_fill_2 FILLER_54_267 ();
 sg13g2_fill_1 FILLER_54_269 ();
 sg13g2_fill_2 FILLER_54_300 ();
 sg13g2_fill_2 FILLER_54_340 ();
 sg13g2_fill_2 FILLER_54_451 ();
 sg13g2_fill_2 FILLER_54_612 ();
 sg13g2_fill_1 FILLER_54_614 ();
 sg13g2_fill_1 FILLER_54_708 ();
 sg13g2_fill_1 FILLER_54_714 ();
 sg13g2_fill_2 FILLER_54_728 ();
 sg13g2_fill_1 FILLER_54_730 ();
 sg13g2_fill_2 FILLER_54_749 ();
 sg13g2_fill_1 FILLER_54_751 ();
 sg13g2_fill_1 FILLER_54_776 ();
 sg13g2_fill_1 FILLER_54_826 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_fill_1 FILLER_55_70 ();
 sg13g2_fill_1 FILLER_55_79 ();
 sg13g2_fill_2 FILLER_55_114 ();
 sg13g2_fill_1 FILLER_55_116 ();
 sg13g2_decap_8 FILLER_55_139 ();
 sg13g2_decap_8 FILLER_55_146 ();
 sg13g2_decap_4 FILLER_55_153 ();
 sg13g2_fill_2 FILLER_55_157 ();
 sg13g2_decap_4 FILLER_55_171 ();
 sg13g2_fill_1 FILLER_55_211 ();
 sg13g2_fill_1 FILLER_55_239 ();
 sg13g2_fill_2 FILLER_55_259 ();
 sg13g2_fill_2 FILLER_55_270 ();
 sg13g2_fill_1 FILLER_55_449 ();
 sg13g2_fill_1 FILLER_55_538 ();
 sg13g2_fill_2 FILLER_55_597 ();
 sg13g2_fill_1 FILLER_55_599 ();
 sg13g2_fill_2 FILLER_55_645 ();
 sg13g2_fill_2 FILLER_55_673 ();
 sg13g2_fill_1 FILLER_55_675 ();
 sg13g2_fill_1 FILLER_55_702 ();
 sg13g2_fill_2 FILLER_55_729 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_fill_2 FILLER_55_766 ();
 sg13g2_fill_1 FILLER_55_768 ();
 sg13g2_fill_2 FILLER_55_816 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_4 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_60 ();
 sg13g2_decap_8 FILLER_56_95 ();
 sg13g2_decap_8 FILLER_56_102 ();
 sg13g2_decap_8 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_116 ();
 sg13g2_fill_1 FILLER_56_118 ();
 sg13g2_fill_1 FILLER_56_168 ();
 sg13g2_fill_2 FILLER_56_174 ();
 sg13g2_fill_1 FILLER_56_176 ();
 sg13g2_fill_1 FILLER_56_186 ();
 sg13g2_fill_1 FILLER_56_213 ();
 sg13g2_fill_1 FILLER_56_307 ();
 sg13g2_fill_2 FILLER_56_317 ();
 sg13g2_fill_2 FILLER_56_360 ();
 sg13g2_fill_2 FILLER_56_469 ();
 sg13g2_decap_4 FILLER_56_481 ();
 sg13g2_decap_4 FILLER_56_530 ();
 sg13g2_fill_2 FILLER_56_578 ();
 sg13g2_fill_1 FILLER_56_624 ();
 sg13g2_fill_2 FILLER_56_655 ();
 sg13g2_fill_1 FILLER_56_657 ();
 sg13g2_fill_2 FILLER_56_778 ();
 sg13g2_fill_1 FILLER_56_784 ();
 sg13g2_fill_1 FILLER_56_794 ();
 sg13g2_fill_2 FILLER_56_833 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_fill_2 FILLER_57_56 ();
 sg13g2_fill_1 FILLER_57_58 ();
 sg13g2_fill_1 FILLER_57_85 ();
 sg13g2_fill_2 FILLER_57_96 ();
 sg13g2_decap_8 FILLER_57_113 ();
 sg13g2_fill_2 FILLER_57_120 ();
 sg13g2_decap_4 FILLER_57_128 ();
 sg13g2_decap_8 FILLER_57_169 ();
 sg13g2_fill_2 FILLER_57_176 ();
 sg13g2_fill_1 FILLER_57_197 ();
 sg13g2_fill_1 FILLER_57_216 ();
 sg13g2_fill_1 FILLER_57_229 ();
 sg13g2_fill_2 FILLER_57_234 ();
 sg13g2_fill_2 FILLER_57_255 ();
 sg13g2_fill_1 FILLER_57_257 ();
 sg13g2_fill_2 FILLER_57_266 ();
 sg13g2_fill_2 FILLER_57_316 ();
 sg13g2_fill_1 FILLER_57_318 ();
 sg13g2_fill_2 FILLER_57_344 ();
 sg13g2_decap_4 FILLER_57_414 ();
 sg13g2_fill_1 FILLER_57_510 ();
 sg13g2_fill_2 FILLER_57_557 ();
 sg13g2_fill_1 FILLER_57_649 ();
 sg13g2_fill_2 FILLER_57_690 ();
 sg13g2_fill_1 FILLER_57_697 ();
 sg13g2_fill_1 FILLER_57_724 ();
 sg13g2_fill_2 FILLER_57_731 ();
 sg13g2_fill_2 FILLER_57_795 ();
 sg13g2_fill_2 FILLER_57_859 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_fill_1 FILLER_58_70 ();
 sg13g2_fill_2 FILLER_58_141 ();
 sg13g2_decap_4 FILLER_58_218 ();
 sg13g2_fill_1 FILLER_58_227 ();
 sg13g2_fill_1 FILLER_58_262 ();
 sg13g2_fill_2 FILLER_58_272 ();
 sg13g2_fill_2 FILLER_58_400 ();
 sg13g2_decap_4 FILLER_58_449 ();
 sg13g2_fill_2 FILLER_58_463 ();
 sg13g2_fill_1 FILLER_58_465 ();
 sg13g2_fill_1 FILLER_58_538 ();
 sg13g2_fill_1 FILLER_58_558 ();
 sg13g2_fill_2 FILLER_58_666 ();
 sg13g2_fill_2 FILLER_58_683 ();
 sg13g2_fill_2 FILLER_58_715 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_4 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_81 ();
 sg13g2_decap_4 FILLER_59_91 ();
 sg13g2_fill_2 FILLER_59_95 ();
 sg13g2_decap_8 FILLER_59_116 ();
 sg13g2_fill_1 FILLER_59_123 ();
 sg13g2_decap_4 FILLER_59_129 ();
 sg13g2_fill_2 FILLER_59_133 ();
 sg13g2_decap_4 FILLER_59_152 ();
 sg13g2_fill_1 FILLER_59_156 ();
 sg13g2_fill_2 FILLER_59_162 ();
 sg13g2_decap_8 FILLER_59_167 ();
 sg13g2_fill_1 FILLER_59_178 ();
 sg13g2_fill_1 FILLER_59_188 ();
 sg13g2_fill_1 FILLER_59_221 ();
 sg13g2_fill_1 FILLER_59_252 ();
 sg13g2_fill_1 FILLER_59_257 ();
 sg13g2_fill_1 FILLER_59_265 ();
 sg13g2_fill_2 FILLER_59_281 ();
 sg13g2_fill_1 FILLER_59_283 ();
 sg13g2_fill_2 FILLER_59_290 ();
 sg13g2_fill_1 FILLER_59_292 ();
 sg13g2_fill_2 FILLER_59_302 ();
 sg13g2_fill_1 FILLER_59_304 ();
 sg13g2_fill_2 FILLER_59_317 ();
 sg13g2_fill_1 FILLER_59_336 ();
 sg13g2_fill_1 FILLER_59_351 ();
 sg13g2_fill_2 FILLER_59_519 ();
 sg13g2_fill_2 FILLER_59_567 ();
 sg13g2_fill_2 FILLER_59_636 ();
 sg13g2_fill_2 FILLER_59_767 ();
 sg13g2_fill_2 FILLER_59_859 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_fill_1 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_113 ();
 sg13g2_fill_2 FILLER_60_120 ();
 sg13g2_decap_8 FILLER_60_130 ();
 sg13g2_decap_8 FILLER_60_137 ();
 sg13g2_decap_4 FILLER_60_144 ();
 sg13g2_fill_2 FILLER_60_153 ();
 sg13g2_decap_4 FILLER_60_186 ();
 sg13g2_decap_4 FILLER_60_195 ();
 sg13g2_fill_1 FILLER_60_199 ();
 sg13g2_fill_2 FILLER_60_219 ();
 sg13g2_fill_1 FILLER_60_221 ();
 sg13g2_fill_2 FILLER_60_227 ();
 sg13g2_fill_2 FILLER_60_353 ();
 sg13g2_fill_1 FILLER_60_384 ();
 sg13g2_fill_1 FILLER_60_454 ();
 sg13g2_fill_2 FILLER_60_464 ();
 sg13g2_fill_1 FILLER_60_528 ();
 sg13g2_fill_1 FILLER_60_537 ();
 sg13g2_fill_1 FILLER_60_552 ();
 sg13g2_decap_4 FILLER_60_562 ();
 sg13g2_fill_2 FILLER_60_594 ();
 sg13g2_fill_1 FILLER_60_596 ();
 sg13g2_fill_1 FILLER_60_611 ();
 sg13g2_fill_1 FILLER_60_656 ();
 sg13g2_fill_1 FILLER_60_697 ();
 sg13g2_fill_2 FILLER_60_715 ();
 sg13g2_fill_1 FILLER_60_740 ();
 sg13g2_fill_1 FILLER_60_750 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_fill_1 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_98 ();
 sg13g2_decap_4 FILLER_61_155 ();
 sg13g2_fill_2 FILLER_61_168 ();
 sg13g2_decap_4 FILLER_61_218 ();
 sg13g2_decap_4 FILLER_61_254 ();
 sg13g2_fill_1 FILLER_61_265 ();
 sg13g2_fill_2 FILLER_61_313 ();
 sg13g2_fill_1 FILLER_61_342 ();
 sg13g2_fill_1 FILLER_61_353 ();
 sg13g2_fill_1 FILLER_61_380 ();
 sg13g2_fill_2 FILLER_61_459 ();
 sg13g2_fill_1 FILLER_61_461 ();
 sg13g2_fill_2 FILLER_61_570 ();
 sg13g2_fill_2 FILLER_61_680 ();
 sg13g2_fill_1 FILLER_61_682 ();
 sg13g2_fill_2 FILLER_61_692 ();
 sg13g2_fill_2 FILLER_61_772 ();
 sg13g2_fill_1 FILLER_61_819 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_fill_2 FILLER_62_99 ();
 sg13g2_decap_8 FILLER_62_127 ();
 sg13g2_decap_8 FILLER_62_134 ();
 sg13g2_decap_4 FILLER_62_141 ();
 sg13g2_fill_2 FILLER_62_156 ();
 sg13g2_fill_1 FILLER_62_158 ();
 sg13g2_fill_1 FILLER_62_165 ();
 sg13g2_fill_2 FILLER_62_191 ();
 sg13g2_fill_1 FILLER_62_193 ();
 sg13g2_fill_1 FILLER_62_207 ();
 sg13g2_decap_8 FILLER_62_220 ();
 sg13g2_fill_2 FILLER_62_227 ();
 sg13g2_fill_1 FILLER_62_229 ();
 sg13g2_fill_1 FILLER_62_239 ();
 sg13g2_fill_2 FILLER_62_295 ();
 sg13g2_fill_1 FILLER_62_390 ();
 sg13g2_fill_2 FILLER_62_421 ();
 sg13g2_fill_2 FILLER_62_438 ();
 sg13g2_fill_1 FILLER_62_446 ();
 sg13g2_fill_2 FILLER_62_456 ();
 sg13g2_fill_2 FILLER_62_494 ();
 sg13g2_fill_2 FILLER_62_585 ();
 sg13g2_fill_1 FILLER_62_587 ();
 sg13g2_fill_2 FILLER_62_598 ();
 sg13g2_fill_1 FILLER_62_696 ();
 sg13g2_fill_1 FILLER_62_712 ();
 sg13g2_fill_2 FILLER_62_728 ();
 sg13g2_fill_2 FILLER_62_747 ();
 sg13g2_fill_1 FILLER_62_749 ();
 sg13g2_fill_2 FILLER_62_764 ();
 sg13g2_fill_2 FILLER_62_818 ();
 sg13g2_fill_1 FILLER_62_825 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_4 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_67 ();
 sg13g2_decap_4 FILLER_63_95 ();
 sg13g2_fill_2 FILLER_63_121 ();
 sg13g2_fill_1 FILLER_63_149 ();
 sg13g2_fill_2 FILLER_63_216 ();
 sg13g2_fill_1 FILLER_63_218 ();
 sg13g2_decap_4 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_239 ();
 sg13g2_fill_2 FILLER_63_243 ();
 sg13g2_fill_1 FILLER_63_256 ();
 sg13g2_fill_2 FILLER_63_263 ();
 sg13g2_fill_2 FILLER_63_288 ();
 sg13g2_fill_1 FILLER_63_290 ();
 sg13g2_fill_1 FILLER_63_306 ();
 sg13g2_fill_1 FILLER_63_335 ();
 sg13g2_fill_2 FILLER_63_341 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_fill_2 FILLER_63_393 ();
 sg13g2_fill_1 FILLER_63_395 ();
 sg13g2_fill_1 FILLER_63_434 ();
 sg13g2_fill_2 FILLER_63_448 ();
 sg13g2_fill_1 FILLER_63_450 ();
 sg13g2_fill_2 FILLER_63_495 ();
 sg13g2_fill_2 FILLER_63_533 ();
 sg13g2_fill_2 FILLER_63_558 ();
 sg13g2_fill_2 FILLER_63_587 ();
 sg13g2_fill_1 FILLER_63_609 ();
 sg13g2_fill_2 FILLER_63_627 ();
 sg13g2_fill_2 FILLER_63_796 ();
 sg13g2_fill_1 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_4 FILLER_64_56 ();
 sg13g2_fill_2 FILLER_64_94 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_2 FILLER_64_122 ();
 sg13g2_fill_1 FILLER_64_124 ();
 sg13g2_decap_4 FILLER_64_151 ();
 sg13g2_decap_8 FILLER_64_164 ();
 sg13g2_fill_1 FILLER_64_171 ();
 sg13g2_fill_1 FILLER_64_175 ();
 sg13g2_fill_2 FILLER_64_258 ();
 sg13g2_decap_8 FILLER_64_295 ();
 sg13g2_decap_4 FILLER_64_302 ();
 sg13g2_fill_1 FILLER_64_306 ();
 sg13g2_fill_2 FILLER_64_319 ();
 sg13g2_fill_1 FILLER_64_321 ();
 sg13g2_fill_2 FILLER_64_382 ();
 sg13g2_fill_1 FILLER_64_384 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_fill_1 FILLER_64_454 ();
 sg13g2_fill_2 FILLER_64_527 ();
 sg13g2_fill_1 FILLER_64_529 ();
 sg13g2_decap_8 FILLER_64_630 ();
 sg13g2_decap_4 FILLER_64_637 ();
 sg13g2_fill_2 FILLER_64_641 ();
 sg13g2_fill_2 FILLER_64_655 ();
 sg13g2_fill_2 FILLER_64_693 ();
 sg13g2_fill_1 FILLER_64_695 ();
 sg13g2_fill_2 FILLER_64_702 ();
 sg13g2_fill_1 FILLER_64_704 ();
 sg13g2_fill_2 FILLER_64_741 ();
 sg13g2_fill_1 FILLER_64_743 ();
 sg13g2_fill_1 FILLER_64_817 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_fill_2 FILLER_65_56 ();
 sg13g2_fill_1 FILLER_65_58 ();
 sg13g2_decap_4 FILLER_65_100 ();
 sg13g2_decap_8 FILLER_65_135 ();
 sg13g2_decap_4 FILLER_65_142 ();
 sg13g2_fill_2 FILLER_65_163 ();
 sg13g2_fill_1 FILLER_65_165 ();
 sg13g2_fill_2 FILLER_65_198 ();
 sg13g2_fill_2 FILLER_65_206 ();
 sg13g2_fill_2 FILLER_65_227 ();
 sg13g2_fill_2 FILLER_65_238 ();
 sg13g2_fill_2 FILLER_65_256 ();
 sg13g2_fill_1 FILLER_65_299 ();
 sg13g2_fill_2 FILLER_65_344 ();
 sg13g2_fill_2 FILLER_65_372 ();
 sg13g2_fill_2 FILLER_65_379 ();
 sg13g2_fill_2 FILLER_65_391 ();
 sg13g2_fill_1 FILLER_65_406 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_fill_1 FILLER_65_450 ();
 sg13g2_fill_1 FILLER_65_565 ();
 sg13g2_fill_2 FILLER_65_580 ();
 sg13g2_fill_2 FILLER_65_588 ();
 sg13g2_fill_2 FILLER_65_604 ();
 sg13g2_fill_1 FILLER_65_606 ();
 sg13g2_fill_1 FILLER_65_722 ();
 sg13g2_fill_1 FILLER_65_738 ();
 sg13g2_fill_1 FILLER_65_744 ();
 sg13g2_fill_2 FILLER_65_793 ();
 sg13g2_fill_1 FILLER_65_811 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_97 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_decap_4 FILLER_66_119 ();
 sg13g2_fill_2 FILLER_66_123 ();
 sg13g2_decap_4 FILLER_66_151 ();
 sg13g2_fill_1 FILLER_66_155 ();
 sg13g2_decap_8 FILLER_66_164 ();
 sg13g2_fill_2 FILLER_66_171 ();
 sg13g2_fill_1 FILLER_66_173 ();
 sg13g2_fill_2 FILLER_66_279 ();
 sg13g2_fill_2 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_417 ();
 sg13g2_fill_2 FILLER_66_424 ();
 sg13g2_fill_2 FILLER_66_528 ();
 sg13g2_fill_1 FILLER_66_530 ();
 sg13g2_fill_2 FILLER_66_580 ();
 sg13g2_fill_1 FILLER_66_582 ();
 sg13g2_fill_2 FILLER_66_593 ();
 sg13g2_fill_1 FILLER_66_595 ();
 sg13g2_decap_8 FILLER_66_639 ();
 sg13g2_decap_8 FILLER_66_646 ();
 sg13g2_decap_4 FILLER_66_657 ();
 sg13g2_fill_1 FILLER_66_699 ();
 sg13g2_fill_2 FILLER_66_749 ();
 sg13g2_fill_2 FILLER_66_791 ();
 sg13g2_fill_1 FILLER_66_793 ();
 sg13g2_fill_1 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_4 FILLER_67_105 ();
 sg13g2_decap_4 FILLER_67_129 ();
 sg13g2_fill_2 FILLER_67_133 ();
 sg13g2_decap_4 FILLER_67_143 ();
 sg13g2_fill_1 FILLER_67_147 ();
 sg13g2_fill_2 FILLER_67_182 ();
 sg13g2_fill_2 FILLER_67_193 ();
 sg13g2_fill_1 FILLER_67_195 ();
 sg13g2_fill_2 FILLER_67_217 ();
 sg13g2_fill_1 FILLER_67_219 ();
 sg13g2_fill_2 FILLER_67_233 ();
 sg13g2_fill_1 FILLER_67_235 ();
 sg13g2_decap_8 FILLER_67_240 ();
 sg13g2_decap_8 FILLER_67_247 ();
 sg13g2_fill_2 FILLER_67_281 ();
 sg13g2_fill_2 FILLER_67_413 ();
 sg13g2_fill_2 FILLER_67_450 ();
 sg13g2_fill_1 FILLER_67_452 ();
 sg13g2_fill_2 FILLER_67_463 ();
 sg13g2_fill_1 FILLER_67_465 ();
 sg13g2_fill_1 FILLER_67_493 ();
 sg13g2_fill_2 FILLER_67_579 ();
 sg13g2_fill_1 FILLER_67_581 ();
 sg13g2_decap_8 FILLER_67_618 ();
 sg13g2_decap_8 FILLER_67_625 ();
 sg13g2_decap_8 FILLER_67_632 ();
 sg13g2_decap_8 FILLER_67_639 ();
 sg13g2_decap_8 FILLER_67_646 ();
 sg13g2_decap_8 FILLER_67_653 ();
 sg13g2_decap_8 FILLER_67_660 ();
 sg13g2_fill_2 FILLER_67_667 ();
 sg13g2_fill_1 FILLER_67_669 ();
 sg13g2_fill_2 FILLER_67_683 ();
 sg13g2_fill_2 FILLER_67_711 ();
 sg13g2_fill_1 FILLER_67_713 ();
 sg13g2_fill_2 FILLER_67_747 ();
 sg13g2_fill_2 FILLER_67_777 ();
 sg13g2_fill_1 FILLER_67_818 ();
 sg13g2_fill_1 FILLER_67_845 ();
 sg13g2_fill_2 FILLER_67_859 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_151 ();
 sg13g2_fill_1 FILLER_68_158 ();
 sg13g2_decap_4 FILLER_68_174 ();
 sg13g2_fill_1 FILLER_68_178 ();
 sg13g2_fill_2 FILLER_68_208 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_fill_2 FILLER_68_235 ();
 sg13g2_fill_2 FILLER_68_242 ();
 sg13g2_fill_2 FILLER_68_257 ();
 sg13g2_fill_1 FILLER_68_259 ();
 sg13g2_fill_1 FILLER_68_271 ();
 sg13g2_fill_1 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_356 ();
 sg13g2_fill_1 FILLER_68_389 ();
 sg13g2_fill_1 FILLER_68_431 ();
 sg13g2_fill_2 FILLER_68_449 ();
 sg13g2_fill_2 FILLER_68_482 ();
 sg13g2_fill_2 FILLER_68_581 ();
 sg13g2_fill_2 FILLER_68_606 ();
 sg13g2_fill_1 FILLER_68_608 ();
 sg13g2_decap_8 FILLER_68_622 ();
 sg13g2_decap_8 FILLER_68_629 ();
 sg13g2_decap_8 FILLER_68_636 ();
 sg13g2_decap_8 FILLER_68_643 ();
 sg13g2_decap_8 FILLER_68_650 ();
 sg13g2_decap_8 FILLER_68_657 ();
 sg13g2_decap_8 FILLER_68_664 ();
 sg13g2_decap_8 FILLER_68_671 ();
 sg13g2_fill_1 FILLER_68_678 ();
 sg13g2_fill_1 FILLER_68_709 ();
 sg13g2_fill_2 FILLER_68_719 ();
 sg13g2_fill_2 FILLER_68_747 ();
 sg13g2_fill_1 FILLER_68_788 ();
 sg13g2_fill_2 FILLER_68_801 ();
 sg13g2_decap_4 FILLER_68_857 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_4 FILLER_69_105 ();
 sg13g2_fill_2 FILLER_69_122 ();
 sg13g2_fill_2 FILLER_69_150 ();
 sg13g2_decap_4 FILLER_69_183 ();
 sg13g2_fill_1 FILLER_69_197 ();
 sg13g2_fill_1 FILLER_69_207 ();
 sg13g2_fill_1 FILLER_69_240 ();
 sg13g2_decap_4 FILLER_69_251 ();
 sg13g2_fill_2 FILLER_69_255 ();
 sg13g2_fill_2 FILLER_69_260 ();
 sg13g2_fill_2 FILLER_69_271 ();
 sg13g2_fill_1 FILLER_69_282 ();
 sg13g2_fill_2 FILLER_69_350 ();
 sg13g2_fill_2 FILLER_69_358 ();
 sg13g2_fill_1 FILLER_69_386 ();
 sg13g2_fill_1 FILLER_69_568 ();
 sg13g2_fill_1 FILLER_69_587 ();
 sg13g2_decap_8 FILLER_69_618 ();
 sg13g2_decap_8 FILLER_69_625 ();
 sg13g2_decap_8 FILLER_69_632 ();
 sg13g2_decap_8 FILLER_69_639 ();
 sg13g2_decap_8 FILLER_69_646 ();
 sg13g2_decap_8 FILLER_69_653 ();
 sg13g2_decap_8 FILLER_69_660 ();
 sg13g2_decap_8 FILLER_69_667 ();
 sg13g2_decap_8 FILLER_69_674 ();
 sg13g2_fill_2 FILLER_69_681 ();
 sg13g2_fill_1 FILLER_69_683 ();
 sg13g2_fill_2 FILLER_69_693 ();
 sg13g2_fill_1 FILLER_69_695 ();
 sg13g2_fill_1 FILLER_69_755 ();
 sg13g2_fill_2 FILLER_69_771 ();
 sg13g2_fill_2 FILLER_69_786 ();
 sg13g2_fill_1 FILLER_69_788 ();
 sg13g2_fill_1 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_69_852 ();
 sg13g2_fill_2 FILLER_69_859 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_4 FILLER_70_112 ();
 sg13g2_fill_1 FILLER_70_150 ();
 sg13g2_fill_2 FILLER_70_214 ();
 sg13g2_decap_4 FILLER_70_246 ();
 sg13g2_fill_1 FILLER_70_250 ();
 sg13g2_fill_2 FILLER_70_282 ();
 sg13g2_fill_1 FILLER_70_336 ();
 sg13g2_fill_2 FILLER_70_364 ();
 sg13g2_fill_1 FILLER_70_411 ();
 sg13g2_fill_2 FILLER_70_421 ();
 sg13g2_fill_2 FILLER_70_465 ();
 sg13g2_fill_1 FILLER_70_467 ();
 sg13g2_fill_2 FILLER_70_482 ();
 sg13g2_fill_1 FILLER_70_484 ();
 sg13g2_fill_2 FILLER_70_508 ();
 sg13g2_decap_8 FILLER_70_631 ();
 sg13g2_decap_8 FILLER_70_638 ();
 sg13g2_decap_8 FILLER_70_645 ();
 sg13g2_decap_8 FILLER_70_652 ();
 sg13g2_decap_8 FILLER_70_659 ();
 sg13g2_decap_8 FILLER_70_666 ();
 sg13g2_decap_8 FILLER_70_673 ();
 sg13g2_decap_8 FILLER_70_680 ();
 sg13g2_decap_8 FILLER_70_687 ();
 sg13g2_decap_4 FILLER_70_694 ();
 sg13g2_fill_1 FILLER_70_702 ();
 sg13g2_fill_2 FILLER_70_722 ();
 sg13g2_fill_2 FILLER_70_732 ();
 sg13g2_fill_1 FILLER_70_734 ();
 sg13g2_fill_1 FILLER_70_765 ();
 sg13g2_fill_2 FILLER_70_792 ();
 sg13g2_fill_1 FILLER_70_794 ();
 sg13g2_decap_8 FILLER_70_842 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_4 FILLER_70_856 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_4 FILLER_71_154 ();
 sg13g2_fill_2 FILLER_71_158 ();
 sg13g2_decap_8 FILLER_71_169 ();
 sg13g2_decap_8 FILLER_71_176 ();
 sg13g2_decap_8 FILLER_71_183 ();
 sg13g2_decap_8 FILLER_71_190 ();
 sg13g2_fill_1 FILLER_71_197 ();
 sg13g2_decap_8 FILLER_71_220 ();
 sg13g2_decap_8 FILLER_71_240 ();
 sg13g2_fill_1 FILLER_71_247 ();
 sg13g2_fill_1 FILLER_71_313 ();
 sg13g2_fill_1 FILLER_71_350 ();
 sg13g2_fill_2 FILLER_71_360 ();
 sg13g2_fill_2 FILLER_71_442 ();
 sg13g2_fill_1 FILLER_71_444 ();
 sg13g2_fill_1 FILLER_71_485 ();
 sg13g2_fill_2 FILLER_71_496 ();
 sg13g2_fill_1 FILLER_71_498 ();
 sg13g2_fill_2 FILLER_71_517 ();
 sg13g2_decap_8 FILLER_71_621 ();
 sg13g2_decap_8 FILLER_71_628 ();
 sg13g2_decap_8 FILLER_71_635 ();
 sg13g2_decap_8 FILLER_71_642 ();
 sg13g2_decap_8 FILLER_71_649 ();
 sg13g2_decap_8 FILLER_71_656 ();
 sg13g2_decap_8 FILLER_71_663 ();
 sg13g2_decap_8 FILLER_71_670 ();
 sg13g2_decap_8 FILLER_71_677 ();
 sg13g2_decap_8 FILLER_71_684 ();
 sg13g2_decap_8 FILLER_71_691 ();
 sg13g2_decap_8 FILLER_71_698 ();
 sg13g2_fill_2 FILLER_71_705 ();
 sg13g2_fill_1 FILLER_71_707 ();
 sg13g2_decap_4 FILLER_71_716 ();
 sg13g2_fill_2 FILLER_71_720 ();
 sg13g2_fill_2 FILLER_71_730 ();
 sg13g2_decap_4 FILLER_71_736 ();
 sg13g2_fill_1 FILLER_71_740 ();
 sg13g2_fill_2 FILLER_71_757 ();
 sg13g2_fill_1 FILLER_71_759 ();
 sg13g2_fill_2 FILLER_71_764 ();
 sg13g2_fill_1 FILLER_71_766 ();
 sg13g2_fill_1 FILLER_71_775 ();
 sg13g2_fill_1 FILLER_71_806 ();
 sg13g2_decap_8 FILLER_71_828 ();
 sg13g2_decap_8 FILLER_71_835 ();
 sg13g2_decap_8 FILLER_71_842 ();
 sg13g2_decap_8 FILLER_71_849 ();
 sg13g2_decap_4 FILLER_71_856 ();
 sg13g2_fill_2 FILLER_71_860 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_fill_2 FILLER_72_238 ();
 sg13g2_fill_1 FILLER_72_240 ();
 sg13g2_fill_1 FILLER_72_267 ();
 sg13g2_fill_1 FILLER_72_377 ();
 sg13g2_fill_2 FILLER_72_432 ();
 sg13g2_fill_1 FILLER_72_434 ();
 sg13g2_decap_4 FILLER_72_471 ();
 sg13g2_decap_8 FILLER_72_606 ();
 sg13g2_decap_8 FILLER_72_613 ();
 sg13g2_decap_8 FILLER_72_620 ();
 sg13g2_decap_8 FILLER_72_627 ();
 sg13g2_decap_8 FILLER_72_634 ();
 sg13g2_decap_8 FILLER_72_641 ();
 sg13g2_decap_8 FILLER_72_648 ();
 sg13g2_decap_8 FILLER_72_655 ();
 sg13g2_decap_8 FILLER_72_662 ();
 sg13g2_decap_8 FILLER_72_669 ();
 sg13g2_decap_8 FILLER_72_676 ();
 sg13g2_decap_8 FILLER_72_683 ();
 sg13g2_decap_8 FILLER_72_690 ();
 sg13g2_decap_8 FILLER_72_697 ();
 sg13g2_decap_8 FILLER_72_704 ();
 sg13g2_decap_8 FILLER_72_711 ();
 sg13g2_decap_8 FILLER_72_718 ();
 sg13g2_decap_8 FILLER_72_725 ();
 sg13g2_decap_8 FILLER_72_732 ();
 sg13g2_decap_8 FILLER_72_739 ();
 sg13g2_decap_8 FILLER_72_746 ();
 sg13g2_decap_8 FILLER_72_753 ();
 sg13g2_decap_8 FILLER_72_760 ();
 sg13g2_decap_8 FILLER_72_767 ();
 sg13g2_fill_2 FILLER_72_774 ();
 sg13g2_decap_4 FILLER_72_780 ();
 sg13g2_fill_2 FILLER_72_788 ();
 sg13g2_fill_1 FILLER_72_790 ();
 sg13g2_fill_2 FILLER_72_795 ();
 sg13g2_fill_1 FILLER_72_797 ();
 sg13g2_fill_1 FILLER_72_804 ();
 sg13g2_decap_8 FILLER_72_818 ();
 sg13g2_decap_8 FILLER_72_825 ();
 sg13g2_decap_8 FILLER_72_832 ();
 sg13g2_decap_8 FILLER_72_839 ();
 sg13g2_decap_8 FILLER_72_846 ();
 sg13g2_decap_8 FILLER_72_853 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_8 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_decap_4 FILLER_73_238 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_fill_1 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_389 ();
 sg13g2_fill_1 FILLER_73_396 ();
 sg13g2_fill_1 FILLER_73_415 ();
 sg13g2_fill_2 FILLER_73_425 ();
 sg13g2_fill_2 FILLER_73_440 ();
 sg13g2_fill_2 FILLER_73_446 ();
 sg13g2_decap_8 FILLER_73_458 ();
 sg13g2_decap_4 FILLER_73_475 ();
 sg13g2_fill_2 FILLER_73_498 ();
 sg13g2_fill_1 FILLER_73_500 ();
 sg13g2_fill_1 FILLER_73_510 ();
 sg13g2_fill_2 FILLER_73_526 ();
 sg13g2_fill_2 FILLER_73_564 ();
 sg13g2_fill_1 FILLER_73_566 ();
 sg13g2_fill_1 FILLER_73_575 ();
 sg13g2_decap_8 FILLER_73_601 ();
 sg13g2_decap_8 FILLER_73_608 ();
 sg13g2_decap_8 FILLER_73_615 ();
 sg13g2_decap_8 FILLER_73_622 ();
 sg13g2_decap_8 FILLER_73_629 ();
 sg13g2_decap_8 FILLER_73_636 ();
 sg13g2_decap_8 FILLER_73_643 ();
 sg13g2_decap_8 FILLER_73_650 ();
 sg13g2_decap_8 FILLER_73_657 ();
 sg13g2_decap_8 FILLER_73_664 ();
 sg13g2_decap_8 FILLER_73_671 ();
 sg13g2_decap_8 FILLER_73_678 ();
 sg13g2_decap_8 FILLER_73_685 ();
 sg13g2_decap_8 FILLER_73_692 ();
 sg13g2_decap_8 FILLER_73_699 ();
 sg13g2_decap_8 FILLER_73_706 ();
 sg13g2_decap_8 FILLER_73_713 ();
 sg13g2_decap_8 FILLER_73_720 ();
 sg13g2_decap_8 FILLER_73_727 ();
 sg13g2_decap_8 FILLER_73_734 ();
 sg13g2_decap_8 FILLER_73_741 ();
 sg13g2_decap_8 FILLER_73_748 ();
 sg13g2_decap_8 FILLER_73_755 ();
 sg13g2_decap_8 FILLER_73_762 ();
 sg13g2_decap_8 FILLER_73_769 ();
 sg13g2_decap_8 FILLER_73_776 ();
 sg13g2_decap_8 FILLER_73_783 ();
 sg13g2_decap_8 FILLER_73_790 ();
 sg13g2_decap_8 FILLER_73_797 ();
 sg13g2_decap_8 FILLER_73_804 ();
 sg13g2_decap_8 FILLER_73_811 ();
 sg13g2_decap_8 FILLER_73_818 ();
 sg13g2_decap_8 FILLER_73_825 ();
 sg13g2_decap_8 FILLER_73_832 ();
 sg13g2_decap_8 FILLER_73_839 ();
 sg13g2_decap_8 FILLER_73_846 ();
 sg13g2_decap_8 FILLER_73_853 ();
 sg13g2_fill_2 FILLER_73_860 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_fill_1 FILLER_74_245 ();
 sg13g2_fill_1 FILLER_74_293 ();
 sg13g2_fill_2 FILLER_74_330 ();
 sg13g2_fill_2 FILLER_74_348 ();
 sg13g2_fill_2 FILLER_74_364 ();
 sg13g2_fill_1 FILLER_74_372 ();
 sg13g2_fill_2 FILLER_74_512 ();
 sg13g2_fill_1 FILLER_74_514 ();
 sg13g2_fill_1 FILLER_74_541 ();
 sg13g2_fill_2 FILLER_74_552 ();
 sg13g2_decap_8 FILLER_74_580 ();
 sg13g2_decap_8 FILLER_74_587 ();
 sg13g2_decap_8 FILLER_74_594 ();
 sg13g2_decap_8 FILLER_74_601 ();
 sg13g2_decap_8 FILLER_74_608 ();
 sg13g2_decap_8 FILLER_74_615 ();
 sg13g2_decap_8 FILLER_74_622 ();
 sg13g2_decap_8 FILLER_74_629 ();
 sg13g2_decap_8 FILLER_74_636 ();
 sg13g2_decap_8 FILLER_74_643 ();
 sg13g2_decap_8 FILLER_74_650 ();
 sg13g2_decap_8 FILLER_74_657 ();
 sg13g2_decap_8 FILLER_74_664 ();
 sg13g2_decap_8 FILLER_74_671 ();
 sg13g2_decap_8 FILLER_74_678 ();
 sg13g2_decap_8 FILLER_74_685 ();
 sg13g2_decap_8 FILLER_74_692 ();
 sg13g2_decap_8 FILLER_74_699 ();
 sg13g2_decap_8 FILLER_74_706 ();
 sg13g2_decap_8 FILLER_74_713 ();
 sg13g2_decap_8 FILLER_74_720 ();
 sg13g2_decap_8 FILLER_74_727 ();
 sg13g2_decap_8 FILLER_74_734 ();
 sg13g2_decap_8 FILLER_74_741 ();
 sg13g2_decap_8 FILLER_74_748 ();
 sg13g2_decap_8 FILLER_74_755 ();
 sg13g2_decap_8 FILLER_74_762 ();
 sg13g2_decap_8 FILLER_74_769 ();
 sg13g2_decap_8 FILLER_74_776 ();
 sg13g2_decap_8 FILLER_74_783 ();
 sg13g2_decap_8 FILLER_74_790 ();
 sg13g2_decap_8 FILLER_74_797 ();
 sg13g2_decap_8 FILLER_74_804 ();
 sg13g2_decap_8 FILLER_74_811 ();
 sg13g2_decap_8 FILLER_74_818 ();
 sg13g2_decap_8 FILLER_74_825 ();
 sg13g2_decap_8 FILLER_74_832 ();
 sg13g2_decap_8 FILLER_74_839 ();
 sg13g2_decap_8 FILLER_74_846 ();
 sg13g2_decap_8 FILLER_74_853 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_4 FILLER_75_238 ();
 sg13g2_fill_1 FILLER_75_242 ();
 sg13g2_fill_2 FILLER_75_269 ();
 sg13g2_fill_2 FILLER_75_302 ();
 sg13g2_fill_2 FILLER_75_332 ();
 sg13g2_fill_2 FILLER_75_350 ();
 sg13g2_fill_2 FILLER_75_415 ();
 sg13g2_fill_1 FILLER_75_422 ();
 sg13g2_fill_1 FILLER_75_458 ();
 sg13g2_fill_1 FILLER_75_530 ();
 sg13g2_decap_8 FILLER_75_563 ();
 sg13g2_decap_8 FILLER_75_570 ();
 sg13g2_decap_8 FILLER_75_577 ();
 sg13g2_decap_8 FILLER_75_584 ();
 sg13g2_decap_8 FILLER_75_591 ();
 sg13g2_decap_8 FILLER_75_598 ();
 sg13g2_decap_8 FILLER_75_605 ();
 sg13g2_decap_8 FILLER_75_612 ();
 sg13g2_decap_8 FILLER_75_619 ();
 sg13g2_decap_8 FILLER_75_626 ();
 sg13g2_decap_8 FILLER_75_633 ();
 sg13g2_decap_8 FILLER_75_640 ();
 sg13g2_decap_8 FILLER_75_647 ();
 sg13g2_decap_8 FILLER_75_654 ();
 sg13g2_decap_8 FILLER_75_661 ();
 sg13g2_decap_8 FILLER_75_668 ();
 sg13g2_decap_8 FILLER_75_675 ();
 sg13g2_decap_8 FILLER_75_682 ();
 sg13g2_decap_8 FILLER_75_689 ();
 sg13g2_decap_8 FILLER_75_696 ();
 sg13g2_decap_8 FILLER_75_703 ();
 sg13g2_decap_8 FILLER_75_710 ();
 sg13g2_decap_8 FILLER_75_717 ();
 sg13g2_decap_8 FILLER_75_724 ();
 sg13g2_decap_8 FILLER_75_731 ();
 sg13g2_decap_8 FILLER_75_738 ();
 sg13g2_decap_8 FILLER_75_745 ();
 sg13g2_decap_8 FILLER_75_752 ();
 sg13g2_decap_8 FILLER_75_759 ();
 sg13g2_decap_8 FILLER_75_766 ();
 sg13g2_decap_8 FILLER_75_773 ();
 sg13g2_decap_8 FILLER_75_780 ();
 sg13g2_decap_8 FILLER_75_787 ();
 sg13g2_decap_8 FILLER_75_794 ();
 sg13g2_decap_8 FILLER_75_801 ();
 sg13g2_decap_8 FILLER_75_808 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_decap_8 FILLER_75_822 ();
 sg13g2_decap_8 FILLER_75_829 ();
 sg13g2_decap_8 FILLER_75_836 ();
 sg13g2_decap_8 FILLER_75_843 ();
 sg13g2_decap_8 FILLER_75_850 ();
 sg13g2_decap_4 FILLER_75_857 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_fill_2 FILLER_76_259 ();
 sg13g2_decap_4 FILLER_76_446 ();
 sg13g2_fill_1 FILLER_76_476 ();
 sg13g2_fill_1 FILLER_76_503 ();
 sg13g2_decap_4 FILLER_76_539 ();
 sg13g2_decap_8 FILLER_76_552 ();
 sg13g2_decap_8 FILLER_76_559 ();
 sg13g2_decap_8 FILLER_76_566 ();
 sg13g2_decap_8 FILLER_76_573 ();
 sg13g2_decap_8 FILLER_76_580 ();
 sg13g2_decap_8 FILLER_76_587 ();
 sg13g2_decap_8 FILLER_76_594 ();
 sg13g2_decap_8 FILLER_76_601 ();
 sg13g2_decap_8 FILLER_76_608 ();
 sg13g2_decap_8 FILLER_76_615 ();
 sg13g2_decap_8 FILLER_76_622 ();
 sg13g2_decap_8 FILLER_76_629 ();
 sg13g2_decap_8 FILLER_76_636 ();
 sg13g2_decap_8 FILLER_76_643 ();
 sg13g2_decap_8 FILLER_76_650 ();
 sg13g2_decap_8 FILLER_76_657 ();
 sg13g2_decap_8 FILLER_76_664 ();
 sg13g2_decap_8 FILLER_76_671 ();
 sg13g2_decap_8 FILLER_76_678 ();
 sg13g2_decap_8 FILLER_76_685 ();
 sg13g2_decap_8 FILLER_76_692 ();
 sg13g2_decap_8 FILLER_76_699 ();
 sg13g2_decap_8 FILLER_76_706 ();
 sg13g2_decap_8 FILLER_76_713 ();
 sg13g2_decap_8 FILLER_76_720 ();
 sg13g2_decap_8 FILLER_76_727 ();
 sg13g2_decap_8 FILLER_76_734 ();
 sg13g2_decap_8 FILLER_76_741 ();
 sg13g2_decap_8 FILLER_76_748 ();
 sg13g2_decap_8 FILLER_76_755 ();
 sg13g2_decap_8 FILLER_76_762 ();
 sg13g2_decap_8 FILLER_76_769 ();
 sg13g2_decap_8 FILLER_76_776 ();
 sg13g2_decap_8 FILLER_76_783 ();
 sg13g2_decap_8 FILLER_76_790 ();
 sg13g2_decap_8 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_804 ();
 sg13g2_decap_8 FILLER_76_811 ();
 sg13g2_decap_8 FILLER_76_818 ();
 sg13g2_decap_8 FILLER_76_825 ();
 sg13g2_decap_8 FILLER_76_832 ();
 sg13g2_decap_8 FILLER_76_839 ();
 sg13g2_decap_8 FILLER_76_846 ();
 sg13g2_decap_8 FILLER_76_853 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_4 FILLER_77_245 ();
 sg13g2_fill_2 FILLER_77_249 ();
 sg13g2_decap_8 FILLER_77_313 ();
 sg13g2_fill_1 FILLER_77_320 ();
 sg13g2_decap_4 FILLER_77_347 ();
 sg13g2_fill_2 FILLER_77_418 ();
 sg13g2_fill_1 FILLER_77_420 ();
 sg13g2_fill_2 FILLER_77_448 ();
 sg13g2_fill_2 FILLER_77_470 ();
 sg13g2_fill_1 FILLER_77_472 ();
 sg13g2_fill_2 FILLER_77_486 ();
 sg13g2_decap_8 FILLER_77_548 ();
 sg13g2_decap_8 FILLER_77_555 ();
 sg13g2_decap_8 FILLER_77_562 ();
 sg13g2_decap_8 FILLER_77_569 ();
 sg13g2_decap_8 FILLER_77_576 ();
 sg13g2_decap_8 FILLER_77_583 ();
 sg13g2_decap_8 FILLER_77_590 ();
 sg13g2_decap_8 FILLER_77_597 ();
 sg13g2_decap_8 FILLER_77_604 ();
 sg13g2_decap_8 FILLER_77_611 ();
 sg13g2_decap_8 FILLER_77_618 ();
 sg13g2_decap_8 FILLER_77_625 ();
 sg13g2_decap_8 FILLER_77_632 ();
 sg13g2_decap_8 FILLER_77_639 ();
 sg13g2_decap_8 FILLER_77_646 ();
 sg13g2_decap_8 FILLER_77_653 ();
 sg13g2_decap_8 FILLER_77_660 ();
 sg13g2_decap_8 FILLER_77_667 ();
 sg13g2_decap_8 FILLER_77_674 ();
 sg13g2_decap_8 FILLER_77_681 ();
 sg13g2_decap_8 FILLER_77_688 ();
 sg13g2_decap_8 FILLER_77_695 ();
 sg13g2_decap_8 FILLER_77_702 ();
 sg13g2_decap_8 FILLER_77_709 ();
 sg13g2_decap_8 FILLER_77_716 ();
 sg13g2_decap_8 FILLER_77_723 ();
 sg13g2_decap_8 FILLER_77_730 ();
 sg13g2_decap_8 FILLER_77_737 ();
 sg13g2_decap_8 FILLER_77_744 ();
 sg13g2_decap_8 FILLER_77_751 ();
 sg13g2_decap_8 FILLER_77_758 ();
 sg13g2_decap_8 FILLER_77_765 ();
 sg13g2_decap_8 FILLER_77_772 ();
 sg13g2_decap_8 FILLER_77_779 ();
 sg13g2_decap_8 FILLER_77_786 ();
 sg13g2_decap_8 FILLER_77_793 ();
 sg13g2_decap_8 FILLER_77_800 ();
 sg13g2_decap_8 FILLER_77_807 ();
 sg13g2_decap_8 FILLER_77_814 ();
 sg13g2_decap_8 FILLER_77_821 ();
 sg13g2_decap_8 FILLER_77_828 ();
 sg13g2_decap_8 FILLER_77_835 ();
 sg13g2_decap_8 FILLER_77_842 ();
 sg13g2_decap_8 FILLER_77_849 ();
 sg13g2_decap_4 FILLER_77_856 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_fill_2 FILLER_78_252 ();
 sg13g2_fill_1 FILLER_78_254 ();
 sg13g2_fill_2 FILLER_78_310 ();
 sg13g2_fill_2 FILLER_78_341 ();
 sg13g2_fill_1 FILLER_78_343 ();
 sg13g2_fill_1 FILLER_78_358 ();
 sg13g2_fill_2 FILLER_78_364 ();
 sg13g2_fill_1 FILLER_78_366 ();
 sg13g2_decap_8 FILLER_78_443 ();
 sg13g2_decap_8 FILLER_78_450 ();
 sg13g2_decap_8 FILLER_78_457 ();
 sg13g2_decap_8 FILLER_78_464 ();
 sg13g2_decap_8 FILLER_78_471 ();
 sg13g2_fill_2 FILLER_78_478 ();
 sg13g2_fill_1 FILLER_78_480 ();
 sg13g2_fill_1 FILLER_78_508 ();
 sg13g2_decap_4 FILLER_78_518 ();
 sg13g2_decap_8 FILLER_78_532 ();
 sg13g2_decap_8 FILLER_78_539 ();
 sg13g2_decap_8 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_553 ();
 sg13g2_decap_8 FILLER_78_560 ();
 sg13g2_decap_8 FILLER_78_567 ();
 sg13g2_decap_8 FILLER_78_574 ();
 sg13g2_decap_8 FILLER_78_581 ();
 sg13g2_decap_8 FILLER_78_588 ();
 sg13g2_decap_8 FILLER_78_595 ();
 sg13g2_decap_8 FILLER_78_602 ();
 sg13g2_decap_8 FILLER_78_609 ();
 sg13g2_decap_8 FILLER_78_616 ();
 sg13g2_decap_8 FILLER_78_623 ();
 sg13g2_decap_8 FILLER_78_630 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_decap_8 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_651 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_decap_8 FILLER_78_672 ();
 sg13g2_decap_8 FILLER_78_679 ();
 sg13g2_decap_8 FILLER_78_686 ();
 sg13g2_decap_8 FILLER_78_693 ();
 sg13g2_decap_8 FILLER_78_700 ();
 sg13g2_decap_8 FILLER_78_707 ();
 sg13g2_decap_8 FILLER_78_714 ();
 sg13g2_decap_8 FILLER_78_721 ();
 sg13g2_decap_8 FILLER_78_728 ();
 sg13g2_decap_8 FILLER_78_735 ();
 sg13g2_decap_8 FILLER_78_742 ();
 sg13g2_decap_8 FILLER_78_749 ();
 sg13g2_decap_8 FILLER_78_756 ();
 sg13g2_decap_8 FILLER_78_763 ();
 sg13g2_decap_8 FILLER_78_770 ();
 sg13g2_decap_8 FILLER_78_777 ();
 sg13g2_decap_8 FILLER_78_784 ();
 sg13g2_decap_8 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_798 ();
 sg13g2_decap_8 FILLER_78_805 ();
 sg13g2_decap_8 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_8 FILLER_78_854 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_fill_1 FILLER_79_280 ();
 sg13g2_fill_2 FILLER_79_286 ();
 sg13g2_decap_8 FILLER_79_306 ();
 sg13g2_fill_2 FILLER_79_313 ();
 sg13g2_fill_1 FILLER_79_315 ();
 sg13g2_decap_4 FILLER_79_350 ();
 sg13g2_fill_1 FILLER_79_354 ();
 sg13g2_fill_2 FILLER_79_379 ();
 sg13g2_fill_1 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_455 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_decap_8 FILLER_79_490 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_decap_8 FILLER_79_504 ();
 sg13g2_decap_4 FILLER_79_511 ();
 sg13g2_fill_2 FILLER_79_515 ();
 sg13g2_decap_8 FILLER_79_522 ();
 sg13g2_decap_8 FILLER_79_529 ();
 sg13g2_decap_8 FILLER_79_536 ();
 sg13g2_decap_8 FILLER_79_543 ();
 sg13g2_decap_8 FILLER_79_550 ();
 sg13g2_decap_8 FILLER_79_557 ();
 sg13g2_decap_8 FILLER_79_564 ();
 sg13g2_decap_8 FILLER_79_571 ();
 sg13g2_decap_8 FILLER_79_578 ();
 sg13g2_decap_8 FILLER_79_585 ();
 sg13g2_decap_8 FILLER_79_592 ();
 sg13g2_decap_8 FILLER_79_599 ();
 sg13g2_decap_8 FILLER_79_606 ();
 sg13g2_decap_8 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_620 ();
 sg13g2_decap_8 FILLER_79_627 ();
 sg13g2_decap_8 FILLER_79_634 ();
 sg13g2_decap_8 FILLER_79_641 ();
 sg13g2_decap_8 FILLER_79_648 ();
 sg13g2_decap_8 FILLER_79_655 ();
 sg13g2_decap_8 FILLER_79_662 ();
 sg13g2_decap_8 FILLER_79_669 ();
 sg13g2_decap_8 FILLER_79_676 ();
 sg13g2_decap_8 FILLER_79_683 ();
 sg13g2_decap_8 FILLER_79_690 ();
 sg13g2_decap_8 FILLER_79_697 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_8 FILLER_79_711 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_decap_8 FILLER_79_725 ();
 sg13g2_decap_8 FILLER_79_732 ();
 sg13g2_decap_8 FILLER_79_739 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_decap_8 FILLER_79_753 ();
 sg13g2_decap_8 FILLER_79_760 ();
 sg13g2_decap_8 FILLER_79_767 ();
 sg13g2_decap_8 FILLER_79_774 ();
 sg13g2_decap_8 FILLER_79_781 ();
 sg13g2_decap_8 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_4 FILLER_79_858 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_8 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_155 ();
 sg13g2_fill_1 FILLER_80_159 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_decap_4 FILLER_80_220 ();
 sg13g2_decap_4 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_4 FILLER_80_250 ();
 sg13g2_fill_2 FILLER_80_254 ();
 sg13g2_decap_4 FILLER_80_260 ();
 sg13g2_decap_4 FILLER_80_268 ();
 sg13g2_decap_8 FILLER_80_276 ();
 sg13g2_decap_8 FILLER_80_283 ();
 sg13g2_decap_8 FILLER_80_290 ();
 sg13g2_decap_8 FILLER_80_297 ();
 sg13g2_decap_8 FILLER_80_304 ();
 sg13g2_decap_4 FILLER_80_311 ();
 sg13g2_fill_1 FILLER_80_315 ();
 sg13g2_fill_2 FILLER_80_324 ();
 sg13g2_fill_1 FILLER_80_335 ();
 sg13g2_fill_2 FILLER_80_341 ();
 sg13g2_fill_1 FILLER_80_343 ();
 sg13g2_decap_8 FILLER_80_349 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_fill_2 FILLER_80_372 ();
 sg13g2_fill_1 FILLER_80_374 ();
 sg13g2_decap_4 FILLER_80_394 ();
 sg13g2_fill_2 FILLER_80_398 ();
 sg13g2_decap_8 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_444 ();
 sg13g2_decap_8 FILLER_80_451 ();
 sg13g2_decap_8 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_decap_8 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_479 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_decap_8 FILLER_80_493 ();
 sg13g2_decap_8 FILLER_80_500 ();
 sg13g2_decap_8 FILLER_80_507 ();
 sg13g2_decap_8 FILLER_80_514 ();
 sg13g2_decap_8 FILLER_80_521 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_decap_8 FILLER_80_535 ();
 sg13g2_decap_8 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_decap_8 FILLER_80_563 ();
 sg13g2_decap_8 FILLER_80_570 ();
 sg13g2_decap_8 FILLER_80_577 ();
 sg13g2_decap_8 FILLER_80_584 ();
 sg13g2_decap_8 FILLER_80_591 ();
 sg13g2_decap_8 FILLER_80_598 ();
 sg13g2_decap_8 FILLER_80_605 ();
 sg13g2_decap_8 FILLER_80_612 ();
 sg13g2_decap_8 FILLER_80_619 ();
 sg13g2_decap_8 FILLER_80_626 ();
 sg13g2_decap_8 FILLER_80_633 ();
 sg13g2_decap_8 FILLER_80_640 ();
 sg13g2_decap_8 FILLER_80_647 ();
 sg13g2_decap_8 FILLER_80_654 ();
 sg13g2_decap_8 FILLER_80_661 ();
 sg13g2_decap_8 FILLER_80_668 ();
 sg13g2_decap_8 FILLER_80_675 ();
 sg13g2_decap_8 FILLER_80_682 ();
 sg13g2_decap_8 FILLER_80_689 ();
 sg13g2_decap_8 FILLER_80_696 ();
 sg13g2_decap_8 FILLER_80_703 ();
 sg13g2_decap_8 FILLER_80_710 ();
 sg13g2_decap_8 FILLER_80_717 ();
 sg13g2_decap_8 FILLER_80_724 ();
 sg13g2_decap_8 FILLER_80_731 ();
 sg13g2_decap_8 FILLER_80_738 ();
 sg13g2_decap_8 FILLER_80_745 ();
 sg13g2_decap_8 FILLER_80_752 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_decap_8 FILLER_80_766 ();
 sg13g2_decap_8 FILLER_80_773 ();
 sg13g2_decap_8 FILLER_80_780 ();
 sg13g2_decap_8 FILLER_80_787 ();
 sg13g2_decap_8 FILLER_80_794 ();
 sg13g2_decap_8 FILLER_80_801 ();
 sg13g2_decap_8 FILLER_80_808 ();
 sg13g2_decap_8 FILLER_80_815 ();
 sg13g2_decap_8 FILLER_80_822 ();
 sg13g2_decap_8 FILLER_80_829 ();
 sg13g2_decap_8 FILLER_80_836 ();
 sg13g2_decap_8 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_850 ();
 sg13g2_decap_4 FILLER_80_857 ();
 sg13g2_fill_1 FILLER_80_861 ();
 assign uio_oe[0] = net541;
 assign uio_oe[1] = net542;
 assign uio_oe[2] = net543;
 assign uio_oe[3] = net544;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net545;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[1] = net18;
 assign uo_out[2] = net19;
 assign uo_out[3] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule

module tt_um_couchand_cora16 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire clk_regs;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire busy;
 wire \cpu_instance.accum[0] ;
 wire \cpu_instance.accum[10] ;
 wire \cpu_instance.accum[11] ;
 wire \cpu_instance.accum[12] ;
 wire \cpu_instance.accum[13] ;
 wire \cpu_instance.accum[14] ;
 wire \cpu_instance.accum[15] ;
 wire \cpu_instance.accum[1] ;
 wire \cpu_instance.accum[2] ;
 wire \cpu_instance.accum[3] ;
 wire \cpu_instance.accum[4] ;
 wire \cpu_instance.accum[5] ;
 wire \cpu_instance.accum[6] ;
 wire \cpu_instance.accum[7] ;
 wire \cpu_instance.accum[8] ;
 wire \cpu_instance.accum[9] ;
 wire \cpu_instance.carry ;
 wire \cpu_instance.dp[0] ;
 wire \cpu_instance.dp[10] ;
 wire \cpu_instance.dp[11] ;
 wire \cpu_instance.dp[12] ;
 wire \cpu_instance.dp[13] ;
 wire \cpu_instance.dp[14] ;
 wire \cpu_instance.dp[15] ;
 wire \cpu_instance.dp[1] ;
 wire \cpu_instance.dp[2] ;
 wire \cpu_instance.dp[3] ;
 wire \cpu_instance.dp[4] ;
 wire \cpu_instance.dp[5] ;
 wire \cpu_instance.dp[6] ;
 wire \cpu_instance.dp[7] ;
 wire \cpu_instance.dp[8] ;
 wire \cpu_instance.dp[9] ;
 wire \cpu_instance.halt ;
 wire \cpu_instance.inst[0] ;
 wire \cpu_instance.inst[10] ;
 wire \cpu_instance.inst[11] ;
 wire \cpu_instance.inst[12] ;
 wire \cpu_instance.inst[13] ;
 wire \cpu_instance.inst[14] ;
 wire \cpu_instance.inst[15] ;
 wire \cpu_instance.inst[1] ;
 wire \cpu_instance.inst[2] ;
 wire \cpu_instance.inst[3] ;
 wire \cpu_instance.inst[4] ;
 wire \cpu_instance.inst[5] ;
 wire \cpu_instance.inst[6] ;
 wire \cpu_instance.inst[7] ;
 wire \cpu_instance.inst[8] ;
 wire \cpu_instance.inst[9] ;
 wire \cpu_instance.neg ;
 wire \cpu_instance.pc[0] ;
 wire \cpu_instance.pc[10] ;
 wire \cpu_instance.pc[11] ;
 wire \cpu_instance.pc[12] ;
 wire \cpu_instance.pc[13] ;
 wire \cpu_instance.pc[14] ;
 wire \cpu_instance.pc[15] ;
 wire \cpu_instance.pc[1] ;
 wire \cpu_instance.pc[2] ;
 wire \cpu_instance.pc[3] ;
 wire \cpu_instance.pc[4] ;
 wire \cpu_instance.pc[5] ;
 wire \cpu_instance.pc[6] ;
 wire \cpu_instance.pc[7] ;
 wire \cpu_instance.pc[8] ;
 wire \cpu_instance.pc[9] ;
 wire \cpu_instance.ram_data_out[0] ;
 wire \cpu_instance.ram_data_out[10] ;
 wire \cpu_instance.ram_data_out[11] ;
 wire \cpu_instance.ram_data_out[12] ;
 wire \cpu_instance.ram_data_out[13] ;
 wire \cpu_instance.ram_data_out[14] ;
 wire \cpu_instance.ram_data_out[15] ;
 wire \cpu_instance.ram_data_out[1] ;
 wire \cpu_instance.ram_data_out[2] ;
 wire \cpu_instance.ram_data_out[3] ;
 wire \cpu_instance.ram_data_out[4] ;
 wire \cpu_instance.ram_data_out[5] ;
 wire \cpu_instance.ram_data_out[6] ;
 wire \cpu_instance.ram_data_out[7] ;
 wire \cpu_instance.ram_data_out[8] ;
 wire \cpu_instance.ram_data_out[9] ;
 wire \cpu_instance.skip ;
 wire \cpu_instance.skipped ;
 wire \cpu_instance.sp[10] ;
 wire \cpu_instance.sp[11] ;
 wire \cpu_instance.sp[12] ;
 wire \cpu_instance.sp[13] ;
 wire \cpu_instance.sp[14] ;
 wire \cpu_instance.sp[15] ;
 wire \cpu_instance.sp[1] ;
 wire \cpu_instance.sp[2] ;
 wire \cpu_instance.sp[3] ;
 wire \cpu_instance.sp[4] ;
 wire \cpu_instance.sp[5] ;
 wire \cpu_instance.sp[6] ;
 wire \cpu_instance.sp[7] ;
 wire \cpu_instance.sp[8] ;
 wire \cpu_instance.sp[9] ;
 wire \cpu_instance.sp_minus_two[1] ;
 wire net155;
 wire \cpu_instance.spi_mosi ;
 wire \cpu_instance.spi_ram.addr[0] ;
 wire \cpu_instance.spi_ram.addr[10] ;
 wire \cpu_instance.spi_ram.addr[11] ;
 wire \cpu_instance.spi_ram.addr[12] ;
 wire \cpu_instance.spi_ram.addr[13] ;
 wire \cpu_instance.spi_ram.addr[14] ;
 wire \cpu_instance.spi_ram.addr[15] ;
 wire \cpu_instance.spi_ram.addr[1] ;
 wire \cpu_instance.spi_ram.addr[2] ;
 wire \cpu_instance.spi_ram.addr[3] ;
 wire \cpu_instance.spi_ram.addr[4] ;
 wire \cpu_instance.spi_ram.addr[5] ;
 wire \cpu_instance.spi_ram.addr[6] ;
 wire \cpu_instance.spi_ram.addr[7] ;
 wire \cpu_instance.spi_ram.addr[8] ;
 wire \cpu_instance.spi_ram.addr[9] ;
 wire \cpu_instance.spi_ram.bits_remaining[0] ;
 wire \cpu_instance.spi_ram.bits_remaining[1] ;
 wire \cpu_instance.spi_ram.bits_remaining[2] ;
 wire \cpu_instance.spi_ram.bits_remaining[3] ;
 wire \cpu_instance.spi_ram.fsm_state[0] ;
 wire \cpu_instance.spi_ram.fsm_state[1] ;
 wire \cpu_instance.spi_ram.spi_miso_buf ;
 wire \cpu_instance.spi_ram.spi_select ;
 wire \cpu_instance.spi_ram.writing ;
 wire \cpu_instance.state[0] ;
 wire \cpu_instance.state[1] ;
 wire \cpu_instance.state[2] ;
 wire \cpu_instance.state[3] ;
 wire \cpu_instance.trap ;
 wire \cpu_instance.zero ;
 wire net12;
 wire net13;
 wire net152;
 wire net153;
 wire net154;
 wire net14;
 wire net15;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;

 sg13g2_inv_1 _2752_ (.Y(_1886_),
    .A(net1282));
 sg13g2_inv_1 _2753_ (.Y(_1887_),
    .A(net296));
 sg13g2_inv_1 _2754_ (.Y(_1888_),
    .A(net293));
 sg13g2_inv_1 _2755_ (.Y(_1889_),
    .A(\cpu_instance.sp[12] ));
 sg13g2_inv_1 _2756_ (.Y(_1890_),
    .A(\cpu_instance.sp[10] ));
 sg13g2_inv_1 _2757_ (.Y(_1891_),
    .A(net239));
 sg13g2_inv_1 _2758_ (.Y(_1892_),
    .A(net301));
 sg13g2_inv_1 _2759_ (.Y(_1893_),
    .A(net189));
 sg13g2_inv_1 _2760_ (.Y(_1894_),
    .A(\cpu_instance.pc[14] ));
 sg13g2_inv_1 _2761_ (.Y(_1895_),
    .A(\cpu_instance.pc[13] ));
 sg13g2_inv_2 _2762_ (.Y(_1896_),
    .A(net304));
 sg13g2_inv_2 _2763_ (.Y(_1897_),
    .A(\cpu_instance.pc[11] ));
 sg13g2_inv_1 _2764_ (.Y(_1898_),
    .A(\cpu_instance.pc[10] ));
 sg13g2_inv_2 _2765_ (.Y(_1899_),
    .A(net314));
 sg13g2_inv_1 _2766_ (.Y(_1900_),
    .A(\cpu_instance.pc[6] ));
 sg13g2_inv_1 _2767_ (.Y(_1901_),
    .A(\cpu_instance.pc[5] ));
 sg13g2_inv_1 _2768_ (.Y(_1902_),
    .A(net312));
 sg13g2_inv_2 _2769_ (.Y(_1903_),
    .A(net171));
 sg13g2_inv_2 _2770_ (.Y(_1904_),
    .A(\cpu_instance.ram_data_out[15] ));
 sg13g2_inv_1 _2771_ (.Y(_1905_),
    .A(net1286));
 sg13g2_inv_4 _2772_ (.A(net276),
    .Y(_1906_));
 sg13g2_inv_1 _2773_ (.Y(_1907_),
    .A(net1288));
 sg13g2_inv_2 _2774_ (.Y(_1908_),
    .A(net281));
 sg13g2_inv_1 _2775_ (.Y(_1909_),
    .A(net1291));
 sg13g2_inv_2 _2776_ (.Y(_1910_),
    .A(net254));
 sg13g2_inv_2 _2777_ (.Y(_1911_),
    .A(net1292));
 sg13g2_inv_2 _2778_ (.Y(_1912_),
    .A(net307));
 sg13g2_inv_4 _2779_ (.A(net1297),
    .Y(_1913_));
 sg13g2_inv_2 _2780_ (.Y(_1914_),
    .A(net248));
 sg13g2_inv_4 _2781_ (.A(net1302),
    .Y(_1915_));
 sg13g2_inv_2 _2782_ (.Y(_1916_),
    .A(net297));
 sg13g2_inv_4 _2783_ (.A(net299),
    .Y(_1917_));
 sg13g2_inv_2 _2784_ (.Y(_1918_),
    .A(net257));
 sg13g2_inv_2 _2785_ (.Y(_1919_),
    .A(\cpu_instance.ram_data_out[5] ));
 sg13g2_inv_2 _2786_ (.Y(_1920_),
    .A(\cpu_instance.ram_data_out[4] ));
 sg13g2_inv_2 _2787_ (.Y(_1921_),
    .A(net309));
 sg13g2_inv_2 _2788_ (.Y(_1922_),
    .A(net300));
 sg13g2_inv_1 _2789_ (.Y(_1923_),
    .A(\cpu_instance.ram_data_out[1] ));
 sg13g2_inv_2 _2790_ (.Y(_1924_),
    .A(net245));
 sg13g2_inv_2 _2791_ (.Y(_1925_),
    .A(\cpu_instance.accum[15] ));
 sg13g2_inv_2 _2792_ (.Y(_1926_),
    .A(\cpu_instance.accum[14] ));
 sg13g2_inv_2 _2793_ (.Y(_1927_),
    .A(net1304));
 sg13g2_inv_1 _2794_ (.Y(_1928_),
    .A(net1305));
 sg13g2_inv_1 _2795_ (.Y(_1929_),
    .A(net1306));
 sg13g2_inv_2 _2796_ (.Y(_1930_),
    .A(net1309));
 sg13g2_inv_2 _2797_ (.Y(_1931_),
    .A(\cpu_instance.accum[7] ));
 sg13g2_inv_4 _2798_ (.A(\cpu_instance.accum[5] ),
    .Y(_1932_));
 sg13g2_inv_1 _2799_ (.Y(_1933_),
    .A(\cpu_instance.accum[4] ));
 sg13g2_inv_2 _2800_ (.Y(_1934_),
    .A(net318));
 sg13g2_inv_4 _2801_ (.A(net313),
    .Y(_1935_));
 sg13g2_inv_4 _2802_ (.A(\cpu_instance.accum[1] ),
    .Y(_1936_));
 sg13g2_inv_1 _2803_ (.Y(_1937_),
    .A(\cpu_instance.accum[0] ));
 sg13g2_inv_1 _2804_ (.Y(_1938_),
    .A(net160));
 sg13g2_inv_1 _2805_ (.Y(_1939_),
    .A(net156));
 sg13g2_inv_1 _2806_ (.Y(_1940_),
    .A(net159));
 sg13g2_inv_1 _2807_ (.Y(_1941_),
    .A(net161));
 sg13g2_inv_1 _2808_ (.Y(_1942_),
    .A(net164));
 sg13g2_inv_2 _2809_ (.Y(_1943_),
    .A(net1319));
 sg13g2_inv_1 _2810_ (.Y(_1944_),
    .A(net268));
 sg13g2_inv_1 _5238__2 (.Y(net155),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _2812_ (.Y(_1945_),
    .A(net197));
 sg13g2_inv_1 _2813_ (.Y(_1946_),
    .A(net174));
 sg13g2_inv_1 _2814_ (.Y(_1947_),
    .A(net2));
 sg13g2_inv_1 _2815_ (.Y(_1948_),
    .A(_0022_));
 sg13g2_inv_1 _2816_ (.Y(_1949_),
    .A(_0038_));
 sg13g2_inv_2 _2817_ (.Y(_1950_),
    .A(_0039_));
 sg13g2_inv_1 _2818_ (.Y(_1951_),
    .A(net157));
 sg13g2_inv_2 _2819_ (.Y(_1952_),
    .A(_0036_));
 sg13g2_inv_4 _2820_ (.A(_0034_),
    .Y(_1953_));
 sg13g2_inv_2 _2821_ (.Y(_1954_),
    .A(_0033_));
 sg13g2_inv_1 _2822_ (.Y(_1955_),
    .A(net165));
 sg13g2_inv_2 _2823_ (.Y(_1956_),
    .A(_0032_));
 sg13g2_inv_1 _2824_ (.Y(_1957_),
    .A(_0031_));
 sg13g2_inv_1 _2825_ (.Y(_1958_),
    .A(_0015_));
 sg13g2_inv_1 _2826_ (.Y(_1959_),
    .A(net172));
 sg13g2_inv_1 _2827_ (.Y(_1960_),
    .A(_0030_));
 sg13g2_inv_1 _2828_ (.Y(_1961_),
    .A(_0029_));
 sg13g2_inv_1 _2829_ (.Y(_1962_),
    .A(net195));
 sg13g2_inv_1 _2830_ (.Y(_1963_),
    .A(_0028_));
 sg13g2_inv_2 _2831_ (.Y(_1964_),
    .A(_0027_));
 sg13g2_inv_1 _2832_ (.Y(_1965_),
    .A(net176));
 sg13g2_inv_1 _2833_ (.Y(_1966_),
    .A(_0026_));
 sg13g2_inv_1 _2834_ (.Y(_1967_),
    .A(_0025_));
 sg13g2_inv_1 _2835_ (.Y(_1968_),
    .A(net169));
 sg13g2_inv_1 _2836_ (.Y(_1969_),
    .A(_0024_));
 sg13g2_inv_1 _2837_ (.Y(_1970_),
    .A(net167));
 sg13g2_inv_1 _2838_ (.Y(_1971_),
    .A(_0052_));
 sg13g2_inv_1 _2839_ (.Y(_1972_),
    .A(_0053_));
 sg13g2_inv_2 _2840_ (.Y(_1973_),
    .A(net1337));
 sg13g2_or2_2 _2841_ (.X(_1974_),
    .B(\cpu_instance.spi_ram.fsm_state[0] ),
    .A(\cpu_instance.spi_ram.fsm_state[1] ));
 sg13g2_inv_2 _2842_ (.Y(\cpu_instance.spi_ram.spi_select ),
    .A(net1277));
 sg13g2_nor2_1 _2843_ (.A(\cpu_instance.state[3] ),
    .B(net1282),
    .Y(_1975_));
 sg13g2_nor2_2 _2844_ (.A(\cpu_instance.state[1] ),
    .B(_1888_),
    .Y(_1976_));
 sg13g2_nand2_1 _2845_ (.Y(_1977_),
    .A(_1887_),
    .B(\cpu_instance.state[0] ));
 sg13g2_nor2b_2 _2846_ (.A(net1282),
    .B_N(\cpu_instance.state[3] ),
    .Y(_1978_));
 sg13g2_nand2b_1 _2847_ (.Y(_1979_),
    .B(\cpu_instance.state[3] ),
    .A_N(net1282));
 sg13g2_nor2_1 _2848_ (.A(_1887_),
    .B(\cpu_instance.state[0] ),
    .Y(_1980_));
 sg13g2_nand2_1 _2849_ (.Y(_1981_),
    .A(\cpu_instance.state[1] ),
    .B(_1888_));
 sg13g2_a22oi_1 _2850_ (.Y(_1982_),
    .B1(_1978_),
    .B2(_1980_),
    .A2(_1976_),
    .A1(_1975_));
 sg13g2_inv_1 _2851_ (.Y(\cpu_instance.halt ),
    .A(_1982_));
 sg13g2_nor4_1 _2852_ (.A(\cpu_instance.spi_ram.bits_remaining[3] ),
    .B(\cpu_instance.spi_ram.bits_remaining[2] ),
    .C(\cpu_instance.spi_ram.bits_remaining[1] ),
    .D(\cpu_instance.spi_ram.fsm_state[1] ),
    .Y(_1983_));
 sg13g2_o21ai_1 _2853_ (.B1(_1983_),
    .Y(_1984_),
    .A1(\cpu_instance.spi_ram.bits_remaining[0] ),
    .A2(_1945_));
 sg13g2_nor2b_2 _2854_ (.A(\cpu_instance.spi_ram.fsm_state[0] ),
    .B_N(\cpu_instance.spi_ram.fsm_state[1] ),
    .Y(_1985_));
 sg13g2_nand2b_2 _2855_ (.Y(_1986_),
    .B(\cpu_instance.spi_ram.fsm_state[1] ),
    .A_N(\cpu_instance.spi_ram.fsm_state[0] ));
 sg13g2_and2_1 _2856_ (.A(\cpu_instance.spi_ram.fsm_state[1] ),
    .B(\cpu_instance.spi_ram.fsm_state[0] ),
    .X(_1987_));
 sg13g2_a22oi_1 _2857_ (.Y(_1988_),
    .B1(net1275),
    .B2(\cpu_instance.ram_data_out[15] ),
    .A2(_1985_),
    .A1(\cpu_instance.spi_ram.addr[15] ));
 sg13g2_a21oi_1 _2858_ (.A1(_1984_),
    .A2(_1988_),
    .Y(\cpu_instance.spi_mosi ),
    .B1(\cpu_instance.spi_ram.spi_select ));
 sg13g2_nor2_1 _2859_ (.A(net1282),
    .B(_1981_),
    .Y(\cpu_instance.trap ));
 sg13g2_nor3_2 _2860_ (.A(\cpu_instance.state[3] ),
    .B(\cpu_instance.state[2] ),
    .C(\cpu_instance.state[0] ),
    .Y(_1989_));
 sg13g2_nor2_1 _2861_ (.A(\cpu_instance.halt ),
    .B(_1989_),
    .Y(busy));
 sg13g2_or2_2 _2862_ (.X(_1990_),
    .B(\cpu_instance.state[0] ),
    .A(\cpu_instance.state[1] ));
 sg13g2_nor2_2 _2863_ (.A(_1979_),
    .B(_1990_),
    .Y(_1991_));
 sg13g2_nor2b_2 _2864_ (.A(\cpu_instance.state[3] ),
    .B_N(net1282),
    .Y(_1992_));
 sg13g2_nand2b_2 _2865_ (.Y(_1993_),
    .B(net1282),
    .A_N(\cpu_instance.state[3] ));
 sg13g2_mux2_1 _2866_ (.A0(_1979_),
    .A1(_1993_),
    .S(_1990_),
    .X(_1994_));
 sg13g2_mux2_1 _2867_ (.A0(_1978_),
    .A1(_1992_),
    .S(_1990_),
    .X(_1995_));
 sg13g2_nor2_2 _2868_ (.A(net1291),
    .B(_1911_),
    .Y(_1996_));
 sg13g2_nand2_1 _2869_ (.Y(_1997_),
    .A(_1909_),
    .B(net1292));
 sg13g2_nor2_2 _2870_ (.A(net1268),
    .B(_1997_),
    .Y(_1998_));
 sg13g2_nand2_2 _2871_ (.Y(_1999_),
    .A(net1264),
    .B(_1996_));
 sg13g2_or2_1 _2872_ (.X(_2000_),
    .B(net1301),
    .A(net1298));
 sg13g2_nor4_1 _2873_ (.A(\cpu_instance.inst[15] ),
    .B(net1287),
    .C(net1288),
    .D(_2000_),
    .Y(_2001_));
 sg13g2_and4_2 _2874_ (.A(net1286),
    .B(net1264),
    .C(_1996_),
    .D(_2001_),
    .X(_2002_));
 sg13g2_nand4_1 _2875_ (.B(net1264),
    .C(_1996_),
    .A(net1286),
    .Y(_2003_),
    .D(_2001_));
 sg13g2_and3_1 _2876_ (.X(_2004_),
    .A(\cpu_instance.inst[15] ),
    .B(_1905_),
    .C(net1264));
 sg13g2_a21oi_1 _2877_ (.A1(net1292),
    .A2(_2004_),
    .Y(_2005_),
    .B1(_2002_));
 sg13g2_a21o_1 _2878_ (.A2(_2004_),
    .A1(net1292),
    .B1(_2002_),
    .X(_2006_));
 sg13g2_nor2_2 _2879_ (.A(net1303),
    .B(net1215),
    .Y(_2007_));
 sg13g2_nand2_2 _2880_ (.Y(_2008_),
    .A(net1291),
    .B(net1265));
 sg13g2_nor2b_1 _2881_ (.A(net1286),
    .B_N(net1287),
    .Y(_2009_));
 sg13g2_nand2b_2 _2882_ (.Y(_2010_),
    .B(net1287),
    .A_N(net1286));
 sg13g2_nor3_2 _2883_ (.A(net1281),
    .B(net1284),
    .C(_2010_),
    .Y(_2011_));
 sg13g2_nand3b_1 _2884_ (.B(_2009_),
    .C(net1288),
    .Y(_2012_),
    .A_N(net1284));
 sg13g2_nor2_1 _2885_ (.A(_2008_),
    .B(_2012_),
    .Y(_2013_));
 sg13g2_o21ai_1 _2886_ (.B1(_2013_),
    .Y(_2014_),
    .A1(_1958_),
    .A2(_2007_));
 sg13g2_a21oi_2 _2887_ (.B1(_2014_),
    .Y(_2015_),
    .A2(_2007_),
    .A1(_0023_));
 sg13g2_nand2_1 _2888_ (.Y(_2016_),
    .A(\cpu_instance.inst[0] ),
    .B(net1213));
 sg13g2_and2_1 _2889_ (.A(_2013_),
    .B(_2016_),
    .X(_2017_));
 sg13g2_and2_2 _2890_ (.A(_1915_),
    .B(_2017_),
    .X(_2018_));
 sg13g2_nand2_1 _2891_ (.Y(_2019_),
    .A(_1915_),
    .B(_2017_));
 sg13g2_nor4_2 _2892_ (.A(net1285),
    .B(net1286),
    .C(net1287),
    .Y(_2020_),
    .D(net1288));
 sg13g2_or4_2 _2893_ (.A(net1285),
    .B(net1286),
    .C(net1287),
    .D(net1288),
    .X(_2021_));
 sg13g2_nand2_2 _2894_ (.Y(_2022_),
    .A(net1298),
    .B(net1302));
 sg13g2_inv_1 _2895_ (.Y(_2023_),
    .A(_2022_));
 sg13g2_nor2_2 _2896_ (.A(_2021_),
    .B(_2022_),
    .Y(_2024_));
 sg13g2_and2_1 _2897_ (.A(_1998_),
    .B(_2024_),
    .X(_2025_));
 sg13g2_nor2_2 _2898_ (.A(_1909_),
    .B(net1293),
    .Y(_2026_));
 sg13g2_nand2_1 _2899_ (.Y(_2027_),
    .A(net1291),
    .B(_1911_));
 sg13g2_nor2_2 _2900_ (.A(net1270),
    .B(_2027_),
    .Y(_2028_));
 sg13g2_and2_1 _2901_ (.A(_2024_),
    .B(_2028_),
    .X(_2029_));
 sg13g2_nand2_2 _2902_ (.Y(_2030_),
    .A(_2024_),
    .B(_2028_));
 sg13g2_nand2b_2 _2903_ (.Y(_2031_),
    .B(_2030_),
    .A_N(net1208));
 sg13g2_nor4_2 _2904_ (.A(\cpu_instance.inst[11] ),
    .B(net1284),
    .C(net1270),
    .Y(_2032_),
    .D(_2010_));
 sg13g2_nor3_2 _2905_ (.A(\cpu_instance.inst[14] ),
    .B(\cpu_instance.inst[13] ),
    .C(net1284),
    .Y(_2033_));
 sg13g2_nor2b_2 _2906_ (.A(_2008_),
    .B_N(_2033_),
    .Y(_2034_));
 sg13g2_nor4_2 _2907_ (.A(net1289),
    .B(net1284),
    .C(_2008_),
    .Y(_2035_),
    .D(_2010_));
 sg13g2_or4_2 _2908_ (.A(net1289),
    .B(net1284),
    .C(_2008_),
    .D(_2010_),
    .X(_2036_));
 sg13g2_nor4_1 _2909_ (.A(_2031_),
    .B(_2032_),
    .C(_2034_),
    .D(net1204),
    .Y(_2037_));
 sg13g2_nand3b_1 _2910_ (.B(_2019_),
    .C(_2037_),
    .Y(_2038_),
    .A_N(net1111));
 sg13g2_inv_2 _2911_ (.Y(_2039_),
    .A(net1067));
 sg13g2_nor2_2 _2912_ (.A(net1290),
    .B(net1293),
    .Y(_2040_));
 sg13g2_nand2_2 _2913_ (.Y(_2041_),
    .A(_1909_),
    .B(_1911_));
 sg13g2_nor2_1 _2914_ (.A(_2000_),
    .B(_2041_),
    .Y(_2042_));
 sg13g2_nor2_1 _2915_ (.A(net1285),
    .B(net1281),
    .Y(_2043_));
 sg13g2_nor4_1 _2916_ (.A(net1286),
    .B(net1287),
    .C(_2000_),
    .D(_2041_),
    .Y(_2044_));
 sg13g2_and2_1 _2917_ (.A(_2043_),
    .B(_2044_),
    .X(_2045_));
 sg13g2_nand2_2 _2918_ (.Y(_2046_),
    .A(net1264),
    .B(_2045_));
 sg13g2_nor2b_2 _2919_ (.A(net1302),
    .B_N(net1299),
    .Y(_2047_));
 sg13g2_nand2_1 _2920_ (.Y(_2048_),
    .A(_2020_),
    .B(_2047_));
 sg13g2_nor4_2 _2921_ (.A(net1285),
    .B(net1281),
    .C(_1911_),
    .Y(_2049_),
    .D(_2010_));
 sg13g2_and4_2 _2922_ (.A(net1290),
    .B(net1263),
    .C(_2023_),
    .D(_2049_),
    .X(_2050_));
 sg13g2_nand4_1 _2923_ (.B(net1263),
    .C(_2023_),
    .A(net1290),
    .Y(_2051_),
    .D(_2049_));
 sg13g2_nand3_1 _2924_ (.B(_2047_),
    .C(_2049_),
    .A(net1290),
    .Y(_2052_));
 sg13g2_nand4_1 _2925_ (.B(net1298),
    .C(net1263),
    .A(net1290),
    .Y(_2053_),
    .D(_2049_));
 sg13g2_o21ai_1 _2926_ (.B1(_2051_),
    .Y(_2054_),
    .A1(net1269),
    .A2(_2052_));
 sg13g2_nor3_2 _2927_ (.A(net1285),
    .B(net1281),
    .C(_2010_),
    .Y(_2055_));
 sg13g2_nand2_2 _2928_ (.Y(_2056_),
    .A(_2009_),
    .B(_2043_));
 sg13g2_nand2_1 _2929_ (.Y(_2057_),
    .A(net1290),
    .B(net1292));
 sg13g2_nand4_1 _2930_ (.B(net1292),
    .C(_2047_),
    .A(net1290),
    .Y(_2058_),
    .D(_2055_));
 sg13g2_nor2_1 _2931_ (.A(net1267),
    .B(_2058_),
    .Y(_2059_));
 sg13g2_nor2_2 _2932_ (.A(net1268),
    .B(_2057_),
    .Y(_2060_));
 sg13g2_nand2b_2 _2933_ (.Y(_2061_),
    .B(net1264),
    .A_N(_2057_));
 sg13g2_nor3_2 _2934_ (.A(_2022_),
    .B(_2056_),
    .C(_2061_),
    .Y(_2062_));
 sg13g2_nand3_1 _2935_ (.B(_2055_),
    .C(_2060_),
    .A(_2023_),
    .Y(_2063_));
 sg13g2_o21ai_1 _2936_ (.B1(_2063_),
    .Y(_2064_),
    .A1(net1269),
    .A2(_2058_));
 sg13g2_nor4_2 _2937_ (.A(_1913_),
    .B(net1301),
    .C(net1267),
    .Y(_2065_),
    .D(_2021_));
 sg13g2_nand2_1 _2938_ (.Y(_2066_),
    .A(_2026_),
    .B(_2065_));
 sg13g2_nor2_2 _2939_ (.A(net1298),
    .B(_2021_),
    .Y(_2067_));
 sg13g2_nand2_2 _2940_ (.Y(_2068_),
    .A(_1913_),
    .B(_2020_));
 sg13g2_nand2_1 _2941_ (.Y(_2069_),
    .A(net1303),
    .B(_2067_));
 sg13g2_nand3_1 _2942_ (.B(_2040_),
    .C(_2067_),
    .A(net1301),
    .Y(_2070_));
 sg13g2_nor2_1 _2943_ (.A(_1999_),
    .B(_2068_),
    .Y(_2071_));
 sg13g2_nand2_1 _2944_ (.Y(_2072_),
    .A(_1998_),
    .B(_2067_));
 sg13g2_nor2_2 _2945_ (.A(net1201),
    .B(net1199),
    .Y(_2073_));
 sg13g2_nor3_1 _2946_ (.A(net1288),
    .B(\cpu_instance.inst[11] ),
    .C(net1270),
    .Y(_2074_));
 sg13g2_a21oi_1 _2947_ (.A1(_2033_),
    .A2(_2074_),
    .Y(_2075_),
    .B1(_2002_));
 sg13g2_a21o_1 _2948_ (.A2(_2074_),
    .A1(_2033_),
    .B1(_2002_),
    .X(_2076_));
 sg13g2_nand2_1 _2949_ (.Y(_2077_),
    .A(_2024_),
    .B(_2040_));
 sg13g2_nand3_1 _2950_ (.B(_2024_),
    .C(_2040_),
    .A(net1263),
    .Y(_2078_));
 sg13g2_nor2_1 _2951_ (.A(_1977_),
    .B(_1993_),
    .Y(_2079_));
 sg13g2_nand2_1 _2952_ (.Y(_2080_),
    .A(_1976_),
    .B(_1992_));
 sg13g2_nor2_2 _2953_ (.A(net1281),
    .B(net1291),
    .Y(_2081_));
 sg13g2_and3_1 _2954_ (.X(_2082_),
    .A(net1263),
    .B(_2033_),
    .C(_2081_));
 sg13g2_nand3_1 _2955_ (.B(_2033_),
    .C(_2081_),
    .A(net1263),
    .Y(_2083_));
 sg13g2_nor2_1 _2956_ (.A(net1268),
    .B(_2021_),
    .Y(_2084_));
 sg13g2_nor4_2 _2957_ (.A(net1298),
    .B(net1267),
    .C(_2021_),
    .Y(_2085_),
    .D(_2041_));
 sg13g2_nand2_2 _2958_ (.Y(_2086_),
    .A(_2040_),
    .B(_2065_));
 sg13g2_inv_1 _2959_ (.Y(_2087_),
    .A(_2086_));
 sg13g2_nand2b_2 _2960_ (.Y(_2088_),
    .B(_2086_),
    .A_N(_2085_));
 sg13g2_nand2b_2 _2961_ (.Y(_2089_),
    .B(net1194),
    .A_N(_2064_));
 sg13g2_nand3_1 _2962_ (.B(_2047_),
    .C(_2084_),
    .A(_2026_),
    .Y(_2090_));
 sg13g2_nand4_1 _2963_ (.B(net1248),
    .C(_2083_),
    .A(net1191),
    .Y(_2091_),
    .D(_2090_));
 sg13g2_a21oi_1 _2964_ (.A1(_0041_),
    .A2(net1067),
    .Y(_2092_),
    .B1(_2091_));
 sg13g2_nand3_1 _2965_ (.B(_2055_),
    .C(_2060_),
    .A(_2047_),
    .Y(_2093_));
 sg13g2_nor3_2 _2966_ (.A(_2022_),
    .B(_2056_),
    .C(_2061_),
    .Y(_2094_));
 sg13g2_nand3_1 _2967_ (.B(_2055_),
    .C(_2060_),
    .A(_2023_),
    .Y(_2095_));
 sg13g2_nand3_1 _2968_ (.B(_2055_),
    .C(_2060_),
    .A(net1298),
    .Y(_2096_));
 sg13g2_nand3_1 _2969_ (.B(_2090_),
    .C(_2096_),
    .A(_2046_),
    .Y(_2097_));
 sg13g2_nor2b_1 _2970_ (.A(_2038_),
    .B_N(_2097_),
    .Y(_2098_));
 sg13g2_nand2_2 _2971_ (.Y(_2099_),
    .A(net1194),
    .B(net1180));
 sg13g2_nor3_1 _2972_ (.A(net1267),
    .B(_2021_),
    .C(_2041_),
    .Y(_2100_));
 sg13g2_nor3_1 _2973_ (.A(_2098_),
    .B(_2099_),
    .C(_2100_),
    .Y(_2101_));
 sg13g2_a21oi_1 _2974_ (.A1(_1911_),
    .A2(_2004_),
    .Y(_2102_),
    .B1(_2031_));
 sg13g2_and2_2 _2975_ (.A(net1278),
    .B(_2102_),
    .X(_2103_));
 sg13g2_nand3_1 _2976_ (.B(_2066_),
    .C(_2078_),
    .A(_2046_),
    .Y(_2104_));
 sg13g2_nor3_2 _2977_ (.A(net1238),
    .B(_2089_),
    .C(_2104_),
    .Y(_2105_));
 sg13g2_nand3_1 _2978_ (.B(net1108),
    .C(_2105_),
    .A(net1067),
    .Y(_2106_));
 sg13g2_nor2_2 _2979_ (.A(_1981_),
    .B(_1993_),
    .Y(_2107_));
 sg13g2_nand2_1 _2980_ (.Y(_2108_),
    .A(_1980_),
    .B(_1992_));
 sg13g2_nor2_1 _2981_ (.A(net1277),
    .B(net1227),
    .Y(_2109_));
 sg13g2_nand2_1 _2982_ (.Y(_2110_),
    .A(net1273),
    .B(net1230));
 sg13g2_nor3_2 _2983_ (.A(net1303),
    .B(_1999_),
    .C(_2068_),
    .Y(_2111_));
 sg13g2_nor4_1 _2984_ (.A(_2007_),
    .B(net1201),
    .C(_2110_),
    .D(_2111_),
    .Y(_2112_));
 sg13g2_nor2_2 _2985_ (.A(_1999_),
    .B(_2069_),
    .Y(_2113_));
 sg13g2_inv_1 _2986_ (.Y(_2114_),
    .A(_2113_));
 sg13g2_nor2_2 _2987_ (.A(_1999_),
    .B(_2048_),
    .Y(_2115_));
 sg13g2_nor2_1 _2988_ (.A(_2113_),
    .B(net1176),
    .Y(_2116_));
 sg13g2_and2_2 _2989_ (.A(_1996_),
    .B(_2065_),
    .X(_2117_));
 sg13g2_nor3_1 _2990_ (.A(net1248),
    .B(_2113_),
    .C(net1178),
    .Y(_2118_));
 sg13g2_nand2_2 _2991_ (.Y(_2119_),
    .A(net1235),
    .B(_2116_));
 sg13g2_nor2_1 _2992_ (.A(_2061_),
    .B(_2069_),
    .Y(_2120_));
 sg13g2_nor2_1 _2993_ (.A(_1905_),
    .B(net1284),
    .Y(_2121_));
 sg13g2_nor4_2 _2994_ (.A(_1905_),
    .B(\cpu_instance.inst[13] ),
    .C(net1291),
    .Y(_2122_),
    .D(net1284));
 sg13g2_and2_2 _2995_ (.A(net1266),
    .B(_2122_),
    .X(_2123_));
 sg13g2_nand2_1 _2996_ (.Y(_2124_),
    .A(net1266),
    .B(_2122_));
 sg13g2_a21oi_1 _2997_ (.A1(net1288),
    .A2(net1223),
    .Y(_2125_),
    .B1(_2120_));
 sg13g2_a21o_1 _2998_ (.A2(net1223),
    .A1(net1288),
    .B1(_2120_),
    .X(_2126_));
 sg13g2_nand3_1 _2999_ (.B(net1166),
    .C(net1163),
    .A(_2112_),
    .Y(_2127_));
 sg13g2_nand2_1 _3000_ (.Y(_2128_),
    .A(\cpu_instance.state[1] ),
    .B(_1989_));
 sg13g2_nand2_1 _3001_ (.Y(_2129_),
    .A(_2026_),
    .B(net1247));
 sg13g2_o21ai_1 _3002_ (.B1(_2128_),
    .Y(_2130_),
    .A1(_2048_),
    .A2(_2129_));
 sg13g2_nor2_2 _3003_ (.A(_1990_),
    .B(_1993_),
    .Y(_2131_));
 sg13g2_nand2b_1 _3004_ (.Y(_2132_),
    .B(_1992_),
    .A_N(_1990_));
 sg13g2_nand2_1 _3005_ (.Y(_2133_),
    .A(_1976_),
    .B(_1978_));
 sg13g2_a21oi_1 _3006_ (.A1(_1976_),
    .A2(_1978_),
    .Y(_2134_),
    .B1(_2131_));
 sg13g2_nand3b_1 _3007_ (.B(\cpu_instance.state[1] ),
    .C(\cpu_instance.state[0] ),
    .Y(_2135_),
    .A_N(\cpu_instance.state[3] ));
 sg13g2_nand2_1 _3008_ (.Y(_2136_),
    .A(_1982_),
    .B(_2132_));
 sg13g2_nand2_1 _3009_ (.Y(_2137_),
    .A(_2133_),
    .B(_2135_));
 sg13g2_a21oi_2 _3010_ (.B1(net1239),
    .Y(_2138_),
    .A2(_2045_),
    .A1(net1264));
 sg13g2_nand2_2 _3011_ (.Y(_2139_),
    .A(_2046_),
    .B(net1250));
 sg13g2_nand2_1 _3012_ (.Y(_2140_),
    .A(_2090_),
    .B(net1159));
 sg13g2_nor2_1 _3013_ (.A(_2077_),
    .B(_2140_),
    .Y(_2141_));
 sg13g2_o21ai_1 _3014_ (.B1(_1974_),
    .Y(_2142_),
    .A1(_1991_),
    .A2(net1230));
 sg13g2_nand2_1 _3015_ (.Y(_2143_),
    .A(net1263),
    .B(_2142_));
 sg13g2_a21oi_1 _3016_ (.A1(_2059_),
    .A2(_2109_),
    .Y(_2144_),
    .B1(_2143_));
 sg13g2_nor4_1 _3017_ (.A(net1301),
    .B(_1997_),
    .C(_2068_),
    .D(net1226),
    .Y(_2145_));
 sg13g2_and2_1 _3018_ (.A(_1887_),
    .B(_1989_),
    .X(_2146_));
 sg13g2_nor2_2 _3019_ (.A(_2039_),
    .B(net1185),
    .Y(_2147_));
 sg13g2_nand2_1 _3020_ (.Y(_2148_),
    .A(net1067),
    .B(net1189));
 sg13g2_nand2_1 _3021_ (.Y(_2149_),
    .A(net1239),
    .B(net1060));
 sg13g2_nor2_1 _3022_ (.A(net1191),
    .B(_2088_),
    .Y(_2150_));
 sg13g2_nor2_1 _3023_ (.A(_2007_),
    .B(net1226),
    .Y(_2151_));
 sg13g2_nor2_2 _3024_ (.A(_2046_),
    .B(net1239),
    .Y(_2152_));
 sg13g2_nor3_1 _3025_ (.A(_2045_),
    .B(net1199),
    .C(net1238),
    .Y(_2153_));
 sg13g2_a22oi_1 _3026_ (.Y(_2154_),
    .B1(_2153_),
    .B2(net1232),
    .A2(_2101_),
    .A1(_2092_));
 sg13g2_nand3_1 _3027_ (.B(net1247),
    .C(_2084_),
    .A(_2042_),
    .Y(_2155_));
 sg13g2_nand2_1 _3028_ (.Y(_2156_),
    .A(_2127_),
    .B(_2155_));
 sg13g2_a21oi_1 _3029_ (.A1(_2070_),
    .A2(_2086_),
    .Y(_2157_),
    .B1(net1238));
 sg13g2_nor3_1 _3030_ (.A(_2136_),
    .B(_2141_),
    .C(_2157_),
    .Y(_2158_));
 sg13g2_nor4_1 _3031_ (.A(_2130_),
    .B(_2137_),
    .C(_2145_),
    .D(_2146_),
    .Y(_2159_));
 sg13g2_a22oi_1 _3032_ (.Y(_2160_),
    .B1(_2109_),
    .B2(_2117_),
    .A2(_2099_),
    .A1(net1247));
 sg13g2_nand4_1 _3033_ (.B(_2158_),
    .C(_2159_),
    .A(_2144_),
    .Y(_2161_),
    .D(_2160_));
 sg13g2_or4_1 _3034_ (.A(_2151_),
    .B(_2152_),
    .C(_2156_),
    .D(_2161_),
    .X(_2162_));
 sg13g2_a21oi_1 _3035_ (.A1(_2105_),
    .A2(_2150_),
    .Y(_2163_),
    .B1(_2162_));
 sg13g2_and4_2 _3036_ (.A(_2106_),
    .B(_2149_),
    .C(_2154_),
    .D(_2163_),
    .X(_2164_));
 sg13g2_nand2b_1 _3037_ (.Y(_2165_),
    .B(net260),
    .A_N(_2164_));
 sg13g2_and2_1 _3038_ (.A(_1907_),
    .B(_2034_),
    .X(_2166_));
 sg13g2_nand2_1 _3039_ (.Y(_2167_),
    .A(_1907_),
    .B(_2034_));
 sg13g2_a21o_1 _3040_ (.A2(_2122_),
    .A1(_0013_),
    .B1(net1270),
    .X(_2168_));
 sg13g2_nor3_1 _3041_ (.A(net1268),
    .B(_2057_),
    .C(_2068_),
    .Y(_2169_));
 sg13g2_nand4_1 _3042_ (.B(net1293),
    .C(net1265),
    .A(net1291),
    .Y(_2170_),
    .D(_2067_));
 sg13g2_nand2_2 _3043_ (.Y(_2171_),
    .A(_2003_),
    .B(_2170_));
 sg13g2_a221oi_1 _3044_ (.B2(_2067_),
    .C1(_2002_),
    .B1(_2060_),
    .A1(_2011_),
    .Y(_2172_),
    .A2(_2028_));
 sg13g2_nand2b_1 _3045_ (.Y(_2173_),
    .B(_0013_),
    .A_N(net1299));
 sg13g2_nand3b_1 _3046_ (.B(net1302),
    .C(_0013_),
    .Y(_2174_),
    .A_N(net1298));
 sg13g2_inv_1 _3047_ (.Y(_2175_),
    .A(_2174_));
 sg13g2_nor2_2 _3048_ (.A(net1293),
    .B(_2022_),
    .Y(_2176_));
 sg13g2_a21oi_1 _3049_ (.A1(net8),
    .A2(_2176_),
    .Y(_2177_),
    .B1(net1262));
 sg13g2_a21oi_2 _3050_ (.B1(_2177_),
    .Y(_2178_),
    .A2(net1262),
    .A1(_0016_));
 sg13g2_a221oi_1 _3051_ (.B2(_2178_),
    .C1(net1224),
    .B1(_2172_),
    .A1(_1969_),
    .Y(_2179_),
    .A2(net1175));
 sg13g2_nor2_2 _3052_ (.A(net1222),
    .B(_2179_),
    .Y(_2180_));
 sg13g2_nand2_2 _3053_ (.Y(_2181_),
    .A(_1904_),
    .B(net1236));
 sg13g2_o21ai_1 _3054_ (.B1(net1244),
    .Y(_2182_),
    .A1(net1222),
    .A2(_2179_));
 sg13g2_nand2_2 _3055_ (.Y(_2183_),
    .A(_2181_),
    .B(_2182_));
 sg13g2_inv_1 _3056_ (.Y(_2184_),
    .A(_2183_));
 sg13g2_nand2_1 _3057_ (.Y(_2185_),
    .A(_1969_),
    .B(_2184_));
 sg13g2_nor2_1 _3058_ (.A(_1969_),
    .B(_2184_),
    .Y(_2186_));
 sg13g2_xnor2_1 _3059_ (.Y(_2187_),
    .A(_0024_),
    .B(_2183_));
 sg13g2_inv_1 _3060_ (.Y(_2188_),
    .A(_2187_));
 sg13g2_a21oi_1 _3061_ (.A1(net7),
    .A2(_2176_),
    .Y(_2189_),
    .B1(net1260));
 sg13g2_a21oi_2 _3062_ (.B1(_2189_),
    .Y(_2190_),
    .A2(net1260),
    .A1(_0017_));
 sg13g2_a221oi_1 _3063_ (.B2(_2190_),
    .C1(net1224),
    .B1(_2172_),
    .A1(_1967_),
    .Y(_2191_),
    .A2(net1175));
 sg13g2_nor2_2 _3064_ (.A(net1221),
    .B(_2191_),
    .Y(_2192_));
 sg13g2_nor3_2 _3065_ (.A(net1236),
    .B(net1221),
    .C(_2191_),
    .Y(_2193_));
 sg13g2_nor2_2 _3066_ (.A(_0043_),
    .B(net1244),
    .Y(_2194_));
 sg13g2_nor2_1 _3067_ (.A(_2193_),
    .B(_2194_),
    .Y(_2195_));
 sg13g2_nor2_1 _3068_ (.A(_1926_),
    .B(_2195_),
    .Y(_2196_));
 sg13g2_nor3_2 _3069_ (.A(\cpu_instance.accum[14] ),
    .B(_2193_),
    .C(_2194_),
    .Y(_2197_));
 sg13g2_nor2_2 _3070_ (.A(_2196_),
    .B(_2197_),
    .Y(_2198_));
 sg13g2_a21oi_1 _3071_ (.A1(net6),
    .A2(_2176_),
    .Y(_2199_),
    .B1(net1260));
 sg13g2_a21oi_2 _3072_ (.B1(_2199_),
    .Y(_2200_),
    .A2(net1261),
    .A1(_0018_));
 sg13g2_a221oi_1 _3073_ (.B2(_2200_),
    .C1(net1224),
    .B1(_2172_),
    .A1(_1966_),
    .Y(_2201_),
    .A2(net1175));
 sg13g2_nor2_2 _3074_ (.A(net1221),
    .B(_2201_),
    .Y(_2202_));
 sg13g2_or2_2 _3075_ (.X(_2203_),
    .B(_2201_),
    .A(net1221));
 sg13g2_nor2_1 _3076_ (.A(_0044_),
    .B(net1243),
    .Y(_2204_));
 sg13g2_a21oi_2 _3077_ (.B1(_2204_),
    .Y(_2205_),
    .A2(_2202_),
    .A1(net1244));
 sg13g2_or2_1 _3078_ (.X(_2206_),
    .B(_2205_),
    .A(net1304));
 sg13g2_nand2_1 _3079_ (.Y(_2207_),
    .A(net1304),
    .B(_2205_));
 sg13g2_a21oi_1 _3080_ (.A1(net5),
    .A2(_2176_),
    .Y(_2208_),
    .B1(net1260));
 sg13g2_a21oi_2 _3081_ (.B1(_2208_),
    .Y(_2209_),
    .A2(net1260),
    .A1(_0019_));
 sg13g2_a221oi_1 _3082_ (.B2(_2209_),
    .C1(net1224),
    .B1(_2172_),
    .A1(_1964_),
    .Y(_2210_),
    .A2(net1175));
 sg13g2_nor2_2 _3083_ (.A(net1222),
    .B(_2210_),
    .Y(_2211_));
 sg13g2_or2_2 _3084_ (.X(_2212_),
    .B(_2210_),
    .A(net1222));
 sg13g2_nor3_2 _3085_ (.A(net1236),
    .B(net1221),
    .C(_2210_),
    .Y(_2213_));
 sg13g2_nor2_2 _3086_ (.A(_0045_),
    .B(net1243),
    .Y(_2214_));
 sg13g2_o21ai_1 _3087_ (.B1(net1305),
    .Y(_2215_),
    .A1(_2213_),
    .A2(_2214_));
 sg13g2_or3_1 _3088_ (.A(net1305),
    .B(_2213_),
    .C(_2214_),
    .X(_2216_));
 sg13g2_and2_2 _3089_ (.A(_2215_),
    .B(_2216_),
    .X(_2217_));
 sg13g2_inv_1 _3090_ (.Y(_2218_),
    .A(_2217_));
 sg13g2_a21oi_1 _3091_ (.A1(net4),
    .A2(_2176_),
    .Y(_2219_),
    .B1(net1260));
 sg13g2_a21oi_2 _3092_ (.B1(_2219_),
    .Y(_2220_),
    .A2(net1261),
    .A1(_0020_));
 sg13g2_a221oi_1 _3093_ (.B2(_2220_),
    .C1(net1224),
    .B1(_2172_),
    .A1(_1963_),
    .Y(_2221_),
    .A2(net1175));
 sg13g2_nor2_2 _3094_ (.A(net1221),
    .B(_2221_),
    .Y(_2222_));
 sg13g2_nor3_2 _3095_ (.A(net1236),
    .B(net1221),
    .C(_2221_),
    .Y(_2223_));
 sg13g2_nor2_1 _3096_ (.A(_0046_),
    .B(net1243),
    .Y(_2224_));
 sg13g2_nor2_1 _3097_ (.A(_2223_),
    .B(_2224_),
    .Y(_2225_));
 sg13g2_nor2_1 _3098_ (.A(net1306),
    .B(_2225_),
    .Y(_2226_));
 sg13g2_a21oi_1 _3099_ (.A1(net3),
    .A2(_2176_),
    .Y(_2227_),
    .B1(net1260));
 sg13g2_a21oi_2 _3100_ (.B1(_2227_),
    .Y(_2228_),
    .A2(net1260),
    .A1(_0021_));
 sg13g2_a221oi_1 _3101_ (.B2(_2228_),
    .C1(net1224),
    .B1(_2172_),
    .A1(_1961_),
    .Y(_2229_),
    .A2(net1175));
 sg13g2_nor2_2 _3102_ (.A(net1221),
    .B(_2229_),
    .Y(_2230_));
 sg13g2_nor2_1 _3103_ (.A(_0047_),
    .B(net1243),
    .Y(_2231_));
 sg13g2_a21oi_2 _3104_ (.B1(_2231_),
    .Y(_2232_),
    .A2(_2230_),
    .A1(net1243));
 sg13g2_nand2b_1 _3105_ (.Y(_2233_),
    .B(net1307),
    .A_N(_2232_));
 sg13g2_inv_1 _3106_ (.Y(_2234_),
    .A(_2233_));
 sg13g2_nor2b_1 _3107_ (.A(net1307),
    .B_N(_2232_),
    .Y(_2235_));
 sg13g2_nor2_2 _3108_ (.A(_2234_),
    .B(_2235_),
    .Y(_2236_));
 sg13g2_a21oi_1 _3109_ (.A1(net2),
    .A2(_2176_),
    .Y(_2237_),
    .B1(net1261));
 sg13g2_a21oi_2 _3110_ (.B1(_2237_),
    .Y(_2238_),
    .A2(net1262),
    .A1(_0022_));
 sg13g2_a221oi_1 _3111_ (.B2(_2238_),
    .C1(net1224),
    .B1(_2172_),
    .A1(_1960_),
    .Y(_2239_),
    .A2(net1175));
 sg13g2_a21o_1 _3112_ (.A2(_2122_),
    .A1(_0014_),
    .B1(net1272),
    .X(_2240_));
 sg13g2_nor2_2 _3113_ (.A(_2239_),
    .B(_2240_),
    .Y(_2241_));
 sg13g2_nand2_2 _3114_ (.Y(_2242_),
    .A(_0048_),
    .B(net1236));
 sg13g2_o21ai_1 _3115_ (.B1(net1246),
    .Y(_2243_),
    .A1(_2239_),
    .A2(_2240_));
 sg13g2_nand2_1 _3116_ (.Y(_2244_),
    .A(_2242_),
    .B(_2243_));
 sg13g2_nand3_1 _3117_ (.B(_2242_),
    .C(_2243_),
    .A(_1930_),
    .Y(_2245_));
 sg13g2_nand2_1 _3118_ (.Y(_2246_),
    .A(net1309),
    .B(_2244_));
 sg13g2_a21oi_1 _3119_ (.A1(net1),
    .A2(_2176_),
    .Y(_2247_),
    .B1(net1262));
 sg13g2_a21oi_2 _3120_ (.B1(_2247_),
    .Y(_2248_),
    .A2(net1262),
    .A1(_0023_));
 sg13g2_a221oi_1 _3121_ (.B2(_2248_),
    .C1(net1224),
    .B1(_2172_),
    .A1(_1957_),
    .Y(_2249_),
    .A2(net1175));
 sg13g2_o21ai_1 _3122_ (.B1(net1265),
    .Y(_2250_),
    .A1(_1958_),
    .A2(_2124_));
 sg13g2_nor2_2 _3123_ (.A(_2249_),
    .B(_2250_),
    .Y(_2251_));
 sg13g2_nor3_2 _3124_ (.A(net1236),
    .B(_2249_),
    .C(_2250_),
    .Y(_2252_));
 sg13g2_nor2_2 _3125_ (.A(_0049_),
    .B(net1244),
    .Y(_2253_));
 sg13g2_nor2_1 _3126_ (.A(_2252_),
    .B(_2253_),
    .Y(_2254_));
 sg13g2_and2_1 _3127_ (.A(net1310),
    .B(_2254_),
    .X(_2255_));
 sg13g2_o21ai_1 _3128_ (.B1(net1311),
    .Y(_2256_),
    .A1(_2252_),
    .A2(_2253_));
 sg13g2_nor3_1 _3129_ (.A(net1310),
    .B(_2252_),
    .C(_2253_),
    .Y(_2257_));
 sg13g2_xnor2_1 _3130_ (.Y(_2258_),
    .A(net1310),
    .B(_2254_));
 sg13g2_and2_1 _3131_ (.A(_0013_),
    .B(_2047_),
    .X(_2259_));
 sg13g2_nand2_1 _3132_ (.Y(_2260_),
    .A(_0013_),
    .B(_2047_));
 sg13g2_nand4_1 _3133_ (.B(net1265),
    .C(_2011_),
    .A(net1299),
    .Y(_2261_),
    .D(_2026_));
 sg13g2_nand2_2 _3134_ (.Y(_2262_),
    .A(_2260_),
    .B(_2261_));
 sg13g2_and3_1 _3135_ (.X(_2263_),
    .A(net1293),
    .B(\cpu_instance.inst[7] ),
    .C(_2173_));
 sg13g2_mux2_1 _3136_ (.A0(_2263_),
    .A1(net8),
    .S(_2262_),
    .X(_2264_));
 sg13g2_nor4_2 _3137_ (.A(net1298),
    .B(net1270),
    .C(_2012_),
    .Y(_2265_),
    .D(_2027_));
 sg13g2_nor3_1 _3138_ (.A(_2002_),
    .B(_2169_),
    .C(_2265_),
    .Y(_2266_));
 sg13g2_nor2b_1 _3139_ (.A(_2122_),
    .B_N(_2266_),
    .Y(_2267_));
 sg13g2_a21oi_1 _3140_ (.A1(_2003_),
    .A2(_2170_),
    .Y(_2268_),
    .B1(_2123_));
 sg13g2_nand2b_1 _3141_ (.Y(_2269_),
    .B(_1915_),
    .A_N(_2173_));
 sg13g2_inv_1 _3142_ (.Y(_2270_),
    .A(_2269_));
 sg13g2_or2_1 _3143_ (.X(_2271_),
    .B(_2265_),
    .A(net1223));
 sg13g2_nor3_2 _3144_ (.A(net1223),
    .B(_2265_),
    .C(_2270_),
    .Y(_2272_));
 sg13g2_or2_1 _3145_ (.X(_2273_),
    .B(_2272_),
    .A(net1174));
 sg13g2_nor3_1 _3146_ (.A(_0016_),
    .B(net1174),
    .C(_2272_),
    .Y(_2274_));
 sg13g2_a221oi_1 _3147_ (.B2(_1956_),
    .C1(_2274_),
    .B1(net1174),
    .A1(_2264_),
    .Y(_2275_),
    .A2(_2267_));
 sg13g2_nor2_2 _3148_ (.A(net1271),
    .B(_2275_),
    .Y(_2276_));
 sg13g2_nor2_1 _3149_ (.A(_0050_),
    .B(net1246),
    .Y(_2277_));
 sg13g2_a21oi_2 _3150_ (.B1(_2277_),
    .Y(_2278_),
    .A2(_2276_),
    .A1(net1246));
 sg13g2_or2_1 _3151_ (.X(_2279_),
    .B(_2278_),
    .A(\cpu_instance.accum[7] ));
 sg13g2_nand2_2 _3152_ (.Y(_2280_),
    .A(\cpu_instance.accum[7] ),
    .B(_2278_));
 sg13g2_nor3_1 _3153_ (.A(_0017_),
    .B(net1174),
    .C(_2272_),
    .Y(_2281_));
 sg13g2_a21oi_2 _3154_ (.B1(_1911_),
    .Y(_2282_),
    .A2(_2022_),
    .A1(_0013_));
 sg13g2_a22oi_1 _3155_ (.Y(_2283_),
    .B1(_2282_),
    .B2(\cpu_instance.inst[6] ),
    .A2(_2262_),
    .A1(net7));
 sg13g2_nand2b_1 _3156_ (.Y(_2284_),
    .B(_2267_),
    .A_N(_2283_));
 sg13g2_a21oi_1 _3157_ (.A1(_1954_),
    .A2(_2268_),
    .Y(_2285_),
    .B1(_2281_));
 sg13g2_a21o_2 _3158_ (.A2(_2285_),
    .A1(_2284_),
    .B1(net1271),
    .X(_2286_));
 sg13g2_mux2_2 _3159_ (.A0(_0051_),
    .A1(_2286_),
    .S(net1246),
    .X(_2287_));
 sg13g2_nor2b_2 _3160_ (.A(_2287_),
    .B_N(net1312),
    .Y(_2288_));
 sg13g2_nand2b_1 _3161_ (.Y(_2289_),
    .B(_2287_),
    .A_N(net1312));
 sg13g2_nor2b_2 _3162_ (.A(_2288_),
    .B_N(_2289_),
    .Y(_2290_));
 sg13g2_nor3_1 _3163_ (.A(_0018_),
    .B(net1174),
    .C(_2272_),
    .Y(_2291_));
 sg13g2_a22oi_1 _3164_ (.Y(_2292_),
    .B1(_2282_),
    .B2(\cpu_instance.inst[5] ),
    .A2(_2262_),
    .A1(net6));
 sg13g2_nand2b_1 _3165_ (.Y(_2293_),
    .B(_2267_),
    .A_N(_2292_));
 sg13g2_a21oi_1 _3166_ (.A1(_1953_),
    .A2(_2268_),
    .Y(_2294_),
    .B1(_2291_));
 sg13g2_a21oi_2 _3167_ (.B1(net1271),
    .Y(_2295_),
    .A2(_2294_),
    .A1(_2293_));
 sg13g2_nor2_1 _3168_ (.A(_1919_),
    .B(net1249),
    .Y(_2296_));
 sg13g2_a21o_2 _3169_ (.A2(net1105),
    .A1(net1249),
    .B1(_2296_),
    .X(_2297_));
 sg13g2_a21oi_2 _3170_ (.B1(_2296_),
    .Y(_2298_),
    .A2(net1105),
    .A1(net1249));
 sg13g2_nand2_1 _3171_ (.Y(_2299_),
    .A(_1953_),
    .B(_2297_));
 sg13g2_o21ai_1 _3172_ (.B1(_2299_),
    .Y(_2300_),
    .A1(\cpu_instance.accum[5] ),
    .A2(_2297_));
 sg13g2_nor2_1 _3173_ (.A(\cpu_instance.ram_data_out[4] ),
    .B(net1249),
    .Y(_2301_));
 sg13g2_a22oi_1 _3174_ (.Y(_2302_),
    .B1(_2282_),
    .B2(\cpu_instance.inst[4] ),
    .A2(_2262_),
    .A1(net5));
 sg13g2_nor2b_1 _3175_ (.A(_2302_),
    .B_N(_2267_),
    .Y(_2303_));
 sg13g2_nand2b_1 _3176_ (.Y(_2304_),
    .B(net1174),
    .A_N(net1313));
 sg13g2_o21ai_1 _3177_ (.B1(_2304_),
    .Y(_2305_),
    .A1(_0019_),
    .A2(_2273_));
 sg13g2_o21ai_1 _3178_ (.B1(net1265),
    .Y(_2306_),
    .A1(_2303_),
    .A2(_2305_));
 sg13g2_a21oi_2 _3179_ (.B1(_2301_),
    .Y(_2307_),
    .A2(_2306_),
    .A1(net1249));
 sg13g2_nor2b_2 _3180_ (.A(net1313),
    .B_N(_2307_),
    .Y(_2308_));
 sg13g2_nand2b_1 _3181_ (.Y(_2309_),
    .B(net1313),
    .A_N(_2307_));
 sg13g2_nor2b_2 _3182_ (.A(_2308_),
    .B_N(_2309_),
    .Y(_2310_));
 sg13g2_nor2_1 _3183_ (.A(_0020_),
    .B(_2273_),
    .Y(_2311_));
 sg13g2_nand2_1 _3184_ (.Y(_2312_),
    .A(net4),
    .B(_2262_));
 sg13g2_a21oi_1 _3185_ (.A1(\cpu_instance.inst[3] ),
    .A2(_2282_),
    .Y(_2313_),
    .B1(_2171_));
 sg13g2_a221oi_1 _3186_ (.B2(_2313_),
    .C1(_2122_),
    .B1(_2312_),
    .A1(_0036_),
    .Y(_2314_),
    .A2(_2171_));
 sg13g2_o21ai_1 _3187_ (.B1(net1265),
    .Y(_2315_),
    .A1(_2311_),
    .A2(_2314_));
 sg13g2_nor2_1 _3188_ (.A(net1239),
    .B(_2315_),
    .Y(_2316_));
 sg13g2_nor2_1 _3189_ (.A(_1921_),
    .B(net1249),
    .Y(_2317_));
 sg13g2_nand2_1 _3190_ (.Y(_2318_),
    .A(\cpu_instance.ram_data_out[3] ),
    .B(net1239));
 sg13g2_nor2_1 _3191_ (.A(_2316_),
    .B(_2317_),
    .Y(_2319_));
 sg13g2_o21ai_1 _3192_ (.B1(_2318_),
    .Y(_2320_),
    .A1(net1239),
    .A2(_2315_));
 sg13g2_nand2_1 _3193_ (.Y(_2321_),
    .A(_1952_),
    .B(net1066));
 sg13g2_xnor2_1 _3194_ (.Y(_2322_),
    .A(_1952_),
    .B(net1066));
 sg13g2_nand2_1 _3195_ (.Y(_2323_),
    .A(\cpu_instance.inst[2] ),
    .B(_2282_));
 sg13g2_o21ai_1 _3196_ (.B1(_2323_),
    .Y(_2324_),
    .A1(_0021_),
    .A2(_2269_));
 sg13g2_a221oi_1 _3197_ (.B2(net3),
    .C1(_2324_),
    .B1(_2262_),
    .A1(net1265),
    .Y(_2325_),
    .A2(_2122_));
 sg13g2_a21o_1 _3198_ (.A2(_2271_),
    .A1(_0021_),
    .B1(net1271),
    .X(_2326_));
 sg13g2_a221oi_1 _3199_ (.B2(_2266_),
    .C1(_2326_),
    .B1(_2325_),
    .A1(_0037_),
    .Y(_2327_),
    .A2(net1174));
 sg13g2_nor2_1 _3200_ (.A(_1922_),
    .B(net1251),
    .Y(_2328_));
 sg13g2_a21o_1 _3201_ (.A2(_2327_),
    .A1(net1251),
    .B1(_2328_),
    .X(_2329_));
 sg13g2_a21oi_1 _3202_ (.A1(net1251),
    .A2(_2327_),
    .Y(_2330_),
    .B1(_2328_));
 sg13g2_nor2_1 _3203_ (.A(_0037_),
    .B(net1098),
    .Y(_2331_));
 sg13g2_nand2b_1 _3204_ (.Y(_2332_),
    .B(net1103),
    .A_N(_0037_));
 sg13g2_nand2_1 _3205_ (.Y(_2333_),
    .A(_1935_),
    .B(net1098));
 sg13g2_nand2_1 _3206_ (.Y(_2334_),
    .A(_2332_),
    .B(_2333_));
 sg13g2_a21o_1 _3207_ (.A2(_2261_),
    .A1(_2260_),
    .B1(_1947_),
    .X(_2335_));
 sg13g2_a22oi_1 _3208_ (.Y(_2336_),
    .B1(_2282_),
    .B2(\cpu_instance.inst[1] ),
    .A2(_2270_),
    .A1(_1948_));
 sg13g2_nand4_1 _3209_ (.B(_2266_),
    .C(_2335_),
    .A(_2124_),
    .Y(_2337_),
    .D(_2336_));
 sg13g2_a221oi_1 _3210_ (.B2(_0022_),
    .C1(net1270),
    .B1(_2271_),
    .A1(_0038_),
    .Y(_2338_),
    .A2(net1174));
 sg13g2_nand2_2 _3211_ (.Y(_2339_),
    .A(_2337_),
    .B(_2338_));
 sg13g2_nand3_1 _3212_ (.B(_2337_),
    .C(_2338_),
    .A(net1251),
    .Y(_2340_));
 sg13g2_nand2_2 _3213_ (.Y(_2341_),
    .A(\cpu_instance.ram_data_out[1] ),
    .B(net1239));
 sg13g2_nand2_1 _3214_ (.Y(_2342_),
    .A(_2340_),
    .B(_2341_));
 sg13g2_and2_1 _3215_ (.A(_2340_),
    .B(_2341_),
    .X(_2343_));
 sg13g2_nand2_1 _3216_ (.Y(_2344_),
    .A(_1949_),
    .B(net1086));
 sg13g2_and2_1 _3217_ (.A(_0023_),
    .B(net1223),
    .X(_2345_));
 sg13g2_nor4_1 _3218_ (.A(_1909_),
    .B(_0013_),
    .C(net1270),
    .D(_2012_),
    .Y(_2346_));
 sg13g2_nor3_1 _3219_ (.A(net1302),
    .B(_0023_),
    .C(_2173_),
    .Y(_2347_));
 sg13g2_a221oi_1 _3220_ (.B2(\cpu_instance.inst[0] ),
    .C1(_2347_),
    .B1(_2282_),
    .A1(net1),
    .Y(_2348_),
    .A2(_2259_));
 sg13g2_nand2b_1 _3221_ (.Y(_2349_),
    .B(net1299),
    .A_N(net1));
 sg13g2_nand4_1 _3222_ (.B(_2011_),
    .C(_2026_),
    .A(net1265),
    .Y(_2350_),
    .D(_2349_));
 sg13g2_o21ai_1 _3223_ (.B1(_2350_),
    .Y(_2351_),
    .A1(_2346_),
    .A2(_2348_));
 sg13g2_a221oi_1 _3224_ (.B2(_0023_),
    .C1(_2002_),
    .B1(_2265_),
    .A1(_2060_),
    .Y(_2352_),
    .A2(_2067_));
 sg13g2_a221oi_1 _3225_ (.B2(_2352_),
    .C1(net1223),
    .B1(_2351_),
    .A1(_1950_),
    .Y(_2353_),
    .A2(_2171_));
 sg13g2_nand2_2 _3226_ (.Y(_2354_),
    .A(_0052_),
    .B(net1240));
 sg13g2_o21ai_1 _3227_ (.B1(net1251),
    .Y(_2355_),
    .A1(_2345_),
    .A2(_2353_));
 sg13g2_nand2_1 _3228_ (.Y(_2356_),
    .A(_2354_),
    .B(_2355_));
 sg13g2_and2_2 _3229_ (.A(_2354_),
    .B(_2355_),
    .X(_2357_));
 sg13g2_nand3_1 _3230_ (.B(_2354_),
    .C(_2355_),
    .A(_0039_),
    .Y(_2358_));
 sg13g2_a21oi_2 _3231_ (.B1(_0038_),
    .Y(_2359_),
    .A2(_2341_),
    .A1(_2340_));
 sg13g2_and3_1 _3232_ (.X(_2360_),
    .A(_1936_),
    .B(_2340_),
    .C(_2341_));
 sg13g2_o21ai_1 _3233_ (.B1(_2358_),
    .Y(_2361_),
    .A1(_2359_),
    .A2(_2360_));
 sg13g2_nand2_1 _3234_ (.Y(_2362_),
    .A(_2344_),
    .B(_2361_));
 sg13g2_a22oi_1 _3235_ (.Y(_2363_),
    .B1(_2344_),
    .B2(_2361_),
    .A2(_2333_),
    .A1(_2332_));
 sg13g2_nand2_1 _3236_ (.Y(_2364_),
    .A(_2334_),
    .B(_2362_));
 sg13g2_nor2_1 _3237_ (.A(_0037_),
    .B(net1103),
    .Y(_2365_));
 sg13g2_o21ai_1 _3238_ (.B1(_2322_),
    .Y(_2366_),
    .A1(_2363_),
    .A2(_2365_));
 sg13g2_nand2_1 _3239_ (.Y(_2367_),
    .A(_1952_),
    .B(net1059));
 sg13g2_a21oi_1 _3240_ (.A1(_2366_),
    .A2(_2367_),
    .Y(_2368_),
    .B1(_2310_));
 sg13g2_nor2_1 _3241_ (.A(net1313),
    .B(_2307_),
    .Y(_2369_));
 sg13g2_o21ai_1 _3242_ (.B1(_2300_),
    .Y(_2370_),
    .A1(_2368_),
    .A2(_2369_));
 sg13g2_nand2_1 _3243_ (.Y(_2371_),
    .A(_1953_),
    .B(_2298_));
 sg13g2_a21oi_2 _3244_ (.B1(_2290_),
    .Y(_2372_),
    .A2(_2371_),
    .A1(_2370_));
 sg13g2_and2_1 _3245_ (.A(net1312),
    .B(_2287_),
    .X(_2373_));
 sg13g2_nor2_1 _3246_ (.A(_2372_),
    .B(_2373_),
    .Y(_2374_));
 sg13g2_o21ai_1 _3247_ (.B1(_2279_),
    .Y(_2375_),
    .A1(_2372_),
    .A2(_2373_));
 sg13g2_a21oi_2 _3248_ (.B1(_2258_),
    .Y(_2376_),
    .A2(_2375_),
    .A1(_2280_));
 sg13g2_nor2_1 _3249_ (.A(_2255_),
    .B(_2376_),
    .Y(_2377_));
 sg13g2_o21ai_1 _3250_ (.B1(_2245_),
    .Y(_2378_),
    .A1(_2255_),
    .A2(_2376_));
 sg13g2_a21oi_2 _3251_ (.B1(_2236_),
    .Y(_2379_),
    .A2(_2378_),
    .A1(_2246_));
 sg13g2_a21oi_1 _3252_ (.A1(net1307),
    .A2(_2232_),
    .Y(_2380_),
    .B1(_2379_));
 sg13g2_a221oi_1 _3253_ (.B2(net1307),
    .C1(_2379_),
    .B1(_2232_),
    .A1(net1306),
    .Y(_2381_),
    .A2(_2225_));
 sg13g2_nor2_1 _3254_ (.A(_2226_),
    .B(_2381_),
    .Y(_2382_));
 sg13g2_nor3_1 _3255_ (.A(_2217_),
    .B(_2226_),
    .C(_2381_),
    .Y(_2383_));
 sg13g2_nor3_1 _3256_ (.A(_1928_),
    .B(_2213_),
    .C(_2214_),
    .Y(_2384_));
 sg13g2_nor2_1 _3257_ (.A(_2383_),
    .B(_2384_),
    .Y(_2385_));
 sg13g2_o21ai_1 _3258_ (.B1(_2206_),
    .Y(_2386_),
    .A1(_2383_),
    .A2(_2384_));
 sg13g2_a21oi_2 _3259_ (.B1(_2198_),
    .Y(_2387_),
    .A2(_2386_),
    .A1(_2207_));
 sg13g2_nor3_1 _3260_ (.A(_1926_),
    .B(_2193_),
    .C(_2194_),
    .Y(_2388_));
 sg13g2_or3_1 _3261_ (.A(_2187_),
    .B(_2387_),
    .C(_2388_),
    .X(_2389_));
 sg13g2_o21ai_1 _3262_ (.B1(_2187_),
    .Y(_2390_),
    .A1(_2387_),
    .A2(_2388_));
 sg13g2_and2_1 _3263_ (.A(net1289),
    .B(_2034_),
    .X(_2391_));
 sg13g2_nand2_2 _3264_ (.Y(_2392_),
    .A(net1289),
    .B(_2034_));
 sg13g2_nand3_1 _3265_ (.B(_2390_),
    .C(net1152),
    .A(_2389_),
    .Y(_2393_));
 sg13g2_nor2_1 _3266_ (.A(_0024_),
    .B(net1205),
    .Y(_2394_));
 sg13g2_and2_2 _3267_ (.A(net1289),
    .B(_2032_),
    .X(_2395_));
 sg13g2_a221oi_1 _3268_ (.B2(net1171),
    .C1(net1203),
    .B1(_2188_),
    .A1(_0024_),
    .Y(_2396_),
    .A2(net1210));
 sg13g2_nor2_2 _3269_ (.A(net1209),
    .B(_2307_),
    .Y(_2397_));
 sg13g2_or2_2 _3270_ (.X(_2398_),
    .B(_2307_),
    .A(net1208));
 sg13g2_a221oi_1 _3271_ (.B2(_2243_),
    .C1(_2231_),
    .B1(_2242_),
    .A1(net1243),
    .Y(_2399_),
    .A2(_2230_));
 sg13g2_nor4_1 _3272_ (.A(_2193_),
    .B(_2194_),
    .C(_2252_),
    .D(_2253_),
    .Y(_2400_));
 sg13g2_nor4_1 _3273_ (.A(_2213_),
    .B(_2214_),
    .C(_2223_),
    .D(_2224_),
    .Y(_2401_));
 sg13g2_a221oi_1 _3274_ (.B2(net1244),
    .C1(_2204_),
    .B1(_2202_),
    .A1(_2181_),
    .Y(_2402_),
    .A2(_2182_));
 sg13g2_and4_1 _3275_ (.A(_2399_),
    .B(_2400_),
    .C(_2401_),
    .D(_2402_),
    .X(_2403_));
 sg13g2_and4_2 _3276_ (.A(_2278_),
    .B(_2287_),
    .C(_2298_),
    .D(_2403_),
    .X(_2404_));
 sg13g2_nand2_2 _3277_ (.Y(_2405_),
    .A(_1960_),
    .B(net1054));
 sg13g2_nand3_1 _3278_ (.B(net1077),
    .C(net1053),
    .A(_1963_),
    .Y(_2406_));
 sg13g2_nand2_1 _3279_ (.Y(_2407_),
    .A(_1961_),
    .B(net1053));
 sg13g2_o21ai_1 _3280_ (.B1(_2406_),
    .Y(_2408_),
    .A1(net1077),
    .A2(_2407_));
 sg13g2_nor2_2 _3281_ (.A(net1109),
    .B(net1065),
    .Y(_2409_));
 sg13g2_nand2_2 _3282_ (.Y(_2410_),
    .A(_2018_),
    .B(net1059));
 sg13g2_nand2_1 _3283_ (.Y(_2411_),
    .A(_1964_),
    .B(net1053));
 sg13g2_nand3_1 _3284_ (.B(net1073),
    .C(net1053),
    .A(_1964_),
    .Y(_2412_));
 sg13g2_nand2_1 _3285_ (.Y(_2413_),
    .A(_1966_),
    .B(net1053));
 sg13g2_nand3_1 _3286_ (.B(net1077),
    .C(net1053),
    .A(_1966_),
    .Y(_2414_));
 sg13g2_and2_1 _3287_ (.A(_2412_),
    .B(_2414_),
    .X(_2415_));
 sg13g2_and2_1 _3288_ (.A(_1969_),
    .B(net1054),
    .X(_2416_));
 sg13g2_nand2_1 _3289_ (.Y(_2417_),
    .A(net1077),
    .B(_2416_));
 sg13g2_nand3_1 _3290_ (.B(net1073),
    .C(net1054),
    .A(_1967_),
    .Y(_2418_));
 sg13g2_nand3_1 _3291_ (.B(_2417_),
    .C(_2418_),
    .A(net1083),
    .Y(_2419_));
 sg13g2_a21oi_1 _3292_ (.A1(net1088),
    .A2(_2415_),
    .Y(_2420_),
    .B1(net1101));
 sg13g2_a21oi_1 _3293_ (.A1(_1957_),
    .A2(net1055),
    .Y(_2421_),
    .B1(net1077));
 sg13g2_a21oi_1 _3294_ (.A1(net1078),
    .A2(_2405_),
    .Y(_2422_),
    .B1(_2421_));
 sg13g2_mux2_1 _3295_ (.A0(_2408_),
    .A1(_2422_),
    .S(net1088),
    .X(_2423_));
 sg13g2_a221oi_1 _3296_ (.B2(net1101),
    .C1(_2410_),
    .B1(_2423_),
    .A1(_2419_),
    .Y(_2424_),
    .A2(_2420_));
 sg13g2_nor2_1 _3297_ (.A(_2398_),
    .B(_2424_),
    .Y(_2425_));
 sg13g2_a21oi_1 _3298_ (.A1(_1952_),
    .A2(net1057),
    .Y(_2426_),
    .B1(net1075));
 sg13g2_nand2b_1 _3299_ (.Y(_2427_),
    .B(net1056),
    .A_N(_0037_));
 sg13g2_a21oi_1 _3300_ (.A1(net1076),
    .A2(_2427_),
    .Y(_2428_),
    .B1(_2426_));
 sg13g2_o21ai_1 _3301_ (.B1(_2358_),
    .Y(_2429_),
    .A1(_1949_),
    .A2(net1076));
 sg13g2_nor2b_1 _3302_ (.A(_2429_),
    .B_N(net1057),
    .Y(_2430_));
 sg13g2_and2_1 _3303_ (.A(net1091),
    .B(_2430_),
    .X(_2431_));
 sg13g2_a21oi_1 _3304_ (.A1(net1085),
    .A2(_2428_),
    .Y(_2432_),
    .B1(_2431_));
 sg13g2_nor3_1 _3305_ (.A(net1110),
    .B(net1096),
    .C(_2432_),
    .Y(_2433_));
 sg13g2_nor2_2 _3306_ (.A(net1110),
    .B(net1102),
    .Y(_2434_));
 sg13g2_nor2_1 _3307_ (.A(net1313),
    .B(net1080),
    .Y(_2435_));
 sg13g2_a21oi_2 _3308_ (.B1(_2435_),
    .Y(_2436_),
    .A2(net1080),
    .A1(_1953_));
 sg13g2_nand2b_1 _3309_ (.Y(_2437_),
    .B(_2404_),
    .A_N(_2436_));
 sg13g2_nand2_2 _3310_ (.Y(_2438_),
    .A(_1956_),
    .B(net1055));
 sg13g2_nand2_2 _3311_ (.Y(_2439_),
    .A(_2015_),
    .B(net1059));
 sg13g2_nor2_1 _3312_ (.A(net1090),
    .B(net1074),
    .Y(_2440_));
 sg13g2_nand2_2 _3313_ (.Y(_2441_),
    .A(net1082),
    .B(net1078));
 sg13g2_nor2_2 _3314_ (.A(net1101),
    .B(net1063),
    .Y(_2442_));
 sg13g2_nand2_1 _3315_ (.Y(_2443_),
    .A(_2416_),
    .B(_2442_));
 sg13g2_a21oi_1 _3316_ (.A1(_1954_),
    .A2(net1057),
    .Y(_2444_),
    .B1(net1080));
 sg13g2_a21oi_2 _3317_ (.B1(_2444_),
    .Y(_2445_),
    .A2(_2438_),
    .A1(net1080));
 sg13g2_nor2_1 _3318_ (.A(net1091),
    .B(_2445_),
    .Y(_2446_));
 sg13g2_a21oi_2 _3319_ (.B1(_2446_),
    .Y(_2447_),
    .A2(_2437_),
    .A1(net1091));
 sg13g2_a21oi_2 _3320_ (.B1(_2433_),
    .Y(_2448_),
    .A2(_2447_),
    .A1(_2434_));
 sg13g2_o21ai_1 _3321_ (.B1(_2448_),
    .Y(_2449_),
    .A1(_2439_),
    .A2(_2443_));
 sg13g2_o21ai_1 _3322_ (.B1(_2425_),
    .Y(_2450_),
    .A1(_2409_),
    .A2(_2449_));
 sg13g2_and2_1 _3323_ (.A(_1907_),
    .B(_2032_),
    .X(_2451_));
 sg13g2_nand2_2 _3324_ (.Y(_2452_),
    .A(net1281),
    .B(_2032_));
 sg13g2_a221oi_1 _3325_ (.B2(_2450_),
    .C1(net1169),
    .B1(_2396_),
    .A1(net1204),
    .Y(_2453_),
    .A2(_2186_));
 sg13g2_nor2_1 _3326_ (.A(_2185_),
    .B(_2452_),
    .Y(_2454_));
 sg13g2_nor3_1 _3327_ (.A(_2394_),
    .B(_2453_),
    .C(_2454_),
    .Y(_2455_));
 sg13g2_a21o_2 _3328_ (.A2(_2455_),
    .A1(_2393_),
    .B1(net1154),
    .X(_2456_));
 sg13g2_nand2_1 _3329_ (.Y(_2457_),
    .A(_1927_),
    .B(_2205_));
 sg13g2_nor2_1 _3330_ (.A(_1927_),
    .B(_2205_),
    .Y(_2458_));
 sg13g2_nor3_2 _3331_ (.A(net1306),
    .B(_2223_),
    .C(_2224_),
    .Y(_2459_));
 sg13g2_nor2_2 _3332_ (.A(_1929_),
    .B(_2225_),
    .Y(_2460_));
 sg13g2_a21oi_2 _3333_ (.B1(net1309),
    .Y(_2461_),
    .A2(_2243_),
    .A1(_2242_));
 sg13g2_nor2_2 _3334_ (.A(_1930_),
    .B(_2244_),
    .Y(_2462_));
 sg13g2_nor2_1 _3335_ (.A(_1931_),
    .B(_2278_),
    .Y(_2463_));
 sg13g2_inv_1 _3336_ (.Y(_2464_),
    .A(_2463_));
 sg13g2_nand2_2 _3337_ (.Y(_2465_),
    .A(_1931_),
    .B(_2278_));
 sg13g2_nand2_1 _3338_ (.Y(_2466_),
    .A(_0034_),
    .B(_2298_));
 sg13g2_and3_1 _3339_ (.X(_2467_),
    .A(\cpu_instance.accum[0] ),
    .B(_2354_),
    .C(_2355_));
 sg13g2_nand3_1 _3340_ (.B(_2340_),
    .C(_2341_),
    .A(_0038_),
    .Y(_2468_));
 sg13g2_nor2b_1 _3341_ (.A(_2359_),
    .B_N(_2468_),
    .Y(_2469_));
 sg13g2_inv_1 _3342_ (.Y(_2470_),
    .A(_2469_));
 sg13g2_a21o_1 _3343_ (.A2(_2468_),
    .A1(_2467_),
    .B1(_2359_),
    .X(_2471_));
 sg13g2_nand2_2 _3344_ (.Y(_2472_),
    .A(_0037_),
    .B(net1098));
 sg13g2_nand2_1 _3345_ (.Y(_2473_),
    .A(_2332_),
    .B(_2472_));
 sg13g2_a21oi_1 _3346_ (.A1(_2471_),
    .A2(_2472_),
    .Y(_2474_),
    .B1(_2331_));
 sg13g2_o21ai_1 _3347_ (.B1(_2321_),
    .Y(_2475_),
    .A1(_2322_),
    .A2(_2474_));
 sg13g2_a21oi_1 _3348_ (.A1(_2310_),
    .A2(_2475_),
    .Y(_2476_),
    .B1(_2308_));
 sg13g2_a221oi_1 _3349_ (.B2(_2475_),
    .C1(_2308_),
    .B1(_2310_),
    .A1(_1953_),
    .Y(_2477_),
    .A2(_2297_));
 sg13g2_a21o_1 _3350_ (.A2(_2298_),
    .A1(_0034_),
    .B1(_2477_),
    .X(_2478_));
 sg13g2_nand3b_1 _3351_ (.B(_2290_),
    .C(_2466_),
    .Y(_2479_),
    .A_N(_2477_));
 sg13g2_nand2b_1 _3352_ (.Y(_2480_),
    .B(_2479_),
    .A_N(_2288_));
 sg13g2_nand3b_1 _3353_ (.B(_2464_),
    .C(_2479_),
    .Y(_2481_),
    .A_N(_2288_));
 sg13g2_nand2_1 _3354_ (.Y(_2482_),
    .A(_2465_),
    .B(_2481_));
 sg13g2_nand3_1 _3355_ (.B(_2465_),
    .C(_2481_),
    .A(_2258_),
    .Y(_2483_));
 sg13g2_nand2_1 _3356_ (.Y(_2484_),
    .A(_2256_),
    .B(_2483_));
 sg13g2_a21oi_1 _3357_ (.A1(_2256_),
    .A2(_2483_),
    .Y(_2485_),
    .B1(_2461_));
 sg13g2_nor2_1 _3358_ (.A(_2462_),
    .B(_2485_),
    .Y(_2486_));
 sg13g2_o21ai_1 _3359_ (.B1(_2236_),
    .Y(_2487_),
    .A1(_2462_),
    .A2(_2485_));
 sg13g2_nand2_1 _3360_ (.Y(_2488_),
    .A(_2233_),
    .B(_2487_));
 sg13g2_a21oi_1 _3361_ (.A1(_2233_),
    .A2(_2487_),
    .Y(_2489_),
    .B1(_2459_));
 sg13g2_nor2_1 _3362_ (.A(_2460_),
    .B(_2489_),
    .Y(_2490_));
 sg13g2_o21ai_1 _3363_ (.B1(_2215_),
    .Y(_2491_),
    .A1(_2218_),
    .A2(_2490_));
 sg13g2_or2_1 _3364_ (.X(_2492_),
    .B(_2491_),
    .A(_2458_));
 sg13g2_nand3_1 _3365_ (.B(_2457_),
    .C(_2492_),
    .A(_2198_),
    .Y(_2493_));
 sg13g2_nand2b_1 _3366_ (.Y(_2494_),
    .B(_2493_),
    .A_N(_2196_));
 sg13g2_xnor2_1 _3367_ (.Y(_2495_),
    .A(_2187_),
    .B(_2494_));
 sg13g2_nand2_2 _3368_ (.Y(_2496_),
    .A(net1154),
    .B(_2495_));
 sg13g2_nand2_1 _3369_ (.Y(_2497_),
    .A(_2456_),
    .B(_2496_));
 sg13g2_a21o_1 _3370_ (.A2(_2492_),
    .A1(_2457_),
    .B1(_2198_),
    .X(_2498_));
 sg13g2_nand2_1 _3371_ (.Y(_2499_),
    .A(_2493_),
    .B(_2498_));
 sg13g2_nand3_1 _3372_ (.B(_2207_),
    .C(_2386_),
    .A(_2198_),
    .Y(_2500_));
 sg13g2_nand3b_1 _3373_ (.B(net1152),
    .C(_2500_),
    .Y(_2501_),
    .A_N(_2387_));
 sg13g2_a221oi_1 _3374_ (.B2(net1171),
    .C1(net1202),
    .B1(_2198_),
    .A1(_0025_),
    .Y(_2502_),
    .A2(net1210));
 sg13g2_nand3_1 _3375_ (.B(net1077),
    .C(net1055),
    .A(_1957_),
    .Y(_2503_));
 sg13g2_o21ai_1 _3376_ (.B1(_2503_),
    .Y(_2504_),
    .A1(net1079),
    .A2(_2438_));
 sg13g2_a21oi_1 _3377_ (.A1(_1961_),
    .A2(net1053),
    .Y(_2505_),
    .B1(net1073));
 sg13g2_a21oi_1 _3378_ (.A1(net1073),
    .A2(_2405_),
    .Y(_2506_),
    .B1(_2505_));
 sg13g2_nor2_1 _3379_ (.A(net1088),
    .B(_2506_),
    .Y(_2507_));
 sg13g2_nor2_1 _3380_ (.A(net1084),
    .B(_2504_),
    .Y(_2508_));
 sg13g2_nor3_1 _3381_ (.A(net1093),
    .B(_2507_),
    .C(_2508_),
    .Y(_2509_));
 sg13g2_a21oi_1 _3382_ (.A1(_1963_),
    .A2(net1053),
    .Y(_2510_),
    .B1(net1077));
 sg13g2_a21oi_1 _3383_ (.A1(net1077),
    .A2(_2411_),
    .Y(_2511_),
    .B1(_2510_));
 sg13g2_inv_1 _3384_ (.Y(_2512_),
    .A(_2511_));
 sg13g2_nand2_1 _3385_ (.Y(_2513_),
    .A(net1073),
    .B(_2413_));
 sg13g2_a21oi_1 _3386_ (.A1(_1967_),
    .A2(net1054),
    .Y(_2514_),
    .B1(net1073));
 sg13g2_nor2_1 _3387_ (.A(net1088),
    .B(_2514_),
    .Y(_2515_));
 sg13g2_a22oi_1 _3388_ (.Y(_2516_),
    .B1(_2513_),
    .B2(_2515_),
    .A2(_2511_),
    .A1(net1088));
 sg13g2_o21ai_1 _3389_ (.B1(_2409_),
    .Y(_2517_),
    .A1(net1101),
    .A2(_2516_));
 sg13g2_o21ai_1 _3390_ (.B1(_2397_),
    .Y(_2518_),
    .A1(_2509_),
    .A2(_2517_));
 sg13g2_nand3_1 _3391_ (.B(net1075),
    .C(net1056),
    .A(_1952_),
    .Y(_2519_));
 sg13g2_nand2b_1 _3392_ (.Y(_2520_),
    .B(net1056),
    .A_N(_0035_));
 sg13g2_nand3b_1 _3393_ (.B(net1080),
    .C(net1056),
    .Y(_2521_),
    .A_N(net1313));
 sg13g2_a21oi_1 _3394_ (.A1(_2519_),
    .A2(_2521_),
    .Y(_2522_),
    .B1(net1085));
 sg13g2_nand3_1 _3395_ (.B(net1075),
    .C(net1056),
    .A(_1953_),
    .Y(_2523_));
 sg13g2_nand3_1 _3396_ (.B(net1080),
    .C(net1057),
    .A(_1954_),
    .Y(_2524_));
 sg13g2_nand2_2 _3397_ (.Y(_2525_),
    .A(_2523_),
    .B(_2524_));
 sg13g2_a21o_1 _3398_ (.A2(_2525_),
    .A1(net1085),
    .B1(_2522_),
    .X(_2526_));
 sg13g2_and2_2 _3399_ (.A(_1950_),
    .B(net1057),
    .X(_2527_));
 sg13g2_nand2_1 _3400_ (.Y(_2528_),
    .A(net1081),
    .B(_2527_));
 sg13g2_nand3_1 _3401_ (.B(net1075),
    .C(net1057),
    .A(_1949_),
    .Y(_2529_));
 sg13g2_nand3b_1 _3402_ (.B(net1081),
    .C(net1056),
    .Y(_2530_),
    .A_N(_0037_));
 sg13g2_nand2_1 _3403_ (.Y(_2531_),
    .A(_2529_),
    .B(_2530_));
 sg13g2_nand2_1 _3404_ (.Y(_2532_),
    .A(net1086),
    .B(_2531_));
 sg13g2_o21ai_1 _3405_ (.B1(_2532_),
    .Y(_2533_),
    .A1(net1085),
    .A2(_2528_));
 sg13g2_mux2_1 _3406_ (.A0(_2526_),
    .A1(_2533_),
    .S(net1102),
    .X(_2534_));
 sg13g2_nor2_1 _3407_ (.A(net1078),
    .B(_2416_),
    .Y(_0190_));
 sg13g2_nand2b_2 _3408_ (.Y(_0191_),
    .B(_2515_),
    .A_N(_0190_));
 sg13g2_nand2b_1 _3409_ (.Y(_0192_),
    .B(net1094),
    .A_N(_0191_));
 sg13g2_o21ai_1 _3410_ (.B1(_2410_),
    .Y(_0193_),
    .A1(_2439_),
    .A2(_0192_));
 sg13g2_a21oi_1 _3411_ (.A1(_2018_),
    .A2(_2534_),
    .Y(_0194_),
    .B1(_0193_));
 sg13g2_or2_1 _3412_ (.X(_0195_),
    .B(_0194_),
    .A(_2518_));
 sg13g2_a22oi_1 _3413_ (.Y(_0196_),
    .B1(_2502_),
    .B2(_0195_),
    .A2(_2197_),
    .A1(net1203));
 sg13g2_a21oi_1 _3414_ (.A1(_2196_),
    .A2(net1169),
    .Y(_0197_),
    .B1(_0196_));
 sg13g2_o21ai_1 _3415_ (.B1(_0197_),
    .Y(_0198_),
    .A1(_0025_),
    .A2(net1205));
 sg13g2_nor2_1 _3416_ (.A(net1154),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_a22oi_1 _3417_ (.Y(_0200_),
    .B1(_2501_),
    .B2(_0199_),
    .A2(_2499_),
    .A1(net1154));
 sg13g2_and2_1 _3418_ (.A(_2206_),
    .B(_2207_),
    .X(_0201_));
 sg13g2_inv_1 _3419_ (.Y(_0202_),
    .A(_0201_));
 sg13g2_a221oi_1 _3420_ (.B2(_0202_),
    .C1(net1202),
    .B1(net1171),
    .A1(_0026_),
    .Y(_0203_),
    .A2(net1210));
 sg13g2_nand2_1 _3421_ (.Y(_0204_),
    .A(net1087),
    .B(_2430_));
 sg13g2_nor3_1 _3422_ (.A(net1110),
    .B(net1096),
    .C(_0204_),
    .Y(_0205_));
 sg13g2_nand2_1 _3423_ (.Y(_0206_),
    .A(net1091),
    .B(_2428_));
 sg13g2_o21ai_1 _3424_ (.B1(_0206_),
    .Y(_0207_),
    .A1(net1091),
    .A2(_2437_));
 sg13g2_a21oi_2 _3425_ (.B1(_0205_),
    .Y(_0208_),
    .A2(_0207_),
    .A1(_2434_));
 sg13g2_nand2_1 _3426_ (.Y(_0209_),
    .A(_2414_),
    .B(_2418_));
 sg13g2_nor2_1 _3427_ (.A(net1088),
    .B(_0209_),
    .Y(_0210_));
 sg13g2_a21oi_2 _3428_ (.B1(_0210_),
    .Y(_0211_),
    .A2(_2417_),
    .A1(net1088));
 sg13g2_nand3_1 _3429_ (.B(net1093),
    .C(_0211_),
    .A(net1111),
    .Y(_0212_));
 sg13g2_a21o_1 _3430_ (.A2(_0212_),
    .A1(net1109),
    .B1(net1065),
    .X(_0213_));
 sg13g2_mux2_1 _3431_ (.A0(_2422_),
    .A1(_2445_),
    .S(net1090),
    .X(_0214_));
 sg13g2_a21oi_1 _3432_ (.A1(net1089),
    .A2(_2408_),
    .Y(_0215_),
    .B1(net1101));
 sg13g2_o21ai_1 _3433_ (.B1(_0215_),
    .Y(_0216_),
    .A1(net1088),
    .A2(_2415_));
 sg13g2_o21ai_1 _3434_ (.B1(_0216_),
    .Y(_0217_),
    .A1(net1093),
    .A2(_0214_));
 sg13g2_a221oi_1 _3435_ (.B2(_2409_),
    .C1(_2398_),
    .B1(_0217_),
    .A1(_0208_),
    .Y(_0218_),
    .A2(_0213_));
 sg13g2_nand2b_1 _3436_ (.Y(_0219_),
    .B(_0203_),
    .A_N(_0218_));
 sg13g2_nand3_1 _3437_ (.B(net1203),
    .C(_2205_),
    .A(_1927_),
    .Y(_0220_));
 sg13g2_nor2_1 _3438_ (.A(_0026_),
    .B(net1205),
    .Y(_0221_));
 sg13g2_xnor2_1 _3439_ (.Y(_0222_),
    .A(_2385_),
    .B(_0201_));
 sg13g2_a221oi_1 _3440_ (.B2(net1152),
    .C1(_0221_),
    .B1(_0222_),
    .A1(net1169),
    .Y(_0223_),
    .A2(_2458_));
 sg13g2_a21oi_1 _3441_ (.A1(_0219_),
    .A2(_0220_),
    .Y(_0224_),
    .B1(net1154));
 sg13g2_xnor2_1 _3442_ (.Y(_0225_),
    .A(_2491_),
    .B(_0202_));
 sg13g2_a22oi_1 _3443_ (.Y(_0226_),
    .B1(_0225_),
    .B2(net1154),
    .A2(_0224_),
    .A1(_0223_));
 sg13g2_xnor2_1 _3444_ (.Y(_0227_),
    .A(_2217_),
    .B(_2490_));
 sg13g2_a21oi_1 _3445_ (.A1(net1083),
    .A2(_2512_),
    .Y(_0228_),
    .B1(net1101));
 sg13g2_o21ai_1 _3446_ (.B1(_0228_),
    .Y(_0229_),
    .A1(net1083),
    .A2(_2506_));
 sg13g2_mux2_1 _3447_ (.A0(_2504_),
    .A1(_2525_),
    .S(net1090),
    .X(_0230_));
 sg13g2_a21oi_1 _3448_ (.A1(net1099),
    .A2(_0230_),
    .Y(_0231_),
    .B1(_2410_));
 sg13g2_a21oi_1 _3449_ (.A1(_0229_),
    .A2(_0231_),
    .Y(_0232_),
    .B1(_2398_));
 sg13g2_nor3_2 _3450_ (.A(net1083),
    .B(_2514_),
    .C(_0190_),
    .Y(_0233_));
 sg13g2_mux2_1 _3451_ (.A0(_2411_),
    .A1(_2413_),
    .S(net1073),
    .X(_0234_));
 sg13g2_nor2_1 _3452_ (.A(net1089),
    .B(_0234_),
    .Y(_0235_));
 sg13g2_nor2_1 _3453_ (.A(_0233_),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_o21ai_1 _3454_ (.B1(net1094),
    .Y(_0237_),
    .A1(_0233_),
    .A2(_0235_));
 sg13g2_a21oi_1 _3455_ (.A1(_2519_),
    .A2(_2521_),
    .Y(_0238_),
    .B1(net1092));
 sg13g2_a21oi_2 _3456_ (.B1(_0238_),
    .Y(_0239_),
    .A2(_2531_),
    .A1(net1091));
 sg13g2_nor2_1 _3457_ (.A(net1110),
    .B(_2441_),
    .Y(_0240_));
 sg13g2_a21oi_1 _3458_ (.A1(_2527_),
    .A2(_0240_),
    .Y(_0241_),
    .B1(_2434_));
 sg13g2_a21o_1 _3459_ (.A2(_0239_),
    .A1(net1096),
    .B1(_0241_),
    .X(_0242_));
 sg13g2_and2_1 _3460_ (.A(_2410_),
    .B(_0242_),
    .X(_0243_));
 sg13g2_o21ai_1 _3461_ (.B1(_0243_),
    .Y(_0244_),
    .A1(_2439_),
    .A2(_0237_));
 sg13g2_nor2_2 _3462_ (.A(net1095),
    .B(_2440_),
    .Y(_0245_));
 sg13g2_a221oi_1 _3463_ (.B2(_2216_),
    .C1(net1155),
    .B1(net1203),
    .A1(_1964_),
    .Y(_0246_),
    .A2(net1207));
 sg13g2_o21ai_1 _3464_ (.B1(_0246_),
    .Y(_0247_),
    .A1(_2215_),
    .A2(_2452_));
 sg13g2_a21o_1 _3465_ (.A2(net1171),
    .A1(_2217_),
    .B1(_0247_),
    .X(_0248_));
 sg13g2_a221oi_1 _3466_ (.B2(_0244_),
    .C1(_0248_),
    .B1(_0232_),
    .A1(_0027_),
    .Y(_0249_),
    .A2(net1210));
 sg13g2_o21ai_1 _3467_ (.B1(net1152),
    .Y(_0250_),
    .A1(_2218_),
    .A2(_2382_));
 sg13g2_o21ai_1 _3468_ (.B1(_0249_),
    .Y(_0251_),
    .A1(_2383_),
    .A2(_0250_));
 sg13g2_o21ai_1 _3469_ (.B1(_0251_),
    .Y(_0252_),
    .A1(net1153),
    .A2(_0227_));
 sg13g2_nor2_2 _3470_ (.A(_2459_),
    .B(_2460_),
    .Y(_0253_));
 sg13g2_xnor2_1 _3471_ (.Y(_0254_),
    .A(_2380_),
    .B(_0253_));
 sg13g2_nand2_1 _3472_ (.Y(_0255_),
    .A(_2406_),
    .B(_2412_));
 sg13g2_mux2_1 _3473_ (.A0(_0209_),
    .A1(_0255_),
    .S(net1082),
    .X(_0256_));
 sg13g2_a21oi_1 _3474_ (.A1(_2416_),
    .A2(_2440_),
    .Y(_0257_),
    .B1(net1093));
 sg13g2_o21ai_1 _3475_ (.B1(net1111),
    .Y(_0258_),
    .A1(net1099),
    .A2(_0256_));
 sg13g2_o21ai_1 _3476_ (.B1(net1109),
    .Y(_0259_),
    .A1(_0257_),
    .A2(_0258_));
 sg13g2_nand2b_1 _3477_ (.Y(_0260_),
    .B(_2434_),
    .A_N(_2432_));
 sg13g2_nand2_1 _3478_ (.Y(_0261_),
    .A(net1094),
    .B(_2423_));
 sg13g2_a21oi_1 _3479_ (.A1(net1100),
    .A2(_2447_),
    .Y(_0262_),
    .B1(_2410_));
 sg13g2_a221oi_1 _3480_ (.B2(_0262_),
    .C1(_2398_),
    .B1(_0261_),
    .A1(net1065),
    .Y(_0263_),
    .A2(_0260_));
 sg13g2_nand2_2 _3481_ (.Y(_0264_),
    .A(_0259_),
    .B(_0263_));
 sg13g2_a221oi_1 _3482_ (.B2(_0253_),
    .C1(net1202),
    .B1(net1171),
    .A1(_0028_),
    .Y(_0265_),
    .A2(net1210));
 sg13g2_a22oi_1 _3483_ (.Y(_0266_),
    .B1(_0264_),
    .B2(_0265_),
    .A2(_2459_),
    .A1(net1202));
 sg13g2_a21oi_1 _3484_ (.A1(net1169),
    .A2(_2460_),
    .Y(_0267_),
    .B1(_0266_));
 sg13g2_o21ai_1 _3485_ (.B1(_0267_),
    .Y(_0268_),
    .A1(_0028_),
    .A2(net1205));
 sg13g2_nor2_1 _3486_ (.A(net1154),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_o21ai_1 _3487_ (.B1(_0269_),
    .Y(_0270_),
    .A1(_2392_),
    .A2(_0254_));
 sg13g2_xor2_1 _3488_ (.B(_0253_),
    .A(_2488_),
    .X(_0271_));
 sg13g2_o21ai_1 _3489_ (.B1(_0270_),
    .Y(_0272_),
    .A1(net1153),
    .A2(_0271_));
 sg13g2_xnor2_1 _3490_ (.Y(_0273_),
    .A(_2322_),
    .B(_2474_));
 sg13g2_a21oi_1 _3491_ (.A1(_1953_),
    .A2(net1056),
    .Y(_0274_),
    .B1(net1075));
 sg13g2_nor2_1 _3492_ (.A(_2444_),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_a21oi_1 _3493_ (.A1(net1075),
    .A2(_2520_),
    .Y(_0276_),
    .B1(_2426_));
 sg13g2_mux2_1 _3494_ (.A0(_0275_),
    .A1(_0276_),
    .S(net1085),
    .X(_0277_));
 sg13g2_a21oi_1 _3495_ (.A1(net1097),
    .A2(_0277_),
    .Y(_0278_),
    .B1(net1066));
 sg13g2_mux2_1 _3496_ (.A0(_2405_),
    .A1(_2407_),
    .S(net1073),
    .X(_0279_));
 sg13g2_a21o_2 _3497_ (.A2(_2438_),
    .A1(net1079),
    .B1(_2421_),
    .X(_0280_));
 sg13g2_mux2_2 _3498_ (.A0(_0279_),
    .A1(_0280_),
    .S(net1084),
    .X(_0281_));
 sg13g2_o21ai_1 _3499_ (.B1(_0278_),
    .Y(_0282_),
    .A1(net1096),
    .A2(_0281_));
 sg13g2_o21ai_1 _3500_ (.B1(_2439_),
    .Y(_0283_),
    .A1(_0257_),
    .A2(_0258_));
 sg13g2_nand3_1 _3501_ (.B(_0282_),
    .C(_0283_),
    .A(net1110),
    .Y(_0284_));
 sg13g2_o21ai_1 _3502_ (.B1(_0284_),
    .Y(_0285_),
    .A1(net1066),
    .A2(_0260_));
 sg13g2_a221oi_1 _3503_ (.B2(_0285_),
    .C1(net1172),
    .B1(_2397_),
    .A1(_0036_),
    .Y(_0286_),
    .A2(net1209));
 sg13g2_a21oi_1 _3504_ (.A1(_2322_),
    .A2(net1172),
    .Y(_0287_),
    .B1(_0286_));
 sg13g2_a21oi_1 _3505_ (.A1(_0036_),
    .A2(net1059),
    .Y(_0288_),
    .B1(_2036_));
 sg13g2_nor3_1 _3506_ (.A(net1170),
    .B(_0287_),
    .C(_0288_),
    .Y(_0289_));
 sg13g2_a21oi_1 _3507_ (.A1(_2321_),
    .A2(net1170),
    .Y(_0290_),
    .B1(_0289_));
 sg13g2_a21oi_1 _3508_ (.A1(_0036_),
    .A2(net1206),
    .Y(_0291_),
    .B1(_2391_));
 sg13g2_o21ai_1 _3509_ (.B1(_0291_),
    .Y(_0292_),
    .A1(net1206),
    .A2(_0290_));
 sg13g2_or3_1 _3510_ (.A(_2322_),
    .B(_2363_),
    .C(_2365_),
    .X(_0293_));
 sg13g2_and2_1 _3511_ (.A(net1151),
    .B(_0293_),
    .X(_0294_));
 sg13g2_a21oi_1 _3512_ (.A1(_2366_),
    .A2(_0294_),
    .Y(_0295_),
    .B1(net1156));
 sg13g2_a22oi_1 _3513_ (.Y(_0296_),
    .B1(_0292_),
    .B2(_0295_),
    .A2(_0273_),
    .A1(net1156));
 sg13g2_or2_1 _3514_ (.X(_0297_),
    .B(_0296_),
    .A(_2039_));
 sg13g2_nor2_2 _3515_ (.A(_2461_),
    .B(_2462_),
    .Y(_0298_));
 sg13g2_xnor2_1 _3516_ (.Y(_0299_),
    .A(_2377_),
    .B(_0298_));
 sg13g2_nor2_1 _3517_ (.A(net1089),
    .B(_0279_),
    .Y(_0300_));
 sg13g2_a21oi_2 _3518_ (.B1(_0300_),
    .Y(_0301_),
    .A2(_0255_),
    .A1(net1089));
 sg13g2_o21ai_1 _3519_ (.B1(net1111),
    .Y(_0302_),
    .A1(net1093),
    .A2(_0211_));
 sg13g2_a21o_1 _3520_ (.A2(_0301_),
    .A1(net1093),
    .B1(_0302_),
    .X(_0303_));
 sg13g2_nand2_1 _3521_ (.Y(_0304_),
    .A(net1109),
    .B(_0303_));
 sg13g2_a21oi_1 _3522_ (.A1(net1102),
    .A2(_0207_),
    .Y(_0305_),
    .B1(_2410_));
 sg13g2_o21ai_1 _3523_ (.B1(_2397_),
    .Y(_0306_),
    .A1(_2018_),
    .A2(net1058));
 sg13g2_nand3_1 _3524_ (.B(net1087),
    .C(_2430_),
    .A(net1096),
    .Y(_0307_));
 sg13g2_nand2_1 _3525_ (.Y(_0308_),
    .A(net1093),
    .B(_0214_));
 sg13g2_a221oi_1 _3526_ (.B2(_0305_),
    .C1(_0306_),
    .B1(_0308_),
    .A1(net1064),
    .Y(_0309_),
    .A2(_0307_));
 sg13g2_a21oi_1 _3527_ (.A1(net1171),
    .A2(_0298_),
    .Y(_0310_),
    .B1(net1202));
 sg13g2_a22oi_1 _3528_ (.Y(_0311_),
    .B1(_0304_),
    .B2(_0309_),
    .A2(net1208),
    .A1(_0030_));
 sg13g2_a221oi_1 _3529_ (.B2(_0311_),
    .C1(net1169),
    .B1(_0310_),
    .A1(net1202),
    .Y(_0312_),
    .A2(_2461_));
 sg13g2_a21oi_1 _3530_ (.A1(_1960_),
    .A2(net1207),
    .Y(_0313_),
    .B1(net1152));
 sg13g2_a21oi_1 _3531_ (.A1(net1169),
    .A2(_2462_),
    .Y(_0314_),
    .B1(_0312_));
 sg13g2_xor2_1 _3532_ (.B(_0298_),
    .A(_2484_),
    .X(_0315_));
 sg13g2_a221oi_1 _3533_ (.B2(_0314_),
    .C1(net1155),
    .B1(_0313_),
    .A1(net1152),
    .Y(_0316_),
    .A2(_0299_));
 sg13g2_a21oi_2 _3534_ (.B1(_0316_),
    .Y(_0317_),
    .A2(_0315_),
    .A1(net1155));
 sg13g2_inv_1 _3535_ (.Y(_0318_),
    .A(_0317_));
 sg13g2_xnor2_1 _3536_ (.Y(_0319_),
    .A(_2467_),
    .B(_2469_));
 sg13g2_a21oi_1 _3537_ (.A1(_0038_),
    .A2(net1209),
    .Y(_0320_),
    .B1(net1173));
 sg13g2_nor3_1 _3538_ (.A(net1102),
    .B(_2410_),
    .C(_0204_),
    .Y(_0321_));
 sg13g2_a21oi_1 _3539_ (.A1(_1949_),
    .A2(net1056),
    .Y(_0322_),
    .B1(net1075));
 sg13g2_nand2_1 _3540_ (.Y(_0323_),
    .A(net1085),
    .B(_0275_));
 sg13g2_o21ai_1 _3541_ (.B1(_0323_),
    .Y(_0324_),
    .A1(net1087),
    .A2(_0280_));
 sg13g2_a21o_1 _3542_ (.A2(_2427_),
    .A1(net1075),
    .B1(net1092),
    .X(_0325_));
 sg13g2_a21oi_1 _3543_ (.A1(net1091),
    .A2(_0276_),
    .Y(_0326_),
    .B1(net1103));
 sg13g2_o21ai_1 _3544_ (.B1(_0326_),
    .Y(_0327_),
    .A1(_0322_),
    .A2(_0325_));
 sg13g2_o21ai_1 _3545_ (.B1(_0327_),
    .Y(_0328_),
    .A1(net1097),
    .A2(_0324_));
 sg13g2_a221oi_1 _3546_ (.B2(net1059),
    .C1(_2018_),
    .B1(_0328_),
    .A1(_2439_),
    .Y(_0329_),
    .A2(_0303_));
 sg13g2_o21ai_1 _3547_ (.B1(_2397_),
    .Y(_0330_),
    .A1(_0321_),
    .A2(_0329_));
 sg13g2_and2_2 _3548_ (.A(net1111),
    .B(net1109),
    .X(_0331_));
 sg13g2_nand2_1 _3549_ (.Y(_0332_),
    .A(net1111),
    .B(net1110));
 sg13g2_a22oi_1 _3550_ (.Y(_0333_),
    .B1(_0320_),
    .B2(_0330_),
    .A2(_2470_),
    .A1(net1172));
 sg13g2_a21oi_1 _3551_ (.A1(_2359_),
    .A2(net1170),
    .Y(_0334_),
    .B1(net1206));
 sg13g2_o21ai_1 _3552_ (.B1(_0334_),
    .Y(_0335_),
    .A1(_2036_),
    .A2(_2360_));
 sg13g2_a21oi_1 _3553_ (.A1(_1936_),
    .A2(net1206),
    .Y(_0336_),
    .B1(net1151));
 sg13g2_o21ai_1 _3554_ (.B1(_0336_),
    .Y(_0337_),
    .A1(_0333_),
    .A2(_0335_));
 sg13g2_or3_1 _3555_ (.A(_2358_),
    .B(_2359_),
    .C(_2360_),
    .X(_0338_));
 sg13g2_and2_1 _3556_ (.A(_2361_),
    .B(_0338_),
    .X(_0339_));
 sg13g2_a21oi_1 _3557_ (.A1(net1151),
    .A2(_0339_),
    .Y(_0340_),
    .B1(net1156));
 sg13g2_a22oi_1 _3558_ (.Y(_0341_),
    .B1(_0337_),
    .B2(_0340_),
    .A2(_0319_),
    .A1(net1157));
 sg13g2_nand2_1 _3559_ (.Y(_0342_),
    .A(net1097),
    .B(_2533_));
 sg13g2_nand2_1 _3560_ (.Y(_0343_),
    .A(_2521_),
    .B(_2523_));
 sg13g2_nand2_1 _3561_ (.Y(_0344_),
    .A(_2519_),
    .B(_2530_));
 sg13g2_o21ai_1 _3562_ (.B1(_2503_),
    .Y(_0345_),
    .A1(net1078),
    .A2(_2405_));
 sg13g2_o21ai_1 _3563_ (.B1(_2524_),
    .Y(_0346_),
    .A1(net1080),
    .A2(_2438_));
 sg13g2_mux2_1 _3564_ (.A0(_0345_),
    .A1(_0346_),
    .S(net1087),
    .X(_0347_));
 sg13g2_nand2_1 _3565_ (.Y(_0348_),
    .A(net1102),
    .B(_0347_));
 sg13g2_mux2_1 _3566_ (.A0(_0343_),
    .A1(_0344_),
    .S(net1085),
    .X(_0349_));
 sg13g2_a21oi_1 _3567_ (.A1(net1097),
    .A2(_0349_),
    .Y(_0350_),
    .B1(net1066));
 sg13g2_nor2_1 _3568_ (.A(_2505_),
    .B(_2510_),
    .Y(_0351_));
 sg13g2_or2_1 _3569_ (.X(_0352_),
    .B(_2510_),
    .A(_2505_));
 sg13g2_mux2_1 _3570_ (.A0(_0234_),
    .A1(_0352_),
    .S(net1082),
    .X(_0353_));
 sg13g2_and2_1 _3571_ (.A(net1093),
    .B(_0353_),
    .X(_0354_));
 sg13g2_a21oi_2 _3572_ (.B1(_0354_),
    .Y(_0355_),
    .A2(_0191_),
    .A1(net1099));
 sg13g2_a21oi_1 _3573_ (.A1(_0348_),
    .A2(_0350_),
    .Y(_0356_),
    .B1(_0332_));
 sg13g2_o21ai_1 _3574_ (.B1(_0356_),
    .Y(_0357_),
    .A1(net1058),
    .A2(_0355_));
 sg13g2_o21ai_1 _3575_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_2410_),
    .A2(_0342_));
 sg13g2_a221oi_1 _3576_ (.B2(_0358_),
    .C1(net1172),
    .B1(_2397_),
    .A1(_0037_),
    .Y(_0359_),
    .A2(net1209));
 sg13g2_a21o_1 _3577_ (.A2(_2473_),
    .A1(net1172),
    .B1(_0359_),
    .X(_0360_));
 sg13g2_a221oi_1 _3578_ (.B2(_2331_),
    .C1(net1207),
    .B1(net1170),
    .A1(net1204),
    .Y(_0361_),
    .A2(_2333_));
 sg13g2_a221oi_1 _3579_ (.B2(_0361_),
    .C1(net1151),
    .B1(_0360_),
    .A1(_1935_),
    .Y(_0362_),
    .A2(net1206));
 sg13g2_o21ai_1 _3580_ (.B1(net1151),
    .Y(_0363_),
    .A1(_2334_),
    .A2(_2362_));
 sg13g2_inv_1 _3581_ (.Y(_0364_),
    .A(_0363_));
 sg13g2_a21oi_1 _3582_ (.A1(_2364_),
    .A2(_0364_),
    .Y(_0365_),
    .B1(_0362_));
 sg13g2_xnor2_1 _3583_ (.Y(_0366_),
    .A(_2471_),
    .B(_2473_));
 sg13g2_nand2_1 _3584_ (.Y(_0367_),
    .A(net1157),
    .B(_0366_));
 sg13g2_o21ai_1 _3585_ (.B1(_0367_),
    .Y(_0368_),
    .A1(net1156),
    .A2(_0365_));
 sg13g2_nor2_1 _3586_ (.A(_0341_),
    .B(_0368_),
    .Y(_0369_));
 sg13g2_xnor2_1 _3587_ (.Y(_0370_),
    .A(_2258_),
    .B(_2482_));
 sg13g2_mux2_1 _3588_ (.A0(_0345_),
    .A1(_0351_),
    .S(net1089),
    .X(_0371_));
 sg13g2_nor2_1 _3589_ (.A(net1100),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_a21oi_1 _3590_ (.A1(net1100),
    .A2(_0236_),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_a21oi_1 _3591_ (.A1(net1111),
    .A2(_0373_),
    .Y(_0374_),
    .B1(_2018_));
 sg13g2_o21ai_1 _3592_ (.B1(_2409_),
    .Y(_0375_),
    .A1(net1096),
    .A2(_0239_));
 sg13g2_a21oi_1 _3593_ (.A1(net1096),
    .A2(_0230_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_a21oi_1 _3594_ (.A1(_2442_),
    .A2(_2527_),
    .Y(_0377_),
    .B1(net1058));
 sg13g2_nor4_2 _3595_ (.A(_0306_),
    .B(_0374_),
    .C(_0376_),
    .Y(_0378_),
    .D(_0377_));
 sg13g2_a21oi_1 _3596_ (.A1(_0031_),
    .A2(net1210),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_a21oi_1 _3597_ (.A1(_2258_),
    .A2(net1171),
    .Y(_0380_),
    .B1(net1204));
 sg13g2_a22oi_1 _3598_ (.Y(_0381_),
    .B1(_0379_),
    .B2(_0380_),
    .A2(_2257_),
    .A1(net1203));
 sg13g2_nor2_1 _3599_ (.A(_2256_),
    .B(_2452_),
    .Y(_0382_));
 sg13g2_o21ai_1 _3600_ (.B1(net1153),
    .Y(_0383_),
    .A1(_0031_),
    .A2(net1205));
 sg13g2_and3_1 _3601_ (.X(_0384_),
    .A(_2258_),
    .B(_2280_),
    .C(_2375_));
 sg13g2_nor3_1 _3602_ (.A(_2376_),
    .B(_2392_),
    .C(_0384_),
    .Y(_0385_));
 sg13g2_or4_1 _3603_ (.A(_0381_),
    .B(_0382_),
    .C(_0383_),
    .D(_0385_),
    .X(_0386_));
 sg13g2_o21ai_1 _3604_ (.B1(_0386_),
    .Y(_0387_),
    .A1(net1153),
    .A2(_0370_));
 sg13g2_nand2_2 _3605_ (.Y(_0388_),
    .A(_2279_),
    .B(_2280_));
 sg13g2_a221oi_1 _3606_ (.B2(_0388_),
    .C1(_2035_),
    .B1(_2395_),
    .A1(_0032_),
    .Y(_0389_),
    .A2(net1208));
 sg13g2_a21o_1 _3607_ (.A2(_2443_),
    .A1(net1064),
    .B1(_2398_),
    .X(_0390_));
 sg13g2_a21oi_1 _3608_ (.A1(net1099),
    .A2(_0256_),
    .Y(_0391_),
    .B1(net1065));
 sg13g2_o21ai_1 _3609_ (.B1(_0391_),
    .Y(_0392_),
    .A1(net1099),
    .A2(_0281_));
 sg13g2_nor2_1 _3610_ (.A(net1064),
    .B(_2448_),
    .Y(_0393_));
 sg13g2_a21oi_1 _3611_ (.A1(_0331_),
    .A2(_0392_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_o21ai_1 _3612_ (.B1(_0389_),
    .Y(_0395_),
    .A1(_0390_),
    .A2(_0394_));
 sg13g2_o21ai_1 _3613_ (.B1(_0395_),
    .Y(_0396_),
    .A1(_2036_),
    .A2(_2465_));
 sg13g2_a221oi_1 _3614_ (.B2(_2463_),
    .C1(net1152),
    .B1(net1169),
    .A1(_1956_),
    .Y(_0397_),
    .A2(net1207));
 sg13g2_xnor2_1 _3615_ (.Y(_0398_),
    .A(_2374_),
    .B(_0388_));
 sg13g2_a22oi_1 _3616_ (.Y(_0399_),
    .B1(_0398_),
    .B2(net1152),
    .A2(_0397_),
    .A1(_0396_));
 sg13g2_xnor2_1 _3617_ (.Y(_0400_),
    .A(_2480_),
    .B(_0388_));
 sg13g2_nand2_1 _3618_ (.Y(_0401_),
    .A(net1155),
    .B(_0400_));
 sg13g2_o21ai_1 _3619_ (.B1(_0401_),
    .Y(_0402_),
    .A1(net1155),
    .A2(_0399_));
 sg13g2_nand4_1 _3620_ (.B(_0369_),
    .C(_0387_),
    .A(_2164_),
    .Y(_0403_),
    .D(_0402_));
 sg13g2_xnor2_1 _3621_ (.Y(_0404_),
    .A(_2236_),
    .B(_2486_));
 sg13g2_and3_1 _3622_ (.X(_0405_),
    .A(_2236_),
    .B(_2246_),
    .C(_2378_));
 sg13g2_nor3_1 _3623_ (.A(_2379_),
    .B(_2392_),
    .C(_0405_),
    .Y(_0406_));
 sg13g2_a21oi_1 _3624_ (.A1(net1102),
    .A2(_2526_),
    .Y(_0407_),
    .B1(_2320_));
 sg13g2_nor4_1 _3625_ (.A(net1109),
    .B(net1099),
    .C(_2507_),
    .D(_2508_),
    .Y(_0408_));
 sg13g2_a21oi_1 _3626_ (.A1(_0331_),
    .A2(_0355_),
    .Y(_0409_),
    .B1(_0408_));
 sg13g2_o21ai_1 _3627_ (.B1(_0409_),
    .Y(_0410_),
    .A1(net1109),
    .A2(_0407_));
 sg13g2_a21oi_1 _3628_ (.A1(net1064),
    .A2(_0342_),
    .Y(_0411_),
    .B1(_0306_));
 sg13g2_a21oi_1 _3629_ (.A1(_2236_),
    .A2(net1171),
    .Y(_0412_),
    .B1(net1202));
 sg13g2_a22oi_1 _3630_ (.Y(_0413_),
    .B1(_0410_),
    .B2(_0411_),
    .A2(net1208),
    .A1(_0029_));
 sg13g2_a22oi_1 _3631_ (.Y(_0414_),
    .B1(_0412_),
    .B2(_0413_),
    .A2(_2235_),
    .A1(net1202));
 sg13g2_a21oi_1 _3632_ (.A1(_2234_),
    .A2(net1169),
    .Y(_0415_),
    .B1(net1154));
 sg13g2_o21ai_1 _3633_ (.B1(_0415_),
    .Y(_0416_),
    .A1(_0029_),
    .A2(net1205));
 sg13g2_or3_1 _3634_ (.A(_0406_),
    .B(_0414_),
    .C(_0416_),
    .X(_0417_));
 sg13g2_o21ai_1 _3635_ (.B1(_0417_),
    .Y(_0418_),
    .A1(net1153),
    .A2(_0404_));
 sg13g2_xnor2_1 _3636_ (.Y(_0419_),
    .A(_2290_),
    .B(_2478_));
 sg13g2_nor2_1 _3637_ (.A(_2167_),
    .B(_0419_),
    .Y(_0420_));
 sg13g2_a21oi_1 _3638_ (.A1(net1099),
    .A2(_0353_),
    .Y(_0421_),
    .B1(net1065));
 sg13g2_o21ai_1 _3639_ (.B1(_0421_),
    .Y(_0422_),
    .A1(net1099),
    .A2(_0347_));
 sg13g2_o21ai_1 _3640_ (.B1(_0422_),
    .Y(_0423_),
    .A1(net1058),
    .A2(_0192_));
 sg13g2_a22oi_1 _3641_ (.Y(_0424_),
    .B1(_0331_),
    .B2(_0423_),
    .A2(_2534_),
    .A1(_2409_));
 sg13g2_a221oi_1 _3642_ (.B2(net1173),
    .C1(net1204),
    .B1(_2290_),
    .A1(_0033_),
    .Y(_0425_),
    .A2(net1208));
 sg13g2_o21ai_1 _3643_ (.B1(_0425_),
    .Y(_0426_),
    .A1(_2398_),
    .A2(_0424_));
 sg13g2_o21ai_1 _3644_ (.B1(_0426_),
    .Y(_0427_),
    .A1(_2036_),
    .A2(_2289_));
 sg13g2_a21oi_1 _3645_ (.A1(_2288_),
    .A2(net1170),
    .Y(_0428_),
    .B1(net1207));
 sg13g2_a221oi_1 _3646_ (.B2(_0428_),
    .C1(net1151),
    .B1(_0427_),
    .A1(_0033_),
    .Y(_0429_),
    .A2(net1207));
 sg13g2_nand3_1 _3647_ (.B(_2370_),
    .C(_2371_),
    .A(_2290_),
    .Y(_0430_));
 sg13g2_nor2_1 _3648_ (.A(_2372_),
    .B(_2392_),
    .Y(_0431_));
 sg13g2_a21oi_1 _3649_ (.A1(_0430_),
    .A2(_0431_),
    .Y(_0432_),
    .B1(_0429_));
 sg13g2_a21o_2 _3650_ (.A2(_0432_),
    .A1(net1153),
    .B1(_0420_),
    .X(_0433_));
 sg13g2_nand2_1 _3651_ (.Y(_0434_),
    .A(_2299_),
    .B(_2466_));
 sg13g2_xor2_1 _3652_ (.B(_0434_),
    .A(_2476_),
    .X(_0435_));
 sg13g2_a21oi_1 _3653_ (.A1(_0034_),
    .A2(net1208),
    .Y(_0436_),
    .B1(net1173));
 sg13g2_nor3_1 _3654_ (.A(_2018_),
    .B(net1058),
    .C(_0212_),
    .Y(_0437_));
 sg13g2_a21oi_1 _3655_ (.A1(net1102),
    .A2(_0301_),
    .Y(_0438_),
    .B1(_0332_));
 sg13g2_o21ai_1 _3656_ (.B1(_0438_),
    .Y(_0439_),
    .A1(net1102),
    .A2(_0324_));
 sg13g2_a21oi_1 _3657_ (.A1(_0208_),
    .A2(_0439_),
    .Y(_0440_),
    .B1(net1064));
 sg13g2_o21ai_1 _3658_ (.B1(_2397_),
    .Y(_0441_),
    .A1(_0437_),
    .A2(_0440_));
 sg13g2_a221oi_1 _3659_ (.B2(_0441_),
    .C1(net1204),
    .B1(_0436_),
    .A1(net1173),
    .Y(_0442_),
    .A2(_0434_));
 sg13g2_o21ai_1 _3660_ (.B1(_2030_),
    .Y(_0443_),
    .A1(_2299_),
    .A2(_2452_));
 sg13g2_a21oi_1 _3661_ (.A1(_1932_),
    .A2(_2298_),
    .Y(_0444_),
    .B1(_2036_));
 sg13g2_or3_1 _3662_ (.A(_0442_),
    .B(_0443_),
    .C(_0444_),
    .X(_0445_));
 sg13g2_o21ai_1 _3663_ (.B1(_0445_),
    .Y(_0446_),
    .A1(\cpu_instance.accum[5] ),
    .A2(net1205));
 sg13g2_or3_1 _3664_ (.A(_2300_),
    .B(_2368_),
    .C(_2369_),
    .X(_0447_));
 sg13g2_nand3_1 _3665_ (.B(net1151),
    .C(_0447_),
    .A(_2370_),
    .Y(_0448_));
 sg13g2_nand3_1 _3666_ (.B(_0446_),
    .C(_0448_),
    .A(net1153),
    .Y(_0449_));
 sg13g2_o21ai_1 _3667_ (.B1(_0449_),
    .Y(_0450_),
    .A1(net1153),
    .A2(_0435_));
 sg13g2_nor2_1 _3668_ (.A(_1950_),
    .B(net1076),
    .Y(_0451_));
 sg13g2_xnor2_1 _3669_ (.Y(_0452_),
    .A(_0039_),
    .B(net1080));
 sg13g2_a21oi_1 _3670_ (.A1(_0039_),
    .A2(net1208),
    .Y(_0453_),
    .B1(net1172));
 sg13g2_mux2_1 _3671_ (.A0(_0343_),
    .A1(_0346_),
    .S(net1091),
    .X(_0454_));
 sg13g2_a21oi_1 _3672_ (.A1(net1103),
    .A2(_0454_),
    .Y(_0455_),
    .B1(net1066));
 sg13g2_nand3_1 _3673_ (.B(_2528_),
    .C(_2529_),
    .A(net1086),
    .Y(_0456_));
 sg13g2_o21ai_1 _3674_ (.B1(_0456_),
    .Y(_0457_),
    .A1(net1085),
    .A2(_0344_));
 sg13g2_o21ai_1 _3675_ (.B1(_0455_),
    .Y(_0458_),
    .A1(net1103),
    .A2(_0457_));
 sg13g2_a21oi_1 _3676_ (.A1(net1111),
    .A2(_0458_),
    .Y(_0459_),
    .B1(_2018_));
 sg13g2_nor3_2 _3677_ (.A(net1064),
    .B(net1100),
    .C(_2441_),
    .Y(_0460_));
 sg13g2_a21oi_1 _3678_ (.A1(_2527_),
    .A2(_0460_),
    .Y(_0461_),
    .B1(net1110));
 sg13g2_nor2_1 _3679_ (.A(net1058),
    .B(_0373_),
    .Y(_0462_));
 sg13g2_or4_1 _3680_ (.A(_2398_),
    .B(_0459_),
    .C(_0461_),
    .D(_0462_),
    .X(_0463_));
 sg13g2_a22oi_1 _3681_ (.Y(_0464_),
    .B1(_0453_),
    .B2(_0463_),
    .A2(_0452_),
    .A1(net1172));
 sg13g2_a21oi_1 _3682_ (.A1(net1170),
    .A2(_2467_),
    .Y(_0465_),
    .B1(net1206));
 sg13g2_nor2_1 _3683_ (.A(_2036_),
    .B(_0451_),
    .Y(_0466_));
 sg13g2_nor2_1 _3684_ (.A(_0464_),
    .B(_0466_),
    .Y(_0467_));
 sg13g2_nor2_1 _3685_ (.A(\cpu_instance.accum[0] ),
    .B(net1205),
    .Y(_0468_));
 sg13g2_a21o_1 _3686_ (.A2(_0467_),
    .A1(_0465_),
    .B1(_0468_),
    .X(_0469_));
 sg13g2_nor3_1 _3687_ (.A(_2392_),
    .B(_2467_),
    .C(_0451_),
    .Y(_0470_));
 sg13g2_nor2_1 _3688_ (.A(net1156),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_a22oi_1 _3689_ (.Y(_0472_),
    .B1(_0469_),
    .B2(_0471_),
    .A2(_0452_),
    .A1(net1156));
 sg13g2_xnor2_1 _3690_ (.Y(_0473_),
    .A(_2310_),
    .B(_2475_));
 sg13g2_a221oi_1 _3691_ (.B2(net1172),
    .C1(net1204),
    .B1(_2310_),
    .A1(net1313),
    .Y(_0474_),
    .A2(net1209));
 sg13g2_mux2_1 _3692_ (.A0(_0371_),
    .A1(_0454_),
    .S(net1096),
    .X(_0475_));
 sg13g2_nand2_1 _3693_ (.Y(_0476_),
    .A(net1058),
    .B(_0475_));
 sg13g2_o21ai_1 _3694_ (.B1(_0476_),
    .Y(_0477_),
    .A1(net1058),
    .A2(_0237_));
 sg13g2_nor2_1 _3695_ (.A(net1064),
    .B(_0242_),
    .Y(_0478_));
 sg13g2_a21oi_1 _3696_ (.A1(_0331_),
    .A2(_0477_),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_o21ai_1 _3697_ (.B1(_0474_),
    .Y(_0480_),
    .A1(_2398_),
    .A2(_0479_));
 sg13g2_o21ai_1 _3698_ (.B1(_0480_),
    .Y(_0481_),
    .A1(_2036_),
    .A2(_2309_));
 sg13g2_a21oi_1 _3699_ (.A1(_2308_),
    .A2(net1170),
    .Y(_0482_),
    .B1(net1206));
 sg13g2_a221oi_1 _3700_ (.B2(_0482_),
    .C1(net1151),
    .B1(_0481_),
    .A1(net1313),
    .Y(_0483_),
    .A2(net1206));
 sg13g2_and3_1 _3701_ (.X(_0484_),
    .A(_2310_),
    .B(_2366_),
    .C(_2367_));
 sg13g2_nor3_1 _3702_ (.A(_2368_),
    .B(_2392_),
    .C(_0484_),
    .Y(_0485_));
 sg13g2_nor3_1 _3703_ (.A(net1156),
    .B(_0483_),
    .C(_0485_),
    .Y(_0486_));
 sg13g2_a21oi_2 _3704_ (.B1(_0486_),
    .Y(_0487_),
    .A2(_0473_),
    .A1(net1156));
 sg13g2_nor2_1 _3705_ (.A(_0472_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_nand4_1 _3706_ (.B(_0433_),
    .C(_0450_),
    .A(_0418_),
    .Y(_0489_),
    .D(_0488_));
 sg13g2_nor4_2 _3707_ (.A(_0297_),
    .B(_0318_),
    .C(_0403_),
    .Y(_0490_),
    .D(_0489_));
 sg13g2_nand3_1 _3708_ (.B(_0272_),
    .C(_0490_),
    .A(_0252_),
    .Y(_0491_));
 sg13g2_or4_2 _3709_ (.A(_2497_),
    .B(_0200_),
    .C(_0226_),
    .D(_0491_),
    .X(_0492_));
 sg13g2_a21oi_1 _3710_ (.A1(_2165_),
    .A2(_0492_),
    .Y(_0055_),
    .B1(net1326));
 sg13g2_nor2_1 _3711_ (.A(net1235),
    .B(net1162),
    .Y(_0493_));
 sg13g2_nand2_1 _3712_ (.Y(_0494_),
    .A(net1242),
    .B(net1161));
 sg13g2_nor2_2 _3713_ (.A(net1237),
    .B(_2093_),
    .Y(_0495_));
 sg13g2_inv_2 _3714_ (.Y(_0496_),
    .A(_0495_));
 sg13g2_nand2_2 _3715_ (.Y(_0497_),
    .A(net1127),
    .B(_0496_));
 sg13g2_or2_2 _3716_ (.X(_0498_),
    .B(_2135_),
    .A(_1886_));
 sg13g2_nand3_1 _3717_ (.B(net1301),
    .C(_2004_),
    .A(net1292),
    .Y(_0499_));
 sg13g2_nor2_2 _3718_ (.A(_0498_),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_nor3_1 _3719_ (.A(_2083_),
    .B(_0498_),
    .C(_0499_),
    .Y(_0501_));
 sg13g2_nand2_2 _3720_ (.Y(_0502_),
    .A(net1248),
    .B(_2111_));
 sg13g2_nand3_1 _3721_ (.B(net1248),
    .C(net1232),
    .A(_2007_),
    .Y(_0503_));
 sg13g2_nor2_2 _3722_ (.A(net1215),
    .B(net1234),
    .Y(_0504_));
 sg13g2_nand2_2 _3723_ (.Y(_0505_),
    .A(net1213),
    .B(net1241));
 sg13g2_and2_2 _3724_ (.A(_0502_),
    .B(_0503_),
    .X(_0506_));
 sg13g2_nand2_1 _3725_ (.Y(_0507_),
    .A(_0502_),
    .B(_0503_));
 sg13g2_nand2b_2 _3726_ (.Y(_0508_),
    .B(_0506_),
    .A_N(net1148));
 sg13g2_or2_1 _3727_ (.X(_0509_),
    .B(_0508_),
    .A(_0497_));
 sg13g2_and3_1 _3728_ (.X(_0510_),
    .A(_0041_),
    .B(net1273),
    .C(_0509_));
 sg13g2_nand3_1 _3729_ (.B(net1273),
    .C(_0509_),
    .A(_0041_),
    .Y(_0511_));
 sg13g2_nor2_2 _3730_ (.A(net1274),
    .B(net1044),
    .Y(_0512_));
 sg13g2_nor2_2 _3731_ (.A(net1285),
    .B(net1267),
    .Y(_0513_));
 sg13g2_nor3_1 _3732_ (.A(net1285),
    .B(_0011_),
    .C(net1267),
    .Y(_0514_));
 sg13g2_xnor2_1 _3733_ (.Y(_0515_),
    .A(_0011_),
    .B(_0513_));
 sg13g2_xor2_1 _3734_ (.B(_0513_),
    .A(_0011_),
    .X(_0516_));
 sg13g2_a22oi_1 _3735_ (.Y(_0517_),
    .B1(_0515_),
    .B2(_0497_),
    .A2(_0508_),
    .A1(\cpu_instance.accum[0] ));
 sg13g2_nor2_1 _3736_ (.A(net1043),
    .B(_0517_),
    .Y(_0518_));
 sg13g2_a221oi_1 _3737_ (.B2(net245),
    .C1(_0518_),
    .B1(_0512_),
    .A1(\cpu_instance.spi_ram.spi_miso_buf ),
    .Y(_0519_),
    .A2(net1275));
 sg13g2_inv_1 _3738_ (.Y(_0056_),
    .A(_0519_));
 sg13g2_a22oi_1 _3739_ (.Y(_0520_),
    .B1(net1027),
    .B2(\cpu_instance.ram_data_out[1] ),
    .A2(net1275),
    .A1(net245));
 sg13g2_xnor2_1 _3740_ (.Y(_0521_),
    .A(_1903_),
    .B(_0514_));
 sg13g2_mux2_1 _3741_ (.A0(_1903_),
    .A1(_0521_),
    .S(_0513_),
    .X(_0522_));
 sg13g2_nand2_1 _3742_ (.Y(_0523_),
    .A(net1131),
    .B(net1145));
 sg13g2_nor2_1 _3743_ (.A(\cpu_instance.accum[1] ),
    .B(_0497_),
    .Y(_0524_));
 sg13g2_o21ai_1 _3744_ (.B1(_0523_),
    .Y(_0525_),
    .A1(_0496_),
    .A2(net1145));
 sg13g2_o21ai_1 _3745_ (.B1(_0510_),
    .Y(_0526_),
    .A1(_0508_),
    .A2(_0525_));
 sg13g2_o21ai_1 _3746_ (.B1(net246),
    .Y(_0057_),
    .A1(_0524_),
    .A2(_0526_));
 sg13g2_a21oi_2 _3747_ (.B1(_1903_),
    .Y(_0527_),
    .A2(_0513_),
    .A1(_0011_));
 sg13g2_nand2_1 _3748_ (.Y(_0528_),
    .A(\cpu_instance.pc[2] ),
    .B(_0527_));
 sg13g2_xor2_1 _3749_ (.B(_0527_),
    .A(\cpu_instance.pc[2] ),
    .X(_0529_));
 sg13g2_inv_2 _3750_ (.Y(_0530_),
    .A(_0529_));
 sg13g2_nand2_2 _3751_ (.Y(_0531_),
    .A(net1145),
    .B(_0529_));
 sg13g2_xor2_1 _3752_ (.B(_0529_),
    .A(net1145),
    .X(_0532_));
 sg13g2_nor2_1 _3753_ (.A(net1131),
    .B(_0532_),
    .Y(_0533_));
 sg13g2_a21oi_1 _3754_ (.A1(net1131),
    .A2(_0530_),
    .Y(_0534_),
    .B1(_0533_));
 sg13g2_a22oi_1 _3755_ (.Y(_0535_),
    .B1(_0534_),
    .B2(_0497_),
    .A2(_0508_),
    .A1(\cpu_instance.accum[2] ));
 sg13g2_nor2_1 _3756_ (.A(net1043),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_a221oi_1 _3757_ (.B2(net300),
    .C1(_0536_),
    .B1(net1027),
    .A1(net290),
    .Y(_0537_),
    .A2(net1275));
 sg13g2_inv_1 _3758_ (.Y(_0058_),
    .A(_0537_));
 sg13g2_nor2_1 _3759_ (.A(\cpu_instance.ram_data_out[3] ),
    .B(net1044),
    .Y(_0538_));
 sg13g2_nand3_1 _3760_ (.B(\cpu_instance.pc[2] ),
    .C(_0527_),
    .A(\cpu_instance.pc[3] ),
    .Y(_0539_));
 sg13g2_xnor2_1 _3761_ (.Y(_0540_),
    .A(\cpu_instance.pc[3] ),
    .B(_0528_));
 sg13g2_xnor2_1 _3762_ (.Y(_0541_),
    .A(_1902_),
    .B(_0528_));
 sg13g2_xnor2_1 _3763_ (.Y(_0542_),
    .A(_0531_),
    .B(_0541_));
 sg13g2_nor2_1 _3764_ (.A(net1127),
    .B(_0540_),
    .Y(_0543_));
 sg13g2_a21oi_1 _3765_ (.A1(net1127),
    .A2(_0542_),
    .Y(_0544_),
    .B1(_0543_));
 sg13g2_a221oi_1 _3766_ (.B2(_0497_),
    .C1(net1043),
    .B1(_0544_),
    .A1(\cpu_instance.accum[3] ),
    .Y(_0545_),
    .A2(_0508_));
 sg13g2_a221oi_1 _3767_ (.B2(_1921_),
    .C1(_0545_),
    .B1(net1027),
    .A1(_1922_),
    .Y(_0059_),
    .A2(net1275));
 sg13g2_nand4_1 _3768_ (.B(\cpu_instance.pc[3] ),
    .C(\cpu_instance.pc[2] ),
    .A(\cpu_instance.pc[4] ),
    .Y(_0546_),
    .D(_0527_));
 sg13g2_xnor2_1 _3769_ (.Y(_0547_),
    .A(\cpu_instance.pc[4] ),
    .B(_0539_));
 sg13g2_xor2_1 _3770_ (.B(_0539_),
    .A(\cpu_instance.pc[4] ),
    .X(_0548_));
 sg13g2_nor3_2 _3771_ (.A(_0531_),
    .B(net1126),
    .C(_0548_),
    .Y(_0549_));
 sg13g2_o21ai_1 _3772_ (.B1(_0548_),
    .Y(_0550_),
    .A1(_0531_),
    .A2(net1126));
 sg13g2_nand2b_2 _3773_ (.Y(_0551_),
    .B(_0550_),
    .A_N(_0549_));
 sg13g2_nor2_1 _3774_ (.A(net1127),
    .B(_0547_),
    .Y(_0552_));
 sg13g2_a21oi_1 _3775_ (.A1(net1127),
    .A2(_0551_),
    .Y(_0553_),
    .B1(_0552_));
 sg13g2_a221oi_1 _3776_ (.B2(_0497_),
    .C1(_0511_),
    .B1(_0553_),
    .A1(\cpu_instance.accum[4] ),
    .Y(_0554_),
    .A2(_0508_));
 sg13g2_nor3_1 _3777_ (.A(net1027),
    .B(_0538_),
    .C(_0554_),
    .Y(_0555_));
 sg13g2_a21o_1 _3778_ (.A2(net1027),
    .A1(net284),
    .B1(_0555_),
    .X(_0060_));
 sg13g2_or2_1 _3779_ (.X(_0556_),
    .B(_0546_),
    .A(_1901_));
 sg13g2_xnor2_1 _3780_ (.Y(_0557_),
    .A(\cpu_instance.pc[5] ),
    .B(_0546_));
 sg13g2_xnor2_1 _3781_ (.Y(_0558_),
    .A(_1901_),
    .B(_0546_));
 sg13g2_a22oi_1 _3782_ (.Y(_0559_),
    .B1(_0557_),
    .B2(net1131),
    .A2(_0508_),
    .A1(\cpu_instance.accum[5] ));
 sg13g2_nand2_1 _3783_ (.Y(_0560_),
    .A(_0549_),
    .B(_0557_));
 sg13g2_xnor2_1 _3784_ (.Y(_0561_),
    .A(_0549_),
    .B(_0558_));
 sg13g2_a21oi_1 _3785_ (.A1(_0495_),
    .A2(_0561_),
    .Y(_0562_),
    .B1(net1042));
 sg13g2_a221oi_1 _3786_ (.B2(_0562_),
    .C1(net1027),
    .B1(_0559_),
    .A1(_1920_),
    .Y(_0563_),
    .A2(net1043));
 sg13g2_a21o_1 _3787_ (.A2(net1027),
    .A1(net283),
    .B1(_0563_),
    .X(_0061_));
 sg13g2_a22oi_1 _3788_ (.Y(_0564_),
    .B1(net1027),
    .B2(net257),
    .A2(net1275),
    .A1(\cpu_instance.ram_data_out[5] ));
 sg13g2_nor2_2 _3789_ (.A(_1900_),
    .B(_0556_),
    .Y(_0565_));
 sg13g2_xnor2_1 _3790_ (.Y(_0566_),
    .A(\cpu_instance.pc[6] ),
    .B(_0556_));
 sg13g2_xnor2_1 _3791_ (.Y(_0567_),
    .A(_1900_),
    .B(_0556_));
 sg13g2_nor2_1 _3792_ (.A(_0560_),
    .B(net1070),
    .Y(_0568_));
 sg13g2_xnor2_1 _3793_ (.Y(_0569_),
    .A(_0560_),
    .B(_0566_));
 sg13g2_a221oi_1 _3794_ (.B2(_0495_),
    .C1(net1131),
    .B1(_0569_),
    .A1(net1312),
    .Y(_0570_),
    .A2(net1148));
 sg13g2_a21oi_1 _3795_ (.A1(net1131),
    .A2(_0567_),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_a21oi_1 _3796_ (.A1(net1312),
    .A2(net1072),
    .Y(_0572_),
    .B1(_0571_));
 sg13g2_o21ai_1 _3797_ (.B1(net258),
    .Y(_0062_),
    .A1(net1043),
    .A2(_0572_));
 sg13g2_a21oi_1 _3798_ (.A1(\cpu_instance.accum[7] ),
    .A2(net1148),
    .Y(_0573_),
    .B1(net1130));
 sg13g2_nand2_1 _3799_ (.Y(_0574_),
    .A(\cpu_instance.pc[7] ),
    .B(_0565_));
 sg13g2_xnor2_1 _3800_ (.Y(_0575_),
    .A(_1899_),
    .B(_0565_));
 sg13g2_xnor2_1 _3801_ (.Y(_0576_),
    .A(\cpu_instance.pc[7] ),
    .B(_0565_));
 sg13g2_nand2_1 _3802_ (.Y(_0577_),
    .A(_0568_),
    .B(_0575_));
 sg13g2_xnor2_1 _3803_ (.Y(_0578_),
    .A(_0568_),
    .B(_0575_));
 sg13g2_o21ai_1 _3804_ (.B1(_0573_),
    .Y(_0579_),
    .A1(_0496_),
    .A2(_0578_));
 sg13g2_a21oi_1 _3805_ (.A1(net1130),
    .A2(_0576_),
    .Y(_0580_),
    .B1(net1072));
 sg13g2_a221oi_1 _3806_ (.B2(_0580_),
    .C1(net1043),
    .B1(_0579_),
    .A1(\cpu_instance.accum[7] ),
    .Y(_0581_),
    .A2(net1072));
 sg13g2_a221oi_1 _3807_ (.B2(_1917_),
    .C1(_0581_),
    .B1(net1026),
    .A1(_1918_),
    .Y(_0063_),
    .A2(net1274));
 sg13g2_a21oi_1 _3808_ (.A1(net1310),
    .A2(net1147),
    .Y(_0582_),
    .B1(net1128));
 sg13g2_nand3_1 _3809_ (.B(\cpu_instance.pc[7] ),
    .C(_0565_),
    .A(\cpu_instance.pc[8] ),
    .Y(_0583_));
 sg13g2_xnor2_1 _3810_ (.Y(_0584_),
    .A(\cpu_instance.pc[8] ),
    .B(_0574_));
 sg13g2_xor2_1 _3811_ (.B(_0574_),
    .A(\cpu_instance.pc[8] ),
    .X(_0585_));
 sg13g2_nor2_1 _3812_ (.A(_0577_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_xnor2_1 _3813_ (.Y(_0587_),
    .A(_0577_),
    .B(_0585_));
 sg13g2_o21ai_1 _3814_ (.B1(_0582_),
    .Y(_0588_),
    .A1(_0496_),
    .A2(_0587_));
 sg13g2_a21oi_1 _3815_ (.A1(net1129),
    .A2(_0585_),
    .Y(_0589_),
    .B1(net1071));
 sg13g2_a221oi_1 _3816_ (.B2(_0589_),
    .C1(net1042),
    .B1(_0588_),
    .A1(net1310),
    .Y(_0590_),
    .A2(net1072));
 sg13g2_a221oi_1 _3817_ (.B2(_1916_),
    .C1(_0590_),
    .B1(net1026),
    .A1(_1917_),
    .Y(_0064_),
    .A2(net1274));
 sg13g2_nand2_1 _3818_ (.Y(_0591_),
    .A(net248),
    .B(net1025));
 sg13g2_nand4_1 _3819_ (.B(\cpu_instance.pc[8] ),
    .C(\cpu_instance.pc[7] ),
    .A(\cpu_instance.pc[9] ),
    .Y(_0592_),
    .D(_0565_));
 sg13g2_xnor2_1 _3820_ (.Y(_0593_),
    .A(\cpu_instance.pc[9] ),
    .B(_0583_));
 sg13g2_and2_1 _3821_ (.A(_0586_),
    .B(net1052),
    .X(_0594_));
 sg13g2_xor2_1 _3822_ (.B(net1051),
    .A(_0586_),
    .X(_0595_));
 sg13g2_a221oi_1 _3823_ (.B2(_0495_),
    .C1(net1130),
    .B1(_0595_),
    .A1(net1309),
    .Y(_0596_),
    .A2(net1147));
 sg13g2_o21ai_1 _3824_ (.B1(_0506_),
    .Y(_0597_),
    .A1(net1127),
    .A2(net1051));
 sg13g2_a21oi_1 _3825_ (.A1(net1309),
    .A2(net1072),
    .Y(_0598_),
    .B1(net1042));
 sg13g2_o21ai_1 _3826_ (.B1(_0598_),
    .Y(_0599_),
    .A1(_0596_),
    .A2(_0597_));
 sg13g2_o21ai_1 _3827_ (.B1(_0599_),
    .Y(_0600_),
    .A1(\cpu_instance.ram_data_out[8] ),
    .A2(net1044));
 sg13g2_o21ai_1 _3828_ (.B1(_0591_),
    .Y(_0065_),
    .A1(net1025),
    .A2(_0600_));
 sg13g2_xnor2_1 _3829_ (.Y(_0601_),
    .A(\cpu_instance.pc[10] ),
    .B(_0592_));
 sg13g2_nand2b_1 _3830_ (.Y(_0602_),
    .B(net1128),
    .A_N(net1049));
 sg13g2_a21oi_1 _3831_ (.A1(net1307),
    .A2(net1147),
    .Y(_0603_),
    .B1(net1128));
 sg13g2_nand2_1 _3832_ (.Y(_0604_),
    .A(_0594_),
    .B(net1050));
 sg13g2_xnor2_1 _3833_ (.Y(_0605_),
    .A(_0594_),
    .B(net1050));
 sg13g2_o21ai_1 _3834_ (.B1(_0603_),
    .Y(_0606_),
    .A1(_0496_),
    .A2(_0605_));
 sg13g2_a221oi_1 _3835_ (.B2(_0606_),
    .C1(net1042),
    .B1(_0602_),
    .A1(net1307),
    .Y(_0607_),
    .A2(net1071));
 sg13g2_a221oi_1 _3836_ (.B2(_1912_),
    .C1(_0607_),
    .B1(net1026),
    .A1(_1914_),
    .Y(_0066_),
    .A2(net1274));
 sg13g2_nand2_1 _3837_ (.Y(_0608_),
    .A(net254),
    .B(net1025));
 sg13g2_or3_2 _3838_ (.A(_1897_),
    .B(_1898_),
    .C(_0592_),
    .X(_0609_));
 sg13g2_o21ai_1 _3839_ (.B1(_1897_),
    .Y(_0610_),
    .A1(_1898_),
    .A2(_0592_));
 sg13g2_and2_1 _3840_ (.A(_0609_),
    .B(_0610_),
    .X(_0611_));
 sg13g2_nor2b_1 _3841_ (.A(_0604_),
    .B_N(net1040),
    .Y(_0612_));
 sg13g2_xnor2_1 _3842_ (.Y(_0613_),
    .A(_0604_),
    .B(net1041));
 sg13g2_a221oi_1 _3843_ (.B2(_0495_),
    .C1(net1129),
    .B1(_0613_),
    .A1(net1306),
    .Y(_0614_),
    .A2(net1147));
 sg13g2_o21ai_1 _3844_ (.B1(_0506_),
    .Y(_0615_),
    .A1(net1127),
    .A2(net1040));
 sg13g2_a21oi_1 _3845_ (.A1(net1306),
    .A2(net1071),
    .Y(_0616_),
    .B1(net1042));
 sg13g2_o21ai_1 _3846_ (.B1(_0616_),
    .Y(_0617_),
    .A1(_0614_),
    .A2(_0615_));
 sg13g2_o21ai_1 _3847_ (.B1(_0617_),
    .Y(_0618_),
    .A1(\cpu_instance.ram_data_out[10] ),
    .A2(net1044));
 sg13g2_o21ai_1 _3848_ (.B1(_0608_),
    .Y(_0067_),
    .A1(net1025),
    .A2(_0618_));
 sg13g2_a22oi_1 _3849_ (.Y(_0619_),
    .B1(net1025),
    .B2(net281),
    .A2(net1274),
    .A1(net254));
 sg13g2_nor2_2 _3850_ (.A(_1896_),
    .B(_0609_),
    .Y(_0620_));
 sg13g2_xnor2_1 _3851_ (.Y(_0621_),
    .A(\cpu_instance.pc[12] ),
    .B(_0609_));
 sg13g2_xnor2_1 _3852_ (.Y(_0622_),
    .A(_1896_),
    .B(_0609_));
 sg13g2_and2_1 _3853_ (.A(_0612_),
    .B(_0621_),
    .X(_0623_));
 sg13g2_xnor2_1 _3854_ (.Y(_0624_),
    .A(_0612_),
    .B(_0622_));
 sg13g2_a221oi_1 _3855_ (.B2(_0495_),
    .C1(net1128),
    .B1(_0624_),
    .A1(net1305),
    .Y(_0625_),
    .A2(net1147));
 sg13g2_a21oi_1 _3856_ (.A1(net1128),
    .A2(_0622_),
    .Y(_0626_),
    .B1(_0625_));
 sg13g2_a21oi_1 _3857_ (.A1(net1305),
    .A2(net1071),
    .Y(_0627_),
    .B1(_0626_));
 sg13g2_o21ai_1 _3858_ (.B1(_0619_),
    .Y(_0068_),
    .A1(net1042),
    .A2(_0627_));
 sg13g2_nand2_1 _3859_ (.Y(_0628_),
    .A(net276),
    .B(net1025));
 sg13g2_a21oi_1 _3860_ (.A1(\cpu_instance.ram_data_out[12] ),
    .A2(net1274),
    .Y(_0629_),
    .B1(net1044));
 sg13g2_a21oi_1 _3861_ (.A1(net1304),
    .A2(net1147),
    .Y(_0630_),
    .B1(net1128));
 sg13g2_nand2_1 _3862_ (.Y(_0631_),
    .A(\cpu_instance.pc[13] ),
    .B(_0620_));
 sg13g2_xnor2_1 _3863_ (.Y(_0632_),
    .A(_1895_),
    .B(_0620_));
 sg13g2_xnor2_1 _3864_ (.Y(_0633_),
    .A(\cpu_instance.pc[13] ),
    .B(_0620_));
 sg13g2_and2_1 _3865_ (.A(_0623_),
    .B(_0632_),
    .X(_0634_));
 sg13g2_xnor2_1 _3866_ (.Y(_0635_),
    .A(_0623_),
    .B(_0632_));
 sg13g2_o21ai_1 _3867_ (.B1(_0630_),
    .Y(_0636_),
    .A1(_0496_),
    .A2(_0635_));
 sg13g2_a21oi_1 _3868_ (.A1(net1128),
    .A2(_0633_),
    .Y(_0637_),
    .B1(net1071));
 sg13g2_a221oi_1 _3869_ (.B2(_0637_),
    .C1(net1042),
    .B1(_0636_),
    .A1(net1304),
    .Y(_0638_),
    .A2(net1071));
 sg13g2_o21ai_1 _3870_ (.B1(_0628_),
    .Y(_0069_),
    .A1(_0629_),
    .A2(_0638_));
 sg13g2_nor3_1 _3871_ (.A(\cpu_instance.ram_data_out[14] ),
    .B(net1274),
    .C(net1044),
    .Y(_0639_));
 sg13g2_nand2b_1 _3872_ (.Y(_0640_),
    .B(_0634_),
    .A_N(_0010_));
 sg13g2_nor2_1 _3873_ (.A(_0010_),
    .B(_0631_),
    .Y(_0641_));
 sg13g2_xor2_1 _3874_ (.B(_0631_),
    .A(_0010_),
    .X(_0642_));
 sg13g2_xnor2_1 _3875_ (.Y(_0643_),
    .A(_0010_),
    .B(_0631_));
 sg13g2_o21ai_1 _3876_ (.B1(_0640_),
    .Y(_0644_),
    .A1(_0634_),
    .A2(_0642_));
 sg13g2_a221oi_1 _3877_ (.B2(net1128),
    .C1(net1071),
    .B1(_0642_),
    .A1(\cpu_instance.accum[14] ),
    .Y(_0645_),
    .A2(net1147));
 sg13g2_o21ai_1 _3878_ (.B1(_0645_),
    .Y(_0646_),
    .A1(_0496_),
    .A2(_0644_));
 sg13g2_o21ai_1 _3879_ (.B1(_0646_),
    .Y(_0647_),
    .A1(\cpu_instance.accum[14] ),
    .A2(_0506_));
 sg13g2_a221oi_1 _3880_ (.B2(_0647_),
    .C1(_0639_),
    .B1(net1044),
    .A1(_1906_),
    .Y(_0070_),
    .A2(net1274));
 sg13g2_nand2_1 _3881_ (.Y(_0648_),
    .A(net278),
    .B(net1025));
 sg13g2_xor2_1 _3882_ (.B(_0641_),
    .A(\cpu_instance.pc[15] ),
    .X(_0649_));
 sg13g2_xnor2_1 _3883_ (.Y(_0650_),
    .A(_0640_),
    .B(net1018));
 sg13g2_a221oi_1 _3884_ (.B2(_0495_),
    .C1(net1129),
    .B1(_0650_),
    .A1(\cpu_instance.accum[15] ),
    .Y(_0651_),
    .A2(net1147));
 sg13g2_o21ai_1 _3885_ (.B1(_0506_),
    .Y(_0652_),
    .A1(net1127),
    .A2(net1017));
 sg13g2_a21oi_1 _3886_ (.A1(\cpu_instance.accum[15] ),
    .A2(net1071),
    .Y(_0653_),
    .B1(net1042));
 sg13g2_o21ai_1 _3887_ (.B1(_0653_),
    .Y(_0654_),
    .A1(_0651_),
    .A2(_0652_));
 sg13g2_o21ai_1 _3888_ (.B1(_0654_),
    .Y(_0655_),
    .A1(\cpu_instance.ram_data_out[14] ),
    .A2(net1044));
 sg13g2_o21ai_1 _3889_ (.B1(_0648_),
    .Y(_0071_),
    .A1(net1025),
    .A2(_0655_));
 sg13g2_nor2_1 _3890_ (.A(net1282),
    .B(_2135_),
    .Y(_0656_));
 sg13g2_nand2b_1 _3891_ (.Y(_0657_),
    .B(_1886_),
    .A_N(_2135_));
 sg13g2_nor2b_2 _3892_ (.A(_0497_),
    .B_N(_0502_),
    .Y(_0658_));
 sg13g2_nand3_1 _3893_ (.B(_0496_),
    .C(_0502_),
    .A(_0494_),
    .Y(_0659_));
 sg13g2_nor2_2 _3894_ (.A(_2051_),
    .B(net1237),
    .Y(_0660_));
 sg13g2_nor3_2 _3895_ (.A(net1269),
    .B(_2052_),
    .C(_0498_),
    .Y(_0661_));
 sg13g2_or2_2 _3896_ (.X(_0662_),
    .B(_0661_),
    .A(_0660_));
 sg13g2_nand2_2 _3897_ (.Y(_0663_),
    .A(_2062_),
    .B(net1242));
 sg13g2_nor3_2 _3898_ (.A(net1269),
    .B(_2058_),
    .C(_0498_),
    .Y(_0664_));
 sg13g2_nor2_1 _3899_ (.A(net1234),
    .B(_2116_),
    .Y(_0665_));
 sg13g2_o21ai_1 _3900_ (.B1(net1241),
    .Y(_0666_),
    .A1(_2113_),
    .A2(net1176));
 sg13g2_or4_2 _3901_ (.A(net1149),
    .B(_0504_),
    .C(_0662_),
    .D(net1124),
    .X(_0667_));
 sg13g2_nor2_1 _3902_ (.A(net1238),
    .B(_2095_),
    .Y(_0668_));
 sg13g2_nor2_2 _3903_ (.A(_2093_),
    .B(_0498_),
    .Y(_0669_));
 sg13g2_o21ai_1 _3904_ (.B1(_0041_),
    .Y(_0670_),
    .A1(_0659_),
    .A2(_0667_));
 sg13g2_nand2_2 _3905_ (.Y(_0671_),
    .A(net1256),
    .B(_0670_));
 sg13g2_a21oi_1 _3906_ (.A1(net1256),
    .A2(_0670_),
    .Y(_0672_),
    .B1(net1277));
 sg13g2_nand2_1 _3907_ (.Y(_0673_),
    .A(net1273),
    .B(_0671_));
 sg13g2_o21ai_1 _3908_ (.B1(net1043),
    .Y(_0072_),
    .A1(_1945_),
    .A2(net1048));
 sg13g2_or2_1 _3909_ (.X(_0674_),
    .B(\cpu_instance.spi_ram.bits_remaining[0] ),
    .A(net181));
 sg13g2_nor2_1 _3910_ (.A(net319),
    .B(_0674_),
    .Y(_0675_));
 sg13g2_nor3_2 _3911_ (.A(net207),
    .B(\cpu_instance.spi_ram.bits_remaining[2] ),
    .C(_0674_),
    .Y(_0676_));
 sg13g2_a21o_1 _3912_ (.A2(_0676_),
    .A1(net1277),
    .B1(net1048),
    .X(_0677_));
 sg13g2_o21ai_1 _3913_ (.B1(net1333),
    .Y(_0678_),
    .A1(net252),
    .A2(_0677_));
 sg13g2_a21oi_1 _3914_ (.A1(net252),
    .A2(_0676_),
    .Y(_0073_),
    .B1(_0678_));
 sg13g2_a21oi_1 _3915_ (.A1(\cpu_instance.spi_ram.fsm_state[0] ),
    .A2(_0676_),
    .Y(_0679_),
    .B1(net220));
 sg13g2_nand2_1 _3916_ (.Y(_0680_),
    .A(net1275),
    .B(_0676_));
 sg13g2_nand2_1 _3917_ (.Y(_0681_),
    .A(net1333),
    .B(_0680_));
 sg13g2_nor2_1 _3918_ (.A(net221),
    .B(_0681_),
    .Y(_0074_));
 sg13g2_o21ai_1 _3919_ (.B1(_0680_),
    .Y(_0682_),
    .A1(net1277),
    .A2(_0671_));
 sg13g2_or2_1 _3920_ (.X(_0683_),
    .B(_0682_),
    .A(net178));
 sg13g2_nand2_1 _3921_ (.Y(_0684_),
    .A(net178),
    .B(net1273));
 sg13g2_a21oi_1 _3922_ (.A1(_0683_),
    .A2(_0684_),
    .Y(_0075_),
    .B1(net1325));
 sg13g2_a21oi_1 _3923_ (.A1(net1277),
    .A2(_0674_),
    .Y(_0685_),
    .B1(_0682_));
 sg13g2_a21oi_1 _3924_ (.A1(net181),
    .A2(_0683_),
    .Y(_0686_),
    .B1(_0685_));
 sg13g2_nor2_1 _3925_ (.A(net1324),
    .B(_0686_),
    .Y(_0076_));
 sg13g2_nor3_1 _3926_ (.A(_1944_),
    .B(net1273),
    .C(_0674_),
    .Y(_0687_));
 sg13g2_o21ai_1 _3927_ (.B1(net1333),
    .Y(_0688_),
    .A1(net268),
    .A2(_0685_));
 sg13g2_nor2_1 _3928_ (.A(_0687_),
    .B(_0688_),
    .Y(_0077_));
 sg13g2_xor2_1 _3929_ (.B(_0675_),
    .A(net207),
    .X(_0689_));
 sg13g2_nand3_1 _3930_ (.B(_0680_),
    .C(_0689_),
    .A(net1277),
    .Y(_0690_));
 sg13g2_nand2_1 _3931_ (.Y(_0691_),
    .A(net207),
    .B(_0682_));
 sg13g2_a21oi_1 _3932_ (.A1(_0690_),
    .A2(_0691_),
    .Y(_0078_),
    .B1(net1324));
 sg13g2_nand2_1 _3933_ (.Y(_0692_),
    .A(net1320),
    .B(net1247));
 sg13g2_nand2_1 _3934_ (.Y(_0693_),
    .A(net262),
    .B(net1239));
 sg13g2_a21oi_1 _3935_ (.A1(_0692_),
    .A2(_0693_),
    .Y(_0079_),
    .B1(net1325));
 sg13g2_nand4_1 _3936_ (.B(net1263),
    .C(_2081_),
    .A(net1287),
    .Y(_0694_),
    .D(_2121_));
 sg13g2_nor2_1 _3937_ (.A(\cpu_instance.inst[3] ),
    .B(_2269_),
    .Y(_0695_));
 sg13g2_nor3_1 _3938_ (.A(\cpu_instance.inst[3] ),
    .B(\cpu_instance.inst[2] ),
    .C(_2269_),
    .Y(_0696_));
 sg13g2_nor4_2 _3939_ (.A(\cpu_instance.inst[7] ),
    .B(\cpu_instance.inst[6] ),
    .C(\cpu_instance.inst[5] ),
    .Y(_0697_),
    .D(\cpu_instance.inst[4] ));
 sg13g2_nor2b_1 _3940_ (.A(\cpu_instance.inst[1] ),
    .B_N(_0697_),
    .Y(_0698_));
 sg13g2_nor2b_1 _3941_ (.A(\cpu_instance.inst[0] ),
    .B_N(_0698_),
    .Y(_0699_));
 sg13g2_a21o_1 _3942_ (.A2(_0699_),
    .A1(_0696_),
    .B1(_0694_),
    .X(_0700_));
 sg13g2_nand3b_1 _3943_ (.B(_0697_),
    .C(\cpu_instance.inst[1] ),
    .Y(_0701_),
    .A_N(\cpu_instance.inst[0] ));
 sg13g2_nand2_1 _3944_ (.Y(_0702_),
    .A(\cpu_instance.inst[0] ),
    .B(_0698_));
 sg13g2_nand2_1 _3945_ (.Y(_0703_),
    .A(_0701_),
    .B(_0702_));
 sg13g2_nand2_1 _3946_ (.Y(_0704_),
    .A(_0695_),
    .B(_0703_));
 sg13g2_nand3_1 _3947_ (.B(\cpu_instance.inst[0] ),
    .C(_0697_),
    .A(\cpu_instance.inst[1] ),
    .Y(_0705_));
 sg13g2_nand2_1 _3948_ (.Y(_0706_),
    .A(\cpu_instance.inst[2] ),
    .B(_0695_));
 sg13g2_o21ai_1 _3949_ (.B1(_0704_),
    .Y(_0707_),
    .A1(_0705_),
    .A2(_0706_));
 sg13g2_nand2b_1 _3950_ (.Y(_0708_),
    .B(_0696_),
    .A_N(_0694_));
 sg13g2_inv_1 _3951_ (.Y(_0709_),
    .A(_0708_));
 sg13g2_nor2_1 _3952_ (.A(_0705_),
    .B(_0708_),
    .Y(_0710_));
 sg13g2_nor2_1 _3953_ (.A(_0694_),
    .B(_0706_),
    .Y(_0711_));
 sg13g2_and2_1 _3954_ (.A(_0699_),
    .B(_0711_),
    .X(_0712_));
 sg13g2_nor4_2 _3955_ (.A(_0700_),
    .B(_0707_),
    .C(_0710_),
    .Y(_0713_),
    .D(_0712_));
 sg13g2_nand2b_1 _3956_ (.Y(_0714_),
    .B(net1247),
    .A_N(_0713_));
 sg13g2_nor2_1 _3957_ (.A(_0701_),
    .B(_0708_),
    .Y(_0715_));
 sg13g2_nand2_1 _3958_ (.Y(_0716_),
    .A(_0703_),
    .B(_0711_));
 sg13g2_or2_1 _3959_ (.X(_0717_),
    .B(_0701_),
    .A(\cpu_instance.carry ));
 sg13g2_o21ai_1 _3960_ (.B1(_0717_),
    .Y(_0718_),
    .A1(_0040_),
    .A2(_0702_));
 sg13g2_a221oi_1 _3961_ (.B2(_0711_),
    .C1(_0712_),
    .B1(_0718_),
    .A1(\cpu_instance.carry ),
    .Y(_0719_),
    .A2(_0716_));
 sg13g2_a21oi_1 _3962_ (.A1(\cpu_instance.neg ),
    .A2(_0712_),
    .Y(_0720_),
    .B1(_0719_));
 sg13g2_nor2_1 _3963_ (.A(_0710_),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_a21oi_1 _3964_ (.A1(_0042_),
    .A2(_0710_),
    .Y(_0722_),
    .B1(_0721_));
 sg13g2_nor2_1 _3965_ (.A(_0702_),
    .B(_0708_),
    .Y(_0723_));
 sg13g2_a21oi_1 _3966_ (.A1(\cpu_instance.skipped ),
    .A2(_0715_),
    .Y(_0724_),
    .B1(_0723_));
 sg13g2_o21ai_1 _3967_ (.B1(_0724_),
    .Y(_0725_),
    .A1(_0715_),
    .A2(_0722_));
 sg13g2_or2_1 _3968_ (.X(_0726_),
    .B(_0694_),
    .A(\cpu_instance.zero ));
 sg13g2_a22oi_1 _3969_ (.Y(_0727_),
    .B1(_0723_),
    .B2(_1972_),
    .A2(_0709_),
    .A1(_0699_));
 sg13g2_a22oi_1 _3970_ (.Y(_0728_),
    .B1(_0727_),
    .B2(_0725_),
    .A2(_0726_),
    .A1(_0700_));
 sg13g2_o21ai_1 _3971_ (.B1(net1333),
    .Y(_0729_),
    .A1(_0714_),
    .A2(_0728_));
 sg13g2_a21oi_1 _3972_ (.A1(net1278),
    .A2(_0714_),
    .Y(_0080_),
    .B1(_0729_));
 sg13g2_o21ai_1 _3973_ (.B1(net1155),
    .Y(_0730_),
    .A1(\cpu_instance.accum[15] ),
    .A2(_2184_));
 sg13g2_a21o_1 _3974_ (.A2(_2497_),
    .A1(_2185_),
    .B1(_0730_),
    .X(_0731_));
 sg13g2_nand2_1 _3975_ (.Y(_0732_),
    .A(_1925_),
    .B(_2184_));
 sg13g2_nand3_1 _3976_ (.B(_2496_),
    .C(_0732_),
    .A(_2456_),
    .Y(_0733_));
 sg13g2_a21oi_1 _3977_ (.A1(\cpu_instance.accum[15] ),
    .A2(_2183_),
    .Y(_0734_),
    .B1(_2392_));
 sg13g2_nor2b_1 _3978_ (.A(_2307_),
    .B_N(_0460_),
    .Y(_0735_));
 sg13g2_xnor2_1 _3979_ (.Y(_0736_),
    .A(_2307_),
    .B(_0460_));
 sg13g2_nor2_2 _3980_ (.A(net1082),
    .B(net1078),
    .Y(_0737_));
 sg13g2_nand2_1 _3981_ (.Y(_0738_),
    .A(net1090),
    .B(_2357_));
 sg13g2_nand2_1 _3982_ (.Y(_0739_),
    .A(net1063),
    .B(_0738_));
 sg13g2_nor2_2 _3983_ (.A(_2442_),
    .B(_0245_),
    .Y(_0740_));
 sg13g2_or2_1 _3984_ (.X(_0741_),
    .B(_0245_),
    .A(_2442_));
 sg13g2_nand2_1 _3985_ (.Y(_0742_),
    .A(_0026_),
    .B(_0741_));
 sg13g2_a21oi_1 _3986_ (.A1(_0030_),
    .A2(_0740_),
    .Y(_0743_),
    .B1(net1074));
 sg13g2_a22oi_1 _3987_ (.Y(_0744_),
    .B1(_0741_),
    .B2(_0027_),
    .A2(net1095),
    .A1(_0031_));
 sg13g2_a22oi_1 _3988_ (.Y(_0745_),
    .B1(_0744_),
    .B2(net1082),
    .A2(_0743_),
    .A1(_0742_));
 sg13g2_a22oi_1 _3989_ (.Y(_0746_),
    .B1(_0740_),
    .B2(_0029_),
    .A2(net1101),
    .A1(_0025_));
 sg13g2_xnor2_1 _3990_ (.Y(_0747_),
    .A(net1064),
    .B(_2442_));
 sg13g2_nand2_1 _3991_ (.Y(_0748_),
    .A(_0024_),
    .B(net1095));
 sg13g2_a21oi_1 _3992_ (.A1(_0028_),
    .A2(net1101),
    .Y(_0749_),
    .B1(net1063));
 sg13g2_a221oi_1 _3993_ (.B2(_0749_),
    .C1(_0747_),
    .B1(_0748_),
    .A1(_0737_),
    .Y(_0750_),
    .A2(_0746_));
 sg13g2_o21ai_1 _3994_ (.B1(_0750_),
    .Y(_0751_),
    .A1(_0739_),
    .A2(_0745_));
 sg13g2_a221oi_1 _3995_ (.B2(_2429_),
    .C1(_0739_),
    .B1(_0740_),
    .A1(net1100),
    .Y(_0752_),
    .A2(_2436_));
 sg13g2_nand2_1 _3996_ (.Y(_0753_),
    .A(_0032_),
    .B(net1095));
 sg13g2_a21oi_1 _3997_ (.A1(_0036_),
    .A2(net1100),
    .Y(_0754_),
    .B1(net1063));
 sg13g2_a21oi_1 _3998_ (.A1(_0033_),
    .A2(net1100),
    .Y(_0755_),
    .B1(_0738_));
 sg13g2_a22oi_1 _3999_ (.Y(_0756_),
    .B1(_0755_),
    .B2(_2472_),
    .A2(_0754_),
    .A1(_0753_));
 sg13g2_nand3b_1 _4000_ (.B(_0756_),
    .C(_0747_),
    .Y(_0757_),
    .A_N(_0752_));
 sg13g2_xnor2_1 _4001_ (.Y(_0758_),
    .A(_2297_),
    .B(_0735_));
 sg13g2_and4_1 _4002_ (.A(_0331_),
    .B(_0751_),
    .C(_0757_),
    .D(_0758_),
    .X(_0759_));
 sg13g2_nand2_1 _4003_ (.Y(_0760_),
    .A(_1931_),
    .B(net1082));
 sg13g2_o21ai_1 _4004_ (.B1(_0760_),
    .Y(_0761_),
    .A1(net1312),
    .A2(net1074));
 sg13g2_nor2_1 _4005_ (.A(\cpu_instance.accum[4] ),
    .B(net1095),
    .Y(_0762_));
 sg13g2_a221oi_1 _4006_ (.B2(net1063),
    .C1(_0762_),
    .B1(_0761_),
    .A1(_1932_),
    .Y(_0763_),
    .A2(_0737_));
 sg13g2_nand2_1 _4007_ (.Y(_0764_),
    .A(\cpu_instance.accum[1] ),
    .B(_0737_));
 sg13g2_a22oi_1 _4008_ (.Y(_0765_),
    .B1(net1079),
    .B2(\cpu_instance.accum[2] ),
    .A2(net1087),
    .A1(\cpu_instance.accum[3] ));
 sg13g2_nand3_1 _4009_ (.B(_0764_),
    .C(_0765_),
    .A(net1063),
    .Y(_0766_));
 sg13g2_a21o_1 _4010_ (.A2(_2442_),
    .A1(\cpu_instance.accum[0] ),
    .B1(_0245_),
    .X(_0767_));
 sg13g2_a221oi_1 _4011_ (.B2(_0767_),
    .C1(_0747_),
    .B1(_0766_),
    .A1(_0740_),
    .Y(_0768_),
    .A2(_0763_));
 sg13g2_nand2_1 _4012_ (.Y(_0769_),
    .A(_1925_),
    .B(net1082));
 sg13g2_o21ai_1 _4013_ (.B1(_0769_),
    .Y(_0770_),
    .A1(\cpu_instance.accum[14] ),
    .A2(net1074));
 sg13g2_nor2_1 _4014_ (.A(\cpu_instance.accum[12] ),
    .B(net1095),
    .Y(_0771_));
 sg13g2_a221oi_1 _4015_ (.B2(net1063),
    .C1(_0771_),
    .B1(_0770_),
    .A1(_1927_),
    .Y(_0772_),
    .A2(_0737_));
 sg13g2_a22oi_1 _4016_ (.Y(_0773_),
    .B1(net1078),
    .B2(net1308),
    .A2(net1082),
    .A1(\cpu_instance.accum[11] ));
 sg13g2_nand2_1 _4017_ (.Y(_0774_),
    .A(net1063),
    .B(_0773_));
 sg13g2_a21oi_1 _4018_ (.A1(net1309),
    .A2(_0737_),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_a21oi_1 _4019_ (.A1(net1311),
    .A2(_2442_),
    .Y(_0776_),
    .B1(_0245_));
 sg13g2_o21ai_1 _4020_ (.B1(_0747_),
    .Y(_0777_),
    .A1(_0775_),
    .A2(_0776_));
 sg13g2_a21oi_1 _4021_ (.A1(_0740_),
    .A2(_0772_),
    .Y(_0778_),
    .B1(_0777_));
 sg13g2_nor4_1 _4022_ (.A(net1109),
    .B(_2297_),
    .C(_0768_),
    .D(_0778_),
    .Y(_0779_));
 sg13g2_o21ai_1 _4023_ (.B1(_0736_),
    .Y(_0780_),
    .A1(_0759_),
    .A2(_0779_));
 sg13g2_nand3b_1 _4024_ (.B(_2164_),
    .C(_0780_),
    .Y(_0781_),
    .A_N(net1210));
 sg13g2_a21oi_1 _4025_ (.A1(_0733_),
    .A2(_0734_),
    .Y(_0782_),
    .B1(_0781_));
 sg13g2_o21ai_1 _4026_ (.B1(net1332),
    .Y(_0783_),
    .A1(net305),
    .A2(_2164_));
 sg13g2_a21oi_2 _4027_ (.B1(_0783_),
    .Y(_0081_),
    .A2(_0782_),
    .A1(_0731_));
 sg13g2_nand3_1 _4028_ (.B(_2456_),
    .C(_2496_),
    .A(_2164_),
    .Y(_0784_));
 sg13g2_o21ai_1 _4029_ (.B1(net1335),
    .Y(_0785_),
    .A1(net267),
    .A2(_2164_));
 sg13g2_nor2b_1 _4030_ (.A(_0785_),
    .B_N(_0784_),
    .Y(_0082_));
 sg13g2_nand3b_1 _4031_ (.B(net1278),
    .C(_1976_),
    .Y(_0786_),
    .A_N(_2090_));
 sg13g2_nor3_2 _4032_ (.A(net1320),
    .B(_1977_),
    .C(_2066_),
    .Y(_0787_));
 sg13g2_o21ai_1 _4033_ (.B1(net1338),
    .Y(_0788_),
    .A1(net191),
    .A2(_0787_));
 sg13g2_a21oi_1 _4034_ (.A1(_1937_),
    .A2(_0787_),
    .Y(_0083_),
    .B1(_0788_));
 sg13g2_o21ai_1 _4035_ (.B1(net1330),
    .Y(_0789_),
    .A1(net185),
    .A2(net1138));
 sg13g2_a21oi_1 _4036_ (.A1(_1936_),
    .A2(net1138),
    .Y(_0084_),
    .B1(_0789_));
 sg13g2_o21ai_1 _4037_ (.B1(net1330),
    .Y(_0790_),
    .A1(net198),
    .A2(net1140));
 sg13g2_a21oi_1 _4038_ (.A1(_1935_),
    .A2(net1140),
    .Y(_0085_),
    .B1(_0790_));
 sg13g2_o21ai_1 _4039_ (.B1(net1328),
    .Y(_0791_),
    .A1(net180),
    .A2(net1139));
 sg13g2_a21oi_1 _4040_ (.A1(_1934_),
    .A2(net1139),
    .Y(_0086_),
    .B1(_0791_));
 sg13g2_o21ai_1 _4041_ (.B1(net1328),
    .Y(_0792_),
    .A1(net182),
    .A2(net1139));
 sg13g2_a21oi_1 _4042_ (.A1(_1933_),
    .A2(net1139),
    .Y(_0087_),
    .B1(_0792_));
 sg13g2_o21ai_1 _4043_ (.B1(net1329),
    .Y(_0793_),
    .A1(net194),
    .A2(net1138));
 sg13g2_a21oi_1 _4044_ (.A1(_1932_),
    .A2(net1138),
    .Y(_0088_),
    .B1(_0793_));
 sg13g2_o21ai_1 _4045_ (.B1(net1328),
    .Y(_0794_),
    .A1(\cpu_instance.accum[6] ),
    .A2(net1141));
 sg13g2_a21oi_1 _4046_ (.A1(_1942_),
    .A2(net1141),
    .Y(_0089_),
    .B1(_0794_));
 sg13g2_o21ai_1 _4047_ (.B1(net1329),
    .Y(_0795_),
    .A1(net186),
    .A2(net1138));
 sg13g2_a21oi_1 _4048_ (.A1(_1931_),
    .A2(net1139),
    .Y(_0090_),
    .B1(_0795_));
 sg13g2_o21ai_1 _4049_ (.B1(net1328),
    .Y(_0796_),
    .A1(net1310),
    .A2(net1141));
 sg13g2_a21oi_1 _4050_ (.A1(_1941_),
    .A2(net1141),
    .Y(_0091_),
    .B1(_0796_));
 sg13g2_o21ai_1 _4051_ (.B1(net1328),
    .Y(_0797_),
    .A1(net184),
    .A2(net1138));
 sg13g2_a21oi_1 _4052_ (.A1(_1930_),
    .A2(net1138),
    .Y(_0092_),
    .B1(_0797_));
 sg13g2_o21ai_1 _4053_ (.B1(net1328),
    .Y(_0798_),
    .A1(net1307),
    .A2(_0786_));
 sg13g2_a21oi_1 _4054_ (.A1(_1940_),
    .A2(net1141),
    .Y(_0093_),
    .B1(_0798_));
 sg13g2_o21ai_1 _4055_ (.B1(net1329),
    .Y(_0799_),
    .A1(net196),
    .A2(net1140));
 sg13g2_a21oi_1 _4056_ (.A1(_1929_),
    .A2(net1140),
    .Y(_0094_),
    .B1(_0799_));
 sg13g2_o21ai_1 _4057_ (.B1(net1328),
    .Y(_0800_),
    .A1(net1305),
    .A2(net1141));
 sg13g2_a21oi_1 _4058_ (.A1(_1939_),
    .A2(net1141),
    .Y(_0095_),
    .B1(_0800_));
 sg13g2_o21ai_1 _4059_ (.B1(net1330),
    .Y(_0801_),
    .A1(net1304),
    .A2(net1141));
 sg13g2_a21oi_1 _4060_ (.A1(_1938_),
    .A2(_0786_),
    .Y(_0096_),
    .B1(_0801_));
 sg13g2_o21ai_1 _4061_ (.B1(net1329),
    .Y(_0802_),
    .A1(net193),
    .A2(net1140));
 sg13g2_a21oi_1 _4062_ (.A1(_1926_),
    .A2(net1140),
    .Y(_0097_),
    .B1(_0802_));
 sg13g2_o21ai_1 _4063_ (.B1(net1328),
    .Y(_0803_),
    .A1(net201),
    .A2(net1139));
 sg13g2_a21oi_1 _4064_ (.A1(_1925_),
    .A2(net1138),
    .Y(_0098_),
    .B1(_0803_));
 sg13g2_nor2_1 _4065_ (.A(net1067),
    .B(net1182),
    .Y(_0804_));
 sg13g2_nand2_2 _4066_ (.Y(_0805_),
    .A(_2039_),
    .B(net1191));
 sg13g2_a21oi_1 _4067_ (.A1(net1253),
    .A2(_2114_),
    .Y(_0806_),
    .B1(net1225));
 sg13g2_o21ai_1 _4068_ (.B1(net1229),
    .Y(_0807_),
    .A1(_2050_),
    .A2(_2113_));
 sg13g2_o21ai_1 _4069_ (.B1(_0807_),
    .Y(_0808_),
    .A1(_1924_),
    .A2(net1192));
 sg13g2_a221oi_1 _4070_ (.B2(\cpu_instance.accum[0] ),
    .C1(_0808_),
    .B1(net1046),
    .A1(_2147_),
    .Y(_0809_),
    .A2(_0472_));
 sg13g2_nor2_1 _4071_ (.A(net1250),
    .B(_0809_),
    .Y(_0810_));
 sg13g2_o21ai_1 _4072_ (.B1(_0810_),
    .Y(_0811_),
    .A1(net245),
    .A2(net1137));
 sg13g2_nor2_1 _4073_ (.A(net1185),
    .B(_0472_),
    .Y(_0812_));
 sg13g2_or3_2 _4074_ (.A(net1270),
    .B(_2345_),
    .C(_2353_),
    .X(_0813_));
 sg13g2_a21oi_1 _4075_ (.A1(net1185),
    .A2(_0813_),
    .Y(_0814_),
    .B1(_0812_));
 sg13g2_nor3_1 _4076_ (.A(_2059_),
    .B(_2110_),
    .C(net1163),
    .Y(_0815_));
 sg13g2_and2_1 _4077_ (.A(_0041_),
    .B(_2102_),
    .X(_0816_));
 sg13g2_or2_1 _4078_ (.X(_0817_),
    .B(_0816_),
    .A(net1320));
 sg13g2_nand3_1 _4079_ (.B(_2150_),
    .C(_0817_),
    .A(_2105_),
    .Y(_0818_));
 sg13g2_nor3_1 _4080_ (.A(_2156_),
    .B(_2161_),
    .C(_0815_),
    .Y(_0819_));
 sg13g2_nand4_1 _4081_ (.B(_2154_),
    .C(_0818_),
    .A(_2106_),
    .Y(_0820_),
    .D(_0819_));
 sg13g2_inv_1 _4082_ (.Y(_0821_),
    .A(net1019));
 sg13g2_a221oi_1 _4083_ (.B2(net1159),
    .C1(net1021),
    .B1(_0814_),
    .A1(\cpu_instance.zero ),
    .Y(_0822_),
    .A2(_2152_));
 sg13g2_a221oi_1 _4084_ (.B2(_0811_),
    .C1(net1325),
    .B1(_0822_),
    .A1(_1937_),
    .Y(_0099_),
    .A2(net1021));
 sg13g2_nand2_1 _4085_ (.Y(_0823_),
    .A(net1192),
    .B(net1137));
 sg13g2_o21ai_1 _4086_ (.B1(net1137),
    .Y(_0824_),
    .A1(_1923_),
    .A2(net1192));
 sg13g2_a221oi_1 _4087_ (.B2(\cpu_instance.accum[1] ),
    .C1(_0824_),
    .B1(net1046),
    .A1(_2147_),
    .Y(_0825_),
    .A2(_0341_));
 sg13g2_nor2_1 _4088_ (.A(net1251),
    .B(_0825_),
    .Y(_0826_));
 sg13g2_o21ai_1 _4089_ (.B1(_0826_),
    .Y(_0827_),
    .A1(\cpu_instance.ram_data_out[1] ),
    .A2(net1137));
 sg13g2_nor2_1 _4090_ (.A(net1184),
    .B(_0341_),
    .Y(_0828_));
 sg13g2_a21oi_1 _4091_ (.A1(net1184),
    .A2(_2339_),
    .Y(_0829_),
    .B1(_0828_));
 sg13g2_a221oi_1 _4092_ (.B2(net1159),
    .C1(net1022),
    .B1(_0829_),
    .A1(net267),
    .Y(_0830_),
    .A2(_2152_));
 sg13g2_a221oi_1 _4093_ (.B2(_0830_),
    .C1(net1325),
    .B1(_0827_),
    .A1(_1936_),
    .Y(_0100_),
    .A2(net1021));
 sg13g2_o21ai_1 _4094_ (.B1(net1137),
    .Y(_0831_),
    .A1(_1922_),
    .A2(net1192));
 sg13g2_a221oi_1 _4095_ (.B2(\cpu_instance.accum[2] ),
    .C1(_0831_),
    .B1(net1046),
    .A1(_2147_),
    .Y(_0832_),
    .A2(_0368_));
 sg13g2_nor2_1 _4096_ (.A(net1250),
    .B(_0832_),
    .Y(_0833_));
 sg13g2_o21ai_1 _4097_ (.B1(_0833_),
    .Y(_0834_),
    .A1(net300),
    .A2(net1137));
 sg13g2_mux2_1 _4098_ (.A0(_2327_),
    .A1(_0368_),
    .S(net1191),
    .X(_0835_));
 sg13g2_a221oi_1 _4099_ (.B2(net1159),
    .C1(net1021),
    .B1(_0835_),
    .A1(net305),
    .Y(_0836_),
    .A2(_2152_));
 sg13g2_a221oi_1 _4100_ (.B2(_0836_),
    .C1(net1325),
    .B1(_0834_),
    .A1(_1935_),
    .Y(_0101_),
    .A2(net1021));
 sg13g2_a221oi_1 _4101_ (.B2(_1934_),
    .C1(_0823_),
    .B1(_2039_),
    .A1(_1976_),
    .Y(_0837_),
    .A2(_1992_));
 sg13g2_a221oi_1 _4102_ (.B2(_0297_),
    .C1(net1021),
    .B1(_0837_),
    .A1(_2317_),
    .Y(_0838_),
    .A2(_0823_));
 sg13g2_a21oi_1 _4103_ (.A1(net1185),
    .A2(_2315_),
    .Y(_0839_),
    .B1(_2139_));
 sg13g2_o21ai_1 _4104_ (.B1(_0839_),
    .Y(_0840_),
    .A1(net1185),
    .A2(_0296_));
 sg13g2_a221oi_1 _4105_ (.B2(_0840_),
    .C1(net1325),
    .B1(_0838_),
    .A1(_1934_),
    .Y(_0102_),
    .A2(net1021));
 sg13g2_a21oi_1 _4106_ (.A1(\cpu_instance.ram_data_out[4] ),
    .A2(net1184),
    .Y(_0841_),
    .B1(net1122));
 sg13g2_a22oi_1 _4107_ (.Y(_0842_),
    .B1(net1047),
    .B2(\cpu_instance.accum[4] ),
    .A2(_0487_),
    .A1(_2147_));
 sg13g2_a221oi_1 _4108_ (.B2(_0842_),
    .C1(net1249),
    .B1(_0841_),
    .A1(_1920_),
    .Y(_0843_),
    .A2(net1122));
 sg13g2_o21ai_1 _4109_ (.B1(net1159),
    .Y(_0844_),
    .A1(net1184),
    .A2(_0487_));
 sg13g2_a21oi_1 _4110_ (.A1(net1184),
    .A2(_2306_),
    .Y(_0845_),
    .B1(_0844_));
 sg13g2_nor3_1 _4111_ (.A(net1022),
    .B(_0843_),
    .C(_0845_),
    .Y(_0846_));
 sg13g2_o21ai_1 _4112_ (.B1(net1332),
    .Y(_0847_),
    .A1(\cpu_instance.accum[4] ),
    .A2(net1016));
 sg13g2_nor2_1 _4113_ (.A(_0846_),
    .B(_0847_),
    .Y(_0103_));
 sg13g2_a221oi_1 _4114_ (.B2(\cpu_instance.accum[5] ),
    .C1(net1122),
    .B1(net1047),
    .A1(\cpu_instance.ram_data_out[5] ),
    .Y(_0848_),
    .A2(net1184));
 sg13g2_o21ai_1 _4115_ (.B1(_0848_),
    .Y(_0849_),
    .A1(net1060),
    .A2(_0450_));
 sg13g2_a21oi_1 _4116_ (.A1(_1919_),
    .A2(net1122),
    .Y(_0850_),
    .B1(net1249));
 sg13g2_nand2_1 _4117_ (.Y(_0851_),
    .A(_0849_),
    .B(_0850_));
 sg13g2_or2_1 _4118_ (.X(_0852_),
    .B(net1105),
    .A(net1191));
 sg13g2_a21oi_1 _4119_ (.A1(net1192),
    .A2(_0450_),
    .Y(_0853_),
    .B1(_2139_));
 sg13g2_a221oi_1 _4120_ (.B2(_0853_),
    .C1(net1021),
    .B1(_0852_),
    .A1(net262),
    .Y(_0854_),
    .A2(_2152_));
 sg13g2_a221oi_1 _4121_ (.B2(_0854_),
    .C1(net1326),
    .B1(_0851_),
    .A1(_1932_),
    .Y(_0104_),
    .A2(net1022));
 sg13g2_a221oi_1 _4122_ (.B2(net1312),
    .C1(_0806_),
    .B1(net1047),
    .A1(\cpu_instance.ram_data_out[6] ),
    .Y(_0855_),
    .A2(net1184));
 sg13g2_o21ai_1 _4123_ (.B1(_0855_),
    .Y(_0856_),
    .A1(_2148_),
    .A2(_0433_));
 sg13g2_a21oi_1 _4124_ (.A1(_1918_),
    .A2(net1122),
    .Y(_0857_),
    .B1(net1246));
 sg13g2_nand2_1 _4125_ (.Y(_0858_),
    .A(net1184),
    .B(_2286_));
 sg13g2_a21oi_1 _4126_ (.A1(net1192),
    .A2(_0433_),
    .Y(_0859_),
    .B1(_2139_));
 sg13g2_a221oi_1 _4127_ (.B2(_0859_),
    .C1(net1022),
    .B1(_0858_),
    .A1(_0856_),
    .Y(_0860_),
    .A2(_0857_));
 sg13g2_o21ai_1 _4128_ (.B1(net1338),
    .Y(_0861_),
    .A1(net1312),
    .A2(net1016));
 sg13g2_nor2_1 _4129_ (.A(_0860_),
    .B(_0861_),
    .Y(_0105_));
 sg13g2_a221oi_1 _4130_ (.B2(\cpu_instance.accum[7] ),
    .C1(net1122),
    .B1(net1047),
    .A1(\cpu_instance.ram_data_out[7] ),
    .Y(_0862_),
    .A2(net1182));
 sg13g2_o21ai_1 _4131_ (.B1(_0862_),
    .Y(_0863_),
    .A1(_2148_),
    .A2(_0402_));
 sg13g2_a21oi_1 _4132_ (.A1(_1917_),
    .A2(net1122),
    .Y(_0864_),
    .B1(net1246));
 sg13g2_nor2_1 _4133_ (.A(net1189),
    .B(_2276_),
    .Y(_0865_));
 sg13g2_a21oi_1 _4134_ (.A1(net1189),
    .A2(_0402_),
    .Y(_0866_),
    .B1(_0865_));
 sg13g2_a221oi_1 _4135_ (.B2(net1158),
    .C1(net1020),
    .B1(_0866_),
    .A1(_0863_),
    .Y(_0867_),
    .A2(_0864_));
 sg13g2_o21ai_1 _4136_ (.B1(net1338),
    .Y(_0868_),
    .A1(\cpu_instance.accum[7] ),
    .A2(net1016));
 sg13g2_nor2_1 _4137_ (.A(_0867_),
    .B(_0868_),
    .Y(_0106_));
 sg13g2_a221oi_1 _4138_ (.B2(net1310),
    .C1(net1120),
    .B1(net1045),
    .A1(\cpu_instance.ram_data_out[8] ),
    .Y(_0869_),
    .A2(net1181));
 sg13g2_o21ai_1 _4139_ (.B1(_0869_),
    .Y(_0870_),
    .A1(net1060),
    .A2(_0387_));
 sg13g2_a21oi_1 _4140_ (.A1(_1916_),
    .A2(net1120),
    .Y(_0871_),
    .B1(net1245));
 sg13g2_nor2_1 _4141_ (.A(net1187),
    .B(_2251_),
    .Y(_0872_));
 sg13g2_a21oi_1 _4142_ (.A1(net1188),
    .A2(_0387_),
    .Y(_0873_),
    .B1(_0872_));
 sg13g2_a221oi_1 _4143_ (.B2(net1158),
    .C1(net1019),
    .B1(_0873_),
    .A1(_0870_),
    .Y(_0874_),
    .A2(_0871_));
 sg13g2_o21ai_1 _4144_ (.B1(net1329),
    .Y(_0875_),
    .A1(net1310),
    .A2(net1016));
 sg13g2_nor2_1 _4145_ (.A(_0874_),
    .B(_0875_),
    .Y(_0107_));
 sg13g2_a221oi_1 _4146_ (.B2(net1309),
    .C1(net1120),
    .B1(net1045),
    .A1(\cpu_instance.ram_data_out[9] ),
    .Y(_0876_),
    .A2(net1182));
 sg13g2_o21ai_1 _4147_ (.B1(_0876_),
    .Y(_0877_),
    .A1(net1060),
    .A2(_0317_));
 sg13g2_a21oi_1 _4148_ (.A1(_1914_),
    .A2(net1121),
    .Y(_0878_),
    .B1(net1245));
 sg13g2_nor2_1 _4149_ (.A(net1188),
    .B(_2241_),
    .Y(_0879_));
 sg13g2_a21oi_1 _4150_ (.A1(net1188),
    .A2(_0317_),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_a221oi_1 _4151_ (.B2(net1158),
    .C1(net1020),
    .B1(_0880_),
    .A1(_0877_),
    .Y(_0881_),
    .A2(_0878_));
 sg13g2_o21ai_1 _4152_ (.B1(net1331),
    .Y(_0882_),
    .A1(net1309),
    .A2(_0821_));
 sg13g2_nor2_1 _4153_ (.A(_0881_),
    .B(_0882_),
    .Y(_0108_));
 sg13g2_a221oi_1 _4154_ (.B2(net1308),
    .C1(net1120),
    .B1(net1045),
    .A1(\cpu_instance.ram_data_out[10] ),
    .Y(_0883_),
    .A2(net1181));
 sg13g2_o21ai_1 _4155_ (.B1(_0883_),
    .Y(_0884_),
    .A1(net1060),
    .A2(_0418_));
 sg13g2_o21ai_1 _4156_ (.B1(_0884_),
    .Y(_0885_),
    .A1(\cpu_instance.ram_data_out[10] ),
    .A2(net1137));
 sg13g2_o21ai_1 _4157_ (.B1(net1158),
    .Y(_0886_),
    .A1(net1187),
    .A2(_2230_));
 sg13g2_a21oi_1 _4158_ (.A1(net1187),
    .A2(_0418_),
    .Y(_0887_),
    .B1(_0886_));
 sg13g2_nor2_1 _4159_ (.A(net1019),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_o21ai_1 _4160_ (.B1(_0888_),
    .Y(_0889_),
    .A1(net1243),
    .A2(_0885_));
 sg13g2_o21ai_1 _4161_ (.B1(_0889_),
    .Y(_0890_),
    .A1(net1307),
    .A2(net1016));
 sg13g2_nor2_1 _4162_ (.A(net1322),
    .B(_0890_),
    .Y(_0109_));
 sg13g2_a221oi_1 _4163_ (.B2(net1306),
    .C1(net1120),
    .B1(net1045),
    .A1(\cpu_instance.ram_data_out[11] ),
    .Y(_0891_),
    .A2(net1181));
 sg13g2_o21ai_1 _4164_ (.B1(_0891_),
    .Y(_0892_),
    .A1(net1060),
    .A2(_0272_));
 sg13g2_a21oi_1 _4165_ (.A1(_1910_),
    .A2(net1120),
    .Y(_0893_),
    .B1(net1245));
 sg13g2_nor2_1 _4166_ (.A(net1187),
    .B(_2222_),
    .Y(_0894_));
 sg13g2_a21oi_1 _4167_ (.A1(net1187),
    .A2(_0272_),
    .Y(_0895_),
    .B1(_0894_));
 sg13g2_a221oi_1 _4168_ (.B2(net1158),
    .C1(net1019),
    .B1(_0895_),
    .A1(_0892_),
    .Y(_0896_),
    .A2(_0893_));
 sg13g2_o21ai_1 _4169_ (.B1(net1331),
    .Y(_0897_),
    .A1(net1306),
    .A2(net1016));
 sg13g2_nor2_1 _4170_ (.A(_0896_),
    .B(_0897_),
    .Y(_0110_));
 sg13g2_a221oi_1 _4171_ (.B2(net1305),
    .C1(net1121),
    .B1(net1045),
    .A1(\cpu_instance.ram_data_out[12] ),
    .Y(_0898_),
    .A2(net1181));
 sg13g2_o21ai_1 _4172_ (.B1(_0898_),
    .Y(_0899_),
    .A1(net1060),
    .A2(_0252_));
 sg13g2_a21oi_1 _4173_ (.A1(_1908_),
    .A2(net1120),
    .Y(_0900_),
    .B1(net1243));
 sg13g2_nor2_1 _4174_ (.A(net1187),
    .B(_2211_),
    .Y(_0901_));
 sg13g2_a21oi_1 _4175_ (.A1(net1187),
    .A2(_0252_),
    .Y(_0902_),
    .B1(_0901_));
 sg13g2_a221oi_1 _4176_ (.B2(net1158),
    .C1(net1019),
    .B1(_0902_),
    .A1(_0899_),
    .Y(_0903_),
    .A2(_0900_));
 sg13g2_o21ai_1 _4177_ (.B1(net1329),
    .Y(_0904_),
    .A1(net1305),
    .A2(net1016));
 sg13g2_nor2_1 _4178_ (.A(_0903_),
    .B(_0904_),
    .Y(_0111_));
 sg13g2_a21oi_1 _4179_ (.A1(\cpu_instance.ram_data_out[13] ),
    .A2(net1181),
    .Y(_0905_),
    .B1(net1120));
 sg13g2_a22oi_1 _4180_ (.Y(_0906_),
    .B1(net1045),
    .B2(net1304),
    .A2(_0226_),
    .A1(_2147_));
 sg13g2_a221oi_1 _4181_ (.B2(_0906_),
    .C1(net1245),
    .B1(_0905_),
    .A1(_1906_),
    .Y(_0907_),
    .A2(net1121));
 sg13g2_o21ai_1 _4182_ (.B1(net1158),
    .Y(_0908_),
    .A1(net1181),
    .A2(_0226_));
 sg13g2_a21oi_1 _4183_ (.A1(net1181),
    .A2(_2203_),
    .Y(_0909_),
    .B1(_0908_));
 sg13g2_nor3_1 _4184_ (.A(net1019),
    .B(_0907_),
    .C(_0909_),
    .Y(_0910_));
 sg13g2_o21ai_1 _4185_ (.B1(net1329),
    .Y(_0911_),
    .A1(net1304),
    .A2(net1016));
 sg13g2_nor2_1 _4186_ (.A(_0910_),
    .B(_0911_),
    .Y(_0112_));
 sg13g2_a21oi_1 _4187_ (.A1(\cpu_instance.ram_data_out[14] ),
    .A2(net1181),
    .Y(_0912_),
    .B1(net1121));
 sg13g2_a22oi_1 _4188_ (.Y(_0913_),
    .B1(net1045),
    .B2(\cpu_instance.accum[14] ),
    .A2(_0200_),
    .A1(_2147_));
 sg13g2_o21ai_1 _4189_ (.B1(net1236),
    .Y(_0914_),
    .A1(\cpu_instance.ram_data_out[14] ),
    .A2(net1137));
 sg13g2_a21o_1 _4190_ (.A2(_0913_),
    .A1(_0912_),
    .B1(_0914_),
    .X(_0915_));
 sg13g2_mux2_1 _4191_ (.A0(_2192_),
    .A1(_0200_),
    .S(net1187),
    .X(_0916_));
 sg13g2_a21oi_1 _4192_ (.A1(net1158),
    .A2(_0916_),
    .Y(_0917_),
    .B1(net1019));
 sg13g2_a221oi_1 _4193_ (.B2(_0917_),
    .C1(net1322),
    .B1(_0915_),
    .A1(_1926_),
    .Y(_0113_),
    .A2(net1019));
 sg13g2_a21oi_1 _4194_ (.A1(_2456_),
    .A2(_2496_),
    .Y(_0918_),
    .B1(net1060));
 sg13g2_a221oi_1 _4195_ (.B2(\cpu_instance.accum[15] ),
    .C1(net1121),
    .B1(net1045),
    .A1(\cpu_instance.ram_data_out[15] ),
    .Y(_0919_),
    .A2(net1182));
 sg13g2_inv_1 _4196_ (.Y(_0920_),
    .A(_0919_));
 sg13g2_a21oi_1 _4197_ (.A1(_1904_),
    .A2(net1121),
    .Y(_0921_),
    .B1(net1246));
 sg13g2_o21ai_1 _4198_ (.B1(_0921_),
    .Y(_0922_),
    .A1(_0918_),
    .A2(_0920_));
 sg13g2_nand3_1 _4199_ (.B(_2456_),
    .C(_2496_),
    .A(net1189),
    .Y(_0923_));
 sg13g2_nor2_1 _4200_ (.A(net1189),
    .B(_2180_),
    .Y(_0924_));
 sg13g2_nor2_1 _4201_ (.A(_2139_),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_a21oi_1 _4202_ (.A1(_0923_),
    .A2(_0925_),
    .Y(_0926_),
    .B1(net1020));
 sg13g2_a221oi_1 _4203_ (.B2(_0926_),
    .C1(net1323),
    .B1(_0922_),
    .A1(_1925_),
    .Y(_0114_),
    .A2(net1020));
 sg13g2_nor2_1 _4204_ (.A(_1974_),
    .B(_2132_),
    .Y(_0927_));
 sg13g2_nand2_1 _4205_ (.Y(_0928_),
    .A(\cpu_instance.spi_ram.spi_select ),
    .B(_2131_));
 sg13g2_o21ai_1 _4206_ (.B1(net1336),
    .Y(_0929_),
    .A1(net275),
    .A2(net1216));
 sg13g2_a21oi_1 _4207_ (.A1(_1924_),
    .A2(net1216),
    .Y(_0115_),
    .B1(_0929_));
 sg13g2_o21ai_1 _4208_ (.B1(net1336),
    .Y(_0930_),
    .A1(net259),
    .A2(net1217));
 sg13g2_a21oi_1 _4209_ (.A1(_1923_),
    .A2(net1217),
    .Y(_0116_),
    .B1(_0930_));
 sg13g2_o21ai_1 _4210_ (.B1(net1335),
    .Y(_0931_),
    .A1(net218),
    .A2(net1218));
 sg13g2_a21oi_1 _4211_ (.A1(_1922_),
    .A2(net1218),
    .Y(_0117_),
    .B1(_0931_));
 sg13g2_o21ai_1 _4212_ (.B1(net1336),
    .Y(_0932_),
    .A1(net250),
    .A2(net1217));
 sg13g2_a21oi_1 _4213_ (.A1(_1921_),
    .A2(net1217),
    .Y(_0118_),
    .B1(_0932_));
 sg13g2_o21ai_1 _4214_ (.B1(net1335),
    .Y(_0933_),
    .A1(net216),
    .A2(net1218));
 sg13g2_a21oi_1 _4215_ (.A1(_1920_),
    .A2(net1218),
    .Y(_0119_),
    .B1(_0933_));
 sg13g2_o21ai_1 _4216_ (.B1(net1334),
    .Y(_0934_),
    .A1(net265),
    .A2(net1218));
 sg13g2_a21oi_1 _4217_ (.A1(_1919_),
    .A2(net1217),
    .Y(_0120_),
    .B1(_0934_));
 sg13g2_o21ai_1 _4218_ (.B1(net1335),
    .Y(_0935_),
    .A1(net222),
    .A2(net1218));
 sg13g2_a21oi_1 _4219_ (.A1(_1918_),
    .A2(net1217),
    .Y(_0121_),
    .B1(_0935_));
 sg13g2_o21ai_1 _4220_ (.B1(net1335),
    .Y(_0936_),
    .A1(net214),
    .A2(net1217));
 sg13g2_a21oi_1 _4221_ (.A1(_1917_),
    .A2(net1217),
    .Y(_0122_),
    .B1(_0936_));
 sg13g2_o21ai_1 _4222_ (.B1(net1332),
    .Y(_0937_),
    .A1(net1303),
    .A2(net1220));
 sg13g2_a21oi_1 _4223_ (.A1(_1916_),
    .A2(net1220),
    .Y(_0123_),
    .B1(_0937_));
 sg13g2_o21ai_1 _4224_ (.B1(net1332),
    .Y(_0938_),
    .A1(net1300),
    .A2(net1220));
 sg13g2_a21oi_1 _4225_ (.A1(_1914_),
    .A2(net1220),
    .Y(_0124_),
    .B1(_0938_));
 sg13g2_o21ai_1 _4226_ (.B1(net1336),
    .Y(_0939_),
    .A1(net1292),
    .A2(net1216));
 sg13g2_a21oi_1 _4227_ (.A1(_1912_),
    .A2(net1216),
    .Y(_0125_),
    .B1(_0939_));
 sg13g2_o21ai_1 _4228_ (.B1(net1336),
    .Y(_0940_),
    .A1(net1290),
    .A2(net1216));
 sg13g2_a21oi_1 _4229_ (.A1(_1910_),
    .A2(net1216),
    .Y(_0126_),
    .B1(_0940_));
 sg13g2_o21ai_1 _4230_ (.B1(net1332),
    .Y(_0941_),
    .A1(net1289),
    .A2(net1220));
 sg13g2_a21oi_1 _4231_ (.A1(_1908_),
    .A2(net1220),
    .Y(_0127_),
    .B1(_0941_));
 sg13g2_o21ai_1 _4232_ (.B1(net1336),
    .Y(_0942_),
    .A1(net1287),
    .A2(net1216));
 sg13g2_a21oi_1 _4233_ (.A1(_1906_),
    .A2(net1216),
    .Y(_0128_),
    .B1(_0942_));
 sg13g2_o21ai_1 _4234_ (.B1(net1333),
    .Y(_0943_),
    .A1(\cpu_instance.ram_data_out[14] ),
    .A2(_0928_));
 sg13g2_a21oi_1 _4235_ (.A1(_1905_),
    .A2(_0928_),
    .Y(_0129_),
    .B1(_0943_));
 sg13g2_o21ai_1 _4236_ (.B1(net1336),
    .Y(_0944_),
    .A1(net1285),
    .A2(net1219));
 sg13g2_a21oi_1 _4237_ (.A1(_1904_),
    .A2(net1219),
    .Y(_0130_),
    .B1(_0944_));
 sg13g2_nor2_2 _4238_ (.A(_2038_),
    .B(net1231),
    .Y(_0945_));
 sg13g2_nand2_2 _4239_ (.Y(_0946_),
    .A(_2039_),
    .B(_2083_));
 sg13g2_nor2_2 _4240_ (.A(net1231),
    .B(_0805_),
    .Y(_0947_));
 sg13g2_nand2_1 _4241_ (.Y(_0948_),
    .A(_2083_),
    .B(net1046));
 sg13g2_nand3b_1 _4242_ (.B(_2090_),
    .C(_2046_),
    .Y(_0949_),
    .A_N(_2100_));
 sg13g2_or2_1 _4243_ (.X(_0950_),
    .B(_0949_),
    .A(net1238));
 sg13g2_nand2_1 _4244_ (.Y(_0951_),
    .A(net1281),
    .B(net1223));
 sg13g2_a22oi_1 _4245_ (.Y(_0952_),
    .B1(_2169_),
    .B2(_1915_),
    .A2(net1223),
    .A1(net1281));
 sg13g2_o21ai_1 _4246_ (.B1(_0951_),
    .Y(_0953_),
    .A1(net1302),
    .A2(_2170_));
 sg13g2_nand2_2 _4247_ (.Y(_0954_),
    .A(_2028_),
    .B(_2067_));
 sg13g2_inv_1 _4248_ (.Y(_0955_),
    .A(_0954_));
 sg13g2_nand2_1 _4249_ (.Y(_0956_),
    .A(_0694_),
    .B(_0954_));
 sg13g2_nand3_1 _4250_ (.B(net1168),
    .C(_0954_),
    .A(_0694_),
    .Y(_0957_));
 sg13g2_nor2_1 _4251_ (.A(net1179),
    .B(_2126_),
    .Y(_0958_));
 sg13g2_nand2b_2 _4252_ (.Y(_0959_),
    .B(net1163),
    .A_N(net1179));
 sg13g2_nor4_1 _4253_ (.A(_2089_),
    .B(_0950_),
    .C(_0957_),
    .D(net1113),
    .Y(_0960_));
 sg13g2_a22oi_1 _4254_ (.Y(_0961_),
    .B1(net1230),
    .B2(_2007_),
    .A2(_2052_),
    .A1(_1991_));
 sg13g2_a21oi_1 _4255_ (.A1(_2033_),
    .A2(_2081_),
    .Y(_0962_),
    .B1(net1277));
 sg13g2_nor2b_1 _4256_ (.A(_0961_),
    .B_N(_0962_),
    .Y(_0963_));
 sg13g2_o21ai_1 _4257_ (.B1(_0947_),
    .Y(_0964_),
    .A1(_0960_),
    .A2(_0963_));
 sg13g2_nand2_1 _4258_ (.Y(_0965_),
    .A(_0041_),
    .B(net1247));
 sg13g2_nor2_1 _4259_ (.A(net1180),
    .B(_0965_),
    .Y(_0966_));
 sg13g2_nor3_1 _4260_ (.A(_2136_),
    .B(_2137_),
    .C(_0966_),
    .Y(_0967_));
 sg13g2_and4_2 _4261_ (.A(_2127_),
    .B(_2144_),
    .C(_0964_),
    .D(_0967_),
    .X(_0968_));
 sg13g2_nand4_1 _4262_ (.B(_2144_),
    .C(_0964_),
    .A(_2127_),
    .Y(_0969_),
    .D(_0967_));
 sg13g2_nor2_1 _4263_ (.A(\cpu_instance.pc[0] ),
    .B(net1319),
    .Y(_0970_));
 sg13g2_a21oi_1 _4264_ (.A1(net1319),
    .A2(_0516_),
    .Y(_0971_),
    .B1(_0970_));
 sg13g2_a21oi_1 _4265_ (.A1(_0516_),
    .A2(net1117),
    .Y(_0972_),
    .B1(net1136));
 sg13g2_o21ai_1 _4266_ (.B1(_0972_),
    .Y(_0973_),
    .A1(net1117),
    .A2(_0971_));
 sg13g2_or4_2 _4267_ (.A(net1267),
    .B(_2345_),
    .C(_2353_),
    .D(_0516_),
    .X(_0974_));
 sg13g2_nor2_1 _4268_ (.A(net1319),
    .B(_0974_),
    .Y(_0975_));
 sg13g2_o21ai_1 _4269_ (.B1(_0516_),
    .Y(_0976_),
    .A1(net1319),
    .A2(_0813_));
 sg13g2_nand2_1 _4270_ (.Y(_0977_),
    .A(_0953_),
    .B(_0976_));
 sg13g2_o21ai_1 _4271_ (.B1(_0973_),
    .Y(_0978_),
    .A1(_0975_),
    .A2(_0977_));
 sg13g2_a22oi_1 _4272_ (.Y(_0979_),
    .B1(_0978_),
    .B2(_0945_),
    .A2(_0971_),
    .A1(net1231));
 sg13g2_nor2_2 _4273_ (.A(_2103_),
    .B(net1046),
    .Y(_0980_));
 sg13g2_nor2b_2 _4274_ (.A(net1046),
    .B_N(net1108),
    .Y(_0981_));
 sg13g2_a22oi_1 _4275_ (.Y(_0982_),
    .B1(_0981_),
    .B2(\cpu_instance.pc[0] ),
    .A2(_0980_),
    .A1(_0515_));
 sg13g2_o21ai_1 _4276_ (.B1(_0982_),
    .Y(_0983_),
    .A1(net1186),
    .A2(_0979_));
 sg13g2_nand2_1 _4277_ (.Y(_0984_),
    .A(net1194),
    .B(_0516_));
 sg13g2_a22oi_1 _4278_ (.Y(_0985_),
    .B1(_0984_),
    .B2(_2099_),
    .A2(_0983_),
    .A1(_2053_));
 sg13g2_nor2_2 _4279_ (.A(_2088_),
    .B(_2104_),
    .Y(_0986_));
 sg13g2_or2_2 _4280_ (.X(_0987_),
    .B(_2104_),
    .A(_2088_));
 sg13g2_o21ai_1 _4281_ (.B1(_0986_),
    .Y(_0988_),
    .A1(net1194),
    .A2(_0971_));
 sg13g2_a21oi_1 _4282_ (.A1(_0515_),
    .A2(net1119),
    .Y(_0989_),
    .B1(net1238));
 sg13g2_o21ai_1 _4283_ (.B1(_0989_),
    .Y(_0990_),
    .A1(_0985_),
    .A2(_0988_));
 sg13g2_nand2_1 _4284_ (.Y(_0991_),
    .A(_0515_),
    .B(net1035));
 sg13g2_a22oi_1 _4285_ (.Y(_0992_),
    .B1(_0516_),
    .B2(net1116),
    .A2(net1179),
    .A1(_1924_));
 sg13g2_a21oi_1 _4286_ (.A1(net1161),
    .A2(_0813_),
    .Y(_0993_),
    .B1(net1227));
 sg13g2_o21ai_1 _4287_ (.B1(_0991_),
    .Y(_0994_),
    .A1(_1924_),
    .A2(net1035));
 sg13g2_a221oi_1 _4288_ (.B2(net1226),
    .C1(net1247),
    .B1(_0994_),
    .A1(_0992_),
    .Y(_0995_),
    .A2(_0993_));
 sg13g2_nor2_1 _4289_ (.A(_0969_),
    .B(_0995_),
    .Y(_0996_));
 sg13g2_a22oi_1 _4290_ (.Y(_0997_),
    .B1(_0990_),
    .B2(_0996_),
    .A2(net1014),
    .A1(net210));
 sg13g2_nor2_1 _4291_ (.A(net1325),
    .B(_0997_),
    .Y(_0131_));
 sg13g2_nand3_1 _4292_ (.B(_2338_),
    .C(net1145),
    .A(_2337_),
    .Y(_0998_));
 sg13g2_a21oi_1 _4293_ (.A1(_2337_),
    .A2(_2338_),
    .Y(_0999_),
    .B1(net1145));
 sg13g2_xnor2_1 _4294_ (.Y(_1000_),
    .A(_2339_),
    .B(net1144));
 sg13g2_xnor2_1 _4295_ (.Y(_1001_),
    .A(_0974_),
    .B(_1000_));
 sg13g2_nand2_1 _4296_ (.Y(_1002_),
    .A(net1279),
    .B(_1001_));
 sg13g2_nand2_1 _4297_ (.Y(_1003_),
    .A(net1319),
    .B(net1144));
 sg13g2_and2_1 _4298_ (.A(_1002_),
    .B(_1003_),
    .X(_1004_));
 sg13g2_o21ai_1 _4299_ (.B1(_1003_),
    .Y(_1005_),
    .A1(_1903_),
    .A2(net1319));
 sg13g2_nand2_1 _4300_ (.Y(_1006_),
    .A(net1144),
    .B(net1116));
 sg13g2_a21oi_1 _4301_ (.A1(net1113),
    .A2(_1005_),
    .Y(_1007_),
    .B1(net1136));
 sg13g2_a221oi_1 _4302_ (.B2(_1007_),
    .C1(net1035),
    .B1(_1006_),
    .A1(net1136),
    .Y(_1008_),
    .A2(_1004_));
 sg13g2_nand2_1 _4303_ (.Y(_1009_),
    .A(net1231),
    .B(_1005_));
 sg13g2_a22oi_1 _4304_ (.Y(_1010_),
    .B1(_0981_),
    .B2(\cpu_instance.pc[1] ),
    .A2(_0980_),
    .A1(net1144));
 sg13g2_nand3_1 _4305_ (.B(_1009_),
    .C(_1010_),
    .A(_2096_),
    .Y(_1011_));
 sg13g2_a21oi_1 _4306_ (.A1(net1201),
    .A2(net1144),
    .Y(_1012_),
    .B1(net1199));
 sg13g2_o21ai_1 _4307_ (.B1(_1012_),
    .Y(_1013_),
    .A1(_1008_),
    .A2(_1011_));
 sg13g2_a21oi_1 _4308_ (.A1(net1199),
    .A2(_1005_),
    .Y(_1014_),
    .B1(net1119));
 sg13g2_nor2_1 _4309_ (.A(net1144),
    .B(_0986_),
    .Y(_1015_));
 sg13g2_a21oi_1 _4310_ (.A1(_1013_),
    .A2(_1014_),
    .Y(_1016_),
    .B1(_1015_));
 sg13g2_nand2_1 _4311_ (.Y(_1017_),
    .A(net1247),
    .B(_1016_));
 sg13g2_nor2_1 _4312_ (.A(\cpu_instance.ram_data_out[1] ),
    .B(net1035),
    .Y(_1018_));
 sg13g2_o21ai_1 _4313_ (.B1(net1226),
    .Y(_1019_),
    .A1(net1144),
    .A2(_0947_));
 sg13g2_and2_1 _4314_ (.A(_2094_),
    .B(net1144),
    .X(_1020_));
 sg13g2_a21oi_1 _4315_ (.A1(_2051_),
    .A2(_1006_),
    .Y(_1021_),
    .B1(_1020_));
 sg13g2_nand2_1 _4316_ (.Y(_1022_),
    .A(\cpu_instance.ram_data_out[1] ),
    .B(net1179));
 sg13g2_o21ai_1 _4317_ (.B1(_1022_),
    .Y(_1023_),
    .A1(net1163),
    .A2(_2339_));
 sg13g2_o21ai_1 _4318_ (.B1(_2107_),
    .Y(_1024_),
    .A1(_1021_),
    .A2(_1023_));
 sg13g2_o21ai_1 _4319_ (.B1(_1024_),
    .Y(_1025_),
    .A1(_1018_),
    .A2(_1019_));
 sg13g2_a21oi_1 _4320_ (.A1(net1238),
    .A2(_1025_),
    .Y(_1026_),
    .B1(net1014));
 sg13g2_a221oi_1 _4321_ (.B2(_1026_),
    .C1(net1324),
    .B1(_1017_),
    .A1(_1903_),
    .Y(_0132_),
    .A2(net1014));
 sg13g2_and2_1 _4322_ (.A(_2327_),
    .B(net1143),
    .X(_1027_));
 sg13g2_nand2b_1 _4323_ (.Y(_1028_),
    .B(_0530_),
    .A_N(_2327_));
 sg13g2_nand2b_1 _4324_ (.Y(_1029_),
    .B(_1028_),
    .A_N(_1027_));
 sg13g2_o21ai_1 _4325_ (.B1(_0998_),
    .Y(_1030_),
    .A1(_0974_),
    .A2(_0999_));
 sg13g2_nand2b_1 _4326_ (.Y(_1031_),
    .B(_1030_),
    .A_N(_1029_));
 sg13g2_nand2b_1 _4327_ (.Y(_1032_),
    .B(_1029_),
    .A_N(_1030_));
 sg13g2_and2_1 _4328_ (.A(net1278),
    .B(_1032_),
    .X(_1033_));
 sg13g2_a22oi_1 _4329_ (.Y(_1034_),
    .B1(_1031_),
    .B2(_1033_),
    .A2(net1143),
    .A1(net1321));
 sg13g2_mux2_1 _4330_ (.A0(\cpu_instance.pc[2] ),
    .A1(net1143),
    .S(net1321),
    .X(_1035_));
 sg13g2_nand2_1 _4331_ (.Y(_1036_),
    .A(net1143),
    .B(net1116));
 sg13g2_a21oi_1 _4332_ (.A1(net1113),
    .A2(_1035_),
    .Y(_1037_),
    .B1(net1136));
 sg13g2_a221oi_1 _4333_ (.B2(_1037_),
    .C1(_0946_),
    .B1(_1036_),
    .A1(net1136),
    .Y(_1038_),
    .A2(_1034_));
 sg13g2_nand2_1 _4334_ (.Y(_1039_),
    .A(\cpu_instance.pc[2] ),
    .B(net1108));
 sg13g2_o21ai_1 _4335_ (.B1(_1039_),
    .Y(_1040_),
    .A1(net1108),
    .A2(_0530_));
 sg13g2_a221oi_1 _4336_ (.B2(_2038_),
    .C1(net1186),
    .B1(_1040_),
    .A1(net1231),
    .Y(_1041_),
    .A2(_1035_));
 sg13g2_nor2b_1 _4337_ (.A(_1038_),
    .B_N(_1041_),
    .Y(_1042_));
 sg13g2_o21ai_1 _4338_ (.B1(_2053_),
    .Y(_1043_),
    .A1(net1191),
    .A2(_1040_));
 sg13g2_a21oi_1 _4339_ (.A1(net1201),
    .A2(_0532_),
    .Y(_1044_),
    .B1(net1199));
 sg13g2_o21ai_1 _4340_ (.B1(_1044_),
    .Y(_1045_),
    .A1(_1042_),
    .A2(_1043_));
 sg13g2_o21ai_1 _4341_ (.B1(net1068),
    .Y(_1046_),
    .A1(net1195),
    .A2(_1035_));
 sg13g2_nand2b_1 _4342_ (.Y(_1047_),
    .B(_1045_),
    .A_N(_1046_));
 sg13g2_nand2_1 _4343_ (.Y(_1048_),
    .A(net1143),
    .B(net1119));
 sg13g2_a21oi_1 _4344_ (.A1(_1047_),
    .A2(_1048_),
    .Y(_1049_),
    .B1(net1237));
 sg13g2_nand2_1 _4345_ (.Y(_1050_),
    .A(\cpu_instance.ram_data_out[2] ),
    .B(net1023));
 sg13g2_a21oi_1 _4346_ (.A1(net1143),
    .A2(net1035),
    .Y(_1051_),
    .B1(net1230));
 sg13g2_nand2_2 _4347_ (.Y(_1052_),
    .A(net1237),
    .B(net1225));
 sg13g2_nor2_1 _4348_ (.A(net1241),
    .B(net1228),
    .Y(_1053_));
 sg13g2_nor2_1 _4349_ (.A(net1143),
    .B(_1020_),
    .Y(_1054_));
 sg13g2_nor2_1 _4350_ (.A(_2063_),
    .B(_0531_),
    .Y(_1055_));
 sg13g2_o21ai_1 _4351_ (.B1(net1116),
    .Y(_1056_),
    .A1(_1054_),
    .A2(_1055_));
 sg13g2_a21oi_1 _4352_ (.A1(_1922_),
    .A2(net1179),
    .Y(_1057_),
    .B1(net1248));
 sg13g2_o21ai_1 _4353_ (.B1(_1057_),
    .Y(_1058_),
    .A1(net1163),
    .A2(_2327_));
 sg13g2_nand2b_1 _4354_ (.Y(_1059_),
    .B(_1056_),
    .A_N(_1058_));
 sg13g2_a22oi_1 _4355_ (.Y(_1060_),
    .B1(_1052_),
    .B2(_1059_),
    .A2(_1051_),
    .A1(_1050_));
 sg13g2_nor3_1 _4356_ (.A(net1014),
    .B(_1049_),
    .C(_1060_),
    .Y(_1061_));
 sg13g2_o21ai_1 _4357_ (.B1(net1332),
    .Y(_1062_),
    .A1(net303),
    .A2(net1015));
 sg13g2_nor2_1 _4358_ (.A(_1061_),
    .B(_1062_),
    .Y(_0133_));
 sg13g2_nand2_1 _4359_ (.Y(_1063_),
    .A(net1321),
    .B(_0540_));
 sg13g2_o21ai_1 _4360_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_1902_),
    .A2(net1321));
 sg13g2_nand2b_1 _4361_ (.Y(_1065_),
    .B(_0540_),
    .A_N(_2315_));
 sg13g2_xnor2_1 _4362_ (.Y(_1066_),
    .A(_2315_),
    .B(net1126));
 sg13g2_a21oi_2 _4363_ (.B1(_1027_),
    .Y(_1067_),
    .A2(_1030_),
    .A1(_1028_));
 sg13g2_or2_1 _4364_ (.X(_1068_),
    .B(_1067_),
    .A(_1066_));
 sg13g2_nand2_1 _4365_ (.Y(_1069_),
    .A(_1066_),
    .B(_1067_));
 sg13g2_nand3_1 _4366_ (.B(_1068_),
    .C(_1069_),
    .A(net1278),
    .Y(_1070_));
 sg13g2_o21ai_1 _4367_ (.B1(net1168),
    .Y(_1071_),
    .A1(net1116),
    .A2(_1064_));
 sg13g2_a21oi_1 _4368_ (.A1(net1126),
    .A2(net1116),
    .Y(_1072_),
    .B1(_1071_));
 sg13g2_nand2_1 _4369_ (.Y(_1073_),
    .A(_1063_),
    .B(_1070_));
 sg13g2_a21o_1 _4370_ (.A2(_1073_),
    .A1(net1136),
    .B1(_1072_),
    .X(_1074_));
 sg13g2_nor2_1 _4371_ (.A(net1108),
    .B(net1126),
    .Y(_1075_));
 sg13g2_a21oi_1 _4372_ (.A1(\cpu_instance.pc[3] ),
    .A2(net1108),
    .Y(_1076_),
    .B1(_1075_));
 sg13g2_a21oi_1 _4373_ (.A1(net1191),
    .A2(_1076_),
    .Y(_1077_),
    .B1(net1046));
 sg13g2_a221oi_1 _4374_ (.B2(_0945_),
    .C1(_1077_),
    .B1(_1074_),
    .A1(net1231),
    .Y(_1078_),
    .A2(_1064_));
 sg13g2_a21o_1 _4375_ (.A2(_1076_),
    .A1(net1186),
    .B1(net1201),
    .X(_1079_));
 sg13g2_a21o_1 _4376_ (.A2(_0542_),
    .A1(net1194),
    .B1(_2073_),
    .X(_1080_));
 sg13g2_o21ai_1 _4377_ (.B1(_1080_),
    .Y(_1081_),
    .A1(_1078_),
    .A2(_1079_));
 sg13g2_o21ai_1 _4378_ (.B1(_1081_),
    .Y(_1082_),
    .A1(net1194),
    .A2(_1064_));
 sg13g2_nand2_1 _4379_ (.Y(_1083_),
    .A(_0986_),
    .B(_1082_));
 sg13g2_a21oi_1 _4380_ (.A1(net1126),
    .A2(net1119),
    .Y(_1084_),
    .B1(net1237));
 sg13g2_nand2_1 _4381_ (.Y(_1085_),
    .A(_1083_),
    .B(_1084_));
 sg13g2_nand2_1 _4382_ (.Y(_1086_),
    .A(\cpu_instance.ram_data_out[3] ),
    .B(net1023));
 sg13g2_a21oi_1 _4383_ (.A1(_0540_),
    .A2(net1035),
    .Y(_1087_),
    .B1(net1230));
 sg13g2_xnor2_1 _4384_ (.Y(_1088_),
    .A(net1126),
    .B(_1055_));
 sg13g2_a221oi_1 _4385_ (.B2(_2315_),
    .C1(net1248),
    .B1(net1161),
    .A1(_1921_),
    .Y(_1089_),
    .A2(net1178));
 sg13g2_o21ai_1 _4386_ (.B1(_1089_),
    .Y(_1090_),
    .A1(net1113),
    .A2(_1088_));
 sg13g2_a22oi_1 _4387_ (.Y(_1091_),
    .B1(_1090_),
    .B2(_1052_),
    .A2(_1087_),
    .A1(_1086_));
 sg13g2_nor2_1 _4388_ (.A(net1014),
    .B(_1091_),
    .Y(_1092_));
 sg13g2_a221oi_1 _4389_ (.B2(_1092_),
    .C1(net1324),
    .B1(_1085_),
    .A1(_1902_),
    .Y(_0134_),
    .A2(net1014));
 sg13g2_nor2_1 _4390_ (.A(net1278),
    .B(_0548_),
    .Y(_1093_));
 sg13g2_nand2_1 _4391_ (.Y(_1094_),
    .A(net1321),
    .B(_0547_));
 sg13g2_nor2_1 _4392_ (.A(_2306_),
    .B(_0548_),
    .Y(_1095_));
 sg13g2_xnor2_1 _4393_ (.Y(_1096_),
    .A(_2306_),
    .B(_0547_));
 sg13g2_o21ai_1 _4394_ (.B1(_1065_),
    .Y(_1097_),
    .A1(_1066_),
    .A2(_1067_));
 sg13g2_a21oi_1 _4395_ (.A1(_1096_),
    .A2(_1097_),
    .Y(_1098_),
    .B1(net1321));
 sg13g2_o21ai_1 _4396_ (.B1(_1098_),
    .Y(_1099_),
    .A1(_1096_),
    .A2(_1097_));
 sg13g2_a21oi_1 _4397_ (.A1(_1094_),
    .A2(_1099_),
    .Y(_1100_),
    .B1(net1168));
 sg13g2_a21oi_1 _4398_ (.A1(\cpu_instance.pc[4] ),
    .A2(net1278),
    .Y(_1101_),
    .B1(_1093_));
 sg13g2_o21ai_1 _4399_ (.B1(net1168),
    .Y(_1102_),
    .A1(_0547_),
    .A2(net1113));
 sg13g2_a21oi_1 _4400_ (.A1(net1113),
    .A2(_1101_),
    .Y(_1103_),
    .B1(_1102_));
 sg13g2_o21ai_1 _4401_ (.B1(net1023),
    .Y(_1104_),
    .A1(_1100_),
    .A2(_1103_));
 sg13g2_o21ai_1 _4402_ (.B1(_2053_),
    .Y(_1105_),
    .A1(_2083_),
    .A2(_1101_));
 sg13g2_a221oi_1 _4403_ (.B2(\cpu_instance.pc[4] ),
    .C1(_1105_),
    .B1(_0981_),
    .A1(_0547_),
    .Y(_1106_),
    .A2(_0980_));
 sg13g2_a221oi_1 _4404_ (.B2(_1106_),
    .C1(net1199),
    .B1(_1104_),
    .A1(net1201),
    .Y(_1107_),
    .A2(_0551_));
 sg13g2_o21ai_1 _4405_ (.B1(net1068),
    .Y(_1108_),
    .A1(net1195),
    .A2(_1101_));
 sg13g2_a21oi_1 _4406_ (.A1(_0548_),
    .A2(net1119),
    .Y(_1109_),
    .B1(net1237));
 sg13g2_o21ai_1 _4407_ (.B1(_1109_),
    .Y(_1110_),
    .A1(_1107_),
    .A2(_1108_));
 sg13g2_nor2_1 _4408_ (.A(net1163),
    .B(_2306_),
    .Y(_1111_));
 sg13g2_nor2_2 _4409_ (.A(_2050_),
    .B(net1113),
    .Y(_1112_));
 sg13g2_a221oi_1 _4410_ (.B2(_1112_),
    .C1(net1226),
    .B1(_0547_),
    .A1(\cpu_instance.ram_data_out[4] ),
    .Y(_1113_),
    .A2(net1178));
 sg13g2_o21ai_1 _4411_ (.B1(_1113_),
    .Y(_1114_),
    .A1(_2095_),
    .A2(_0551_));
 sg13g2_nor2_1 _4412_ (.A(_1111_),
    .B(_1114_),
    .Y(_1115_));
 sg13g2_o21ai_1 _4413_ (.B1(net1226),
    .Y(_1116_),
    .A1(_0548_),
    .A2(net1023));
 sg13g2_a21oi_1 _4414_ (.A1(\cpu_instance.ram_data_out[4] ),
    .A2(net1023),
    .Y(_1117_),
    .B1(_1116_));
 sg13g2_nor3_1 _4415_ (.A(net1248),
    .B(_1115_),
    .C(_1117_),
    .Y(_1118_));
 sg13g2_nor2_1 _4416_ (.A(net1014),
    .B(_1118_),
    .Y(_1119_));
 sg13g2_o21ai_1 _4417_ (.B1(net1332),
    .Y(_1120_),
    .A1(net308),
    .A2(_0968_));
 sg13g2_a21oi_1 _4418_ (.A1(_1110_),
    .A2(_1119_),
    .Y(_0135_),
    .B1(_1120_));
 sg13g2_nand2_1 _4419_ (.Y(_1121_),
    .A(net1318),
    .B(_0557_));
 sg13g2_a21oi_1 _4420_ (.A1(_1096_),
    .A2(_1097_),
    .Y(_1122_),
    .B1(_1095_));
 sg13g2_nand2b_1 _4421_ (.Y(_1123_),
    .B(_0558_),
    .A_N(_2295_));
 sg13g2_inv_1 _4422_ (.Y(_1124_),
    .A(_1123_));
 sg13g2_xnor2_1 _4423_ (.Y(_1125_),
    .A(net1105),
    .B(_0557_));
 sg13g2_o21ai_1 _4424_ (.B1(net1280),
    .Y(_1126_),
    .A1(_1122_),
    .A2(_1125_));
 sg13g2_a21oi_1 _4425_ (.A1(_1122_),
    .A2(_1125_),
    .Y(_1127_),
    .B1(_1126_));
 sg13g2_a21oi_1 _4426_ (.A1(net1318),
    .A2(_0557_),
    .Y(_1128_),
    .B1(_1127_));
 sg13g2_o21ai_1 _4427_ (.B1(_1121_),
    .Y(_1129_),
    .A1(_1901_),
    .A2(net1318));
 sg13g2_a21oi_1 _4428_ (.A1(_0558_),
    .A2(net1115),
    .Y(_1130_),
    .B1(net1136));
 sg13g2_o21ai_1 _4429_ (.B1(_1130_),
    .Y(_1131_),
    .A1(net1115),
    .A2(_1129_));
 sg13g2_o21ai_1 _4430_ (.B1(_1131_),
    .Y(_1132_),
    .A1(net1167),
    .A2(_1128_));
 sg13g2_nand2_1 _4431_ (.Y(_1133_),
    .A(\cpu_instance.pc[5] ),
    .B(net1108));
 sg13g2_o21ai_1 _4432_ (.B1(_1133_),
    .Y(_1134_),
    .A1(net1108),
    .A2(_0558_));
 sg13g2_a21oi_1 _4433_ (.A1(net1067),
    .A2(_1134_),
    .Y(_1135_),
    .B1(net1186));
 sg13g2_a22oi_1 _4434_ (.Y(_1136_),
    .B1(_1132_),
    .B2(_0945_),
    .A2(_1129_),
    .A1(net1232));
 sg13g2_o21ai_1 _4435_ (.B1(_2053_),
    .Y(_1137_),
    .A1(net1191),
    .A2(_1134_));
 sg13g2_a21oi_1 _4436_ (.A1(_1135_),
    .A2(_1136_),
    .Y(_1138_),
    .B1(_1137_));
 sg13g2_a21oi_1 _4437_ (.A1(net1200),
    .A2(_0561_),
    .Y(_1139_),
    .B1(_1138_));
 sg13g2_a21oi_1 _4438_ (.A1(net1198),
    .A2(_1129_),
    .Y(_1140_),
    .B1(net1118));
 sg13g2_o21ai_1 _4439_ (.B1(_1140_),
    .Y(_1141_),
    .A1(net1199),
    .A2(_1139_));
 sg13g2_a21oi_1 _4440_ (.A1(_0558_),
    .A2(net1118),
    .Y(_1142_),
    .B1(net1237));
 sg13g2_a21oi_1 _4441_ (.A1(_0558_),
    .A2(_0948_),
    .Y(_1143_),
    .B1(net1229));
 sg13g2_o21ai_1 _4442_ (.B1(_1143_),
    .Y(_1144_),
    .A1(\cpu_instance.ram_data_out[5] ),
    .A2(net1035));
 sg13g2_nand2b_1 _4443_ (.Y(_1145_),
    .B(_2050_),
    .A_N(_0561_));
 sg13g2_a21oi_1 _4444_ (.A1(_2095_),
    .A2(_0558_),
    .Y(_1146_),
    .B1(net1178));
 sg13g2_a221oi_1 _4445_ (.B2(_1146_),
    .C1(net1161),
    .B1(_1145_),
    .A1(\cpu_instance.ram_data_out[5] ),
    .Y(_1147_),
    .A2(net1178));
 sg13g2_o21ai_1 _4446_ (.B1(net1229),
    .Y(_1148_),
    .A1(net1162),
    .A2(net1105));
 sg13g2_o21ai_1 _4447_ (.B1(_1144_),
    .Y(_1149_),
    .A1(_1147_),
    .A2(_1148_));
 sg13g2_a221oi_1 _4448_ (.B2(net1237),
    .C1(net1014),
    .B1(_1149_),
    .A1(_1141_),
    .Y(_1150_),
    .A2(_1142_));
 sg13g2_o21ai_1 _4449_ (.B1(net1332),
    .Y(_1151_),
    .A1(net244),
    .A2(net1015));
 sg13g2_nor2_1 _4450_ (.A(_1150_),
    .B(_1151_),
    .Y(_0136_));
 sg13g2_nand2_1 _4451_ (.Y(_1152_),
    .A(net1318),
    .B(_0566_));
 sg13g2_nor2_1 _4452_ (.A(_2286_),
    .B(net1070),
    .Y(_1153_));
 sg13g2_xnor2_1 _4453_ (.Y(_1154_),
    .A(_2286_),
    .B(net1070));
 sg13g2_a221oi_1 _4454_ (.B2(_1097_),
    .C1(_1095_),
    .B1(_1096_),
    .A1(net1105),
    .Y(_1155_),
    .A2(_0557_));
 sg13g2_nor2_1 _4455_ (.A(_1124_),
    .B(_1155_),
    .Y(_1156_));
 sg13g2_nor3_2 _4456_ (.A(_1124_),
    .B(_1154_),
    .C(_1155_),
    .Y(_1157_));
 sg13g2_xor2_1 _4457_ (.B(_1156_),
    .A(_1154_),
    .X(_1158_));
 sg13g2_o21ai_1 _4458_ (.B1(_1152_),
    .Y(_1159_),
    .A1(net1318),
    .A2(_1158_));
 sg13g2_o21ai_1 _4459_ (.B1(_1152_),
    .Y(_1160_),
    .A1(_1900_),
    .A2(net1318));
 sg13g2_nand2b_1 _4460_ (.Y(_1161_),
    .B(net1112),
    .A_N(_1160_));
 sg13g2_a21oi_1 _4461_ (.A1(net1070),
    .A2(net1115),
    .Y(_1162_),
    .B1(net1135));
 sg13g2_a22oi_1 _4462_ (.Y(_1163_),
    .B1(_1161_),
    .B2(_1162_),
    .A2(_1159_),
    .A1(net1135));
 sg13g2_a21o_1 _4463_ (.A2(_0980_),
    .A1(_0566_),
    .B1(_2064_),
    .X(_1164_));
 sg13g2_a221oi_1 _4464_ (.B2(net1233),
    .C1(_1164_),
    .B1(_1160_),
    .A1(\cpu_instance.pc[6] ),
    .Y(_1165_),
    .A2(_0981_));
 sg13g2_o21ai_1 _4465_ (.B1(_1165_),
    .Y(_1166_),
    .A1(net1034),
    .A2(_1163_));
 sg13g2_o21ai_1 _4466_ (.B1(net1196),
    .Y(_1167_),
    .A1(_2053_),
    .A2(_0569_));
 sg13g2_nand2b_1 _4467_ (.Y(_1168_),
    .B(_1166_),
    .A_N(_1167_));
 sg13g2_a21oi_1 _4468_ (.A1(net1198),
    .A2(_1160_),
    .Y(_1169_),
    .B1(net1119));
 sg13g2_a22oi_1 _4469_ (.Y(_1170_),
    .B1(_1168_),
    .B2(_1169_),
    .A2(_0987_),
    .A1(net1070));
 sg13g2_nand2_1 _4470_ (.Y(_1171_),
    .A(net1242),
    .B(_1170_));
 sg13g2_a21oi_1 _4471_ (.A1(\cpu_instance.ram_data_out[6] ),
    .A2(net1178),
    .Y(_1172_),
    .B1(net1161));
 sg13g2_a21oi_1 _4472_ (.A1(net1253),
    .A2(net1070),
    .Y(_1173_),
    .B1(net1177));
 sg13g2_o21ai_1 _4473_ (.B1(_1173_),
    .Y(_1174_),
    .A1(net1253),
    .A2(_0569_));
 sg13g2_a221oi_1 _4474_ (.B2(_1174_),
    .C1(net1227),
    .B1(_1172_),
    .A1(net1161),
    .Y(_1175_),
    .A2(_2286_));
 sg13g2_o21ai_1 _4475_ (.B1(net1227),
    .Y(_1176_),
    .A1(\cpu_instance.ram_data_out[6] ),
    .A2(net1034));
 sg13g2_a21oi_1 _4476_ (.A1(net1070),
    .A2(net1034),
    .Y(_1177_),
    .B1(_1176_));
 sg13g2_o21ai_1 _4477_ (.B1(net1235),
    .Y(_1178_),
    .A1(_1175_),
    .A2(_1177_));
 sg13g2_and2_1 _4478_ (.A(_0968_),
    .B(_1178_),
    .X(_1179_));
 sg13g2_a221oi_1 _4479_ (.B2(_1179_),
    .C1(net1326),
    .B1(_1171_),
    .A1(_1900_),
    .Y(_0137_),
    .A2(net1013));
 sg13g2_nor2_1 _4480_ (.A(net1106),
    .B(_0576_),
    .Y(_1180_));
 sg13g2_a21oi_1 _4481_ (.A1(\cpu_instance.pc[7] ),
    .A2(net1106),
    .Y(_1181_),
    .B1(_1180_));
 sg13g2_nor2_1 _4482_ (.A(_1153_),
    .B(_1157_),
    .Y(_1182_));
 sg13g2_nand2_1 _4483_ (.Y(_1183_),
    .A(_2276_),
    .B(_0575_));
 sg13g2_nand2b_1 _4484_ (.Y(_1184_),
    .B(_0576_),
    .A_N(_2276_));
 sg13g2_nand2_1 _4485_ (.Y(_1185_),
    .A(_1183_),
    .B(_1184_));
 sg13g2_xnor2_1 _4486_ (.Y(_1186_),
    .A(_1182_),
    .B(_1185_));
 sg13g2_nand2_1 _4487_ (.Y(_1187_),
    .A(net1314),
    .B(_0575_));
 sg13g2_a21oi_1 _4488_ (.A1(net1314),
    .A2(_0575_),
    .Y(_1188_),
    .B1(net1167));
 sg13g2_o21ai_1 _4489_ (.B1(_1188_),
    .Y(_1189_),
    .A1(net1314),
    .A2(_1186_));
 sg13g2_o21ai_1 _4490_ (.B1(_1187_),
    .Y(_1190_),
    .A1(_1899_),
    .A2(net1314));
 sg13g2_a21oi_1 _4491_ (.A1(net1112),
    .A2(_1190_),
    .Y(_1191_),
    .B1(net1135));
 sg13g2_o21ai_1 _4492_ (.B1(_1191_),
    .Y(_1192_),
    .A1(_0576_),
    .A2(net1112));
 sg13g2_nand3_1 _4493_ (.B(_1189_),
    .C(_1192_),
    .A(_0945_),
    .Y(_1193_));
 sg13g2_nand2_1 _4494_ (.Y(_1194_),
    .A(net1190),
    .B(_1181_));
 sg13g2_a22oi_1 _4495_ (.Y(_1195_),
    .B1(_1194_),
    .B2(_0805_),
    .A2(_1190_),
    .A1(net1233));
 sg13g2_a22oi_1 _4496_ (.Y(_1196_),
    .B1(_1193_),
    .B2(_1195_),
    .A2(_1181_),
    .A1(net1183));
 sg13g2_a21oi_1 _4497_ (.A1(net1200),
    .A2(_0578_),
    .Y(_1197_),
    .B1(net1197));
 sg13g2_o21ai_1 _4498_ (.B1(_1197_),
    .Y(_1198_),
    .A1(_2064_),
    .A2(_1196_));
 sg13g2_a21oi_1 _4499_ (.A1(net1197),
    .A2(_1190_),
    .Y(_1199_),
    .B1(net1118));
 sg13g2_a22oi_1 _4500_ (.Y(_1200_),
    .B1(_1198_),
    .B2(_1199_),
    .A2(_0987_),
    .A1(_0576_));
 sg13g2_nand2_1 _4501_ (.Y(_1201_),
    .A(net1241),
    .B(_1200_));
 sg13g2_a21oi_1 _4502_ (.A1(_1917_),
    .A2(net1024),
    .Y(_1202_),
    .B1(net1229));
 sg13g2_o21ai_1 _4503_ (.B1(_1202_),
    .Y(_1203_),
    .A1(_0575_),
    .A2(net1024));
 sg13g2_nand2_1 _4504_ (.Y(_1204_),
    .A(_2050_),
    .B(_0578_));
 sg13g2_a21oi_1 _4505_ (.A1(net1253),
    .A2(_0576_),
    .Y(_1205_),
    .B1(net1177));
 sg13g2_a221oi_1 _4506_ (.B2(_1205_),
    .C1(net1160),
    .B1(_1204_),
    .A1(\cpu_instance.ram_data_out[7] ),
    .Y(_1206_),
    .A2(net1177));
 sg13g2_o21ai_1 _4507_ (.B1(net1228),
    .Y(_1207_),
    .A1(net1162),
    .A2(_2276_));
 sg13g2_o21ai_1 _4508_ (.B1(_1203_),
    .Y(_1208_),
    .A1(_1206_),
    .A2(_1207_));
 sg13g2_a21oi_1 _4509_ (.A1(net1234),
    .A2(_1208_),
    .Y(_1209_),
    .B1(net1012));
 sg13g2_a221oi_1 _4510_ (.B2(_1209_),
    .C1(net1322),
    .B1(_1201_),
    .A1(_1899_),
    .Y(_0138_),
    .A2(net1012));
 sg13g2_mux2_1 _4511_ (.A0(\cpu_instance.pc[8] ),
    .A1(_0584_),
    .S(net1314),
    .X(_1210_));
 sg13g2_o21ai_1 _4512_ (.B1(net1167),
    .Y(_1211_),
    .A1(net1114),
    .A2(_1210_));
 sg13g2_a21oi_1 _4513_ (.A1(_0585_),
    .A2(net1114),
    .Y(_1212_),
    .B1(_1211_));
 sg13g2_nand2_1 _4514_ (.Y(_1213_),
    .A(_2251_),
    .B(_0584_));
 sg13g2_xnor2_1 _4515_ (.Y(_1214_),
    .A(_2251_),
    .B(_0584_));
 sg13g2_o21ai_1 _4516_ (.B1(_1184_),
    .Y(_1215_),
    .A1(_1153_),
    .A2(_1157_));
 sg13g2_nand2_1 _4517_ (.Y(_1216_),
    .A(_1183_),
    .B(_1215_));
 sg13g2_a21o_1 _4518_ (.A2(_1215_),
    .A1(_1183_),
    .B1(_1214_),
    .X(_1217_));
 sg13g2_xnor2_1 _4519_ (.Y(_1218_),
    .A(_1214_),
    .B(_1216_));
 sg13g2_mux2_1 _4520_ (.A0(_0584_),
    .A1(_1218_),
    .S(net1280),
    .X(_1219_));
 sg13g2_a21oi_1 _4521_ (.A1(net1134),
    .A2(_1219_),
    .Y(_1220_),
    .B1(_1212_));
 sg13g2_nor2_1 _4522_ (.A(net1034),
    .B(_1220_),
    .Y(_1221_));
 sg13g2_nand2_1 _4523_ (.Y(_1222_),
    .A(net1233),
    .B(_1210_));
 sg13g2_a22oi_1 _4524_ (.Y(_1223_),
    .B1(_0981_),
    .B2(\cpu_instance.pc[8] ),
    .A2(_0980_),
    .A1(_0584_));
 sg13g2_nand3_1 _4525_ (.B(_1222_),
    .C(_1223_),
    .A(net1180),
    .Y(_1224_));
 sg13g2_a21oi_1 _4526_ (.A1(net1200),
    .A2(_0587_),
    .Y(_1225_),
    .B1(net1197));
 sg13g2_o21ai_1 _4527_ (.B1(_1225_),
    .Y(_1226_),
    .A1(_1221_),
    .A2(_1224_));
 sg13g2_a21oi_1 _4528_ (.A1(net1197),
    .A2(_1210_),
    .Y(_1227_),
    .B1(net1118));
 sg13g2_a22oi_1 _4529_ (.Y(_1228_),
    .B1(_1226_),
    .B2(_1227_),
    .A2(_0987_),
    .A1(_0585_));
 sg13g2_nand2_1 _4530_ (.Y(_1229_),
    .A(net1241),
    .B(_1228_));
 sg13g2_a21oi_1 _4531_ (.A1(_0585_),
    .A2(net1032),
    .Y(_1230_),
    .B1(net1228));
 sg13g2_o21ai_1 _4532_ (.B1(_1230_),
    .Y(_1231_),
    .A1(\cpu_instance.ram_data_out[8] ),
    .A2(net1032));
 sg13g2_o21ai_1 _4533_ (.B1(net1228),
    .Y(_1232_),
    .A1(net1162),
    .A2(_2251_));
 sg13g2_nand2_1 _4534_ (.Y(_1233_),
    .A(_2050_),
    .B(_0587_));
 sg13g2_a21oi_1 _4535_ (.A1(net1253),
    .A2(_0585_),
    .Y(_1234_),
    .B1(net1177));
 sg13g2_a221oi_1 _4536_ (.B2(_1234_),
    .C1(net1160),
    .B1(_1233_),
    .A1(\cpu_instance.ram_data_out[8] ),
    .Y(_1235_),
    .A2(net1177));
 sg13g2_o21ai_1 _4537_ (.B1(_1231_),
    .Y(_1236_),
    .A1(_1232_),
    .A2(_1235_));
 sg13g2_a21oi_1 _4538_ (.A1(net1234),
    .A2(_1236_),
    .Y(_1237_),
    .B1(net1012));
 sg13g2_o21ai_1 _4539_ (.B1(net1331),
    .Y(_1238_),
    .A1(net295),
    .A2(net1015));
 sg13g2_a21oi_1 _4540_ (.A1(_1229_),
    .A2(_1237_),
    .Y(_0139_),
    .B1(_1238_));
 sg13g2_nor2_1 _4541_ (.A(_2241_),
    .B(net1052),
    .Y(_1239_));
 sg13g2_nand2_1 _4542_ (.Y(_1240_),
    .A(_2241_),
    .B(net1052));
 sg13g2_nand2b_1 _4543_ (.Y(_1241_),
    .B(_1240_),
    .A_N(_1239_));
 sg13g2_nand2_1 _4544_ (.Y(_1242_),
    .A(_1213_),
    .B(_1217_));
 sg13g2_xor2_1 _4545_ (.B(_1242_),
    .A(_1241_),
    .X(_1243_));
 sg13g2_a21oi_1 _4546_ (.A1(net1315),
    .A2(net1052),
    .Y(_1244_),
    .B1(net1167));
 sg13g2_o21ai_1 _4547_ (.B1(_1244_),
    .Y(_1245_),
    .A1(net1314),
    .A2(_1243_));
 sg13g2_mux2_1 _4548_ (.A0(\cpu_instance.pc[9] ),
    .A1(net1051),
    .S(net1318),
    .X(_1246_));
 sg13g2_inv_1 _4549_ (.Y(_1247_),
    .A(_1246_));
 sg13g2_a21oi_1 _4550_ (.A1(net1051),
    .A2(net1115),
    .Y(_1248_),
    .B1(net1135));
 sg13g2_o21ai_1 _4551_ (.B1(_1248_),
    .Y(_1249_),
    .A1(net1115),
    .A2(_1247_));
 sg13g2_nand3_1 _4552_ (.B(_1245_),
    .C(_1249_),
    .A(_0945_),
    .Y(_1250_));
 sg13g2_nor2b_1 _4553_ (.A(net1107),
    .B_N(net1051),
    .Y(_1251_));
 sg13g2_a21oi_1 _4554_ (.A1(\cpu_instance.pc[9] ),
    .A2(net1107),
    .Y(_1252_),
    .B1(_1251_));
 sg13g2_nand2_1 _4555_ (.Y(_1253_),
    .A(net1190),
    .B(_1252_));
 sg13g2_a22oi_1 _4556_ (.Y(_1254_),
    .B1(_1253_),
    .B2(_0805_),
    .A2(_1246_),
    .A1(net1233));
 sg13g2_a221oi_1 _4557_ (.B2(_1250_),
    .C1(net1200),
    .B1(_1254_),
    .A1(net1183),
    .Y(_1255_),
    .A2(_1252_));
 sg13g2_a221oi_1 _4558_ (.B2(net1200),
    .C1(_1255_),
    .B1(_0595_),
    .A1(_1998_),
    .Y(_1256_),
    .A2(_2067_));
 sg13g2_o21ai_1 _4559_ (.B1(net1068),
    .Y(_1257_),
    .A1(net1196),
    .A2(_1246_));
 sg13g2_a21oi_1 _4560_ (.A1(net1051),
    .A2(_0987_),
    .Y(_1258_),
    .B1(net1235));
 sg13g2_o21ai_1 _4561_ (.B1(_1258_),
    .Y(_1259_),
    .A1(_1256_),
    .A2(_1257_));
 sg13g2_a22oi_1 _4562_ (.Y(_1260_),
    .B1(net1160),
    .B2(_2241_),
    .A2(_2117_),
    .A1(\cpu_instance.ram_data_out[9] ));
 sg13g2_a22oi_1 _4563_ (.Y(_1261_),
    .B1(_1112_),
    .B2(net1051),
    .A2(_0595_),
    .A1(_2062_));
 sg13g2_nand3_1 _4564_ (.B(_1260_),
    .C(_1261_),
    .A(net1235),
    .Y(_1262_));
 sg13g2_nor2_1 _4565_ (.A(net1051),
    .B(net1024),
    .Y(_1263_));
 sg13g2_a21oi_1 _4566_ (.A1(_1914_),
    .A2(net1024),
    .Y(_1264_),
    .B1(_1263_));
 sg13g2_a22oi_1 _4567_ (.Y(_1265_),
    .B1(_1264_),
    .B2(net1225),
    .A2(_1262_),
    .A1(_1052_));
 sg13g2_nor2_1 _4568_ (.A(net1013),
    .B(_1265_),
    .Y(_1266_));
 sg13g2_a22oi_1 _4569_ (.Y(_1267_),
    .B1(_1259_),
    .B2(_1266_),
    .A2(net1013),
    .A1(net289));
 sg13g2_nor2_1 _4570_ (.A(net1326),
    .B(_1267_),
    .Y(_0140_));
 sg13g2_nand2_1 _4571_ (.Y(_1268_),
    .A(net1315),
    .B(net1049));
 sg13g2_o21ai_1 _4572_ (.B1(_1268_),
    .Y(_1269_),
    .A1(_1898_),
    .A2(net1315));
 sg13g2_nor2_1 _4573_ (.A(net1049),
    .B(net1112),
    .Y(_1270_));
 sg13g2_o21ai_1 _4574_ (.B1(net1167),
    .Y(_1271_),
    .A1(net1114),
    .A2(_1269_));
 sg13g2_nor2_1 _4575_ (.A(_1270_),
    .B(_1271_),
    .Y(_1272_));
 sg13g2_nand2_1 _4576_ (.Y(_1273_),
    .A(_2230_),
    .B(net1050));
 sg13g2_xnor2_1 _4577_ (.Y(_1274_),
    .A(_2230_),
    .B(net1050));
 sg13g2_and2_1 _4578_ (.A(_1213_),
    .B(_1240_),
    .X(_1275_));
 sg13g2_a21o_1 _4579_ (.A2(_1275_),
    .A1(_1217_),
    .B1(_1239_),
    .X(_1276_));
 sg13g2_a21oi_1 _4580_ (.A1(_1217_),
    .A2(_1275_),
    .Y(_1277_),
    .B1(_1239_));
 sg13g2_xnor2_1 _4581_ (.Y(_1278_),
    .A(_1274_),
    .B(_1276_));
 sg13g2_o21ai_1 _4582_ (.B1(_1268_),
    .Y(_1279_),
    .A1(net1315),
    .A2(_1278_));
 sg13g2_a21oi_1 _4583_ (.A1(net1134),
    .A2(_1279_),
    .Y(_1280_),
    .B1(_1272_));
 sg13g2_nor2_1 _4584_ (.A(net1034),
    .B(_1280_),
    .Y(_1281_));
 sg13g2_a22oi_1 _4585_ (.Y(_1282_),
    .B1(_0981_),
    .B2(\cpu_instance.pc[10] ),
    .A2(_0980_),
    .A1(net1049));
 sg13g2_nand2_1 _4586_ (.Y(_1283_),
    .A(net1233),
    .B(_1269_));
 sg13g2_nand3_1 _4587_ (.B(_1282_),
    .C(_1283_),
    .A(net1180),
    .Y(_1284_));
 sg13g2_a21oi_1 _4588_ (.A1(net1200),
    .A2(_0605_),
    .Y(_1285_),
    .B1(net1198));
 sg13g2_o21ai_1 _4589_ (.B1(_1285_),
    .Y(_1286_),
    .A1(_1281_),
    .A2(_1284_));
 sg13g2_a21oi_1 _4590_ (.A1(net1197),
    .A2(_1269_),
    .Y(_1287_),
    .B1(net1118));
 sg13g2_nor2_1 _4591_ (.A(net1049),
    .B(net1068),
    .Y(_1288_));
 sg13g2_a21oi_1 _4592_ (.A1(_1286_),
    .A2(_1287_),
    .Y(_1289_),
    .B1(_1288_));
 sg13g2_nor3_1 _4593_ (.A(net1162),
    .B(net1222),
    .C(_2229_),
    .Y(_1290_));
 sg13g2_a221oi_1 _4594_ (.B2(_1112_),
    .C1(_1290_),
    .B1(net1049),
    .A1(\cpu_instance.ram_data_out[10] ),
    .Y(_1291_),
    .A2(net1176));
 sg13g2_o21ai_1 _4595_ (.B1(_1291_),
    .Y(_1292_),
    .A1(_2063_),
    .A2(_0605_));
 sg13g2_nor2_1 _4596_ (.A(net1049),
    .B(net1024),
    .Y(_1293_));
 sg13g2_o21ai_1 _4597_ (.B1(_1053_),
    .Y(_1294_),
    .A1(\cpu_instance.ram_data_out[10] ),
    .A2(net1032));
 sg13g2_o21ai_1 _4598_ (.B1(net1015),
    .Y(_1295_),
    .A1(_1293_),
    .A2(_1294_));
 sg13g2_a221oi_1 _4599_ (.B2(net1228),
    .C1(_1295_),
    .B1(_1292_),
    .A1(net1241),
    .Y(_1296_),
    .A2(_1289_));
 sg13g2_o21ai_1 _4600_ (.B1(net1331),
    .Y(_1297_),
    .A1(net288),
    .A2(net1015));
 sg13g2_nor2_1 _4601_ (.A(_1296_),
    .B(_1297_),
    .Y(_0141_));
 sg13g2_nor2b_1 _4602_ (.A(net1106),
    .B_N(net1040),
    .Y(_1298_));
 sg13g2_a21oi_1 _4603_ (.A1(\cpu_instance.pc[11] ),
    .A2(net1106),
    .Y(_1299_),
    .B1(_1298_));
 sg13g2_nand2_1 _4604_ (.Y(_1300_),
    .A(_2222_),
    .B(net1041));
 sg13g2_nor2_1 _4605_ (.A(_2222_),
    .B(net1041),
    .Y(_1301_));
 sg13g2_xnor2_1 _4606_ (.Y(_1302_),
    .A(_2222_),
    .B(net1041));
 sg13g2_o21ai_1 _4607_ (.B1(_1273_),
    .Y(_1303_),
    .A1(_1274_),
    .A2(_1276_));
 sg13g2_xor2_1 _4608_ (.B(_1303_),
    .A(_1302_),
    .X(_1304_));
 sg13g2_a21oi_1 _4609_ (.A1(net1315),
    .A2(net1041),
    .Y(_1305_),
    .B1(net1167));
 sg13g2_o21ai_1 _4610_ (.B1(_1305_),
    .Y(_1306_),
    .A1(net1315),
    .A2(_1304_));
 sg13g2_nor2_1 _4611_ (.A(_1897_),
    .B(net1314),
    .Y(_1307_));
 sg13g2_a21oi_1 _4612_ (.A1(net1314),
    .A2(net1040),
    .Y(_1308_),
    .B1(_1307_));
 sg13g2_inv_1 _4613_ (.Y(_1309_),
    .A(_1308_));
 sg13g2_a21oi_1 _4614_ (.A1(net1040),
    .A2(net1114),
    .Y(_1310_),
    .B1(net1134));
 sg13g2_o21ai_1 _4615_ (.B1(_1310_),
    .Y(_1311_),
    .A1(net1114),
    .A2(_1308_));
 sg13g2_nand3_1 _4616_ (.B(_1306_),
    .C(_1311_),
    .A(_0945_),
    .Y(_1312_));
 sg13g2_nand2_1 _4617_ (.Y(_1313_),
    .A(net1190),
    .B(_1299_));
 sg13g2_a22oi_1 _4618_ (.Y(_1314_),
    .B1(_1313_),
    .B2(_0805_),
    .A2(_1309_),
    .A1(net1233));
 sg13g2_a22oi_1 _4619_ (.Y(_1315_),
    .B1(_1312_),
    .B2(_1314_),
    .A2(_1299_),
    .A1(net1183));
 sg13g2_nor2_1 _4620_ (.A(net1200),
    .B(_1315_),
    .Y(_1316_));
 sg13g2_o21ai_1 _4621_ (.B1(net1196),
    .Y(_1317_),
    .A1(net1180),
    .A2(_0613_));
 sg13g2_a21oi_1 _4622_ (.A1(net1197),
    .A2(_1309_),
    .Y(_1318_),
    .B1(_0987_));
 sg13g2_o21ai_1 _4623_ (.B1(_1318_),
    .Y(_1319_),
    .A1(_1316_),
    .A2(_1317_));
 sg13g2_o21ai_1 _4624_ (.B1(_1319_),
    .Y(_1320_),
    .A1(net1040),
    .A2(net1068));
 sg13g2_a22oi_1 _4625_ (.Y(_1321_),
    .B1(net1160),
    .B2(_2222_),
    .A2(_2117_),
    .A1(\cpu_instance.ram_data_out[11] ));
 sg13g2_a22oi_1 _4626_ (.Y(_1322_),
    .B1(_1112_),
    .B2(net1040),
    .A2(_0613_),
    .A1(_2094_));
 sg13g2_nand3_1 _4627_ (.B(_1321_),
    .C(_1322_),
    .A(net1228),
    .Y(_1323_));
 sg13g2_o21ai_1 _4628_ (.B1(net1225),
    .Y(_1324_),
    .A1(_1910_),
    .A2(net1033));
 sg13g2_a21oi_1 _4629_ (.A1(net1040),
    .A2(net1033),
    .Y(_1325_),
    .B1(_1324_));
 sg13g2_nor2_1 _4630_ (.A(net1241),
    .B(_1325_),
    .Y(_1326_));
 sg13g2_a21oi_1 _4631_ (.A1(_1323_),
    .A2(_1326_),
    .Y(_1327_),
    .B1(net1012));
 sg13g2_o21ai_1 _4632_ (.B1(_1327_),
    .Y(_1328_),
    .A1(net1234),
    .A2(_1320_));
 sg13g2_o21ai_1 _4633_ (.B1(net1331),
    .Y(_1329_),
    .A1(net208),
    .A2(net1015));
 sg13g2_nor2b_1 _4634_ (.A(_1329_),
    .B_N(_1328_),
    .Y(_0142_));
 sg13g2_nand2_1 _4635_ (.Y(_1330_),
    .A(net1317),
    .B(_0621_));
 sg13g2_o21ai_1 _4636_ (.B1(_1330_),
    .Y(_1331_),
    .A1(_1896_),
    .A2(net1317));
 sg13g2_o21ai_1 _4637_ (.B1(net1167),
    .Y(_1332_),
    .A1(net1115),
    .A2(_1331_));
 sg13g2_a21oi_1 _4638_ (.A1(_0622_),
    .A2(net1114),
    .Y(_1333_),
    .B1(_1332_));
 sg13g2_nand2_1 _4639_ (.Y(_1334_),
    .A(_2211_),
    .B(_0621_));
 sg13g2_xnor2_1 _4640_ (.Y(_1335_),
    .A(_2211_),
    .B(_0621_));
 sg13g2_nor2_1 _4641_ (.A(_1274_),
    .B(_1302_),
    .Y(_1336_));
 sg13g2_a21oi_1 _4642_ (.A1(_1273_),
    .A2(_1300_),
    .Y(_1337_),
    .B1(_1301_));
 sg13g2_a21oi_2 _4643_ (.B1(_1337_),
    .Y(_1338_),
    .A2(_1336_),
    .A1(_1277_));
 sg13g2_xnor2_1 _4644_ (.Y(_1339_),
    .A(_1335_),
    .B(_1338_));
 sg13g2_o21ai_1 _4645_ (.B1(_1330_),
    .Y(_1340_),
    .A1(net1317),
    .A2(_1339_));
 sg13g2_a21o_1 _4646_ (.A2(_1340_),
    .A1(net1134),
    .B1(_1333_),
    .X(_1341_));
 sg13g2_a22oi_1 _4647_ (.Y(_1342_),
    .B1(_0981_),
    .B2(\cpu_instance.pc[12] ),
    .A2(_0980_),
    .A1(_0621_));
 sg13g2_nand2b_1 _4648_ (.Y(_1343_),
    .B(_1342_),
    .A_N(_2064_));
 sg13g2_a221oi_1 _4649_ (.B2(net1024),
    .C1(_1343_),
    .B1(_1341_),
    .A1(net1233),
    .Y(_1344_),
    .A2(_1331_));
 sg13g2_o21ai_1 _4650_ (.B1(net1196),
    .Y(_1345_),
    .A1(net1180),
    .A2(_0624_));
 sg13g2_a21oi_1 _4651_ (.A1(net1198),
    .A2(_1331_),
    .Y(_1346_),
    .B1(_0987_));
 sg13g2_o21ai_1 _4652_ (.B1(_1346_),
    .Y(_1347_),
    .A1(_1344_),
    .A2(_1345_));
 sg13g2_a21oi_1 _4653_ (.A1(_0622_),
    .A2(net1118),
    .Y(_1348_),
    .B1(net1234));
 sg13g2_nand2_1 _4654_ (.Y(_1349_),
    .A(_1347_),
    .B(_1348_));
 sg13g2_a21oi_1 _4655_ (.A1(\cpu_instance.ram_data_out[12] ),
    .A2(net1176),
    .Y(_1350_),
    .B1(net1160));
 sg13g2_a21oi_1 _4656_ (.A1(net1253),
    .A2(_0622_),
    .Y(_1351_),
    .B1(net1176));
 sg13g2_o21ai_1 _4657_ (.B1(_1351_),
    .Y(_1352_),
    .A1(net1253),
    .A2(_0624_));
 sg13g2_a221oi_1 _4658_ (.B2(_1352_),
    .C1(net1225),
    .B1(_1350_),
    .A1(net1160),
    .Y(_1353_),
    .A2(_2212_));
 sg13g2_o21ai_1 _4659_ (.B1(_1053_),
    .Y(_1354_),
    .A1(\cpu_instance.ram_data_out[12] ),
    .A2(net1032));
 sg13g2_a21oi_1 _4660_ (.A1(_0622_),
    .A2(net1033),
    .Y(_1355_),
    .B1(_1354_));
 sg13g2_nor3_1 _4661_ (.A(net1012),
    .B(_1353_),
    .C(_1355_),
    .Y(_1356_));
 sg13g2_a221oi_1 _4662_ (.B2(_1356_),
    .C1(net1323),
    .B1(_1349_),
    .A1(_1896_),
    .Y(_0143_),
    .A2(net1012));
 sg13g2_nor2_1 _4663_ (.A(net1280),
    .B(_0633_),
    .Y(_1357_));
 sg13g2_xnor2_1 _4664_ (.Y(_1358_),
    .A(_2202_),
    .B(_0632_));
 sg13g2_o21ai_1 _4665_ (.B1(_1334_),
    .Y(_1359_),
    .A1(_1335_),
    .A2(_1338_));
 sg13g2_xnor2_1 _4666_ (.Y(_1360_),
    .A(_1358_),
    .B(_1359_));
 sg13g2_a21o_1 _4667_ (.A2(_1360_),
    .A1(net1280),
    .B1(_1357_),
    .X(_1361_));
 sg13g2_a21oi_1 _4668_ (.A1(\cpu_instance.pc[13] ),
    .A2(net1280),
    .Y(_1362_),
    .B1(_1357_));
 sg13g2_nand2_1 _4669_ (.Y(_1363_),
    .A(_0633_),
    .B(net1114));
 sg13g2_a21oi_1 _4670_ (.A1(net1112),
    .A2(_1362_),
    .Y(_1364_),
    .B1(net1135));
 sg13g2_a22oi_1 _4671_ (.Y(_1365_),
    .B1(_1363_),
    .B2(_1364_),
    .A2(_1361_),
    .A1(net1134));
 sg13g2_nand2_1 _4672_ (.Y(_1366_),
    .A(\cpu_instance.pc[13] ),
    .B(net1107));
 sg13g2_o21ai_1 _4673_ (.B1(_1366_),
    .Y(_1367_),
    .A1(net1106),
    .A2(_0633_));
 sg13g2_o21ai_1 _4674_ (.B1(net1190),
    .Y(_1368_),
    .A1(_2083_),
    .A2(_1362_));
 sg13g2_a21oi_1 _4675_ (.A1(net1067),
    .A2(_1367_),
    .Y(_1369_),
    .B1(_1368_));
 sg13g2_o21ai_1 _4676_ (.B1(_1369_),
    .Y(_1370_),
    .A1(_0946_),
    .A2(_1365_));
 sg13g2_o21ai_1 _4677_ (.B1(_2053_),
    .Y(_1371_),
    .A1(net1190),
    .A2(_1367_));
 sg13g2_nor2b_1 _4678_ (.A(_1371_),
    .B_N(_1370_),
    .Y(_1372_));
 sg13g2_o21ai_1 _4679_ (.B1(net1196),
    .Y(_1373_),
    .A1(net1180),
    .A2(_0635_));
 sg13g2_a21oi_1 _4680_ (.A1(net1197),
    .A2(_1362_),
    .Y(_1374_),
    .B1(_0987_));
 sg13g2_o21ai_1 _4681_ (.B1(_1374_),
    .Y(_1375_),
    .A1(_1372_),
    .A2(_1373_));
 sg13g2_a21oi_1 _4682_ (.A1(_0632_),
    .A2(net1118),
    .Y(_1376_),
    .B1(net1235));
 sg13g2_nor2_1 _4683_ (.A(net1162),
    .B(_2203_),
    .Y(_1377_));
 sg13g2_a221oi_1 _4684_ (.B2(_1112_),
    .C1(_1377_),
    .B1(_0632_),
    .A1(\cpu_instance.ram_data_out[13] ),
    .Y(_1378_),
    .A2(net1176));
 sg13g2_o21ai_1 _4685_ (.B1(_1378_),
    .Y(_1379_),
    .A1(_2095_),
    .A2(_0635_));
 sg13g2_nand2_1 _4686_ (.Y(_1380_),
    .A(net1229),
    .B(_1379_));
 sg13g2_o21ai_1 _4687_ (.B1(net1225),
    .Y(_1381_),
    .A1(\cpu_instance.ram_data_out[13] ),
    .A2(net1032));
 sg13g2_a21oi_1 _4688_ (.A1(_0633_),
    .A2(net1032),
    .Y(_1382_),
    .B1(_1381_));
 sg13g2_nor2_1 _4689_ (.A(net1241),
    .B(_1382_),
    .Y(_1383_));
 sg13g2_a221oi_1 _4690_ (.B2(_1383_),
    .C1(net1013),
    .B1(_1380_),
    .A1(_1375_),
    .Y(_1384_),
    .A2(_1376_));
 sg13g2_a21oi_1 _4691_ (.A1(net272),
    .A2(net1012),
    .Y(_1385_),
    .B1(_1384_));
 sg13g2_nor2_1 _4692_ (.A(net1323),
    .B(_1385_),
    .Y(_0144_));
 sg13g2_nand2_1 _4693_ (.Y(_1386_),
    .A(\cpu_instance.pc[14] ),
    .B(net1106));
 sg13g2_o21ai_1 _4694_ (.B1(_1386_),
    .Y(_1387_),
    .A1(net1106),
    .A2(_0643_));
 sg13g2_nor2_1 _4695_ (.A(net1280),
    .B(_0643_),
    .Y(_1388_));
 sg13g2_or2_1 _4696_ (.X(_1389_),
    .B(_1358_),
    .A(_1335_));
 sg13g2_a21oi_1 _4697_ (.A1(_2203_),
    .A2(_0633_),
    .Y(_1390_),
    .B1(_1334_));
 sg13g2_a21oi_1 _4698_ (.A1(_2202_),
    .A2(_0632_),
    .Y(_1391_),
    .B1(_1390_));
 sg13g2_o21ai_1 _4699_ (.B1(_1391_),
    .Y(_1392_),
    .A1(_1338_),
    .A2(_1389_));
 sg13g2_and2_1 _4700_ (.A(_2192_),
    .B(_0642_),
    .X(_1393_));
 sg13g2_nand2b_1 _4701_ (.Y(_1394_),
    .B(_0643_),
    .A_N(_2192_));
 sg13g2_nand2b_1 _4702_ (.Y(_1395_),
    .B(_1394_),
    .A_N(_1393_));
 sg13g2_xnor2_1 _4703_ (.Y(_1396_),
    .A(_1392_),
    .B(_1395_));
 sg13g2_a21o_1 _4704_ (.A2(_1396_),
    .A1(net1280),
    .B1(_1388_),
    .X(_1397_));
 sg13g2_a21oi_2 _4705_ (.B1(_1388_),
    .Y(_1398_),
    .A2(net1280),
    .A1(\cpu_instance.pc[14] ));
 sg13g2_nand2_1 _4706_ (.Y(_1399_),
    .A(_0643_),
    .B(net1114));
 sg13g2_a21oi_1 _4707_ (.A1(net1112),
    .A2(_1398_),
    .Y(_1400_),
    .B1(net1134));
 sg13g2_a22oi_1 _4708_ (.Y(_1401_),
    .B1(_1399_),
    .B2(_1400_),
    .A2(_1397_),
    .A1(net1134));
 sg13g2_nand2b_1 _4709_ (.Y(_1402_),
    .B(net1233),
    .A_N(_1398_));
 sg13g2_o21ai_1 _4710_ (.B1(_1402_),
    .Y(_1403_),
    .A1(_0946_),
    .A2(_1401_));
 sg13g2_o21ai_1 _4711_ (.B1(_1403_),
    .Y(_1404_),
    .A1(net1190),
    .A2(_1387_));
 sg13g2_a21oi_1 _4712_ (.A1(_0805_),
    .A2(_1387_),
    .Y(_1405_),
    .B1(net1200));
 sg13g2_nand2_1 _4713_ (.Y(_1406_),
    .A(_1404_),
    .B(_1405_));
 sg13g2_a21oi_1 _4714_ (.A1(_2064_),
    .A2(_0644_),
    .Y(_1407_),
    .B1(net1197));
 sg13g2_o21ai_1 _4715_ (.B1(net1068),
    .Y(_1408_),
    .A1(net1196),
    .A2(_1398_));
 sg13g2_a21o_1 _4716_ (.A2(_1407_),
    .A1(_1406_),
    .B1(_1408_),
    .X(_1409_));
 sg13g2_a21oi_1 _4717_ (.A1(_0643_),
    .A2(net1118),
    .Y(_1410_),
    .B1(net1234));
 sg13g2_a21oi_1 _4718_ (.A1(_0643_),
    .A2(net1032),
    .Y(_1411_),
    .B1(net1228));
 sg13g2_o21ai_1 _4719_ (.B1(_1411_),
    .Y(_1412_),
    .A1(\cpu_instance.ram_data_out[14] ),
    .A2(net1032));
 sg13g2_o21ai_1 _4720_ (.B1(net1228),
    .Y(_1413_),
    .A1(net1162),
    .A2(_2192_));
 sg13g2_nand2_1 _4721_ (.Y(_1414_),
    .A(_2050_),
    .B(_0644_));
 sg13g2_a21oi_1 _4722_ (.A1(net1253),
    .A2(_0643_),
    .Y(_1415_),
    .B1(net1176));
 sg13g2_a221oi_1 _4723_ (.B2(_1415_),
    .C1(net1160),
    .B1(_1414_),
    .A1(\cpu_instance.ram_data_out[14] ),
    .Y(_1416_),
    .A2(net1176));
 sg13g2_o21ai_1 _4724_ (.B1(_1412_),
    .Y(_1417_),
    .A1(_1413_),
    .A2(_1416_));
 sg13g2_a221oi_1 _4725_ (.B2(net1234),
    .C1(net1012),
    .B1(_1417_),
    .A1(_1409_),
    .Y(_1418_),
    .A2(_1410_));
 sg13g2_o21ai_1 _4726_ (.B1(net1331),
    .Y(_1419_),
    .A1(net274),
    .A2(net1015));
 sg13g2_nor2_1 _4727_ (.A(_1418_),
    .B(_1419_),
    .Y(_0145_));
 sg13g2_mux2_1 _4728_ (.A0(net1017),
    .A1(\cpu_instance.pc[15] ),
    .S(net1106),
    .X(_1420_));
 sg13g2_nand2_1 _4729_ (.Y(_1421_),
    .A(net1317),
    .B(net1018));
 sg13g2_nor2b_1 _4730_ (.A(net1316),
    .B_N(\cpu_instance.pc[15] ),
    .Y(_1422_));
 sg13g2_a21oi_2 _4731_ (.B1(_1422_),
    .Y(_1423_),
    .A2(net1017),
    .A1(net1316));
 sg13g2_o21ai_1 _4732_ (.B1(net1167),
    .Y(_1424_),
    .A1(net1017),
    .A2(net1112));
 sg13g2_a21oi_1 _4733_ (.A1(net1112),
    .A2(_1423_),
    .Y(_1425_),
    .B1(_1424_));
 sg13g2_a21oi_1 _4734_ (.A1(_1392_),
    .A2(_1394_),
    .Y(_1426_),
    .B1(_1393_));
 sg13g2_xnor2_1 _4735_ (.Y(_1427_),
    .A(_2180_),
    .B(net1017));
 sg13g2_xnor2_1 _4736_ (.Y(_1428_),
    .A(_1426_),
    .B(_1427_));
 sg13g2_o21ai_1 _4737_ (.B1(_1421_),
    .Y(_1429_),
    .A1(net1317),
    .A2(_1428_));
 sg13g2_a21oi_1 _4738_ (.A1(net1134),
    .A2(_1429_),
    .Y(_1430_),
    .B1(_1425_));
 sg13g2_o21ai_1 _4739_ (.B1(net1190),
    .Y(_1431_),
    .A1(_2083_),
    .A2(_1423_));
 sg13g2_a21oi_1 _4740_ (.A1(net1067),
    .A2(_1420_),
    .Y(_1432_),
    .B1(_1431_));
 sg13g2_o21ai_1 _4741_ (.B1(_1432_),
    .Y(_1433_),
    .A1(_0946_),
    .A2(_1430_));
 sg13g2_o21ai_1 _4742_ (.B1(_1433_),
    .Y(_1434_),
    .A1(net1190),
    .A2(_1420_));
 sg13g2_o21ai_1 _4743_ (.B1(net1196),
    .Y(_1435_),
    .A1(_2053_),
    .A2(_0650_));
 sg13g2_a21oi_1 _4744_ (.A1(net1180),
    .A2(_1434_),
    .Y(_1436_),
    .B1(_1435_));
 sg13g2_o21ai_1 _4745_ (.B1(net1068),
    .Y(_1437_),
    .A1(net1196),
    .A2(_1423_));
 sg13g2_nor2_1 _4746_ (.A(_1436_),
    .B(_1437_),
    .Y(_1438_));
 sg13g2_nor2_1 _4747_ (.A(net1017),
    .B(net1068),
    .Y(_1439_));
 sg13g2_o21ai_1 _4748_ (.B1(net1242),
    .Y(_1440_),
    .A1(_1438_),
    .A2(_1439_));
 sg13g2_a22oi_1 _4749_ (.Y(_1441_),
    .B1(net1160),
    .B2(_2180_),
    .A2(net1177),
    .A1(\cpu_instance.ram_data_out[15] ));
 sg13g2_inv_1 _4750_ (.Y(_1442_),
    .A(_1441_));
 sg13g2_a221oi_1 _4751_ (.B2(net1017),
    .C1(_1442_),
    .B1(_1112_),
    .A1(_2050_),
    .Y(_1443_),
    .A2(_0650_));
 sg13g2_o21ai_1 _4752_ (.B1(net1225),
    .Y(_1444_),
    .A1(net1017),
    .A2(net1024));
 sg13g2_nand2_1 _4753_ (.Y(_1445_),
    .A(net1235),
    .B(_1444_));
 sg13g2_o21ai_1 _4754_ (.B1(_1445_),
    .Y(_1446_),
    .A1(_2181_),
    .A2(net1033));
 sg13g2_o21ai_1 _4755_ (.B1(_1446_),
    .Y(_1447_),
    .A1(net1225),
    .A2(_1443_));
 sg13g2_and2_1 _4756_ (.A(net1015),
    .B(_1447_),
    .X(_1448_));
 sg13g2_a22oi_1 _4757_ (.Y(_1449_),
    .B1(_1440_),
    .B2(_1448_),
    .A2(net1013),
    .A1(net270));
 sg13g2_nor2_1 _4758_ (.A(net1323),
    .B(_1449_),
    .Y(_0146_));
 sg13g2_nor2_2 _4759_ (.A(net1301),
    .B(_0954_),
    .Y(_1450_));
 sg13g2_nand2_2 _4760_ (.Y(_1451_),
    .A(_1915_),
    .B(_0955_));
 sg13g2_nor2_1 _4761_ (.A(net1301),
    .B(_0041_),
    .Y(_1452_));
 sg13g2_a21oi_1 _4762_ (.A1(net1302),
    .A2(net1320),
    .Y(_1453_),
    .B1(_1452_));
 sg13g2_and4_2 _4763_ (.A(_0012_),
    .B(_1976_),
    .C(_0955_),
    .D(_1453_),
    .X(_1454_));
 sg13g2_nand4_1 _4764_ (.B(_1976_),
    .C(_0955_),
    .A(_0012_),
    .Y(_1455_),
    .D(_1453_));
 sg13g2_o21ai_1 _4765_ (.B1(net1334),
    .Y(_1456_),
    .A1(net224),
    .A2(_1454_));
 sg13g2_nand2_1 _4766_ (.Y(_1457_),
    .A(\cpu_instance.accum[0] ),
    .B(_1450_));
 sg13g2_a21oi_1 _4767_ (.A1(net1311),
    .A2(_1451_),
    .Y(_1458_),
    .B1(_1455_));
 sg13g2_a21oi_1 _4768_ (.A1(_1457_),
    .A2(_1458_),
    .Y(_0147_),
    .B1(net225));
 sg13g2_o21ai_1 _4769_ (.B1(net1334),
    .Y(_1459_),
    .A1(net227),
    .A2(_1454_));
 sg13g2_nand2_1 _4770_ (.Y(_1460_),
    .A(\cpu_instance.accum[1] ),
    .B(_1450_));
 sg13g2_a21oi_1 _4771_ (.A1(\cpu_instance.accum[9] ),
    .A2(_1451_),
    .Y(_1461_),
    .B1(_1455_));
 sg13g2_a21oi_1 _4772_ (.A1(_1460_),
    .A2(_1461_),
    .Y(_0148_),
    .B1(net228));
 sg13g2_o21ai_1 _4773_ (.B1(net1334),
    .Y(_1462_),
    .A1(net230),
    .A2(_1454_));
 sg13g2_nand2_1 _4774_ (.Y(_1463_),
    .A(\cpu_instance.accum[2] ),
    .B(_1450_));
 sg13g2_a21oi_1 _4775_ (.A1(net1308),
    .A2(_1451_),
    .Y(_1464_),
    .B1(_1455_));
 sg13g2_a21oi_1 _4776_ (.A1(_1463_),
    .A2(_1464_),
    .Y(_0149_),
    .B1(net231));
 sg13g2_o21ai_1 _4777_ (.B1(net1334),
    .Y(_1465_),
    .A1(net236),
    .A2(_1454_));
 sg13g2_nand2_1 _4778_ (.Y(_1466_),
    .A(\cpu_instance.accum[3] ),
    .B(_1450_));
 sg13g2_a21oi_1 _4779_ (.A1(\cpu_instance.accum[11] ),
    .A2(_1451_),
    .Y(_1467_),
    .B1(_1455_));
 sg13g2_a21oi_1 _4780_ (.A1(_1466_),
    .A2(_1467_),
    .Y(_0150_),
    .B1(net237));
 sg13g2_o21ai_1 _4781_ (.B1(net1334),
    .Y(_1468_),
    .A1(net233),
    .A2(_1454_));
 sg13g2_nand2_1 _4782_ (.Y(_1469_),
    .A(\cpu_instance.accum[4] ),
    .B(_1450_));
 sg13g2_a21oi_1 _4783_ (.A1(\cpu_instance.accum[12] ),
    .A2(_1451_),
    .Y(_1470_),
    .B1(_1455_));
 sg13g2_a21oi_1 _4784_ (.A1(_1469_),
    .A2(_1470_),
    .Y(_0151_),
    .B1(net234));
 sg13g2_o21ai_1 _4785_ (.B1(net1334),
    .Y(_1471_),
    .A1(net241),
    .A2(_1454_));
 sg13g2_nand2_1 _4786_ (.Y(_1472_),
    .A(\cpu_instance.accum[5] ),
    .B(_1450_));
 sg13g2_a21oi_1 _4787_ (.A1(\cpu_instance.accum[13] ),
    .A2(_1451_),
    .Y(_1473_),
    .B1(_1455_));
 sg13g2_a21oi_1 _4788_ (.A1(_1472_),
    .A2(_1473_),
    .Y(_0152_),
    .B1(net242));
 sg13g2_o21ai_1 _4789_ (.B1(net1334),
    .Y(_1474_),
    .A1(net211),
    .A2(_1454_));
 sg13g2_nand2_1 _4790_ (.Y(_1475_),
    .A(\cpu_instance.accum[6] ),
    .B(_1450_));
 sg13g2_a21oi_1 _4791_ (.A1(\cpu_instance.accum[14] ),
    .A2(_1451_),
    .Y(_1476_),
    .B1(_1455_));
 sg13g2_a21oi_1 _4792_ (.A1(_1475_),
    .A2(_1476_),
    .Y(_0153_),
    .B1(net212));
 sg13g2_o21ai_1 _4793_ (.B1(net1333),
    .Y(_1477_),
    .A1(net204),
    .A2(_1454_));
 sg13g2_nand2_1 _4794_ (.Y(_1478_),
    .A(\cpu_instance.accum[7] ),
    .B(_1450_));
 sg13g2_a21oi_1 _4795_ (.A1(\cpu_instance.accum[15] ),
    .A2(_1451_),
    .Y(_1479_),
    .B1(_1455_));
 sg13g2_a21oi_1 _4796_ (.A1(_1478_),
    .A2(_1479_),
    .Y(_0154_),
    .B1(net205));
 sg13g2_nand4_1 _4797_ (.B(_2093_),
    .C(_2109_),
    .A(net1195),
    .Y(_1480_),
    .D(net1116));
 sg13g2_o21ai_1 _4798_ (.B1(_1052_),
    .Y(_1481_),
    .A1(net1273),
    .A2(net1226));
 sg13g2_or2_1 _4799_ (.X(_1482_),
    .B(_0692_),
    .A(_2077_));
 sg13g2_nor3_1 _4800_ (.A(_2130_),
    .B(_2152_),
    .C(_1481_),
    .Y(_1483_));
 sg13g2_nand3_1 _4801_ (.B(_1482_),
    .C(_1483_),
    .A(_2155_),
    .Y(_1484_));
 sg13g2_nor2_1 _4802_ (.A(_2157_),
    .B(_1484_),
    .Y(_1485_));
 sg13g2_and3_2 _4803_ (.X(_1486_),
    .A(_0950_),
    .B(_1480_),
    .C(_1485_));
 sg13g2_nand3_1 _4804_ (.B(_1480_),
    .C(_1485_),
    .A(_0950_),
    .Y(_1487_));
 sg13g2_o21ai_1 _4805_ (.B1(net1327),
    .Y(_1488_),
    .A1(net1283),
    .A2(net1031));
 sg13g2_a21oi_1 _4806_ (.A1(_1893_),
    .A2(net1031),
    .Y(_0155_),
    .B1(_1488_));
 sg13g2_xnor2_1 _4807_ (.Y(_1489_),
    .A(\cpu_instance.sp[2] ),
    .B(net1283));
 sg13g2_xor2_1 _4808_ (.B(_1489_),
    .A(net1166),
    .X(_1490_));
 sg13g2_o21ai_1 _4809_ (.B1(net1327),
    .Y(_1491_),
    .A1(net316),
    .A2(net1031));
 sg13g2_a21oi_1 _4810_ (.A1(net1031),
    .A2(_1490_),
    .Y(_0156_),
    .B1(_1491_));
 sg13g2_nor3_2 _4811_ (.A(\cpu_instance.sp[3] ),
    .B(\cpu_instance.sp[2] ),
    .C(net1283),
    .Y(_1492_));
 sg13g2_o21ai_1 _4812_ (.B1(\cpu_instance.sp[3] ),
    .Y(_1493_),
    .A1(\cpu_instance.sp[2] ),
    .A2(net1283));
 sg13g2_nor2b_1 _4813_ (.A(_1492_),
    .B_N(_1493_),
    .Y(_1494_));
 sg13g2_nand3_1 _4814_ (.B(\cpu_instance.sp[2] ),
    .C(net1283),
    .A(\cpu_instance.sp[3] ),
    .Y(_1495_));
 sg13g2_a21o_1 _4815_ (.A2(net1283),
    .A1(\cpu_instance.sp[2] ),
    .B1(\cpu_instance.sp[3] ),
    .X(_1496_));
 sg13g2_and2_1 _4816_ (.A(_1495_),
    .B(_1496_),
    .X(_1497_));
 sg13g2_nand2_1 _4817_ (.Y(_1498_),
    .A(net1164),
    .B(_1494_));
 sg13g2_o21ai_1 _4818_ (.B1(_1498_),
    .Y(_1499_),
    .A1(net1165),
    .A2(_1497_));
 sg13g2_o21ai_1 _4819_ (.B1(net1327),
    .Y(_1500_),
    .A1(net302),
    .A2(net1030));
 sg13g2_a21oi_1 _4820_ (.A1(net1030),
    .A2(_1499_),
    .Y(_0157_),
    .B1(_1500_));
 sg13g2_nand4_1 _4821_ (.B(\cpu_instance.sp[3] ),
    .C(\cpu_instance.sp[2] ),
    .A(\cpu_instance.sp[4] ),
    .Y(_1501_),
    .D(net1283));
 sg13g2_inv_1 _4822_ (.Y(_1502_),
    .A(_1501_));
 sg13g2_nor2b_1 _4823_ (.A(net280),
    .B_N(_1495_),
    .Y(_1503_));
 sg13g2_nor2b_2 _4824_ (.A(\cpu_instance.sp[4] ),
    .B_N(_1492_),
    .Y(_1504_));
 sg13g2_xor2_1 _4825_ (.B(_1492_),
    .A(\cpu_instance.sp[4] ),
    .X(_1505_));
 sg13g2_nor3_1 _4826_ (.A(net1164),
    .B(_1502_),
    .C(_1503_),
    .Y(_1506_));
 sg13g2_a21oi_1 _4827_ (.A1(net1164),
    .A2(_1505_),
    .Y(_1507_),
    .B1(_1506_));
 sg13g2_o21ai_1 _4828_ (.B1(net1327),
    .Y(_1508_),
    .A1(net280),
    .A2(net1031));
 sg13g2_a21oi_1 _4829_ (.A1(net1031),
    .A2(_1507_),
    .Y(_0158_),
    .B1(_1508_));
 sg13g2_xor2_1 _4830_ (.B(_1501_),
    .A(\cpu_instance.sp[5] ),
    .X(_1509_));
 sg13g2_nand2_1 _4831_ (.Y(_1510_),
    .A(_0007_),
    .B(_1504_));
 sg13g2_xnor2_1 _4832_ (.Y(_1511_),
    .A(_0007_),
    .B(_1504_));
 sg13g2_nor2_1 _4833_ (.A(net1164),
    .B(_1509_),
    .Y(_1512_));
 sg13g2_a21oi_1 _4834_ (.A1(net1164),
    .A2(_1511_),
    .Y(_1513_),
    .B1(_1512_));
 sg13g2_o21ai_1 _4835_ (.B1(net1327),
    .Y(_1514_),
    .A1(net291),
    .A2(net1030));
 sg13g2_a21oi_1 _4836_ (.A1(net1030),
    .A2(_1513_),
    .Y(_0159_),
    .B1(_1514_));
 sg13g2_xor2_1 _4837_ (.B(_1510_),
    .A(\cpu_instance.sp[6] ),
    .X(_1515_));
 sg13g2_nor2_1 _4838_ (.A(_0007_),
    .B(_1501_),
    .Y(_1516_));
 sg13g2_xor2_1 _4839_ (.B(_1516_),
    .A(\cpu_instance.sp[6] ),
    .X(_1517_));
 sg13g2_nand2_1 _4840_ (.Y(_1518_),
    .A(net1164),
    .B(_1515_));
 sg13g2_o21ai_1 _4841_ (.B1(_1518_),
    .Y(_1519_),
    .A1(net1164),
    .A2(_1517_));
 sg13g2_o21ai_1 _4842_ (.B1(net1327),
    .Y(_1520_),
    .A1(net287),
    .A2(net1030));
 sg13g2_a21oi_1 _4843_ (.A1(net1030),
    .A2(_1519_),
    .Y(_0160_),
    .B1(_1520_));
 sg13g2_nor2_1 _4844_ (.A(\cpu_instance.sp[6] ),
    .B(\cpu_instance.sp[5] ),
    .Y(_1521_));
 sg13g2_and2_1 _4845_ (.A(_1504_),
    .B(_1521_),
    .X(_1522_));
 sg13g2_nor2b_1 _4846_ (.A(\cpu_instance.sp[7] ),
    .B_N(_1522_),
    .Y(_1523_));
 sg13g2_xnor2_1 _4847_ (.Y(_1524_),
    .A(\cpu_instance.sp[7] ),
    .B(_1522_));
 sg13g2_and3_1 _4848_ (.X(_1525_),
    .A(\cpu_instance.sp[6] ),
    .B(\cpu_instance.sp[5] ),
    .C(_1502_));
 sg13g2_a21oi_1 _4849_ (.A1(\cpu_instance.sp[7] ),
    .A2(_1525_),
    .Y(_1526_),
    .B1(net1164));
 sg13g2_o21ai_1 _4850_ (.B1(_1526_),
    .Y(_1527_),
    .A1(\cpu_instance.sp[7] ),
    .A2(_1525_));
 sg13g2_o21ai_1 _4851_ (.B1(_1527_),
    .Y(_1528_),
    .A1(net1132),
    .A2(_1524_));
 sg13g2_nor2_1 _4852_ (.A(net1029),
    .B(_1528_),
    .Y(_1529_));
 sg13g2_nor2_1 _4853_ (.A(net286),
    .B(net1030),
    .Y(_1530_));
 sg13g2_nor3_1 _4854_ (.A(net1322),
    .B(_1529_),
    .C(_1530_),
    .Y(_0161_));
 sg13g2_o21ai_1 _4855_ (.B1(_1892_),
    .Y(_1531_),
    .A1(net1029),
    .A2(_1526_));
 sg13g2_nand3_1 _4856_ (.B(\cpu_instance.sp[7] ),
    .C(_1525_),
    .A(\cpu_instance.sp[8] ),
    .Y(_1532_));
 sg13g2_a21o_1 _4857_ (.A2(_1532_),
    .A1(net1132),
    .B1(net1029),
    .X(_1533_));
 sg13g2_and2_1 _4858_ (.A(_1892_),
    .B(_1523_),
    .X(_1534_));
 sg13g2_xnor2_1 _4859_ (.Y(_1535_),
    .A(_1892_),
    .B(_1523_));
 sg13g2_a21oi_1 _4860_ (.A1(net1166),
    .A2(_1535_),
    .Y(_1536_),
    .B1(_1533_));
 sg13g2_nand2_1 _4861_ (.Y(_1537_),
    .A(net1330),
    .B(_1531_));
 sg13g2_nor2_1 _4862_ (.A(_1536_),
    .B(_1537_),
    .Y(_0162_));
 sg13g2_nor2_1 _4863_ (.A(_1891_),
    .B(_1532_),
    .Y(_1538_));
 sg13g2_o21ai_1 _4864_ (.B1(net1030),
    .Y(_1539_),
    .A1(net1165),
    .A2(_1538_));
 sg13g2_nand2_1 _4865_ (.Y(_1540_),
    .A(_0004_),
    .B(_1534_));
 sg13g2_xnor2_1 _4866_ (.Y(_1541_),
    .A(_0004_),
    .B(_1534_));
 sg13g2_and2_1 _4867_ (.A(net1165),
    .B(_1541_),
    .X(_1542_));
 sg13g2_o21ai_1 _4868_ (.B1(net1327),
    .Y(_1543_),
    .A1(_1539_),
    .A2(_1542_));
 sg13g2_a21oi_1 _4869_ (.A1(_1891_),
    .A2(_1533_),
    .Y(_0163_),
    .B1(_1543_));
 sg13g2_a21oi_1 _4870_ (.A1(net263),
    .A2(net1132),
    .Y(_1544_),
    .B1(_1533_));
 sg13g2_xnor2_1 _4871_ (.Y(_1545_),
    .A(_1890_),
    .B(_1540_));
 sg13g2_nor2_1 _4872_ (.A(net1132),
    .B(_1545_),
    .Y(_1546_));
 sg13g2_a21oi_1 _4873_ (.A1(_1890_),
    .A2(net1133),
    .Y(_1547_),
    .B1(_1546_));
 sg13g2_o21ai_1 _4874_ (.B1(net1327),
    .Y(_1548_),
    .A1(\cpu_instance.sp[10] ),
    .A2(_1544_));
 sg13g2_a21oi_1 _4875_ (.A1(_1544_),
    .A2(_1547_),
    .Y(_0164_),
    .B1(_1548_));
 sg13g2_a21oi_1 _4876_ (.A1(_1890_),
    .A2(net1133),
    .Y(_1549_),
    .B1(_1539_));
 sg13g2_nand3_1 _4877_ (.B(\cpu_instance.sp[10] ),
    .C(_1538_),
    .A(\cpu_instance.sp[11] ),
    .Y(_1550_));
 sg13g2_a21oi_1 _4878_ (.A1(net1133),
    .A2(_1550_),
    .Y(_1551_),
    .B1(net1029));
 sg13g2_and3_1 _4879_ (.X(_1552_),
    .A(_1890_),
    .B(_1891_),
    .C(_1534_));
 sg13g2_nor2b_1 _4880_ (.A(\cpu_instance.sp[11] ),
    .B_N(_1552_),
    .Y(_1553_));
 sg13g2_xnor2_1 _4881_ (.Y(_1554_),
    .A(\cpu_instance.sp[11] ),
    .B(_1552_));
 sg13g2_o21ai_1 _4882_ (.B1(_1551_),
    .Y(_1555_),
    .A1(net1132),
    .A2(_1554_));
 sg13g2_o21ai_1 _4883_ (.B1(_1555_),
    .Y(_1556_),
    .A1(net311),
    .A2(_1549_));
 sg13g2_nor2_1 _4884_ (.A(net1322),
    .B(_1556_),
    .Y(_0165_));
 sg13g2_nor2_1 _4885_ (.A(_1889_),
    .B(_1550_),
    .Y(_1557_));
 sg13g2_or2_1 _4886_ (.X(_1558_),
    .B(_1550_),
    .A(_1889_));
 sg13g2_a21oi_1 _4887_ (.A1(net1133),
    .A2(_1558_),
    .Y(_1559_),
    .B1(net1029));
 sg13g2_and2_1 _4888_ (.A(_1889_),
    .B(_1553_),
    .X(_1560_));
 sg13g2_inv_1 _4889_ (.Y(_1561_),
    .A(_1560_));
 sg13g2_xnor2_1 _4890_ (.Y(_1562_),
    .A(\cpu_instance.sp[12] ),
    .B(_1553_));
 sg13g2_o21ai_1 _4891_ (.B1(_1559_),
    .Y(_1563_),
    .A1(net1132),
    .A2(_1562_));
 sg13g2_o21ai_1 _4892_ (.B1(_1563_),
    .Y(_1564_),
    .A1(net261),
    .A2(_1551_));
 sg13g2_nor2_1 _4893_ (.A(net1322),
    .B(_1564_),
    .Y(_0166_));
 sg13g2_nand2_1 _4894_ (.Y(_1565_),
    .A(_0001_),
    .B(_1560_));
 sg13g2_xor2_1 _4895_ (.B(_1560_),
    .A(_0001_),
    .X(_1566_));
 sg13g2_inv_1 _4896_ (.Y(_1567_),
    .A(_1566_));
 sg13g2_a21oi_1 _4897_ (.A1(net256),
    .A2(_1557_),
    .Y(_1568_),
    .B1(net1165));
 sg13g2_a21oi_1 _4898_ (.A1(net1165),
    .A2(_1567_),
    .Y(_1569_),
    .B1(_1568_));
 sg13g2_o21ai_1 _4899_ (.B1(net1330),
    .Y(_1570_),
    .A1(net256),
    .A2(_1559_));
 sg13g2_a21oi_1 _4900_ (.A1(net1031),
    .A2(_1569_),
    .Y(_0167_),
    .B1(_1570_));
 sg13g2_nor2_1 _4901_ (.A(_0001_),
    .B(_1558_),
    .Y(_1571_));
 sg13g2_xnor2_1 _4902_ (.Y(_1572_),
    .A(\cpu_instance.sp[14] ),
    .B(_1571_));
 sg13g2_xor2_1 _4903_ (.B(_1565_),
    .A(\cpu_instance.sp[14] ),
    .X(_1573_));
 sg13g2_nand2_1 _4904_ (.Y(_1574_),
    .A(net1165),
    .B(_1573_));
 sg13g2_a21oi_1 _4905_ (.A1(net1132),
    .A2(_1572_),
    .Y(_1575_),
    .B1(net1029));
 sg13g2_a22oi_1 _4906_ (.Y(_1576_),
    .B1(_1574_),
    .B2(_1575_),
    .A2(net1029),
    .A1(net273));
 sg13g2_nor2_1 _4907_ (.A(net1322),
    .B(_1576_),
    .Y(_0168_));
 sg13g2_nand3_1 _4908_ (.B(\cpu_instance.sp[13] ),
    .C(_1557_),
    .A(\cpu_instance.sp[14] ),
    .Y(_1577_));
 sg13g2_xor2_1 _4909_ (.B(_1577_),
    .A(\cpu_instance.sp[15] ),
    .X(_1578_));
 sg13g2_nor3_1 _4910_ (.A(\cpu_instance.sp[14] ),
    .B(\cpu_instance.sp[13] ),
    .C(_1561_),
    .Y(_1579_));
 sg13g2_xnor2_1 _4911_ (.Y(_1580_),
    .A(\cpu_instance.sp[15] ),
    .B(_1579_));
 sg13g2_nand2_1 _4912_ (.Y(_1581_),
    .A(net1165),
    .B(_1580_));
 sg13g2_a21oi_1 _4913_ (.A1(net1132),
    .A2(_1578_),
    .Y(_1582_),
    .B1(net1029));
 sg13g2_a22oi_1 _4914_ (.Y(_1583_),
    .B1(_1581_),
    .B2(_1582_),
    .A2(_1487_),
    .A1(net279));
 sg13g2_nor2_1 _4915_ (.A(net1322),
    .B(_1583_),
    .Y(_0169_));
 sg13g2_nor2_1 _4916_ (.A(_1985_),
    .B(net1048),
    .Y(_1584_));
 sg13g2_nand2_2 _4917_ (.Y(_1585_),
    .A(net1276),
    .B(net1036));
 sg13g2_nand3_1 _4918_ (.B(\cpu_instance.dp[0] ),
    .C(net1213),
    .A(_1913_),
    .Y(_1586_));
 sg13g2_nor4_2 _4919_ (.A(net1269),
    .B(_2345_),
    .C(_2353_),
    .Y(_1587_),
    .D(_1586_));
 sg13g2_nor2b_1 _4920_ (.A(net1297),
    .B_N(\cpu_instance.dp[1] ),
    .Y(_1588_));
 sg13g2_a21oi_1 _4921_ (.A1(\cpu_instance.sp[1] ),
    .A2(net1297),
    .Y(_1589_),
    .B1(_1588_));
 sg13g2_nor2_2 _4922_ (.A(net1214),
    .B(_1589_),
    .Y(_1590_));
 sg13g2_and3_1 _4923_ (.X(_1591_),
    .A(_2337_),
    .B(_2338_),
    .C(_1590_));
 sg13g2_a21o_1 _4924_ (.A2(_2338_),
    .A1(_2337_),
    .B1(_1590_),
    .X(_1592_));
 sg13g2_nor2b_1 _4925_ (.A(_1591_),
    .B_N(_1592_),
    .Y(_1593_));
 sg13g2_a21oi_1 _4926_ (.A1(_1587_),
    .A2(_1593_),
    .Y(_1594_),
    .B1(_0505_));
 sg13g2_o21ai_1 _4927_ (.B1(_1594_),
    .Y(_1595_),
    .A1(_1587_),
    .A2(_1593_));
 sg13g2_a221oi_1 _4928_ (.B2(_0662_),
    .C1(net1125),
    .B1(net1145),
    .A1(\cpu_instance.ram_data_out[1] ),
    .Y(_1596_),
    .A2(net1150));
 sg13g2_o21ai_1 _4929_ (.B1(net1062),
    .Y(_1597_),
    .A1(net1283),
    .A2(_0666_));
 sg13g2_a21oi_1 _4930_ (.A1(_1595_),
    .A2(_1596_),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_a21oi_1 _4931_ (.A1(\cpu_instance.pc[1] ),
    .A2(net1259),
    .Y(_1599_),
    .B1(net1039));
 sg13g2_a21oi_1 _4932_ (.A1(\cpu_instance.sp_minus_two[1] ),
    .A2(_0659_),
    .Y(_1600_),
    .B1(_1598_));
 sg13g2_a21oi_1 _4933_ (.A1(net162),
    .A2(_1985_),
    .Y(_1601_),
    .B1(_0672_));
 sg13g2_a21oi_1 _4934_ (.A1(_1599_),
    .A2(_1600_),
    .Y(_1602_),
    .B1(_1601_));
 sg13g2_a21o_1 _4935_ (.A2(net1028),
    .A1(net157),
    .B1(_1602_),
    .X(_0170_));
 sg13g2_a21o_2 _4936_ (.A2(_1592_),
    .A1(_1587_),
    .B1(_1591_),
    .X(_1603_));
 sg13g2_nand2_1 _4937_ (.Y(_1604_),
    .A(_1913_),
    .B(\cpu_instance.dp[2] ));
 sg13g2_nand2b_1 _4938_ (.Y(_1605_),
    .B(net1297),
    .A_N(_0009_));
 sg13g2_a21oi_1 _4939_ (.A1(_1604_),
    .A2(_1605_),
    .Y(_1606_),
    .B1(net1214));
 sg13g2_and2_1 _4940_ (.A(_2327_),
    .B(_1606_),
    .X(_1607_));
 sg13g2_xor2_1 _4941_ (.B(_1606_),
    .A(_2327_),
    .X(_1608_));
 sg13g2_and2_1 _4942_ (.A(_1603_),
    .B(_1608_),
    .X(_1609_));
 sg13g2_o21ai_1 _4943_ (.B1(_0504_),
    .Y(_1610_),
    .A1(_1603_),
    .A2(_1608_));
 sg13g2_a221oi_1 _4944_ (.B2(_0664_),
    .C1(_0668_),
    .B1(net1143),
    .A1(\cpu_instance.ram_data_out[2] ),
    .Y(_1611_),
    .A2(net1150));
 sg13g2_o21ai_1 _4945_ (.B1(_1611_),
    .Y(_1612_),
    .A1(_1609_),
    .A2(_1610_));
 sg13g2_a21oi_1 _4946_ (.A1(_0530_),
    .A2(net1142),
    .Y(_1613_),
    .B1(net1125));
 sg13g2_a221oi_1 _4947_ (.B2(_1613_),
    .C1(_0659_),
    .B1(_1612_),
    .A1(\cpu_instance.sp[2] ),
    .Y(_1614_),
    .A2(net1125));
 sg13g2_o21ai_1 _4948_ (.B1(net1254),
    .Y(_1615_),
    .A1(net1062),
    .A2(_1489_));
 sg13g2_a21oi_1 _4949_ (.A1(\cpu_instance.pc[2] ),
    .A2(net1259),
    .Y(_1616_),
    .B1(net1039));
 sg13g2_o21ai_1 _4950_ (.B1(_1616_),
    .Y(_1617_),
    .A1(_1614_),
    .A2(_1615_));
 sg13g2_o21ai_1 _4951_ (.B1(_1617_),
    .Y(_1618_),
    .A1(\cpu_instance.spi_ram.addr[2] ),
    .A2(_1585_));
 sg13g2_a21oi_1 _4952_ (.A1(_1951_),
    .A2(_1985_),
    .Y(_0171_),
    .B1(_1618_));
 sg13g2_a21o_1 _4953_ (.A2(_1608_),
    .A1(_1603_),
    .B1(_1607_),
    .X(_1619_));
 sg13g2_mux2_1 _4954_ (.A0(\cpu_instance.dp[3] ),
    .A1(\cpu_instance.sp[3] ),
    .S(net1297),
    .X(_1620_));
 sg13g2_nand2_2 _4955_ (.Y(_1621_),
    .A(net1211),
    .B(_1620_));
 sg13g2_nor2_1 _4956_ (.A(_2315_),
    .B(_1621_),
    .Y(_1622_));
 sg13g2_xor2_1 _4957_ (.B(_1621_),
    .A(_2315_),
    .X(_1623_));
 sg13g2_a21oi_1 _4958_ (.A1(_1619_),
    .A2(_1623_),
    .Y(_1624_),
    .B1(_0505_));
 sg13g2_o21ai_1 _4959_ (.B1(_1624_),
    .Y(_1625_),
    .A1(_1619_),
    .A2(_1623_));
 sg13g2_a22oi_1 _4960_ (.Y(_1626_),
    .B1(_0540_),
    .B2(_0664_),
    .A2(net1150),
    .A1(\cpu_instance.ram_data_out[3] ));
 sg13g2_nand3_1 _4961_ (.B(_1625_),
    .C(_1626_),
    .A(_0663_),
    .Y(_1627_));
 sg13g2_nand2_1 _4962_ (.Y(_1628_),
    .A(net1126),
    .B(net1142));
 sg13g2_a21oi_1 _4963_ (.A1(\cpu_instance.sp[3] ),
    .A2(net1123),
    .Y(_1629_),
    .B1(net1257));
 sg13g2_o21ai_1 _4964_ (.B1(_1629_),
    .Y(_1630_),
    .A1(net1061),
    .A2(_1494_));
 sg13g2_a21oi_1 _4965_ (.A1(_1627_),
    .A2(_1628_),
    .Y(_1631_),
    .B1(_1630_));
 sg13g2_o21ai_1 _4966_ (.B1(net1048),
    .Y(_1632_),
    .A1(\cpu_instance.pc[3] ),
    .A2(net1256));
 sg13g2_o21ai_1 _4967_ (.B1(net1039),
    .Y(_1633_),
    .A1(\cpu_instance.spi_ram.addr[2] ),
    .A2(_1986_));
 sg13g2_o21ai_1 _4968_ (.B1(_1633_),
    .Y(_1634_),
    .A1(_1631_),
    .A2(_1632_));
 sg13g2_o21ai_1 _4969_ (.B1(_1634_),
    .Y(_1635_),
    .A1(net187),
    .A2(_1585_));
 sg13g2_inv_1 _4970_ (.Y(_0172_),
    .A(net188));
 sg13g2_a21o_1 _4971_ (.A2(_1623_),
    .A1(_1619_),
    .B1(_1622_),
    .X(_1636_));
 sg13g2_nor2b_1 _4972_ (.A(net1297),
    .B_N(\cpu_instance.dp[4] ),
    .Y(_1637_));
 sg13g2_nor2_1 _4973_ (.A(_1913_),
    .B(_0008_),
    .Y(_1638_));
 sg13g2_o21ai_1 _4974_ (.B1(net1211),
    .Y(_1639_),
    .A1(_1637_),
    .A2(_1638_));
 sg13g2_nor2_1 _4975_ (.A(_2306_),
    .B(_1639_),
    .Y(_1640_));
 sg13g2_xor2_1 _4976_ (.B(_1639_),
    .A(_2306_),
    .X(_1641_));
 sg13g2_o21ai_1 _4977_ (.B1(net1146),
    .Y(_1642_),
    .A1(_1636_),
    .A2(_1641_));
 sg13g2_a21oi_2 _4978_ (.B1(_1642_),
    .Y(_1643_),
    .A2(_1641_),
    .A1(_1636_));
 sg13g2_a22oi_1 _4979_ (.Y(_1644_),
    .B1(_0547_),
    .B2(_0664_),
    .A2(net1150),
    .A1(\cpu_instance.ram_data_out[4] ));
 sg13g2_nand2_1 _4980_ (.Y(_1645_),
    .A(_0663_),
    .B(_1644_));
 sg13g2_a21oi_1 _4981_ (.A1(_0548_),
    .A2(_0660_),
    .Y(_1646_),
    .B1(net1125));
 sg13g2_o21ai_1 _4982_ (.B1(_1646_),
    .Y(_1647_),
    .A1(_1643_),
    .A2(_1645_));
 sg13g2_a221oi_1 _4983_ (.B2(net1069),
    .C1(net1257),
    .B1(_1505_),
    .A1(\cpu_instance.sp[4] ),
    .Y(_1648_),
    .A2(net1123));
 sg13g2_nand2_1 _4984_ (.Y(_1649_),
    .A(_1647_),
    .B(_1648_));
 sg13g2_o21ai_1 _4985_ (.B1(_1649_),
    .Y(_1650_),
    .A1(\cpu_instance.pc[4] ),
    .A2(net1256));
 sg13g2_o21ai_1 _4986_ (.B1(_0673_),
    .Y(_1651_),
    .A1(net187),
    .A2(_1986_));
 sg13g2_o21ai_1 _4987_ (.B1(_1651_),
    .Y(_1652_),
    .A1(net1039),
    .A2(_1650_));
 sg13g2_o21ai_1 _4988_ (.B1(_1652_),
    .Y(_1653_),
    .A1(net203),
    .A2(_1585_));
 sg13g2_inv_1 _4989_ (.Y(_0173_),
    .A(_1653_));
 sg13g2_a21oi_1 _4990_ (.A1(net1069),
    .A2(_1511_),
    .Y(_1654_),
    .B1(net1257));
 sg13g2_o21ai_1 _4991_ (.B1(net1062),
    .Y(_1655_),
    .A1(\cpu_instance.sp[5] ),
    .A2(_0666_));
 sg13g2_a21o_1 _4992_ (.A2(_1641_),
    .A1(_1636_),
    .B1(_1640_),
    .X(_1656_));
 sg13g2_mux2_1 _4993_ (.A0(\cpu_instance.dp[5] ),
    .A1(\cpu_instance.sp[5] ),
    .S(net1295),
    .X(_1657_));
 sg13g2_and3_1 _4994_ (.X(_1658_),
    .A(net1211),
    .B(net1105),
    .C(_1657_));
 sg13g2_a21oi_1 _4995_ (.A1(net1211),
    .A2(_1657_),
    .Y(_1659_),
    .B1(net1105));
 sg13g2_inv_1 _4996_ (.Y(_1660_),
    .A(_1659_));
 sg13g2_nor2_1 _4997_ (.A(_1658_),
    .B(_1659_),
    .Y(_1661_));
 sg13g2_o21ai_1 _4998_ (.B1(net1146),
    .Y(_1662_),
    .A1(_1656_),
    .A2(_1661_));
 sg13g2_a21oi_1 _4999_ (.A1(_1656_),
    .A2(_1661_),
    .Y(_1663_),
    .B1(_1662_));
 sg13g2_a221oi_1 _5000_ (.B2(_0662_),
    .C1(net1125),
    .B1(_0557_),
    .A1(\cpu_instance.ram_data_out[5] ),
    .Y(_1664_),
    .A2(_0500_));
 sg13g2_nor2b_1 _5001_ (.A(_1663_),
    .B_N(_1664_),
    .Y(_1665_));
 sg13g2_o21ai_1 _5002_ (.B1(_1654_),
    .Y(_1666_),
    .A1(_1655_),
    .A2(_1665_));
 sg13g2_a21oi_2 _5003_ (.B1(net1039),
    .Y(_1667_),
    .A2(net1259),
    .A1(_1901_));
 sg13g2_a221oi_1 _5004_ (.B2(_1667_),
    .C1(_1584_),
    .B1(_1666_),
    .A1(\cpu_instance.spi_ram.addr[4] ),
    .Y(_1668_),
    .A2(net1038));
 sg13g2_a21oi_1 _5005_ (.A1(_1955_),
    .A2(net1028),
    .Y(_0174_),
    .B1(_1668_));
 sg13g2_nand2_1 _5006_ (.Y(_1669_),
    .A(net1294),
    .B(_0006_));
 sg13g2_o21ai_1 _5007_ (.B1(_1669_),
    .Y(_1670_),
    .A1(net1294),
    .A2(\cpu_instance.dp[6] ));
 sg13g2_nor2_1 _5008_ (.A(net1214),
    .B(_1670_),
    .Y(_1671_));
 sg13g2_nor2b_1 _5009_ (.A(_2286_),
    .B_N(_1671_),
    .Y(_1672_));
 sg13g2_xnor2_1 _5010_ (.Y(_1673_),
    .A(_2286_),
    .B(_1671_));
 sg13g2_a21o_1 _5011_ (.A2(_1660_),
    .A1(_1656_),
    .B1(_1658_),
    .X(_1674_));
 sg13g2_nand2_1 _5012_ (.Y(_1675_),
    .A(_1673_),
    .B(_1674_));
 sg13g2_nor2_1 _5013_ (.A(_1673_),
    .B(_1674_),
    .Y(_1676_));
 sg13g2_nand3b_1 _5014_ (.B(net1146),
    .C(_1675_),
    .Y(_1677_),
    .A_N(_1676_));
 sg13g2_a22oi_1 _5015_ (.Y(_1678_),
    .B1(_0566_),
    .B2(_0664_),
    .A2(_0500_),
    .A1(\cpu_instance.ram_data_out[6] ));
 sg13g2_nand3_1 _5016_ (.B(_1677_),
    .C(_1678_),
    .A(_0663_),
    .Y(_1679_));
 sg13g2_a21oi_1 _5017_ (.A1(net1070),
    .A2(net1142),
    .Y(_1680_),
    .B1(net1124));
 sg13g2_o21ai_1 _5018_ (.B1(net1254),
    .Y(_1681_),
    .A1(net1061),
    .A2(_1515_));
 sg13g2_a221oi_1 _5019_ (.B2(_1680_),
    .C1(_1681_),
    .B1(_1679_),
    .A1(\cpu_instance.sp[6] ),
    .Y(_1682_),
    .A2(net1123));
 sg13g2_o21ai_1 _5020_ (.B1(net1048),
    .Y(_1683_),
    .A1(\cpu_instance.pc[6] ),
    .A2(net1255));
 sg13g2_o21ai_1 _5021_ (.B1(net1037),
    .Y(_1684_),
    .A1(net165),
    .A2(net1276));
 sg13g2_o21ai_1 _5022_ (.B1(_1684_),
    .Y(_1685_),
    .A1(_1682_),
    .A2(_1683_));
 sg13g2_o21ai_1 _5023_ (.B1(_1685_),
    .Y(_1686_),
    .A1(net200),
    .A2(_1585_));
 sg13g2_inv_1 _5024_ (.Y(_0175_),
    .A(_1686_));
 sg13g2_a21oi_2 _5025_ (.B1(_1672_),
    .Y(_1687_),
    .A2(_1674_),
    .A1(_1673_));
 sg13g2_mux2_1 _5026_ (.A0(\cpu_instance.dp[7] ),
    .A1(\cpu_instance.sp[7] ),
    .S(net1295),
    .X(_1688_));
 sg13g2_and3_1 _5027_ (.X(_1689_),
    .A(net1211),
    .B(_2276_),
    .C(_1688_));
 sg13g2_nand3_1 _5028_ (.B(_2276_),
    .C(_1688_),
    .A(net1211),
    .Y(_1690_));
 sg13g2_a21oi_1 _5029_ (.A1(net1211),
    .A2(_1688_),
    .Y(_1691_),
    .B1(_2276_));
 sg13g2_or2_1 _5030_ (.X(_1692_),
    .B(_1691_),
    .A(_1689_));
 sg13g2_a21oi_1 _5031_ (.A1(_1687_),
    .A2(_1692_),
    .Y(_1693_),
    .B1(_0505_));
 sg13g2_o21ai_1 _5032_ (.B1(_1693_),
    .Y(_1694_),
    .A1(_1687_),
    .A2(_1692_));
 sg13g2_a221oi_1 _5033_ (.B2(_0662_),
    .C1(net1125),
    .B1(_0575_),
    .A1(\cpu_instance.ram_data_out[7] ),
    .Y(_1695_),
    .A2(net1150));
 sg13g2_o21ai_1 _5034_ (.B1(net1061),
    .Y(_1696_),
    .A1(\cpu_instance.sp[7] ),
    .A2(_0666_));
 sg13g2_a21oi_1 _5035_ (.A1(_1694_),
    .A2(_1695_),
    .Y(_1697_),
    .B1(_1696_));
 sg13g2_o21ai_1 _5036_ (.B1(net1254),
    .Y(_1698_),
    .A1(net1061),
    .A2(_1524_));
 sg13g2_a21oi_1 _5037_ (.A1(_1899_),
    .A2(net1257),
    .Y(_1699_),
    .B1(net1037));
 sg13g2_o21ai_1 _5038_ (.B1(_1699_),
    .Y(_1700_),
    .A1(_1697_),
    .A2(_1698_));
 sg13g2_o21ai_1 _5039_ (.B1(net1036),
    .Y(_1701_),
    .A1(\cpu_instance.spi_ram.addr[6] ),
    .A2(net1276));
 sg13g2_a22oi_1 _5040_ (.Y(_0176_),
    .B1(_1700_),
    .B2(_1701_),
    .A2(net1028),
    .A1(_1959_));
 sg13g2_nor2_1 _5041_ (.A(net179),
    .B(_1585_),
    .Y(_1702_));
 sg13g2_nand2_1 _5042_ (.Y(_1703_),
    .A(net1294),
    .B(_0005_));
 sg13g2_o21ai_1 _5043_ (.B1(_1703_),
    .Y(_1704_),
    .A1(net1294),
    .A2(\cpu_instance.dp[8] ));
 sg13g2_nor2_1 _5044_ (.A(net1214),
    .B(_1704_),
    .Y(_1705_));
 sg13g2_and2_1 _5045_ (.A(_2251_),
    .B(_1705_),
    .X(_1706_));
 sg13g2_xnor2_1 _5046_ (.Y(_1707_),
    .A(_2251_),
    .B(_1705_));
 sg13g2_inv_1 _5047_ (.Y(_1708_),
    .A(_1707_));
 sg13g2_a21oi_2 _5048_ (.B1(_1691_),
    .Y(_1709_),
    .A2(_1690_),
    .A1(_1687_));
 sg13g2_o21ai_1 _5049_ (.B1(net1146),
    .Y(_1710_),
    .A1(_1708_),
    .A2(_1709_));
 sg13g2_a21o_1 _5050_ (.A2(_1709_),
    .A1(_1708_),
    .B1(_1710_),
    .X(_1711_));
 sg13g2_a221oi_1 _5051_ (.B2(_0662_),
    .C1(net1124),
    .B1(_0584_),
    .A1(\cpu_instance.ram_data_out[8] ),
    .Y(_1712_),
    .A2(net1149));
 sg13g2_nand2_1 _5052_ (.Y(_1713_),
    .A(_1711_),
    .B(_1712_));
 sg13g2_a21oi_1 _5053_ (.A1(_1892_),
    .A2(net1123),
    .Y(_1714_),
    .B1(net1069));
 sg13g2_a221oi_1 _5054_ (.B2(_1714_),
    .C1(net1257),
    .B1(_1713_),
    .A1(net1069),
    .Y(_1715_),
    .A2(_1535_));
 sg13g2_o21ai_1 _5055_ (.B1(net1048),
    .Y(_1716_),
    .A1(\cpu_instance.pc[8] ),
    .A2(net1255));
 sg13g2_nor2_1 _5056_ (.A(_1715_),
    .B(_1716_),
    .Y(_1717_));
 sg13g2_a21oi_1 _5057_ (.A1(net172),
    .A2(net1036),
    .Y(_1718_),
    .B1(_1717_));
 sg13g2_a21oi_1 _5058_ (.A1(_1585_),
    .A2(_1718_),
    .Y(_0177_),
    .B1(_1702_));
 sg13g2_a21oi_2 _5059_ (.B1(_1706_),
    .Y(_1719_),
    .A2(_1709_),
    .A1(_1708_));
 sg13g2_mux2_1 _5060_ (.A0(\cpu_instance.dp[9] ),
    .A1(\cpu_instance.sp[9] ),
    .S(net1294),
    .X(_1720_));
 sg13g2_nand3_1 _5061_ (.B(_2241_),
    .C(_1720_),
    .A(net1211),
    .Y(_1721_));
 sg13g2_a21oi_1 _5062_ (.A1(net1212),
    .A2(_1720_),
    .Y(_1722_),
    .B1(_2241_));
 sg13g2_inv_1 _5063_ (.Y(_1723_),
    .A(_1722_));
 sg13g2_nand2_1 _5064_ (.Y(_1724_),
    .A(_1721_),
    .B(_1723_));
 sg13g2_a21oi_1 _5065_ (.A1(_1719_),
    .A2(_1724_),
    .Y(_1725_),
    .B1(_0505_));
 sg13g2_o21ai_1 _5066_ (.B1(_1725_),
    .Y(_1726_),
    .A1(_1719_),
    .A2(_1724_));
 sg13g2_a221oi_1 _5067_ (.B2(_0662_),
    .C1(net1124),
    .B1(net1052),
    .A1(\cpu_instance.ram_data_out[9] ),
    .Y(_1727_),
    .A2(net1149));
 sg13g2_nand2_1 _5068_ (.Y(_1728_),
    .A(_1726_),
    .B(_1727_));
 sg13g2_a21oi_1 _5069_ (.A1(_1891_),
    .A2(net1123),
    .Y(_1729_),
    .B1(net1069));
 sg13g2_a22oi_1 _5070_ (.Y(_1730_),
    .B1(_1728_),
    .B2(_1729_),
    .A2(_1541_),
    .A1(net1069));
 sg13g2_o21ai_1 _5071_ (.B1(net1048),
    .Y(_1731_),
    .A1(\cpu_instance.pc[9] ),
    .A2(net1255));
 sg13g2_a21o_1 _5072_ (.A2(_1730_),
    .A1(net1254),
    .B1(_1731_),
    .X(_1732_));
 sg13g2_o21ai_1 _5073_ (.B1(net1036),
    .Y(_1733_),
    .A1(net179),
    .A2(net1276));
 sg13g2_a22oi_1 _5074_ (.Y(_0178_),
    .B1(_1732_),
    .B2(_1733_),
    .A2(net1028),
    .A1(_1962_));
 sg13g2_o21ai_1 _5075_ (.B1(net1036),
    .Y(_1734_),
    .A1(net195),
    .A2(net1276));
 sg13g2_nand2_1 _5076_ (.Y(_1735_),
    .A(net1294),
    .B(_0003_));
 sg13g2_o21ai_1 _5077_ (.B1(_1735_),
    .Y(_1736_),
    .A1(net1294),
    .A2(\cpu_instance.dp[10] ));
 sg13g2_nor2_1 _5078_ (.A(net1214),
    .B(_1736_),
    .Y(_1737_));
 sg13g2_and2_1 _5079_ (.A(_2230_),
    .B(_1737_),
    .X(_1738_));
 sg13g2_xnor2_1 _5080_ (.Y(_1739_),
    .A(_2230_),
    .B(_1737_));
 sg13g2_inv_1 _5081_ (.Y(_1740_),
    .A(_1739_));
 sg13g2_a21oi_1 _5082_ (.A1(_1719_),
    .A2(_1721_),
    .Y(_1741_),
    .B1(_1722_));
 sg13g2_and2_1 _5083_ (.A(_1740_),
    .B(_1741_),
    .X(_1742_));
 sg13g2_o21ai_1 _5084_ (.B1(net1146),
    .Y(_1743_),
    .A1(_1740_),
    .A2(_1741_));
 sg13g2_a22oi_1 _5085_ (.Y(_1744_),
    .B1(net1049),
    .B2(_0669_),
    .A2(net1150),
    .A1(\cpu_instance.ram_data_out[10] ));
 sg13g2_o21ai_1 _5086_ (.B1(_1744_),
    .Y(_1745_),
    .A1(_1742_),
    .A2(_1743_));
 sg13g2_o21ai_1 _5087_ (.B1(net1254),
    .Y(_1746_),
    .A1(net1061),
    .A2(_1545_));
 sg13g2_a221oi_1 _5088_ (.B2(net1050),
    .C1(_1746_),
    .B1(net1142),
    .A1(\cpu_instance.sp[10] ),
    .Y(_1747_),
    .A2(net1124));
 sg13g2_nand2b_1 _5089_ (.Y(_1748_),
    .B(_1747_),
    .A_N(_1745_));
 sg13g2_o21ai_1 _5090_ (.B1(_1748_),
    .Y(_1749_),
    .A1(\cpu_instance.pc[10] ),
    .A2(net1254));
 sg13g2_o21ai_1 _5091_ (.B1(_1734_),
    .Y(_1750_),
    .A1(net1036),
    .A2(_1749_));
 sg13g2_o21ai_1 _5092_ (.B1(_1750_),
    .Y(_1751_),
    .A1(net209),
    .A2(_1585_));
 sg13g2_inv_1 _5093_ (.Y(_0179_),
    .A(_1751_));
 sg13g2_nor2_1 _5094_ (.A(_1738_),
    .B(_1742_),
    .Y(_1752_));
 sg13g2_mux2_1 _5095_ (.A0(\cpu_instance.dp[11] ),
    .A1(\cpu_instance.sp[11] ),
    .S(net1300),
    .X(_1753_));
 sg13g2_nand3_1 _5096_ (.B(_2222_),
    .C(_1753_),
    .A(net1212),
    .Y(_1754_));
 sg13g2_inv_1 _5097_ (.Y(_1755_),
    .A(_1754_));
 sg13g2_a21oi_2 _5098_ (.B1(_2222_),
    .Y(_1756_),
    .A2(_1753_),
    .A1(net1212));
 sg13g2_nor2_1 _5099_ (.A(_1755_),
    .B(_1756_),
    .Y(_1757_));
 sg13g2_nand2_1 _5100_ (.Y(_1758_),
    .A(net1041),
    .B(net1142));
 sg13g2_a221oi_1 _5101_ (.B2(_0664_),
    .C1(_0504_),
    .B1(net1041),
    .A1(\cpu_instance.ram_data_out[11] ),
    .Y(_1759_),
    .A2(net1149));
 sg13g2_xor2_1 _5102_ (.B(_1757_),
    .A(_1752_),
    .X(_1760_));
 sg13g2_a21oi_1 _5103_ (.A1(net1146),
    .A2(_1760_),
    .Y(_1761_),
    .B1(_1759_));
 sg13g2_nor2_1 _5104_ (.A(net1124),
    .B(_1761_),
    .Y(_1762_));
 sg13g2_o21ai_1 _5105_ (.B1(net1062),
    .Y(_1763_),
    .A1(\cpu_instance.sp[11] ),
    .A2(_0666_));
 sg13g2_a21oi_1 _5106_ (.A1(_1758_),
    .A2(_1762_),
    .Y(_1764_),
    .B1(_1763_));
 sg13g2_o21ai_1 _5107_ (.B1(net1254),
    .Y(_1765_),
    .A1(net1062),
    .A2(_1554_));
 sg13g2_a21oi_1 _5108_ (.A1(_1897_),
    .A2(net1257),
    .Y(_1766_),
    .B1(net1037));
 sg13g2_o21ai_1 _5109_ (.B1(_1766_),
    .Y(_1767_),
    .A1(_1764_),
    .A2(_1765_));
 sg13g2_o21ai_1 _5110_ (.B1(net1036),
    .Y(_1768_),
    .A1(\cpu_instance.spi_ram.addr[10] ),
    .A2(net1276));
 sg13g2_a22oi_1 _5111_ (.Y(_0180_),
    .B1(_1767_),
    .B2(_1768_),
    .A2(net1028),
    .A1(_1965_));
 sg13g2_nor2_1 _5112_ (.A(net1296),
    .B(\cpu_instance.dp[12] ),
    .Y(_1769_));
 sg13g2_a21oi_1 _5113_ (.A1(net1296),
    .A2(_0002_),
    .Y(_1770_),
    .B1(_1769_));
 sg13g2_nand2_1 _5114_ (.Y(_1771_),
    .A(net1212),
    .B(_1770_));
 sg13g2_nor2_1 _5115_ (.A(_2212_),
    .B(_1771_),
    .Y(_1772_));
 sg13g2_xnor2_1 _5116_ (.Y(_1773_),
    .A(_2212_),
    .B(_1771_));
 sg13g2_nor3_1 _5117_ (.A(_1738_),
    .B(_1742_),
    .C(_1755_),
    .Y(_1774_));
 sg13g2_o21ai_1 _5118_ (.B1(_1754_),
    .Y(_1775_),
    .A1(_1752_),
    .A2(_1756_));
 sg13g2_o21ai_1 _5119_ (.B1(_1773_),
    .Y(_1776_),
    .A1(_1756_),
    .A2(_1774_));
 sg13g2_nor3_1 _5120_ (.A(_1756_),
    .B(_1773_),
    .C(_1774_),
    .Y(_1777_));
 sg13g2_nand2b_1 _5121_ (.Y(_1778_),
    .B(_1775_),
    .A_N(_1773_));
 sg13g2_nand3_1 _5122_ (.B(_1776_),
    .C(_1778_),
    .A(net1146),
    .Y(_1779_));
 sg13g2_a22oi_1 _5123_ (.Y(_1780_),
    .B1(_0621_),
    .B2(_0664_),
    .A2(net1149),
    .A1(\cpu_instance.ram_data_out[12] ));
 sg13g2_nand3_1 _5124_ (.B(_1779_),
    .C(_1780_),
    .A(_0663_),
    .Y(_1781_));
 sg13g2_nand2_1 _5125_ (.Y(_1782_),
    .A(_0622_),
    .B(net1142));
 sg13g2_a21oi_1 _5126_ (.A1(\cpu_instance.sp[12] ),
    .A2(net1123),
    .Y(_1783_),
    .B1(net1257));
 sg13g2_o21ai_1 _5127_ (.B1(_1783_),
    .Y(_1784_),
    .A1(net1061),
    .A2(_1562_));
 sg13g2_a21oi_1 _5128_ (.A1(_1781_),
    .A2(_1782_),
    .Y(_1785_),
    .B1(_1784_));
 sg13g2_o21ai_1 _5129_ (.B1(net1048),
    .Y(_1786_),
    .A1(\cpu_instance.pc[12] ),
    .A2(net1255));
 sg13g2_o21ai_1 _5130_ (.B1(net1036),
    .Y(_1787_),
    .A1(net176),
    .A2(net1276));
 sg13g2_o21ai_1 _5131_ (.B1(_1787_),
    .Y(_1788_),
    .A1(_1785_),
    .A2(_1786_));
 sg13g2_o21ai_1 _5132_ (.B1(_1788_),
    .Y(_1789_),
    .A1(net202),
    .A2(_1585_));
 sg13g2_inv_1 _5133_ (.Y(_0181_),
    .A(_1789_));
 sg13g2_nand2_1 _5134_ (.Y(_1790_),
    .A(net1295),
    .B(_0001_));
 sg13g2_o21ai_1 _5135_ (.B1(_1790_),
    .Y(_1791_),
    .A1(net1295),
    .A2(\cpu_instance.dp[13] ));
 sg13g2_nand3b_1 _5136_ (.B(net1213),
    .C(_2202_),
    .Y(_1792_),
    .A_N(_1791_));
 sg13g2_o21ai_1 _5137_ (.B1(_2203_),
    .Y(_1793_),
    .A1(net1214),
    .A2(_1791_));
 sg13g2_nand2_1 _5138_ (.Y(_1794_),
    .A(_1792_),
    .B(_1793_));
 sg13g2_nand3b_1 _5139_ (.B(_1778_),
    .C(_1794_),
    .Y(_1795_),
    .A_N(_1772_));
 sg13g2_o21ai_1 _5140_ (.B1(_1793_),
    .Y(_1796_),
    .A1(_1772_),
    .A2(_1777_));
 sg13g2_nand2b_1 _5141_ (.Y(_1797_),
    .B(_1792_),
    .A_N(_1796_));
 sg13g2_nand3_1 _5142_ (.B(_1795_),
    .C(_1797_),
    .A(net1146),
    .Y(_1798_));
 sg13g2_a221oi_1 _5143_ (.B2(_0662_),
    .C1(net1124),
    .B1(_0632_),
    .A1(\cpu_instance.ram_data_out[13] ),
    .Y(_1799_),
    .A2(net1149));
 sg13g2_o21ai_1 _5144_ (.B1(net1061),
    .Y(_1800_),
    .A1(\cpu_instance.sp[13] ),
    .A2(_0666_));
 sg13g2_a21oi_1 _5145_ (.A1(_1798_),
    .A2(_1799_),
    .Y(_1801_),
    .B1(_1800_));
 sg13g2_o21ai_1 _5146_ (.B1(net1254),
    .Y(_1802_),
    .A1(net1062),
    .A2(_1566_));
 sg13g2_a21oi_1 _5147_ (.A1(_1895_),
    .A2(net1258),
    .Y(_1803_),
    .B1(net1037));
 sg13g2_o21ai_1 _5148_ (.B1(_1803_),
    .Y(_1804_),
    .A1(_1801_),
    .A2(_1802_));
 sg13g2_o21ai_1 _5149_ (.B1(net1037),
    .Y(_1805_),
    .A1(\cpu_instance.spi_ram.addr[12] ),
    .A2(net1276));
 sg13g2_a22oi_1 _5150_ (.Y(_0182_),
    .B1(_1804_),
    .B2(_1805_),
    .A2(net1028),
    .A1(_1968_));
 sg13g2_nand2_1 _5151_ (.Y(_1806_),
    .A(_1913_),
    .B(\cpu_instance.dp[14] ));
 sg13g2_nand2b_1 _5152_ (.Y(_1807_),
    .B(net1294),
    .A_N(_0000_));
 sg13g2_a21oi_1 _5153_ (.A1(_1806_),
    .A2(_1807_),
    .Y(_1808_),
    .B1(net1214));
 sg13g2_and2_1 _5154_ (.A(_2192_),
    .B(_1808_),
    .X(_1809_));
 sg13g2_xnor2_1 _5155_ (.Y(_1810_),
    .A(_2192_),
    .B(_1808_));
 sg13g2_nand2_1 _5156_ (.Y(_1811_),
    .A(_1792_),
    .B(_1796_));
 sg13g2_a21oi_1 _5157_ (.A1(_1792_),
    .A2(_1796_),
    .Y(_1812_),
    .B1(_1810_));
 sg13g2_xor2_1 _5158_ (.B(_1811_),
    .A(_1810_),
    .X(_1813_));
 sg13g2_a22oi_1 _5159_ (.Y(_1814_),
    .B1(_0642_),
    .B2(_0661_),
    .A2(net1149),
    .A1(\cpu_instance.ram_data_out[14] ));
 sg13g2_o21ai_1 _5160_ (.B1(_1814_),
    .Y(_1815_),
    .A1(_0505_),
    .A2(_1813_));
 sg13g2_a21oi_1 _5161_ (.A1(\cpu_instance.sp[14] ),
    .A2(net1123),
    .Y(_1816_),
    .B1(net1257));
 sg13g2_o21ai_1 _5162_ (.B1(_1816_),
    .Y(_1817_),
    .A1(net1061),
    .A2(_1573_));
 sg13g2_a21oi_1 _5163_ (.A1(_0642_),
    .A2(_0660_),
    .Y(_1818_),
    .B1(_1817_));
 sg13g2_nand2b_1 _5164_ (.Y(_1819_),
    .B(_1818_),
    .A_N(_1815_));
 sg13g2_a21oi_1 _5165_ (.A1(_1894_),
    .A2(net1258),
    .Y(_1820_),
    .B1(net1038));
 sg13g2_a221oi_1 _5166_ (.B2(_1820_),
    .C1(net1028),
    .B1(_1819_),
    .A1(\cpu_instance.spi_ram.addr[13] ),
    .Y(_1821_),
    .A2(net1038));
 sg13g2_a21oi_1 _5167_ (.A1(_1970_),
    .A2(net1028),
    .Y(_0183_),
    .B1(_1821_));
 sg13g2_a22oi_1 _5168_ (.Y(_1822_),
    .B1(net1018),
    .B2(_0664_),
    .A2(net1149),
    .A1(\cpu_instance.ram_data_out[15] ));
 sg13g2_nor2b_1 _5169_ (.A(net1296),
    .B_N(\cpu_instance.dp[15] ),
    .Y(_1823_));
 sg13g2_a21oi_1 _5170_ (.A1(\cpu_instance.sp[15] ),
    .A2(net1297),
    .Y(_1824_),
    .B1(_1823_));
 sg13g2_nor2_1 _5171_ (.A(net1214),
    .B(_1824_),
    .Y(_1825_));
 sg13g2_xnor2_1 _5172_ (.Y(_1826_),
    .A(_2180_),
    .B(_1825_));
 sg13g2_nor3_1 _5173_ (.A(_1809_),
    .B(_1812_),
    .C(_1826_),
    .Y(_1827_));
 sg13g2_o21ai_1 _5174_ (.B1(_1826_),
    .Y(_1828_),
    .A1(_1809_),
    .A2(_1812_));
 sg13g2_nor2_1 _5175_ (.A(_0505_),
    .B(_1827_),
    .Y(_1829_));
 sg13g2_a22oi_1 _5176_ (.Y(_1830_),
    .B1(_1828_),
    .B2(_1829_),
    .A2(_1822_),
    .A1(_0505_));
 sg13g2_or2_1 _5177_ (.X(_1831_),
    .B(_0663_),
    .A(net1018));
 sg13g2_o21ai_1 _5178_ (.B1(_1831_),
    .Y(_1832_),
    .A1(net1142),
    .A2(_1830_));
 sg13g2_a21oi_1 _5179_ (.A1(\cpu_instance.sp[15] ),
    .A2(net1123),
    .Y(_1833_),
    .B1(net1069));
 sg13g2_a22oi_1 _5180_ (.Y(_1834_),
    .B1(_1832_),
    .B2(_1833_),
    .A2(_1580_),
    .A1(net1069));
 sg13g2_a21oi_1 _5181_ (.A1(\cpu_instance.pc[15] ),
    .A2(net1258),
    .Y(_1835_),
    .B1(net1038));
 sg13g2_nor2b_1 _5182_ (.A(_1834_),
    .B_N(_1835_),
    .Y(_1836_));
 sg13g2_a221oi_1 _5183_ (.B2(_1946_),
    .C1(_1836_),
    .B1(_1584_),
    .A1(_1970_),
    .Y(_0184_),
    .A2(_1985_));
 sg13g2_xnor2_1 _5184_ (.Y(_1837_),
    .A(_0813_),
    .B(_1586_));
 sg13g2_a221oi_1 _5185_ (.B2(_0669_),
    .C1(net1142),
    .B1(_0515_),
    .A1(_1971_),
    .Y(_1838_),
    .A2(net1150));
 sg13g2_o21ai_1 _5186_ (.B1(_1838_),
    .Y(_1839_),
    .A1(_0505_),
    .A2(_1837_));
 sg13g2_a21oi_1 _5187_ (.A1(_0516_),
    .A2(_0660_),
    .Y(_1840_),
    .B1(net1259));
 sg13g2_a22oi_1 _5188_ (.Y(_1841_),
    .B1(_1839_),
    .B2(_1840_),
    .A2(net1259),
    .A1(\cpu_instance.pc[0] ));
 sg13g2_nand3_1 _5189_ (.B(_1986_),
    .C(net1039),
    .A(net162),
    .Y(_1842_));
 sg13g2_o21ai_1 _5190_ (.B1(_1842_),
    .Y(_0185_),
    .A1(net1039),
    .A2(_1841_));
 sg13g2_nor3_1 _5191_ (.A(net1267),
    .B(_2070_),
    .C(_0965_),
    .Y(_1843_));
 sg13g2_nor3_1 _5192_ (.A(_1989_),
    .B(_2131_),
    .C(_1843_),
    .Y(_1844_));
 sg13g2_a21oi_1 _5193_ (.A1(_2093_),
    .A2(_0499_),
    .Y(_1845_),
    .B1(net1226));
 sg13g2_nand2_1 _5194_ (.Y(_1846_),
    .A(net10),
    .B(_2133_));
 sg13g2_o21ai_1 _5195_ (.B1(_1846_),
    .Y(_1847_),
    .A1(net10),
    .A2(_1989_));
 sg13g2_nand2_1 _5196_ (.Y(_1848_),
    .A(_1974_),
    .B(_2131_));
 sg13g2_nand4_1 _5197_ (.B(_2142_),
    .C(_1847_),
    .A(_1982_),
    .Y(_1849_),
    .D(_1848_));
 sg13g2_nor2_1 _5198_ (.A(_1845_),
    .B(_1849_),
    .Y(_1850_));
 sg13g2_a221oi_1 _5199_ (.B2(_1844_),
    .C1(net1324),
    .B1(_1850_),
    .A1(_1888_),
    .Y(_0186_),
    .A2(_1849_));
 sg13g2_nor2_1 _5200_ (.A(_2146_),
    .B(_1849_),
    .Y(_1851_));
 sg13g2_a21oi_1 _5201_ (.A1(net1279),
    .A2(net1178),
    .Y(_1852_),
    .B1(net1161));
 sg13g2_o21ai_1 _5202_ (.B1(_1852_),
    .Y(_1853_),
    .A1(net1178),
    .A2(_0956_));
 sg13g2_nor2_1 _5203_ (.A(net1279),
    .B(net1163),
    .Y(_1854_));
 sg13g2_nor3_1 _5204_ (.A(net1232),
    .B(net1136),
    .C(_1854_),
    .Y(_1855_));
 sg13g2_nor2_1 _5205_ (.A(net1278),
    .B(_2073_),
    .Y(_1856_));
 sg13g2_nor2_1 _5206_ (.A(net1046),
    .B(_0816_),
    .Y(_1857_));
 sg13g2_a221oi_1 _5207_ (.B2(_1855_),
    .C1(_0805_),
    .B1(_1853_),
    .A1(net1279),
    .Y(_1858_),
    .A2(net1231));
 sg13g2_nor3_1 _5208_ (.A(_2089_),
    .B(_1857_),
    .C(_1858_),
    .Y(_1859_));
 sg13g2_a21oi_1 _5209_ (.A1(net1279),
    .A2(_2089_),
    .Y(_1860_),
    .B1(_1859_));
 sg13g2_o21ai_1 _5210_ (.B1(_2086_),
    .Y(_1861_),
    .A1(_2104_),
    .A2(_1860_));
 sg13g2_a21oi_1 _5211_ (.A1(net1319),
    .A2(_2087_),
    .Y(_1862_),
    .B1(_2085_));
 sg13g2_a21oi_1 _5212_ (.A1(_1861_),
    .A2(_1862_),
    .Y(_1863_),
    .B1(_0714_));
 sg13g2_nand2_1 _5213_ (.Y(_1864_),
    .A(_2093_),
    .B(_0947_));
 sg13g2_nand2_1 _5214_ (.Y(_1865_),
    .A(net1194),
    .B(_1112_));
 sg13g2_a21o_1 _5215_ (.A2(net1230),
    .A1(_2007_),
    .B1(_1991_),
    .X(_1866_));
 sg13g2_a22oi_1 _5216_ (.Y(_1867_),
    .B1(_1866_),
    .B2(_1864_),
    .A2(_1865_),
    .A1(net1230));
 sg13g2_nand4_1 _5217_ (.B(_2134_),
    .C(_2135_),
    .A(_2128_),
    .Y(_1868_),
    .D(_1867_));
 sg13g2_or2_1 _5218_ (.X(_1869_),
    .B(_1868_),
    .A(_1863_));
 sg13g2_a221oi_1 _5219_ (.B2(_1869_),
    .C1(net1324),
    .B1(_1851_),
    .A1(_1887_),
    .Y(_0187_),
    .A2(_1849_));
 sg13g2_nor3_1 _5220_ (.A(net1320),
    .B(net1215),
    .C(net1023),
    .Y(_1870_));
 sg13g2_o21ai_1 _5221_ (.B1(net1023),
    .Y(_1871_),
    .A1(_0041_),
    .A2(net1162));
 sg13g2_o21ai_1 _5222_ (.B1(_2073_),
    .Y(_1872_),
    .A1(_1852_),
    .A2(_1871_));
 sg13g2_nor4_1 _5223_ (.A(_2088_),
    .B(_2140_),
    .C(_0713_),
    .D(_1856_),
    .Y(_1873_));
 sg13g2_o21ai_1 _5224_ (.B1(_1873_),
    .Y(_1874_),
    .A1(_1870_),
    .A2(_1872_));
 sg13g2_nor4_1 _5225_ (.A(_2131_),
    .B(net1259),
    .C(_1845_),
    .D(_1849_),
    .Y(_1875_));
 sg13g2_a221oi_1 _5226_ (.B2(_1875_),
    .C1(net1324),
    .B1(_1874_),
    .A1(_1886_),
    .Y(_0188_),
    .A2(_1849_));
 sg13g2_a21o_1 _5227_ (.A2(net1231),
    .A1(net1279),
    .B1(_0981_),
    .X(_1876_));
 sg13g2_nor2_1 _5228_ (.A(_0957_),
    .B(net1113),
    .Y(_1877_));
 sg13g2_a22oi_1 _5229_ (.Y(_1878_),
    .B1(_1877_),
    .B2(net1023),
    .A2(_1876_),
    .A1(net1215));
 sg13g2_nor3_1 _5230_ (.A(_2099_),
    .B(net1119),
    .C(_1878_),
    .Y(_1879_));
 sg13g2_or2_1 _5231_ (.X(_1880_),
    .B(_1879_),
    .A(_0714_));
 sg13g2_o21ai_1 _5232_ (.B1(net1213),
    .Y(_1881_),
    .A1(net1301),
    .A2(_1864_));
 sg13g2_nand4_1 _5233_ (.B(_2096_),
    .C(net1116),
    .A(net1194),
    .Y(_1882_),
    .D(_1881_));
 sg13g2_nand3_1 _5234_ (.B(net1256),
    .C(_1880_),
    .A(_2134_),
    .Y(_1883_));
 sg13g2_a221oi_1 _5235_ (.B2(net1230),
    .C1(_1883_),
    .B1(_1882_),
    .A1(_1991_),
    .Y(_1884_),
    .A2(_1864_));
 sg13g2_a22oi_1 _5236_ (.Y(_1885_),
    .B1(_1851_),
    .B2(_1884_),
    .A2(_1849_),
    .A1(net271));
 sg13g2_nor2_1 _5237_ (.A(net1324),
    .B(_1885_),
    .Y(_0189_));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _5239_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net99),
    .D(_0055_),
    .Q_N(_0053_),
    .Q(\cpu_instance.zero ));
 sg13g2_dfrbp_1 _5240_ (.CLK(net155),
    .RESET_B(net32),
    .D(net9),
    .Q_N(_2615_),
    .Q(\cpu_instance.spi_ram.spi_miso_buf ));
 sg13g2_dfrbp_1 _5241_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net31),
    .D(_0056_),
    .Q_N(_0052_),
    .Q(\cpu_instance.ram_data_out[0] ));
 sg13g2_dfrbp_1 _5242_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net30),
    .D(net247),
    .Q_N(_2614_),
    .Q(\cpu_instance.ram_data_out[1] ));
 sg13g2_dfrbp_1 _5243_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net29),
    .D(_0058_),
    .Q_N(_2613_),
    .Q(\cpu_instance.ram_data_out[2] ));
 sg13g2_dfrbp_1 _5244_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net28),
    .D(net310),
    .Q_N(_2612_),
    .Q(\cpu_instance.ram_data_out[3] ));
 sg13g2_dfrbp_1 _5245_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net27),
    .D(net285),
    .Q_N(_2611_),
    .Q(\cpu_instance.ram_data_out[4] ));
 sg13g2_dfrbp_1 _5246_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net26),
    .D(_0061_),
    .Q_N(_2610_),
    .Q(\cpu_instance.ram_data_out[5] ));
 sg13g2_dfrbp_1 _5247_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net25),
    .D(_0062_),
    .Q_N(_0051_),
    .Q(\cpu_instance.ram_data_out[6] ));
 sg13g2_dfrbp_1 _5248_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net24),
    .D(_0063_),
    .Q_N(_0050_),
    .Q(\cpu_instance.ram_data_out[7] ));
 sg13g2_dfrbp_1 _5249_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net23),
    .D(_0064_),
    .Q_N(_0049_),
    .Q(\cpu_instance.ram_data_out[8] ));
 sg13g2_dfrbp_1 _5250_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net22),
    .D(net249),
    .Q_N(_0048_),
    .Q(\cpu_instance.ram_data_out[9] ));
 sg13g2_dfrbp_1 _5251_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net21),
    .D(_0066_),
    .Q_N(_0047_),
    .Q(\cpu_instance.ram_data_out[10] ));
 sg13g2_dfrbp_1 _5252_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net20),
    .D(net255),
    .Q_N(_0046_),
    .Q(\cpu_instance.ram_data_out[11] ));
 sg13g2_dfrbp_1 _5253_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net19),
    .D(_0068_),
    .Q_N(_0045_),
    .Q(\cpu_instance.ram_data_out[12] ));
 sg13g2_dfrbp_1 _5254_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net18),
    .D(net277),
    .Q_N(_0044_),
    .Q(\cpu_instance.ram_data_out[13] ));
 sg13g2_dfrbp_1 _5255_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net17),
    .D(_0070_),
    .Q_N(_0043_),
    .Q(\cpu_instance.ram_data_out[14] ));
 sg13g2_dfrbp_1 _5256_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net16),
    .D(_0071_),
    .Q_N(_2609_),
    .Q(\cpu_instance.ram_data_out[15] ));
 sg13g2_dfrbp_1 _5257_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net15),
    .D(_0072_),
    .Q_N(_2608_),
    .Q(\cpu_instance.spi_ram.writing ));
 sg13g2_dfrbp_1 _5258_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net150),
    .D(net253),
    .Q_N(_2607_),
    .Q(\cpu_instance.spi_ram.fsm_state[0] ));
 sg13g2_dfrbp_1 _5259_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net148),
    .D(_0074_),
    .Q_N(_2606_),
    .Q(\cpu_instance.spi_ram.fsm_state[1] ));
 sg13g2_dfrbp_1 _5260_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net146),
    .D(_0075_),
    .Q_N(_2605_),
    .Q(\cpu_instance.spi_ram.bits_remaining[0] ));
 sg13g2_dfrbp_1 _5261_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net144),
    .D(_0076_),
    .Q_N(_2604_),
    .Q(\cpu_instance.spi_ram.bits_remaining[1] ));
 sg13g2_dfrbp_1 _5262_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net142),
    .D(net269),
    .Q_N(_2603_),
    .Q(\cpu_instance.spi_ram.bits_remaining[2] ));
 sg13g2_dfrbp_1 _5263_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net140),
    .D(_0078_),
    .Q_N(_2602_),
    .Q(\cpu_instance.spi_ram.bits_remaining[3] ));
 sg13g2_dfrbp_1 _5264_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net138),
    .D(_0079_),
    .Q_N(_0042_),
    .Q(\cpu_instance.skipped ));
 sg13g2_dfrbp_1 _5265_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net136),
    .D(_0080_),
    .Q_N(_0041_),
    .Q(\cpu_instance.skip ));
 sg13g2_dfrbp_1 _5266_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net134),
    .D(_0081_),
    .Q_N(_2601_),
    .Q(\cpu_instance.carry ));
 sg13g2_dfrbp_1 _5267_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net132),
    .D(_0082_),
    .Q_N(_0040_),
    .Q(\cpu_instance.neg ));
 sg13g2_dfrbp_1 _5268_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net130),
    .D(net192),
    .Q_N(_2600_),
    .Q(\cpu_instance.dp[0] ));
 sg13g2_dfrbp_1 _5269_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net128),
    .D(_0084_),
    .Q_N(_2599_),
    .Q(\cpu_instance.dp[1] ));
 sg13g2_dfrbp_1 _5270_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net126),
    .D(net199),
    .Q_N(_2598_),
    .Q(\cpu_instance.dp[2] ));
 sg13g2_dfrbp_1 _5271_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net124),
    .D(_0086_),
    .Q_N(_2597_),
    .Q(\cpu_instance.dp[3] ));
 sg13g2_dfrbp_1 _5272_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net122),
    .D(net183),
    .Q_N(_2596_),
    .Q(\cpu_instance.dp[4] ));
 sg13g2_dfrbp_1 _5273_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net120),
    .D(_0088_),
    .Q_N(_2595_),
    .Q(\cpu_instance.dp[5] ));
 sg13g2_dfrbp_1 _5274_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net118),
    .D(_0089_),
    .Q_N(_2594_),
    .Q(\cpu_instance.dp[6] ));
 sg13g2_dfrbp_1 _5275_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net116),
    .D(_0090_),
    .Q_N(_2593_),
    .Q(\cpu_instance.dp[7] ));
 sg13g2_dfrbp_1 _5276_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net114),
    .D(_0091_),
    .Q_N(_2592_),
    .Q(\cpu_instance.dp[8] ));
 sg13g2_dfrbp_1 _5277_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net112),
    .D(_0092_),
    .Q_N(_2591_),
    .Q(\cpu_instance.dp[9] ));
 sg13g2_dfrbp_1 _5278_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net110),
    .D(_0093_),
    .Q_N(_2590_),
    .Q(\cpu_instance.dp[10] ));
 sg13g2_dfrbp_1 _5279_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net108),
    .D(_0094_),
    .Q_N(_2589_),
    .Q(\cpu_instance.dp[11] ));
 sg13g2_dfrbp_1 _5280_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net106),
    .D(_0095_),
    .Q_N(_2588_),
    .Q(\cpu_instance.dp[12] ));
 sg13g2_dfrbp_1 _5281_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net104),
    .D(_0096_),
    .Q_N(_2587_),
    .Q(\cpu_instance.dp[13] ));
 sg13g2_dfrbp_1 _5282_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net102),
    .D(_0097_),
    .Q_N(_2586_),
    .Q(\cpu_instance.dp[14] ));
 sg13g2_dfrbp_1 _5283_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net100),
    .D(_0098_),
    .Q_N(_2585_),
    .Q(\cpu_instance.dp[15] ));
 sg13g2_dfrbp_1 _5284_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net98),
    .D(_0099_),
    .Q_N(_0039_),
    .Q(\cpu_instance.accum[0] ));
 sg13g2_dfrbp_1 _5285_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net96),
    .D(_0100_),
    .Q_N(_0038_),
    .Q(\cpu_instance.accum[1] ));
 sg13g2_dfrbp_1 _5286_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net94),
    .D(_0101_),
    .Q_N(_0037_),
    .Q(\cpu_instance.accum[2] ));
 sg13g2_dfrbp_1 _5287_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net92),
    .D(_0102_),
    .Q_N(_0036_),
    .Q(\cpu_instance.accum[3] ));
 sg13g2_dfrbp_1 _5288_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net90),
    .D(_0103_),
    .Q_N(_0035_),
    .Q(\cpu_instance.accum[4] ));
 sg13g2_dfrbp_1 _5289_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net88),
    .D(_0104_),
    .Q_N(_0034_),
    .Q(\cpu_instance.accum[5] ));
 sg13g2_dfrbp_1 _5290_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net86),
    .D(_0105_),
    .Q_N(_0033_),
    .Q(\cpu_instance.accum[6] ));
 sg13g2_dfrbp_1 _5291_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net84),
    .D(_0106_),
    .Q_N(_0032_),
    .Q(\cpu_instance.accum[7] ));
 sg13g2_dfrbp_1 _5292_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net82),
    .D(_0107_),
    .Q_N(_0031_),
    .Q(\cpu_instance.accum[8] ));
 sg13g2_dfrbp_1 _5293_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net80),
    .D(_0108_),
    .Q_N(_0030_),
    .Q(\cpu_instance.accum[9] ));
 sg13g2_dfrbp_1 _5294_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net78),
    .D(_0109_),
    .Q_N(_0029_),
    .Q(\cpu_instance.accum[10] ));
 sg13g2_dfrbp_1 _5295_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net76),
    .D(_0110_),
    .Q_N(_0028_),
    .Q(\cpu_instance.accum[11] ));
 sg13g2_dfrbp_1 _5296_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net74),
    .D(_0111_),
    .Q_N(_0027_),
    .Q(\cpu_instance.accum[12] ));
 sg13g2_dfrbp_1 _5297_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net72),
    .D(_0112_),
    .Q_N(_0026_),
    .Q(\cpu_instance.accum[13] ));
 sg13g2_dfrbp_1 _5298_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net70),
    .D(_0113_),
    .Q_N(_0025_),
    .Q(\cpu_instance.accum[14] ));
 sg13g2_dfrbp_1 _5299_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net68),
    .D(_0114_),
    .Q_N(_0024_),
    .Q(\cpu_instance.accum[15] ));
 sg13g2_dfrbp_1 _5300_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net66),
    .D(_0115_),
    .Q_N(_0023_),
    .Q(\cpu_instance.inst[0] ));
 sg13g2_dfrbp_1 _5301_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net64),
    .D(_0116_),
    .Q_N(_0022_),
    .Q(\cpu_instance.inst[1] ));
 sg13g2_dfrbp_1 _5302_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net62),
    .D(net219),
    .Q_N(_0021_),
    .Q(\cpu_instance.inst[2] ));
 sg13g2_dfrbp_1 _5303_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net60),
    .D(net251),
    .Q_N(_0020_),
    .Q(\cpu_instance.inst[3] ));
 sg13g2_dfrbp_1 _5304_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net58),
    .D(net217),
    .Q_N(_0019_),
    .Q(\cpu_instance.inst[4] ));
 sg13g2_dfrbp_1 _5305_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net56),
    .D(net266),
    .Q_N(_0018_),
    .Q(\cpu_instance.inst[5] ));
 sg13g2_dfrbp_1 _5306_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net54),
    .D(net223),
    .Q_N(_0017_),
    .Q(\cpu_instance.inst[6] ));
 sg13g2_dfrbp_1 _5307_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net52),
    .D(net215),
    .Q_N(_0016_),
    .Q(\cpu_instance.inst[7] ));
 sg13g2_dfrbp_1 _5308_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net50),
    .D(net298),
    .Q_N(_0015_),
    .Q(\cpu_instance.inst[8] ));
 sg13g2_dfrbp_1 _5309_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net48),
    .D(_0124_),
    .Q_N(_0014_),
    .Q(\cpu_instance.inst[9] ));
 sg13g2_dfrbp_1 _5310_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net46),
    .D(_0125_),
    .Q_N(_0013_),
    .Q(\cpu_instance.inst[10] ));
 sg13g2_dfrbp_1 _5311_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net44),
    .D(_0126_),
    .Q_N(_2584_),
    .Q(\cpu_instance.inst[11] ));
 sg13g2_dfrbp_1 _5312_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net42),
    .D(net282),
    .Q_N(_2583_),
    .Q(\cpu_instance.inst[12] ));
 sg13g2_dfrbp_1 _5313_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net40),
    .D(_0128_),
    .Q_N(_2582_),
    .Q(\cpu_instance.inst[13] ));
 sg13g2_dfrbp_1 _5314_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net38),
    .D(_0129_),
    .Q_N(_2581_),
    .Q(\cpu_instance.inst[14] ));
 sg13g2_dfrbp_1 _5315_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net36),
    .D(_0130_),
    .Q_N(_0012_),
    .Q(\cpu_instance.inst[15] ));
 sg13g2_dfrbp_1 _5316_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net34),
    .D(_0131_),
    .Q_N(_0011_),
    .Q(\cpu_instance.pc[0] ));
 sg13g2_dfrbp_1 _5317_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net149),
    .D(_0132_),
    .Q_N(_2580_),
    .Q(\cpu_instance.pc[1] ));
 sg13g2_dfrbp_1 _5318_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net145),
    .D(_0133_),
    .Q_N(_2579_),
    .Q(\cpu_instance.pc[2] ));
 sg13g2_dfrbp_1 _5319_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net141),
    .D(_0134_),
    .Q_N(_2578_),
    .Q(\cpu_instance.pc[3] ));
 sg13g2_dfrbp_1 _5320_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net137),
    .D(_0135_),
    .Q_N(_2577_),
    .Q(\cpu_instance.pc[4] ));
 sg13g2_dfrbp_1 _5321_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net133),
    .D(_0136_),
    .Q_N(_2576_),
    .Q(\cpu_instance.pc[5] ));
 sg13g2_dfrbp_1 _5322_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net129),
    .D(_0137_),
    .Q_N(_2575_),
    .Q(\cpu_instance.pc[6] ));
 sg13g2_dfrbp_1 _5323_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net125),
    .D(_0138_),
    .Q_N(_2574_),
    .Q(\cpu_instance.pc[7] ));
 sg13g2_dfrbp_1 _5324_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net121),
    .D(_0139_),
    .Q_N(_2573_),
    .Q(\cpu_instance.pc[8] ));
 sg13g2_dfrbp_1 _5325_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net117),
    .D(_0140_),
    .Q_N(_2572_),
    .Q(\cpu_instance.pc[9] ));
 sg13g2_dfrbp_1 _5326_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net113),
    .D(_0141_),
    .Q_N(_2571_),
    .Q(\cpu_instance.pc[10] ));
 sg13g2_dfrbp_1 _5327_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net109),
    .D(_0142_),
    .Q_N(_2570_),
    .Q(\cpu_instance.pc[11] ));
 sg13g2_dfrbp_1 _5328_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net105),
    .D(_0143_),
    .Q_N(_2569_),
    .Q(\cpu_instance.pc[12] ));
 sg13g2_dfrbp_1 _5329_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net101),
    .D(_0144_),
    .Q_N(_2568_),
    .Q(\cpu_instance.pc[13] ));
 sg13g2_dfrbp_1 _5330_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net97),
    .D(_0145_),
    .Q_N(_0010_),
    .Q(\cpu_instance.pc[14] ));
 sg13g2_dfrbp_1 _5331_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net93),
    .D(_0146_),
    .Q_N(_2567_),
    .Q(\cpu_instance.pc[15] ));
 sg13g2_dfrbp_1 _5332_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net89),
    .D(net226),
    .Q_N(_2566_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _5333_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net85),
    .D(net229),
    .Q_N(_2565_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _5334_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net81),
    .D(net232),
    .Q_N(_2564_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _5335_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net77),
    .D(net238),
    .Q_N(_2563_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _5336_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net73),
    .D(net235),
    .Q_N(_2562_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _5337_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net69),
    .D(net243),
    .Q_N(_2561_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _5338_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net65),
    .D(net213),
    .Q_N(_2560_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _5339_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net61),
    .D(net206),
    .Q_N(_2559_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _5340_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net57),
    .D(net190),
    .Q_N(\cpu_instance.sp_minus_two[1] ),
    .Q(\cpu_instance.sp[1] ));
 sg13g2_dfrbp_1 _5341_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net53),
    .D(_0156_),
    .Q_N(_0009_),
    .Q(\cpu_instance.sp[2] ));
 sg13g2_dfrbp_1 _5342_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net49),
    .D(_0157_),
    .Q_N(_2558_),
    .Q(\cpu_instance.sp[3] ));
 sg13g2_dfrbp_1 _5343_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net45),
    .D(_0158_),
    .Q_N(_0008_),
    .Q(\cpu_instance.sp[4] ));
 sg13g2_dfrbp_1 _5344_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net41),
    .D(net292),
    .Q_N(_0007_),
    .Q(\cpu_instance.sp[5] ));
 sg13g2_dfrbp_1 _5345_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net37),
    .D(_0160_),
    .Q_N(_0006_),
    .Q(\cpu_instance.sp[6] ));
 sg13g2_dfrbp_1 _5346_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net33),
    .D(_0161_),
    .Q_N(_2557_),
    .Q(\cpu_instance.sp[7] ));
 sg13g2_dfrbp_1 _5347_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net143),
    .D(_0162_),
    .Q_N(_0005_),
    .Q(\cpu_instance.sp[8] ));
 sg13g2_dfrbp_1 _5348_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net135),
    .D(net240),
    .Q_N(_0004_),
    .Q(\cpu_instance.sp[9] ));
 sg13g2_dfrbp_1 _5349_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net127),
    .D(net264),
    .Q_N(_0003_),
    .Q(\cpu_instance.sp[10] ));
 sg13g2_dfrbp_1 _5350_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net119),
    .D(_0165_),
    .Q_N(_2556_),
    .Q(\cpu_instance.sp[11] ));
 sg13g2_dfrbp_1 _5351_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net111),
    .D(_0166_),
    .Q_N(_0002_),
    .Q(\cpu_instance.sp[12] ));
 sg13g2_dfrbp_1 _5352_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net103),
    .D(_0167_),
    .Q_N(_0001_),
    .Q(\cpu_instance.sp[13] ));
 sg13g2_dfrbp_1 _5353_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net95),
    .D(_0168_),
    .Q_N(_0000_),
    .Q(\cpu_instance.sp[14] ));
 sg13g2_dfrbp_1 _5354_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net87),
    .D(_0169_),
    .Q_N(_2555_),
    .Q(\cpu_instance.sp[15] ));
 sg13g2_dfrbp_1 _5355_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net79),
    .D(_0170_),
    .Q_N(_2554_),
    .Q(\cpu_instance.spi_ram.addr[1] ));
 sg13g2_dfrbp_1 _5356_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net75),
    .D(net158),
    .Q_N(_2553_),
    .Q(\cpu_instance.spi_ram.addr[2] ));
 sg13g2_dfrbp_1 _5357_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net71),
    .D(_0172_),
    .Q_N(_2552_),
    .Q(\cpu_instance.spi_ram.addr[3] ));
 sg13g2_dfrbp_1 _5358_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net67),
    .D(_0173_),
    .Q_N(_2551_),
    .Q(\cpu_instance.spi_ram.addr[4] ));
 sg13g2_dfrbp_1 _5359_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net63),
    .D(net166),
    .Q_N(_2550_),
    .Q(\cpu_instance.spi_ram.addr[5] ));
 sg13g2_dfrbp_1 _5360_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net59),
    .D(_0175_),
    .Q_N(_2549_),
    .Q(\cpu_instance.spi_ram.addr[6] ));
 sg13g2_dfrbp_1 _5361_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net55),
    .D(net173),
    .Q_N(_2548_),
    .Q(\cpu_instance.spi_ram.addr[7] ));
 sg13g2_dfrbp_1 _5362_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net51),
    .D(_0177_),
    .Q_N(_2547_),
    .Q(\cpu_instance.spi_ram.addr[8] ));
 sg13g2_dfrbp_1 _5363_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net47),
    .D(_0178_),
    .Q_N(_2546_),
    .Q(\cpu_instance.spi_ram.addr[9] ));
 sg13g2_dfrbp_1 _5364_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net43),
    .D(_0179_),
    .Q_N(_2545_),
    .Q(\cpu_instance.spi_ram.addr[10] ));
 sg13g2_dfrbp_1 _5365_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net39),
    .D(net177),
    .Q_N(_2544_),
    .Q(\cpu_instance.spi_ram.addr[11] ));
 sg13g2_dfrbp_1 _5366_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net35),
    .D(_0181_),
    .Q_N(_2543_),
    .Q(\cpu_instance.spi_ram.addr[12] ));
 sg13g2_dfrbp_1 _5367_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net147),
    .D(net170),
    .Q_N(_2542_),
    .Q(\cpu_instance.spi_ram.addr[13] ));
 sg13g2_dfrbp_1 _5368_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net139),
    .D(net168),
    .Q_N(_2541_),
    .Q(\cpu_instance.spi_ram.addr[14] ));
 sg13g2_dfrbp_1 _5369_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net131),
    .D(net175),
    .Q_N(_2540_),
    .Q(\cpu_instance.spi_ram.addr[15] ));
 sg13g2_dfrbp_1 _5370_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net123),
    .D(net163),
    .Q_N(_2539_),
    .Q(\cpu_instance.spi_ram.addr[0] ));
 sg13g2_dfrbp_1 _5371_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net107),
    .D(net294),
    .Q_N(_2538_),
    .Q(\cpu_instance.state[0] ));
 sg13g2_dfrbp_1 _5372_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net91),
    .D(_0187_),
    .Q_N(_2537_),
    .Q(\cpu_instance.state[1] ));
 sg13g2_dfrbp_1 _5373_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net115),
    .D(_0188_),
    .Q_N(_2536_),
    .Q(\cpu_instance.state[2] ));
 sg13g2_dfrbp_1 _5374_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net83),
    .D(_0189_),
    .Q_N(_2535_),
    .Q(\cpu_instance.state[3] ));
 sg13g2_tiehi _5256__16 (.L_HI(net16));
 sg13g2_tiehi _5255__17 (.L_HI(net17));
 sg13g2_tiehi _5254__18 (.L_HI(net18));
 sg13g2_tiehi _5253__19 (.L_HI(net19));
 sg13g2_tiehi _5252__20 (.L_HI(net20));
 sg13g2_tiehi _5251__21 (.L_HI(net21));
 sg13g2_tiehi _5250__22 (.L_HI(net22));
 sg13g2_tiehi _5249__23 (.L_HI(net23));
 sg13g2_tiehi _5248__24 (.L_HI(net24));
 sg13g2_tiehi _5247__25 (.L_HI(net25));
 sg13g2_tiehi _5246__26 (.L_HI(net26));
 sg13g2_tiehi _5245__27 (.L_HI(net27));
 sg13g2_tiehi _5244__28 (.L_HI(net28));
 sg13g2_tiehi _5243__29 (.L_HI(net29));
 sg13g2_tiehi _5242__30 (.L_HI(net30));
 sg13g2_tiehi _5241__31 (.L_HI(net31));
 sg13g2_tiehi _5240__32 (.L_HI(net32));
 sg13g2_tiehi _5346__33 (.L_HI(net33));
 sg13g2_tiehi _5316__34 (.L_HI(net34));
 sg13g2_tiehi _5366__35 (.L_HI(net35));
 sg13g2_tiehi _5315__36 (.L_HI(net36));
 sg13g2_tiehi _5345__37 (.L_HI(net37));
 sg13g2_tiehi _5314__38 (.L_HI(net38));
 sg13g2_tiehi _5365__39 (.L_HI(net39));
 sg13g2_tiehi _5313__40 (.L_HI(net40));
 sg13g2_tiehi _5344__41 (.L_HI(net41));
 sg13g2_tiehi _5312__42 (.L_HI(net42));
 sg13g2_tiehi _5364__43 (.L_HI(net43));
 sg13g2_tiehi _5311__44 (.L_HI(net44));
 sg13g2_tiehi _5343__45 (.L_HI(net45));
 sg13g2_tiehi _5310__46 (.L_HI(net46));
 sg13g2_tiehi _5363__47 (.L_HI(net47));
 sg13g2_tiehi _5309__48 (.L_HI(net48));
 sg13g2_tiehi _5342__49 (.L_HI(net49));
 sg13g2_tiehi _5308__50 (.L_HI(net50));
 sg13g2_tiehi _5362__51 (.L_HI(net51));
 sg13g2_tiehi _5307__52 (.L_HI(net52));
 sg13g2_tiehi _5341__53 (.L_HI(net53));
 sg13g2_tiehi _5306__54 (.L_HI(net54));
 sg13g2_tiehi _5361__55 (.L_HI(net55));
 sg13g2_tiehi _5305__56 (.L_HI(net56));
 sg13g2_tiehi _5340__57 (.L_HI(net57));
 sg13g2_tiehi _5304__58 (.L_HI(net58));
 sg13g2_tiehi _5360__59 (.L_HI(net59));
 sg13g2_tiehi _5303__60 (.L_HI(net60));
 sg13g2_tiehi _5339__61 (.L_HI(net61));
 sg13g2_tiehi _5302__62 (.L_HI(net62));
 sg13g2_tiehi _5359__63 (.L_HI(net63));
 sg13g2_tiehi _5301__64 (.L_HI(net64));
 sg13g2_tiehi _5338__65 (.L_HI(net65));
 sg13g2_tiehi _5300__66 (.L_HI(net66));
 sg13g2_tiehi _5358__67 (.L_HI(net67));
 sg13g2_tiehi _5299__68 (.L_HI(net68));
 sg13g2_tiehi _5337__69 (.L_HI(net69));
 sg13g2_tiehi _5298__70 (.L_HI(net70));
 sg13g2_tiehi _5357__71 (.L_HI(net71));
 sg13g2_tiehi _5297__72 (.L_HI(net72));
 sg13g2_tiehi _5336__73 (.L_HI(net73));
 sg13g2_tiehi _5296__74 (.L_HI(net74));
 sg13g2_tiehi _5356__75 (.L_HI(net75));
 sg13g2_tiehi _5295__76 (.L_HI(net76));
 sg13g2_tiehi _5335__77 (.L_HI(net77));
 sg13g2_tiehi _5294__78 (.L_HI(net78));
 sg13g2_tiehi _5355__79 (.L_HI(net79));
 sg13g2_tiehi _5293__80 (.L_HI(net80));
 sg13g2_tiehi _5334__81 (.L_HI(net81));
 sg13g2_tiehi _5292__82 (.L_HI(net82));
 sg13g2_tiehi _5374__83 (.L_HI(net83));
 sg13g2_tiehi _5291__84 (.L_HI(net84));
 sg13g2_tiehi _5333__85 (.L_HI(net85));
 sg13g2_tiehi _5290__86 (.L_HI(net86));
 sg13g2_tiehi _5354__87 (.L_HI(net87));
 sg13g2_tiehi _5289__88 (.L_HI(net88));
 sg13g2_tiehi _5332__89 (.L_HI(net89));
 sg13g2_tiehi _5288__90 (.L_HI(net90));
 sg13g2_tiehi _5372__91 (.L_HI(net91));
 sg13g2_tiehi _5287__92 (.L_HI(net92));
 sg13g2_tiehi _5331__93 (.L_HI(net93));
 sg13g2_tiehi _5286__94 (.L_HI(net94));
 sg13g2_tiehi _5353__95 (.L_HI(net95));
 sg13g2_tiehi _5285__96 (.L_HI(net96));
 sg13g2_tiehi _5330__97 (.L_HI(net97));
 sg13g2_tiehi _5284__98 (.L_HI(net98));
 sg13g2_tiehi _5239__99 (.L_HI(net99));
 sg13g2_tiehi _5283__100 (.L_HI(net100));
 sg13g2_tiehi _5329__101 (.L_HI(net101));
 sg13g2_tiehi _5282__102 (.L_HI(net102));
 sg13g2_tiehi _5352__103 (.L_HI(net103));
 sg13g2_tiehi _5281__104 (.L_HI(net104));
 sg13g2_tiehi _5328__105 (.L_HI(net105));
 sg13g2_tiehi _5280__106 (.L_HI(net106));
 sg13g2_tiehi _5371__107 (.L_HI(net107));
 sg13g2_tiehi _5279__108 (.L_HI(net108));
 sg13g2_tiehi _5327__109 (.L_HI(net109));
 sg13g2_tiehi _5278__110 (.L_HI(net110));
 sg13g2_tiehi _5351__111 (.L_HI(net111));
 sg13g2_tiehi _5277__112 (.L_HI(net112));
 sg13g2_tiehi _5326__113 (.L_HI(net113));
 sg13g2_tiehi _5276__114 (.L_HI(net114));
 sg13g2_tiehi _5373__115 (.L_HI(net115));
 sg13g2_tiehi _5275__116 (.L_HI(net116));
 sg13g2_tiehi _5325__117 (.L_HI(net117));
 sg13g2_tiehi _5274__118 (.L_HI(net118));
 sg13g2_tiehi _5350__119 (.L_HI(net119));
 sg13g2_tiehi _5273__120 (.L_HI(net120));
 sg13g2_tiehi _5324__121 (.L_HI(net121));
 sg13g2_tiehi _5272__122 (.L_HI(net122));
 sg13g2_tiehi _5370__123 (.L_HI(net123));
 sg13g2_tiehi _5271__124 (.L_HI(net124));
 sg13g2_tiehi _5323__125 (.L_HI(net125));
 sg13g2_tiehi _5270__126 (.L_HI(net126));
 sg13g2_tiehi _5349__127 (.L_HI(net127));
 sg13g2_tiehi _5269__128 (.L_HI(net128));
 sg13g2_tiehi _5322__129 (.L_HI(net129));
 sg13g2_tiehi _5268__130 (.L_HI(net130));
 sg13g2_tiehi _5369__131 (.L_HI(net131));
 sg13g2_tiehi _5267__132 (.L_HI(net132));
 sg13g2_tiehi _5321__133 (.L_HI(net133));
 sg13g2_tiehi _5266__134 (.L_HI(net134));
 sg13g2_tiehi _5348__135 (.L_HI(net135));
 sg13g2_tiehi _5265__136 (.L_HI(net136));
 sg13g2_tiehi _5320__137 (.L_HI(net137));
 sg13g2_tiehi _5264__138 (.L_HI(net138));
 sg13g2_tiehi _5368__139 (.L_HI(net139));
 sg13g2_tiehi _5263__140 (.L_HI(net140));
 sg13g2_tiehi _5319__141 (.L_HI(net141));
 sg13g2_tiehi _5262__142 (.L_HI(net142));
 sg13g2_tiehi _5347__143 (.L_HI(net143));
 sg13g2_tiehi _5261__144 (.L_HI(net144));
 sg13g2_tiehi _5318__145 (.L_HI(net145));
 sg13g2_tiehi _5260__146 (.L_HI(net146));
 sg13g2_tiehi _5367__147 (.L_HI(net147));
 sg13g2_tiehi _5259__148 (.L_HI(net148));
 sg13g2_tiehi _5317__149 (.L_HI(net149));
 sg13g2_tiehi _5258__150 (.L_HI(net150));
 sg13g2_tiehi tt_um_couchand_cora16_151 (.L_HI(net151));
 sg13g2_tiehi tt_um_couchand_cora16_152 (.L_HI(net152));
 sg13g2_tiehi tt_um_couchand_cora16_153 (.L_HI(net153));
 sg13g2_inv_1 _2811__1 (.Y(net154),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_couchand_cora16_12 (.L_LO(net12));
 sg13g2_tielo tt_um_couchand_cora16_13 (.L_LO(net13));
 sg13g2_tielo tt_um_couchand_cora16_14 (.L_LO(net14));
 sg13g2_tiehi _5257__15 (.L_HI(net15));
 sg13g2_buf_1 _5518_ (.A(net1337),
    .X(uio_oe[0]));
 sg13g2_buf_1 _5519_ (.A(net1333),
    .X(uio_oe[1]));
 sg13g2_buf_1 _5520_ (.A(net1333),
    .X(uio_oe[2]));
 sg13g2_buf_2 _5521_ (.A(\cpu_instance.spi_mosi ),
    .X(uio_out[0]));
 sg13g2_buf_2 _5522_ (.A(net1273),
    .X(uio_out[1]));
 sg13g2_buf_1 _5523_ (.A(net154),
    .X(uio_out[2]));
 sg13g2_buf_1 _5524_ (.A(busy),
    .X(uio_out[5]));
 sg13g2_buf_1 _5525_ (.A(\cpu_instance.halt ),
    .X(uio_out[6]));
 sg13g2_buf_1 _5526_ (.A(\cpu_instance.trap ),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout1012 (.A(net1013),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_0969_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_0969_),
    .X(net1014));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(_0968_));
 sg13g2_buf_4 fanout1016 (.X(net1016),
    .A(_0821_));
 sg13g2_buf_4 fanout1017 (.X(net1017),
    .A(net1018));
 sg13g2_buf_2 fanout1018 (.A(_0649_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_0820_),
    .X(net1019));
 sg13g2_buf_1 fanout1020 (.A(_0820_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_0820_),
    .X(net1022));
 sg13g2_buf_4 fanout1023 (.X(net1023),
    .A(net1024));
 sg13g2_buf_4 fanout1024 (.X(net1024),
    .A(_0947_));
 sg13g2_buf_2 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_buf_1 fanout1026 (.A(_0512_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_0512_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_1584_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_1487_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_1486_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net1033),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(net1035),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_0948_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(net1037),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(net1038),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_0673_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(net1041),
    .X(net1040));
 sg13g2_buf_4 fanout1041 (.X(net1041),
    .A(_0611_));
 sg13g2_buf_2 fanout1042 (.A(net1043),
    .X(net1042));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(_0511_));
 sg13g2_buf_4 fanout1044 (.X(net1044),
    .A(_0510_));
 sg13g2_buf_2 fanout1045 (.A(net1047),
    .X(net1045));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(net1047));
 sg13g2_buf_2 fanout1047 (.A(_0804_),
    .X(net1047));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(_0672_));
 sg13g2_buf_2 fanout1049 (.A(net1050),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_0601_),
    .X(net1050));
 sg13g2_buf_4 fanout1051 (.X(net1051),
    .A(net1052));
 sg13g2_buf_2 fanout1052 (.A(_0593_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(net1054),
    .X(net1053));
 sg13g2_buf_1 fanout1054 (.A(net1055),
    .X(net1054));
 sg13g2_buf_1 fanout1055 (.A(_2404_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(net1057),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_2404_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(net1059),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_2319_),
    .X(net1059));
 sg13g2_buf_4 fanout1060 (.X(net1060),
    .A(_2148_));
 sg13g2_buf_2 fanout1061 (.A(net1062),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_0658_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_2441_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(net1066),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(net1066),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_2320_),
    .X(net1066));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(_2038_));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(_0986_));
 sg13g2_buf_2 fanout1069 (.A(_0659_),
    .X(net1069));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(_0567_));
 sg13g2_buf_2 fanout1071 (.A(net1072),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_0507_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_2357_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_1 fanout1076 (.A(_2357_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(net1078),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(net1081),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_1 fanout1081 (.A(_2356_),
    .X(net1081));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(net1084));
 sg13g2_buf_1 fanout1083 (.A(net1084),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_2343_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_1 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_2343_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(net1089),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(net1090),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(net1092),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_1 fanout1092 (.A(_2342_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_1 fanout1094 (.A(net1095),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_2330_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(net1098),
    .X(net1096));
 sg13g2_buf_1 fanout1097 (.A(net1098),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_2330_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(net1100),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(net1104),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(net1104),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(net1104),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_buf_1 fanout1104 (.A(_2329_),
    .X(net1104));
 sg13g2_buf_4 fanout1105 (.X(net1105),
    .A(_2295_));
 sg13g2_buf_2 fanout1106 (.A(net1107),
    .X(net1106));
 sg13g2_buf_1 fanout1107 (.A(_2103_),
    .X(net1107));
 sg13g2_buf_4 fanout1108 (.X(net1108),
    .A(_2103_));
 sg13g2_buf_2 fanout1109 (.A(_2019_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_2019_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_2015_),
    .X(net1111));
 sg13g2_buf_4 fanout1112 (.X(net1112),
    .A(_0959_));
 sg13g2_buf_4 fanout1113 (.X(net1113),
    .A(_0959_));
 sg13g2_buf_2 fanout1114 (.A(net1115),
    .X(net1114));
 sg13g2_buf_4 fanout1115 (.X(net1115),
    .A(net1117));
 sg13g2_buf_4 fanout1116 (.X(net1116),
    .A(net1117));
 sg13g2_buf_2 fanout1117 (.A(_0958_),
    .X(net1117));
 sg13g2_buf_4 fanout1118 (.X(net1118),
    .A(net1119));
 sg13g2_buf_4 fanout1119 (.X(net1119),
    .A(_0949_));
 sg13g2_buf_2 fanout1120 (.A(net1121),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_0806_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(net1124),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(net1125),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_0665_),
    .X(net1125));
 sg13g2_buf_4 fanout1126 (.X(net1126),
    .A(_0541_));
 sg13g2_buf_4 fanout1127 (.X(net1127),
    .A(_0494_));
 sg13g2_buf_2 fanout1128 (.A(net1129),
    .X(net1128));
 sg13g2_buf_1 fanout1129 (.A(net1130),
    .X(net1129));
 sg13g2_buf_1 fanout1130 (.A(net1131),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_0493_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(_2119_),
    .X(net1132));
 sg13g2_buf_1 fanout1133 (.A(_2119_),
    .X(net1133));
 sg13g2_buf_2 fanout1134 (.A(net1135),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(_0953_),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(_0953_),
    .X(net1136));
 sg13g2_buf_4 fanout1137 (.X(net1137),
    .A(_0807_));
 sg13g2_buf_2 fanout1138 (.A(net1139),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(_0787_),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(_0786_),
    .X(net1141));
 sg13g2_buf_4 fanout1142 (.X(net1142),
    .A(_0668_));
 sg13g2_buf_2 fanout1143 (.A(_0529_),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(net1145),
    .X(net1144));
 sg13g2_buf_4 fanout1145 (.X(net1145),
    .A(_0522_));
 sg13g2_buf_2 fanout1146 (.A(_0504_),
    .X(net1146));
 sg13g2_buf_2 fanout1147 (.A(net1148),
    .X(net1147));
 sg13g2_buf_1 fanout1148 (.A(_0501_),
    .X(net1148));
 sg13g2_buf_2 fanout1149 (.A(net1150),
    .X(net1149));
 sg13g2_buf_4 fanout1150 (.X(net1150),
    .A(_0500_));
 sg13g2_buf_2 fanout1151 (.A(_2391_),
    .X(net1151));
 sg13g2_buf_4 fanout1152 (.X(net1152),
    .A(_2391_));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(_2167_));
 sg13g2_buf_2 fanout1154 (.A(net1155),
    .X(net1154));
 sg13g2_buf_2 fanout1155 (.A(net1157),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(_2166_),
    .X(net1157));
 sg13g2_buf_2 fanout1158 (.A(_2138_),
    .X(net1158));
 sg13g2_buf_2 fanout1159 (.A(_2138_),
    .X(net1159));
 sg13g2_buf_2 fanout1160 (.A(net1161),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(_2126_),
    .X(net1161));
 sg13g2_buf_4 fanout1162 (.X(net1162),
    .A(_2125_));
 sg13g2_buf_2 fanout1163 (.A(_2125_),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(net1165),
    .X(net1164));
 sg13g2_buf_2 fanout1165 (.A(net1166),
    .X(net1165));
 sg13g2_buf_4 fanout1166 (.X(net1166),
    .A(_2118_));
 sg13g2_buf_4 fanout1167 (.X(net1167),
    .A(_0952_));
 sg13g2_buf_2 fanout1168 (.A(_0952_),
    .X(net1168));
 sg13g2_buf_2 fanout1169 (.A(_2451_),
    .X(net1169));
 sg13g2_buf_2 fanout1170 (.A(_2451_),
    .X(net1170));
 sg13g2_buf_2 fanout1171 (.A(_2395_),
    .X(net1171));
 sg13g2_buf_2 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_2 fanout1173 (.A(_2395_),
    .X(net1173));
 sg13g2_buf_2 fanout1174 (.A(_2268_),
    .X(net1174));
 sg13g2_buf_2 fanout1175 (.A(_2171_),
    .X(net1175));
 sg13g2_buf_2 fanout1176 (.A(net1177),
    .X(net1176));
 sg13g2_buf_2 fanout1177 (.A(_2115_),
    .X(net1177));
 sg13g2_buf_2 fanout1178 (.A(_2115_),
    .X(net1178));
 sg13g2_buf_1 fanout1179 (.A(_2115_),
    .X(net1179));
 sg13g2_buf_4 fanout1180 (.X(net1180),
    .A(_2096_));
 sg13g2_buf_2 fanout1181 (.A(net1182),
    .X(net1181));
 sg13g2_buf_2 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_2 fanout1183 (.A(_2076_),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(net1186),
    .X(net1184));
 sg13g2_buf_1 fanout1185 (.A(net1186),
    .X(net1185));
 sg13g2_buf_2 fanout1186 (.A(_2076_),
    .X(net1186));
 sg13g2_buf_2 fanout1187 (.A(net1188),
    .X(net1187));
 sg13g2_buf_1 fanout1188 (.A(net1189),
    .X(net1188));
 sg13g2_buf_2 fanout1189 (.A(net1193),
    .X(net1189));
 sg13g2_buf_4 fanout1190 (.X(net1190),
    .A(net1193));
 sg13g2_buf_4 fanout1191 (.X(net1191),
    .A(net1193));
 sg13g2_buf_2 fanout1192 (.A(net1193),
    .X(net1192));
 sg13g2_buf_2 fanout1193 (.A(_2075_),
    .X(net1193));
 sg13g2_buf_4 fanout1194 (.X(net1194),
    .A(net1195));
 sg13g2_buf_2 fanout1195 (.A(_2072_),
    .X(net1195));
 sg13g2_buf_2 fanout1196 (.A(_2072_),
    .X(net1196));
 sg13g2_buf_2 fanout1197 (.A(net1198),
    .X(net1197));
 sg13g2_buf_2 fanout1198 (.A(net1199),
    .X(net1198));
 sg13g2_buf_4 fanout1199 (.X(net1199),
    .A(_2071_));
 sg13g2_buf_2 fanout1200 (.A(_2054_),
    .X(net1200));
 sg13g2_buf_2 fanout1201 (.A(_2054_),
    .X(net1201));
 sg13g2_buf_2 fanout1202 (.A(net1203),
    .X(net1202));
 sg13g2_buf_2 fanout1203 (.A(net1204),
    .X(net1203));
 sg13g2_buf_4 fanout1204 (.X(net1204),
    .A(_2035_));
 sg13g2_buf_4 fanout1205 (.X(net1205),
    .A(_2030_));
 sg13g2_buf_2 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_4 fanout1207 (.X(net1207),
    .A(_2029_));
 sg13g2_buf_4 fanout1208 (.X(net1208),
    .A(_2025_));
 sg13g2_buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_4 fanout1210 (.X(net1210),
    .A(_2025_));
 sg13g2_buf_2 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_2 fanout1212 (.A(net1213),
    .X(net1212));
 sg13g2_buf_4 fanout1213 (.X(net1213),
    .A(_2006_));
 sg13g2_buf_2 fanout1214 (.A(net1215),
    .X(net1214));
 sg13g2_buf_4 fanout1215 (.X(net1215),
    .A(_2005_));
 sg13g2_buf_2 fanout1216 (.A(net1219),
    .X(net1216));
 sg13g2_buf_2 fanout1217 (.A(net1219),
    .X(net1217));
 sg13g2_buf_2 fanout1218 (.A(net1219),
    .X(net1218));
 sg13g2_buf_2 fanout1219 (.A(net1220),
    .X(net1219));
 sg13g2_buf_4 fanout1220 (.X(net1220),
    .A(_0927_));
 sg13g2_buf_4 fanout1221 (.X(net1221),
    .A(net1222));
 sg13g2_buf_2 fanout1222 (.A(_2168_),
    .X(net1222));
 sg13g2_buf_2 fanout1223 (.A(_2123_),
    .X(net1223));
 sg13g2_buf_2 fanout1224 (.A(_2123_),
    .X(net1224));
 sg13g2_buf_4 fanout1225 (.X(net1225),
    .A(net1227));
 sg13g2_buf_2 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_buf_4 fanout1227 (.X(net1227),
    .A(_2108_));
 sg13g2_buf_2 fanout1228 (.A(net1229),
    .X(net1228));
 sg13g2_buf_2 fanout1229 (.A(_2107_),
    .X(net1229));
 sg13g2_buf_2 fanout1230 (.A(_2107_),
    .X(net1230));
 sg13g2_buf_4 fanout1231 (.X(net1231),
    .A(net1232));
 sg13g2_buf_2 fanout1232 (.A(_2082_),
    .X(net1232));
 sg13g2_buf_4 fanout1233 (.X(net1233),
    .A(_2082_));
 sg13g2_buf_2 fanout1234 (.A(net1235),
    .X(net1234));
 sg13g2_buf_4 fanout1235 (.X(net1235),
    .A(net1236));
 sg13g2_buf_4 fanout1236 (.X(net1236),
    .A(net1240));
 sg13g2_buf_4 fanout1237 (.X(net1237),
    .A(net1238));
 sg13g2_buf_4 fanout1238 (.X(net1238),
    .A(net1240));
 sg13g2_buf_4 fanout1239 (.X(net1239),
    .A(net1240));
 sg13g2_buf_2 fanout1240 (.A(_2080_),
    .X(net1240));
 sg13g2_buf_4 fanout1241 (.X(net1241),
    .A(net1252));
 sg13g2_buf_2 fanout1242 (.A(net1252),
    .X(net1242));
 sg13g2_buf_2 fanout1243 (.A(net1244),
    .X(net1243));
 sg13g2_buf_2 fanout1244 (.A(net1245),
    .X(net1244));
 sg13g2_buf_1 fanout1245 (.A(net1246),
    .X(net1245));
 sg13g2_buf_2 fanout1246 (.A(net1252),
    .X(net1246));
 sg13g2_buf_2 fanout1247 (.A(net1248),
    .X(net1247));
 sg13g2_buf_4 fanout1248 (.X(net1248),
    .A(net1252));
 sg13g2_buf_2 fanout1249 (.A(net1250),
    .X(net1249));
 sg13g2_buf_1 fanout1250 (.A(net1251),
    .X(net1250));
 sg13g2_buf_2 fanout1251 (.A(net1252),
    .X(net1251));
 sg13g2_buf_4 fanout1252 (.X(net1252),
    .A(_2079_));
 sg13g2_buf_2 fanout1253 (.A(_2051_),
    .X(net1253));
 sg13g2_buf_2 fanout1254 (.A(net1256),
    .X(net1254));
 sg13g2_buf_1 fanout1255 (.A(net1256),
    .X(net1255));
 sg13g2_buf_4 fanout1256 (.X(net1256),
    .A(_0657_));
 sg13g2_buf_2 fanout1257 (.A(net1258),
    .X(net1257));
 sg13g2_buf_2 fanout1258 (.A(net1259),
    .X(net1258));
 sg13g2_buf_4 fanout1259 (.X(net1259),
    .A(_0656_));
 sg13g2_buf_2 fanout1260 (.A(net1261),
    .X(net1260));
 sg13g2_buf_1 fanout1261 (.A(net1262),
    .X(net1261));
 sg13g2_buf_2 fanout1262 (.A(_2175_),
    .X(net1262));
 sg13g2_buf_2 fanout1263 (.A(net1266),
    .X(net1263));
 sg13g2_buf_4 fanout1264 (.X(net1264),
    .A(net1266));
 sg13g2_buf_2 fanout1265 (.A(net1266),
    .X(net1265));
 sg13g2_buf_2 fanout1266 (.A(_1995_),
    .X(net1266));
 sg13g2_buf_4 fanout1267 (.X(net1267),
    .A(net1269));
 sg13g2_buf_2 fanout1268 (.A(net1269),
    .X(net1268));
 sg13g2_buf_4 fanout1269 (.X(net1269),
    .A(net1272));
 sg13g2_buf_2 fanout1270 (.A(net1272),
    .X(net1270));
 sg13g2_buf_1 fanout1271 (.A(net1272),
    .X(net1271));
 sg13g2_buf_2 fanout1272 (.A(_1994_),
    .X(net1272));
 sg13g2_buf_4 fanout1273 (.X(net1273),
    .A(\cpu_instance.spi_ram.spi_select ));
 sg13g2_buf_2 fanout1274 (.A(net1275),
    .X(net1274));
 sg13g2_buf_4 fanout1275 (.X(net1275),
    .A(_1987_));
 sg13g2_buf_2 fanout1276 (.A(_1986_),
    .X(net1276));
 sg13g2_buf_4 fanout1277 (.X(net1277),
    .A(_1974_));
 sg13g2_buf_4 fanout1278 (.X(net1278),
    .A(_1943_));
 sg13g2_buf_2 fanout1279 (.A(_1943_),
    .X(net1279));
 sg13g2_buf_4 fanout1280 (.X(net1280),
    .A(_1943_));
 sg13g2_buf_4 fanout1281 (.X(net1281),
    .A(_1907_));
 sg13g2_buf_2 fanout1282 (.A(net317),
    .X(net1282));
 sg13g2_buf_2 fanout1283 (.A(\cpu_instance.sp[1] ),
    .X(net1283));
 sg13g2_buf_4 fanout1284 (.X(net1284),
    .A(_0012_));
 sg13g2_buf_4 fanout1285 (.X(net1285),
    .A(net315));
 sg13g2_buf_2 fanout1286 (.A(\cpu_instance.inst[14] ),
    .X(net1286));
 sg13g2_buf_2 fanout1287 (.A(\cpu_instance.inst[13] ),
    .X(net1287));
 sg13g2_buf_4 fanout1288 (.X(net1288),
    .A(\cpu_instance.inst[12] ));
 sg13g2_buf_2 fanout1289 (.A(\cpu_instance.inst[12] ),
    .X(net1289));
 sg13g2_buf_2 fanout1290 (.A(net1291),
    .X(net1290));
 sg13g2_buf_4 fanout1291 (.X(net1291),
    .A(\cpu_instance.inst[11] ));
 sg13g2_buf_2 fanout1292 (.A(net1293),
    .X(net1292));
 sg13g2_buf_2 fanout1293 (.A(\cpu_instance.inst[10] ),
    .X(net1293));
 sg13g2_buf_2 fanout1294 (.A(net1296),
    .X(net1294));
 sg13g2_buf_1 fanout1295 (.A(net1296),
    .X(net1295));
 sg13g2_buf_1 fanout1296 (.A(net1297),
    .X(net1296));
 sg13g2_buf_2 fanout1297 (.A(net1300),
    .X(net1297));
 sg13g2_buf_4 fanout1298 (.X(net1298),
    .A(net1300));
 sg13g2_buf_1 fanout1299 (.A(net1300),
    .X(net1299));
 sg13g2_buf_4 fanout1300 (.X(net1300),
    .A(net306));
 sg13g2_buf_2 fanout1301 (.A(net1302),
    .X(net1301));
 sg13g2_buf_4 fanout1302 (.X(net1302),
    .A(net1303));
 sg13g2_buf_2 fanout1303 (.A(\cpu_instance.inst[8] ),
    .X(net1303));
 sg13g2_buf_4 fanout1304 (.X(net1304),
    .A(\cpu_instance.accum[13] ));
 sg13g2_buf_4 fanout1305 (.X(net1305),
    .A(\cpu_instance.accum[12] ));
 sg13g2_buf_2 fanout1306 (.A(\cpu_instance.accum[11] ),
    .X(net1306));
 sg13g2_buf_4 fanout1307 (.X(net1307),
    .A(net1308));
 sg13g2_buf_4 fanout1308 (.X(net1308),
    .A(\cpu_instance.accum[10] ));
 sg13g2_buf_4 fanout1309 (.X(net1309),
    .A(\cpu_instance.accum[9] ));
 sg13g2_buf_4 fanout1310 (.X(net1310),
    .A(net1311));
 sg13g2_buf_4 fanout1311 (.X(net1311),
    .A(\cpu_instance.accum[8] ));
 sg13g2_buf_2 fanout1312 (.A(\cpu_instance.accum[6] ),
    .X(net1312));
 sg13g2_buf_2 fanout1313 (.A(_0035_),
    .X(net1313));
 sg13g2_buf_2 fanout1314 (.A(net1316),
    .X(net1314));
 sg13g2_buf_1 fanout1315 (.A(net1316),
    .X(net1315));
 sg13g2_buf_1 fanout1316 (.A(net1317),
    .X(net1316));
 sg13g2_buf_2 fanout1317 (.A(net1318),
    .X(net1317));
 sg13g2_buf_2 fanout1318 (.A(\cpu_instance.skip ),
    .X(net1318));
 sg13g2_buf_2 fanout1319 (.A(net1321),
    .X(net1319));
 sg13g2_buf_2 fanout1320 (.A(net1321),
    .X(net1320));
 sg13g2_buf_4 fanout1321 (.X(net1321),
    .A(\cpu_instance.skip ));
 sg13g2_buf_4 fanout1322 (.X(net1322),
    .A(_1973_));
 sg13g2_buf_2 fanout1323 (.A(_1973_),
    .X(net1323));
 sg13g2_buf_4 fanout1324 (.X(net1324),
    .A(net1325));
 sg13g2_buf_4 fanout1325 (.X(net1325),
    .A(net1326));
 sg13g2_buf_4 fanout1326 (.X(net1326),
    .A(_1973_));
 sg13g2_buf_2 fanout1327 (.A(net1330),
    .X(net1327));
 sg13g2_buf_2 fanout1328 (.A(net1329),
    .X(net1328));
 sg13g2_buf_2 fanout1329 (.A(net1330),
    .X(net1329));
 sg13g2_buf_2 fanout1330 (.A(net1331),
    .X(net1330));
 sg13g2_buf_4 fanout1331 (.X(net1331),
    .A(rst_n));
 sg13g2_buf_4 fanout1332 (.X(net1332),
    .A(net1338));
 sg13g2_buf_4 fanout1333 (.X(net1333),
    .A(net1337));
 sg13g2_buf_2 fanout1334 (.A(net1337),
    .X(net1334));
 sg13g2_buf_2 fanout1335 (.A(net1336),
    .X(net1335));
 sg13g2_buf_4 fanout1336 (.X(net1336),
    .A(net1337));
 sg13g2_buf_4 fanout1337 (.X(net1337),
    .A(net1338));
 sg13g2_buf_2 fanout1338 (.A(rst_n),
    .X(net1338));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_tielo tt_um_couchand_cora16_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_9__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_17__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_21__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cpu_instance.dp[12] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold2 (.A(\cpu_instance.spi_ram.addr[1] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0171_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold4 (.A(\cpu_instance.dp[10] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cpu_instance.dp[13] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold6 (.A(\cpu_instance.dp[8] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cpu_instance.spi_ram.addr[0] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0185_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cpu_instance.dp[6] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cpu_instance.spi_ram.addr[5] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0174_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cpu_instance.spi_ram.addr[14] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0183_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cpu_instance.spi_ram.addr[13] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0182_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cpu_instance.pc[1] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold17 (.A(\cpu_instance.spi_ram.addr[7] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0176_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold19 (.A(\cpu_instance.spi_ram.addr[15] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0184_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cpu_instance.spi_ram.addr[11] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0180_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold23 (.A(\cpu_instance.spi_ram.bits_remaining[0] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cpu_instance.spi_ram.addr[8] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold25 (.A(\cpu_instance.dp[3] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold26 (.A(\cpu_instance.spi_ram.bits_remaining[1] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cpu_instance.dp[4] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0087_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cpu_instance.dp[9] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cpu_instance.dp[1] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cpu_instance.dp[7] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cpu_instance.spi_ram.addr[3] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold33 (.A(_1635_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu_instance.sp_minus_two[1] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0155_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cpu_instance.dp[0] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0083_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cpu_instance.dp[14] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cpu_instance.dp[5] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cpu_instance.spi_ram.addr[9] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cpu_instance.dp[11] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold42 (.A(\cpu_instance.spi_ram.writing ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu_instance.dp[2] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0085_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold45 (.A(\cpu_instance.spi_ram.addr[6] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cpu_instance.dp[15] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cpu_instance.spi_ram.addr[12] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cpu_instance.spi_ram.addr[4] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold49 (.A(uo_out[7]),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold50 (.A(_1477_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0154_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cpu_instance.spi_ram.bits_remaining[3] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold53 (.A(\cpu_instance.pc[11] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu_instance.spi_ram.addr[10] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu_instance.pc[0] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold56 (.A(uo_out[6]),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold57 (.A(_1474_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0153_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cpu_instance.inst[7] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0122_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cpu_instance.inst[4] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0119_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu_instance.inst[2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0117_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cpu_instance.spi_ram.fsm_state[1] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0679_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cpu_instance.inst[6] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0121_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold69 (.A(uo_out[0]),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold70 (.A(_1456_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0147_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold72 (.A(uo_out[1]),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold73 (.A(_1459_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0148_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold75 (.A(uo_out[2]),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold76 (.A(_1462_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0149_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold78 (.A(uo_out[4]),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold79 (.A(_1468_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0151_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold81 (.A(uo_out[3]),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold82 (.A(_1465_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0150_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cpu_instance.sp[9] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0163_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold86 (.A(uo_out[5]),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold87 (.A(_1471_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0152_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cpu_instance.pc[5] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cpu_instance.ram_data_out[0] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0520_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0057_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu_instance.ram_data_out[9] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0065_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu_instance.inst[3] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0118_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu_instance.spi_ram.fsm_state[0] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0073_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cpu_instance.ram_data_out[11] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0067_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cpu_instance.sp[13] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cpu_instance.ram_data_out[6] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0564_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu_instance.inst[1] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cpu_instance.zero ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cpu_instance.sp[12] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cpu_instance.skipped ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0004_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0164_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cpu_instance.inst[5] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0120_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cpu_instance.neg ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cpu_instance.spi_ram.bits_remaining[2] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0077_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cpu_instance.pc[15] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold116 (.A(\cpu_instance.state[3] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cpu_instance.pc[13] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cpu_instance.sp[14] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cpu_instance.pc[14] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cpu_instance.inst[0] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold121 (.A(\cpu_instance.ram_data_out[13] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0069_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cpu_instance.ram_data_out[15] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cpu_instance.sp[15] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cpu_instance.sp[4] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu_instance.ram_data_out[12] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0127_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cpu_instance.ram_data_out[5] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cpu_instance.ram_data_out[4] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0060_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold131 (.A(\cpu_instance.sp[7] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cpu_instance.sp[6] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold133 (.A(\cpu_instance.pc[10] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cpu_instance.pc[9] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold135 (.A(\cpu_instance.ram_data_out[1] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold136 (.A(\cpu_instance.sp[5] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0159_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cpu_instance.state[0] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0186_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cpu_instance.pc[8] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cpu_instance.state[1] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu_instance.ram_data_out[8] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0123_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu_instance.ram_data_out[7] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cpu_instance.ram_data_out[2] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cpu_instance.sp[8] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cpu_instance.sp[3] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold148 (.A(\cpu_instance.pc[2] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu_instance.pc[12] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cpu_instance.carry ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cpu_instance.inst[9] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cpu_instance.ram_data_out[10] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cpu_instance.pc[4] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cpu_instance.ram_data_out[3] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0059_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cpu_instance.sp[11] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold157 (.A(\cpu_instance.pc[3] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cpu_instance.accum[2] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold159 (.A(\cpu_instance.pc[7] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold160 (.A(\cpu_instance.inst[15] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold161 (.A(\cpu_instance.sp[2] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cpu_instance.state[2] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cpu_instance.accum[3] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu_instance.spi_ram.bits_remaining[2] ),
    .X(net319));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_fill_1 FILLER_0_105 ();
 sg13g2_fill_2 FILLER_0_134 ();
 sg13g2_fill_1 FILLER_0_136 ();
 sg13g2_fill_2 FILLER_0_153 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_4 FILLER_0_189 ();
 sg13g2_fill_1 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_219 ();
 sg13g2_decap_8 FILLER_0_226 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_decap_8 FILLER_0_240 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_4 FILLER_1_98 ();
 sg13g2_fill_1 FILLER_1_102 ();
 sg13g2_fill_2 FILLER_1_146 ();
 sg13g2_fill_1 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_209 ();
 sg13g2_decap_8 FILLER_1_216 ();
 sg13g2_decap_8 FILLER_1_223 ();
 sg13g2_decap_8 FILLER_1_230 ();
 sg13g2_decap_8 FILLER_1_237 ();
 sg13g2_decap_8 FILLER_1_244 ();
 sg13g2_decap_8 FILLER_1_251 ();
 sg13g2_decap_8 FILLER_1_258 ();
 sg13g2_decap_8 FILLER_1_265 ();
 sg13g2_decap_8 FILLER_1_272 ();
 sg13g2_decap_8 FILLER_1_279 ();
 sg13g2_decap_8 FILLER_1_286 ();
 sg13g2_decap_8 FILLER_1_293 ();
 sg13g2_decap_8 FILLER_1_300 ();
 sg13g2_decap_8 FILLER_1_307 ();
 sg13g2_decap_8 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_4 FILLER_2_91 ();
 sg13g2_fill_2 FILLER_2_174 ();
 sg13g2_fill_2 FILLER_2_181 ();
 sg13g2_fill_1 FILLER_2_183 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_fill_2 FILLER_3_77 ();
 sg13g2_fill_2 FILLER_3_152 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_fill_1 FILLER_4_77 ();
 sg13g2_fill_1 FILLER_4_121 ();
 sg13g2_fill_1 FILLER_4_127 ();
 sg13g2_fill_2 FILLER_4_151 ();
 sg13g2_fill_1 FILLER_4_182 ();
 sg13g2_fill_2 FILLER_4_204 ();
 sg13g2_fill_1 FILLER_4_206 ();
 sg13g2_decap_8 FILLER_4_215 ();
 sg13g2_decap_8 FILLER_4_222 ();
 sg13g2_decap_8 FILLER_4_229 ();
 sg13g2_decap_8 FILLER_4_236 ();
 sg13g2_decap_8 FILLER_4_243 ();
 sg13g2_decap_8 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_257 ();
 sg13g2_decap_8 FILLER_4_264 ();
 sg13g2_decap_8 FILLER_4_271 ();
 sg13g2_decap_8 FILLER_4_278 ();
 sg13g2_decap_8 FILLER_4_285 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_decap_8 FILLER_4_299 ();
 sg13g2_decap_8 FILLER_4_306 ();
 sg13g2_decap_8 FILLER_4_313 ();
 sg13g2_decap_8 FILLER_4_320 ();
 sg13g2_decap_8 FILLER_4_327 ();
 sg13g2_decap_8 FILLER_4_334 ();
 sg13g2_decap_8 FILLER_4_341 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_4 FILLER_5_77 ();
 sg13g2_fill_1 FILLER_5_81 ();
 sg13g2_fill_2 FILLER_5_95 ();
 sg13g2_fill_1 FILLER_5_110 ();
 sg13g2_fill_2 FILLER_5_118 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_fill_1 FILLER_5_195 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_8 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_decap_8 FILLER_5_251 ();
 sg13g2_decap_8 FILLER_5_258 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_300 ();
 sg13g2_decap_8 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_fill_1 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_97 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_fill_1 FILLER_6_146 ();
 sg13g2_fill_1 FILLER_6_161 ();
 sg13g2_fill_2 FILLER_6_220 ();
 sg13g2_fill_2 FILLER_6_251 ();
 sg13g2_fill_1 FILLER_6_253 ();
 sg13g2_decap_8 FILLER_6_258 ();
 sg13g2_decap_8 FILLER_6_265 ();
 sg13g2_decap_8 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_279 ();
 sg13g2_decap_8 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_293 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_fill_1 FILLER_7_84 ();
 sg13g2_fill_2 FILLER_7_133 ();
 sg13g2_fill_2 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_195 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_271 ();
 sg13g2_decap_8 FILLER_7_278 ();
 sg13g2_decap_8 FILLER_7_285 ();
 sg13g2_decap_8 FILLER_7_292 ();
 sg13g2_decap_8 FILLER_7_299 ();
 sg13g2_decap_8 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_decap_8 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_decap_8 FILLER_7_348 ();
 sg13g2_decap_8 FILLER_7_355 ();
 sg13g2_decap_8 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_369 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_fill_2 FILLER_8_70 ();
 sg13g2_fill_2 FILLER_8_107 ();
 sg13g2_fill_1 FILLER_8_109 ();
 sg13g2_fill_1 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_156 ();
 sg13g2_fill_1 FILLER_8_166 ();
 sg13g2_decap_8 FILLER_8_190 ();
 sg13g2_decap_4 FILLER_8_201 ();
 sg13g2_fill_1 FILLER_8_209 ();
 sg13g2_fill_1 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_288 ();
 sg13g2_decap_8 FILLER_8_295 ();
 sg13g2_decap_8 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_309 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_decap_8 FILLER_8_323 ();
 sg13g2_decap_8 FILLER_8_330 ();
 sg13g2_decap_8 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_fill_1 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_68 ();
 sg13g2_decap_4 FILLER_9_75 ();
 sg13g2_fill_2 FILLER_9_92 ();
 sg13g2_fill_1 FILLER_9_94 ();
 sg13g2_decap_8 FILLER_9_134 ();
 sg13g2_fill_2 FILLER_9_141 ();
 sg13g2_decap_4 FILLER_9_152 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_decap_8 FILLER_9_183 ();
 sg13g2_fill_2 FILLER_9_190 ();
 sg13g2_fill_1 FILLER_9_208 ();
 sg13g2_fill_2 FILLER_9_219 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_fill_1 FILLER_10_49 ();
 sg13g2_decap_4 FILLER_10_151 ();
 sg13g2_fill_1 FILLER_10_155 ();
 sg13g2_decap_4 FILLER_10_180 ();
 sg13g2_fill_1 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_1 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_285 ();
 sg13g2_decap_8 FILLER_10_292 ();
 sg13g2_decap_8 FILLER_10_299 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_125 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_fill_2 FILLER_11_171 ();
 sg13g2_fill_2 FILLER_11_201 ();
 sg13g2_fill_1 FILLER_11_203 ();
 sg13g2_fill_1 FILLER_11_223 ();
 sg13g2_fill_1 FILLER_11_244 ();
 sg13g2_fill_1 FILLER_11_260 ();
 sg13g2_fill_1 FILLER_11_271 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_4 FILLER_12_28 ();
 sg13g2_fill_1 FILLER_12_58 ();
 sg13g2_fill_2 FILLER_12_123 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_153 ();
 sg13g2_fill_1 FILLER_12_169 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_fill_2 FILLER_12_219 ();
 sg13g2_fill_1 FILLER_12_221 ();
 sg13g2_fill_1 FILLER_12_253 ();
 sg13g2_decap_4 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_decap_8 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_21 ();
 sg13g2_fill_1 FILLER_13_23 ();
 sg13g2_fill_2 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_87 ();
 sg13g2_fill_1 FILLER_13_108 ();
 sg13g2_fill_2 FILLER_13_114 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_fill_1 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_151 ();
 sg13g2_fill_2 FILLER_13_156 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_164 ();
 sg13g2_fill_1 FILLER_13_166 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_fill_2 FILLER_13_268 ();
 sg13g2_fill_1 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_4 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_25 ();
 sg13g2_fill_2 FILLER_14_65 ();
 sg13g2_fill_1 FILLER_14_76 ();
 sg13g2_fill_2 FILLER_14_82 ();
 sg13g2_fill_2 FILLER_14_89 ();
 sg13g2_decap_8 FILLER_14_110 ();
 sg13g2_decap_8 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_fill_2 FILLER_14_131 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_152 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_240 ();
 sg13g2_decap_8 FILLER_14_295 ();
 sg13g2_decap_8 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_309 ();
 sg13g2_decap_8 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_323 ();
 sg13g2_decap_8 FILLER_14_330 ();
 sg13g2_decap_8 FILLER_14_337 ();
 sg13g2_decap_8 FILLER_14_344 ();
 sg13g2_decap_8 FILLER_14_351 ();
 sg13g2_decap_8 FILLER_14_358 ();
 sg13g2_decap_8 FILLER_14_365 ();
 sg13g2_decap_8 FILLER_14_372 ();
 sg13g2_decap_8 FILLER_14_379 ();
 sg13g2_decap_8 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_fill_2 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_23 ();
 sg13g2_fill_2 FILLER_15_90 ();
 sg13g2_fill_1 FILLER_15_92 ();
 sg13g2_fill_2 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_107 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_187 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_fill_1 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_216 ();
 sg13g2_fill_2 FILLER_15_229 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_30 ();
 sg13g2_fill_2 FILLER_16_57 ();
 sg13g2_fill_1 FILLER_16_73 ();
 sg13g2_fill_1 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_133 ();
 sg13g2_fill_1 FILLER_16_170 ();
 sg13g2_decap_8 FILLER_16_176 ();
 sg13g2_fill_1 FILLER_16_183 ();
 sg13g2_fill_2 FILLER_16_216 ();
 sg13g2_fill_1 FILLER_16_218 ();
 sg13g2_fill_1 FILLER_16_227 ();
 sg13g2_fill_1 FILLER_16_264 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_46 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_decap_4 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_decap_4 FILLER_17_206 ();
 sg13g2_fill_1 FILLER_17_227 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_fill_2 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_264 ();
 sg13g2_decap_4 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_fill_2 FILLER_18_88 ();
 sg13g2_fill_1 FILLER_18_90 ();
 sg13g2_fill_1 FILLER_18_100 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_4 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_4 FILLER_18_158 ();
 sg13g2_fill_2 FILLER_18_162 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_decap_8 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_decap_4 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_4 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_67 ();
 sg13g2_fill_2 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_decap_4 FILLER_19_117 ();
 sg13g2_fill_1 FILLER_19_121 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_fill_2 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_fill_2 FILLER_20_66 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_116 ();
 sg13g2_fill_1 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_186 ();
 sg13g2_fill_2 FILLER_20_209 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_2 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_fill_2 FILLER_20_309 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_37 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_fill_1 FILLER_21_74 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_fill_2 FILLER_21_137 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_decap_8 FILLER_21_160 ();
 sg13g2_fill_2 FILLER_21_167 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_fill_2 FILLER_21_190 ();
 sg13g2_fill_1 FILLER_21_192 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_fill_1 FILLER_21_205 ();
 sg13g2_decap_8 FILLER_21_220 ();
 sg13g2_decap_4 FILLER_21_227 ();
 sg13g2_fill_2 FILLER_21_267 ();
 sg13g2_decap_4 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_92 ();
 sg13g2_fill_1 FILLER_22_96 ();
 sg13g2_fill_2 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_fill_1 FILLER_22_116 ();
 sg13g2_decap_4 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_222 ();
 sg13g2_fill_1 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_30 ();
 sg13g2_fill_2 FILLER_23_107 ();
 sg13g2_fill_1 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_118 ();
 sg13g2_decap_4 FILLER_23_125 ();
 sg13g2_decap_8 FILLER_23_138 ();
 sg13g2_decap_4 FILLER_23_145 ();
 sg13g2_fill_2 FILLER_23_159 ();
 sg13g2_fill_2 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_172 ();
 sg13g2_decap_4 FILLER_23_185 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_255 ();
 sg13g2_fill_2 FILLER_23_272 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_decap_4 FILLER_23_305 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_decap_4 FILLER_24_109 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_decap_4 FILLER_24_160 ();
 sg13g2_fill_1 FILLER_24_164 ();
 sg13g2_fill_2 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_2 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_226 ();
 sg13g2_fill_2 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_decap_4 FILLER_24_290 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_302 ();
 sg13g2_decap_4 FILLER_24_330 ();
 sg13g2_fill_2 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_fill_1 FILLER_25_88 ();
 sg13g2_fill_2 FILLER_25_93 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_123 ();
 sg13g2_decap_4 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_2 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_37 ();
 sg13g2_fill_2 FILLER_26_64 ();
 sg13g2_fill_2 FILLER_26_103 ();
 sg13g2_fill_2 FILLER_26_115 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_decap_8 FILLER_26_128 ();
 sg13g2_decap_4 FILLER_26_135 ();
 sg13g2_fill_2 FILLER_26_139 ();
 sg13g2_fill_2 FILLER_26_156 ();
 sg13g2_fill_1 FILLER_26_182 ();
 sg13g2_decap_4 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_203 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_fill_2 FILLER_26_276 ();
 sg13g2_fill_1 FILLER_26_278 ();
 sg13g2_decap_8 FILLER_26_289 ();
 sg13g2_fill_2 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_fill_2 FILLER_27_79 ();
 sg13g2_fill_2 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_129 ();
 sg13g2_fill_2 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_157 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_247 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_decap_4 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_296 ();
 sg13g2_decap_8 FILLER_27_303 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_340 ();
 sg13g2_fill_2 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_86 ();
 sg13g2_fill_1 FILLER_28_99 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_122 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_decap_4 FILLER_28_220 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_decap_4 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_323 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_156 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_decap_4 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_decap_4 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_decap_4 FILLER_29_313 ();
 sg13g2_fill_1 FILLER_29_317 ();
 sg13g2_fill_2 FILLER_29_323 ();
 sg13g2_fill_1 FILLER_29_325 ();
 sg13g2_decap_8 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_95 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_121 ();
 sg13g2_fill_1 FILLER_30_132 ();
 sg13g2_decap_4 FILLER_30_148 ();
 sg13g2_fill_2 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_decap_8 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_191 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_decap_4 FILLER_30_226 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_decap_4 FILLER_30_235 ();
 sg13g2_decap_4 FILLER_30_279 ();
 sg13g2_decap_4 FILLER_30_291 ();
 sg13g2_fill_2 FILLER_30_308 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_fill_1 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_47 ();
 sg13g2_fill_2 FILLER_31_116 ();
 sg13g2_fill_2 FILLER_31_127 ();
 sg13g2_fill_1 FILLER_31_129 ();
 sg13g2_decap_8 FILLER_31_134 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_decap_4 FILLER_31_149 ();
 sg13g2_decap_4 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_decap_4 FILLER_31_195 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_decap_4 FILLER_31_217 ();
 sg13g2_decap_4 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_366 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_4 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_fill_2 FILLER_32_54 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_68 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_fill_1 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_fill_1 FILLER_32_116 ();
 sg13g2_decap_4 FILLER_32_121 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_decap_4 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_221 ();
 sg13g2_fill_1 FILLER_32_315 ();
 sg13g2_fill_2 FILLER_32_325 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_4 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_374 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_80 ();
 sg13g2_fill_2 FILLER_33_139 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_153 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_decap_4 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_184 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_2 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_decap_4 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_2 FILLER_33_276 ();
 sg13g2_fill_2 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_291 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_decap_8 FILLER_33_334 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_52 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_fill_2 FILLER_34_113 ();
 sg13g2_fill_2 FILLER_34_143 ();
 sg13g2_fill_1 FILLER_34_158 ();
 sg13g2_fill_2 FILLER_34_174 ();
 sg13g2_decap_8 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_4 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_decap_4 FILLER_34_229 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_4 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_fill_1 FILLER_34_269 ();
 sg13g2_decap_8 FILLER_34_276 ();
 sg13g2_decap_4 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_4 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_93 ();
 sg13g2_fill_2 FILLER_35_128 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_153 ();
 sg13g2_fill_1 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_204 ();
 sg13g2_fill_1 FILLER_35_211 ();
 sg13g2_fill_2 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_219 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_decap_4 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_fill_1 FILLER_35_253 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_4 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_4 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_61 ();
 sg13g2_decap_8 FILLER_36_81 ();
 sg13g2_fill_2 FILLER_36_88 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_decap_8 FILLER_36_139 ();
 sg13g2_decap_4 FILLER_36_150 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_decap_4 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_207 ();
 sg13g2_fill_2 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_229 ();
 sg13g2_fill_1 FILLER_36_234 ();
 sg13g2_decap_4 FILLER_36_310 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_2 FILLER_36_325 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_decap_8 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_82 ();
 sg13g2_fill_2 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_decap_4 FILLER_37_106 ();
 sg13g2_fill_1 FILLER_37_110 ();
 sg13g2_fill_1 FILLER_37_141 ();
 sg13g2_decap_4 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_184 ();
 sg13g2_fill_2 FILLER_37_200 ();
 sg13g2_decap_4 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_245 ();
 sg13g2_fill_2 FILLER_37_254 ();
 sg13g2_fill_1 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_293 ();
 sg13g2_decap_8 FILLER_37_299 ();
 sg13g2_decap_8 FILLER_37_310 ();
 sg13g2_decap_8 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_324 ();
 sg13g2_decap_4 FILLER_37_331 ();
 sg13g2_fill_2 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_37_366 ();
 sg13g2_decap_8 FILLER_37_373 ();
 sg13g2_fill_2 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_56 ();
 sg13g2_fill_1 FILLER_38_81 ();
 sg13g2_fill_1 FILLER_38_101 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_138 ();
 sg13g2_decap_4 FILLER_38_145 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_162 ();
 sg13g2_decap_4 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_fill_1 FILLER_38_186 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_233 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_283 ();
 sg13g2_decap_4 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_2 FILLER_38_311 ();
 sg13g2_decap_4 FILLER_38_317 ();
 sg13g2_fill_2 FILLER_38_321 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_367 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_fill_2 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_fill_1 FILLER_39_84 ();
 sg13g2_fill_2 FILLER_39_120 ();
 sg13g2_fill_1 FILLER_39_122 ();
 sg13g2_decap_8 FILLER_39_127 ();
 sg13g2_decap_4 FILLER_39_134 ();
 sg13g2_fill_2 FILLER_39_138 ();
 sg13g2_decap_4 FILLER_39_144 ();
 sg13g2_fill_2 FILLER_39_148 ();
 sg13g2_fill_1 FILLER_39_190 ();
 sg13g2_decap_8 FILLER_39_211 ();
 sg13g2_fill_2 FILLER_39_218 ();
 sg13g2_fill_1 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_226 ();
 sg13g2_decap_8 FILLER_39_233 ();
 sg13g2_fill_2 FILLER_39_240 ();
 sg13g2_fill_2 FILLER_39_255 ();
 sg13g2_fill_1 FILLER_39_257 ();
 sg13g2_decap_4 FILLER_39_275 ();
 sg13g2_fill_1 FILLER_39_279 ();
 sg13g2_fill_1 FILLER_39_348 ();
 sg13g2_fill_2 FILLER_39_365 ();
 sg13g2_fill_2 FILLER_39_376 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_fill_2 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_fill_2 FILLER_40_64 ();
 sg13g2_fill_2 FILLER_40_71 ();
 sg13g2_fill_2 FILLER_40_90 ();
 sg13g2_fill_2 FILLER_40_97 ();
 sg13g2_decap_8 FILLER_40_108 ();
 sg13g2_fill_2 FILLER_40_115 ();
 sg13g2_fill_1 FILLER_40_117 ();
 sg13g2_decap_4 FILLER_40_123 ();
 sg13g2_fill_1 FILLER_40_127 ();
 sg13g2_decap_4 FILLER_40_138 ();
 sg13g2_fill_1 FILLER_40_142 ();
 sg13g2_decap_4 FILLER_40_155 ();
 sg13g2_fill_1 FILLER_40_159 ();
 sg13g2_fill_2 FILLER_40_168 ();
 sg13g2_fill_2 FILLER_40_242 ();
 sg13g2_fill_1 FILLER_40_244 ();
 sg13g2_fill_2 FILLER_40_250 ();
 sg13g2_fill_2 FILLER_40_266 ();
 sg13g2_fill_2 FILLER_40_349 ();
 sg13g2_fill_2 FILLER_40_357 ();
 sg13g2_fill_1 FILLER_40_359 ();
 sg13g2_fill_1 FILLER_40_363 ();
 sg13g2_fill_2 FILLER_40_374 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_75 ();
 sg13g2_fill_1 FILLER_41_85 ();
 sg13g2_fill_2 FILLER_41_117 ();
 sg13g2_fill_1 FILLER_41_133 ();
 sg13g2_fill_2 FILLER_41_154 ();
 sg13g2_decap_4 FILLER_41_198 ();
 sg13g2_fill_2 FILLER_41_251 ();
 sg13g2_decap_4 FILLER_41_261 ();
 sg13g2_fill_2 FILLER_41_281 ();
 sg13g2_fill_2 FILLER_41_303 ();
 sg13g2_fill_1 FILLER_41_305 ();
 sg13g2_decap_4 FILLER_41_311 ();
 sg13g2_fill_2 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_341 ();
 sg13g2_fill_2 FILLER_41_348 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_decap_4 FILLER_41_354 ();
 sg13g2_fill_1 FILLER_41_358 ();
 sg13g2_decap_4 FILLER_41_362 ();
 sg13g2_fill_1 FILLER_41_366 ();
 sg13g2_fill_2 FILLER_41_392 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_53 ();
 sg13g2_decap_8 FILLER_42_64 ();
 sg13g2_fill_1 FILLER_42_71 ();
 sg13g2_fill_1 FILLER_42_77 ();
 sg13g2_fill_2 FILLER_42_122 ();
 sg13g2_fill_1 FILLER_42_124 ();
 sg13g2_fill_2 FILLER_42_138 ();
 sg13g2_fill_1 FILLER_42_158 ();
 sg13g2_fill_2 FILLER_42_169 ();
 sg13g2_fill_1 FILLER_42_171 ();
 sg13g2_fill_1 FILLER_42_189 ();
 sg13g2_decap_4 FILLER_42_199 ();
 sg13g2_fill_2 FILLER_42_203 ();
 sg13g2_fill_2 FILLER_42_217 ();
 sg13g2_fill_1 FILLER_42_219 ();
 sg13g2_fill_1 FILLER_42_241 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_4 FILLER_42_281 ();
 sg13g2_decap_8 FILLER_42_290 ();
 sg13g2_fill_2 FILLER_42_309 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_fill_2 FILLER_42_318 ();
 sg13g2_fill_1 FILLER_42_320 ();
 sg13g2_fill_1 FILLER_42_331 ();
 sg13g2_decap_4 FILLER_42_337 ();
 sg13g2_decap_4 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_4 FILLER_43_56 ();
 sg13g2_decap_4 FILLER_43_73 ();
 sg13g2_fill_2 FILLER_43_81 ();
 sg13g2_fill_2 FILLER_43_96 ();
 sg13g2_fill_1 FILLER_43_103 ();
 sg13g2_decap_4 FILLER_43_117 ();
 sg13g2_fill_1 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_148 ();
 sg13g2_decap_4 FILLER_43_155 ();
 sg13g2_fill_2 FILLER_43_167 ();
 sg13g2_fill_2 FILLER_43_174 ();
 sg13g2_decap_8 FILLER_43_206 ();
 sg13g2_decap_4 FILLER_43_213 ();
 sg13g2_fill_2 FILLER_43_217 ();
 sg13g2_fill_2 FILLER_43_223 ();
 sg13g2_decap_4 FILLER_43_269 ();
 sg13g2_decap_8 FILLER_43_278 ();
 sg13g2_decap_8 FILLER_43_285 ();
 sg13g2_decap_4 FILLER_43_292 ();
 sg13g2_fill_1 FILLER_43_296 ();
 sg13g2_decap_8 FILLER_43_331 ();
 sg13g2_fill_1 FILLER_43_338 ();
 sg13g2_fill_2 FILLER_43_380 ();
 sg13g2_fill_1 FILLER_43_391 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_fill_2 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_44 ();
 sg13g2_fill_1 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_79 ();
 sg13g2_fill_2 FILLER_44_90 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_fill_2 FILLER_44_96 ();
 sg13g2_fill_1 FILLER_44_98 ();
 sg13g2_decap_4 FILLER_44_109 ();
 sg13g2_fill_1 FILLER_44_113 ();
 sg13g2_decap_4 FILLER_44_124 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_4 FILLER_44_149 ();
 sg13g2_fill_1 FILLER_44_158 ();
 sg13g2_fill_2 FILLER_44_180 ();
 sg13g2_fill_1 FILLER_44_182 ();
 sg13g2_fill_2 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_238 ();
 sg13g2_fill_1 FILLER_44_247 ();
 sg13g2_fill_1 FILLER_44_262 ();
 sg13g2_decap_8 FILLER_44_275 ();
 sg13g2_decap_8 FILLER_44_282 ();
 sg13g2_decap_4 FILLER_44_289 ();
 sg13g2_fill_2 FILLER_44_306 ();
 sg13g2_decap_8 FILLER_44_312 ();
 sg13g2_decap_8 FILLER_44_319 ();
 sg13g2_fill_2 FILLER_44_336 ();
 sg13g2_fill_1 FILLER_44_354 ();
 sg13g2_fill_1 FILLER_44_396 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_4 FILLER_45_28 ();
 sg13g2_fill_2 FILLER_45_32 ();
 sg13g2_decap_4 FILLER_45_105 ();
 sg13g2_fill_1 FILLER_45_114 ();
 sg13g2_decap_8 FILLER_45_125 ();
 sg13g2_fill_2 FILLER_45_132 ();
 sg13g2_decap_8 FILLER_45_142 ();
 sg13g2_fill_2 FILLER_45_176 ();
 sg13g2_fill_1 FILLER_45_178 ();
 sg13g2_fill_2 FILLER_45_185 ();
 sg13g2_fill_1 FILLER_45_187 ();
 sg13g2_fill_2 FILLER_45_201 ();
 sg13g2_fill_1 FILLER_45_203 ();
 sg13g2_decap_4 FILLER_45_254 ();
 sg13g2_fill_1 FILLER_45_286 ();
 sg13g2_decap_8 FILLER_45_302 ();
 sg13g2_decap_8 FILLER_45_309 ();
 sg13g2_fill_1 FILLER_45_316 ();
 sg13g2_fill_2 FILLER_45_340 ();
 sg13g2_fill_1 FILLER_45_342 ();
 sg13g2_fill_2 FILLER_45_348 ();
 sg13g2_fill_2 FILLER_45_355 ();
 sg13g2_fill_1 FILLER_45_375 ();
 sg13g2_fill_1 FILLER_45_386 ();
 sg13g2_fill_2 FILLER_45_395 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_35 ();
 sg13g2_fill_2 FILLER_46_64 ();
 sg13g2_fill_1 FILLER_46_66 ();
 sg13g2_fill_2 FILLER_46_81 ();
 sg13g2_fill_1 FILLER_46_83 ();
 sg13g2_fill_2 FILLER_46_128 ();
 sg13g2_fill_1 FILLER_46_130 ();
 sg13g2_decap_4 FILLER_46_163 ();
 sg13g2_fill_2 FILLER_46_184 ();
 sg13g2_fill_1 FILLER_46_186 ();
 sg13g2_fill_2 FILLER_46_208 ();
 sg13g2_decap_4 FILLER_46_245 ();
 sg13g2_fill_2 FILLER_46_249 ();
 sg13g2_decap_4 FILLER_46_256 ();
 sg13g2_fill_2 FILLER_46_268 ();
 sg13g2_fill_1 FILLER_46_275 ();
 sg13g2_fill_2 FILLER_46_334 ();
 sg13g2_fill_1 FILLER_46_336 ();
 sg13g2_fill_2 FILLER_46_345 ();
 sg13g2_decap_8 FILLER_46_352 ();
 sg13g2_fill_1 FILLER_46_359 ();
 sg13g2_decap_4 FILLER_46_374 ();
 sg13g2_fill_2 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_fill_2 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_70 ();
 sg13g2_fill_2 FILLER_47_77 ();
 sg13g2_fill_2 FILLER_47_89 ();
 sg13g2_fill_2 FILLER_47_96 ();
 sg13g2_fill_1 FILLER_47_98 ();
 sg13g2_fill_2 FILLER_47_125 ();
 sg13g2_fill_2 FILLER_47_137 ();
 sg13g2_fill_1 FILLER_47_139 ();
 sg13g2_decap_8 FILLER_47_164 ();
 sg13g2_fill_2 FILLER_47_175 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_fill_1 FILLER_47_210 ();
 sg13g2_decap_4 FILLER_47_245 ();
 sg13g2_fill_2 FILLER_47_257 ();
 sg13g2_decap_4 FILLER_47_311 ();
 sg13g2_fill_2 FILLER_47_315 ();
 sg13g2_fill_2 FILLER_47_340 ();
 sg13g2_fill_1 FILLER_47_342 ();
 sg13g2_decap_8 FILLER_47_352 ();
 sg13g2_decap_8 FILLER_47_359 ();
 sg13g2_decap_4 FILLER_47_405 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_60 ();
 sg13g2_fill_2 FILLER_48_70 ();
 sg13g2_fill_1 FILLER_48_72 ();
 sg13g2_fill_2 FILLER_48_85 ();
 sg13g2_fill_1 FILLER_48_92 ();
 sg13g2_decap_4 FILLER_48_97 ();
 sg13g2_fill_1 FILLER_48_101 ();
 sg13g2_decap_4 FILLER_48_107 ();
 sg13g2_fill_1 FILLER_48_111 ();
 sg13g2_fill_1 FILLER_48_117 ();
 sg13g2_decap_8 FILLER_48_136 ();
 sg13g2_fill_2 FILLER_48_148 ();
 sg13g2_decap_8 FILLER_48_155 ();
 sg13g2_fill_2 FILLER_48_162 ();
 sg13g2_fill_1 FILLER_48_164 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_fill_2 FILLER_48_198 ();
 sg13g2_fill_1 FILLER_48_206 ();
 sg13g2_fill_2 FILLER_48_217 ();
 sg13g2_fill_2 FILLER_48_228 ();
 sg13g2_decap_4 FILLER_48_290 ();
 sg13g2_fill_1 FILLER_48_320 ();
 sg13g2_fill_1 FILLER_48_381 ();
 sg13g2_decap_4 FILLER_48_391 ();
 sg13g2_decap_4 FILLER_48_405 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_4 FILLER_49_49 ();
 sg13g2_fill_1 FILLER_49_99 ();
 sg13g2_decap_4 FILLER_49_110 ();
 sg13g2_decap_8 FILLER_49_128 ();
 sg13g2_fill_2 FILLER_49_135 ();
 sg13g2_decap_4 FILLER_49_142 ();
 sg13g2_fill_1 FILLER_49_146 ();
 sg13g2_decap_4 FILLER_49_152 ();
 sg13g2_fill_2 FILLER_49_156 ();
 sg13g2_decap_4 FILLER_49_180 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_fill_2 FILLER_49_254 ();
 sg13g2_fill_1 FILLER_49_299 ();
 sg13g2_decap_4 FILLER_49_340 ();
 sg13g2_fill_2 FILLER_49_344 ();
 sg13g2_decap_8 FILLER_49_352 ();
 sg13g2_fill_2 FILLER_49_359 ();
 sg13g2_fill_1 FILLER_49_361 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_fill_2 FILLER_50_42 ();
 sg13g2_fill_1 FILLER_50_44 ();
 sg13g2_fill_2 FILLER_50_92 ();
 sg13g2_fill_1 FILLER_50_94 ();
 sg13g2_decap_4 FILLER_50_125 ();
 sg13g2_fill_2 FILLER_50_170 ();
 sg13g2_fill_2 FILLER_50_186 ();
 sg13g2_fill_2 FILLER_50_202 ();
 sg13g2_fill_2 FILLER_50_237 ();
 sg13g2_fill_1 FILLER_50_239 ();
 sg13g2_fill_2 FILLER_50_244 ();
 sg13g2_fill_2 FILLER_50_255 ();
 sg13g2_fill_1 FILLER_50_276 ();
 sg13g2_fill_1 FILLER_50_282 ();
 sg13g2_fill_1 FILLER_50_288 ();
 sg13g2_fill_2 FILLER_50_303 ();
 sg13g2_fill_1 FILLER_50_305 ();
 sg13g2_fill_2 FILLER_50_320 ();
 sg13g2_fill_2 FILLER_50_379 ();
 sg13g2_fill_1 FILLER_50_381 ();
 sg13g2_decap_4 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_fill_2 FILLER_51_42 ();
 sg13g2_fill_1 FILLER_51_44 ();
 sg13g2_fill_2 FILLER_51_71 ();
 sg13g2_fill_1 FILLER_51_73 ();
 sg13g2_fill_2 FILLER_51_87 ();
 sg13g2_fill_1 FILLER_51_89 ();
 sg13g2_fill_1 FILLER_51_114 ();
 sg13g2_decap_4 FILLER_51_148 ();
 sg13g2_fill_1 FILLER_51_166 ();
 sg13g2_fill_2 FILLER_51_171 ();
 sg13g2_decap_8 FILLER_51_177 ();
 sg13g2_fill_1 FILLER_51_218 ();
 sg13g2_fill_1 FILLER_51_232 ();
 sg13g2_fill_2 FILLER_51_253 ();
 sg13g2_fill_1 FILLER_51_261 ();
 sg13g2_fill_2 FILLER_51_270 ();
 sg13g2_fill_2 FILLER_51_315 ();
 sg13g2_fill_2 FILLER_51_325 ();
 sg13g2_fill_1 FILLER_51_327 ();
 sg13g2_decap_4 FILLER_51_333 ();
 sg13g2_fill_2 FILLER_51_337 ();
 sg13g2_fill_1 FILLER_51_349 ();
 sg13g2_fill_1 FILLER_51_369 ();
 sg13g2_decap_4 FILLER_51_405 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_fill_2 FILLER_52_42 ();
 sg13g2_fill_1 FILLER_52_70 ();
 sg13g2_fill_2 FILLER_52_79 ();
 sg13g2_fill_1 FILLER_52_81 ();
 sg13g2_fill_2 FILLER_52_92 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_fill_2 FILLER_52_143 ();
 sg13g2_fill_1 FILLER_52_145 ();
 sg13g2_decap_8 FILLER_52_163 ();
 sg13g2_decap_8 FILLER_52_170 ();
 sg13g2_decap_4 FILLER_52_182 ();
 sg13g2_fill_2 FILLER_52_194 ();
 sg13g2_decap_4 FILLER_52_319 ();
 sg13g2_fill_1 FILLER_52_323 ();
 sg13g2_decap_8 FILLER_52_333 ();
 sg13g2_fill_2 FILLER_52_340 ();
 sg13g2_fill_1 FILLER_52_342 ();
 sg13g2_fill_1 FILLER_52_357 ();
 sg13g2_fill_2 FILLER_52_372 ();
 sg13g2_fill_1 FILLER_52_374 ();
 sg13g2_fill_1 FILLER_52_379 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_fill_2 FILLER_53_42 ();
 sg13g2_fill_2 FILLER_53_71 ();
 sg13g2_fill_2 FILLER_53_81 ();
 sg13g2_fill_2 FILLER_53_97 ();
 sg13g2_fill_1 FILLER_53_99 ();
 sg13g2_fill_1 FILLER_53_136 ();
 sg13g2_fill_2 FILLER_53_168 ();
 sg13g2_decap_4 FILLER_53_190 ();
 sg13g2_fill_1 FILLER_53_211 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_fill_1 FILLER_53_255 ();
 sg13g2_decap_4 FILLER_53_311 ();
 sg13g2_fill_2 FILLER_53_319 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_decap_4 FILLER_53_346 ();
 sg13g2_fill_2 FILLER_53_368 ();
 sg13g2_decap_4 FILLER_53_375 ();
 sg13g2_fill_2 FILLER_53_379 ();
 sg13g2_decap_4 FILLER_53_386 ();
 sg13g2_fill_2 FILLER_53_390 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_4 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_39 ();
 sg13g2_fill_2 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_fill_2 FILLER_54_100 ();
 sg13g2_fill_1 FILLER_54_102 ();
 sg13g2_fill_2 FILLER_54_115 ();
 sg13g2_fill_1 FILLER_54_117 ();
 sg13g2_decap_4 FILLER_54_122 ();
 sg13g2_fill_2 FILLER_54_126 ();
 sg13g2_fill_1 FILLER_54_136 ();
 sg13g2_fill_2 FILLER_54_150 ();
 sg13g2_fill_2 FILLER_54_158 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_fill_1 FILLER_54_174 ();
 sg13g2_decap_4 FILLER_54_234 ();
 sg13g2_fill_2 FILLER_54_249 ();
 sg13g2_fill_1 FILLER_54_255 ();
 sg13g2_fill_2 FILLER_54_261 ();
 sg13g2_fill_1 FILLER_54_263 ();
 sg13g2_fill_1 FILLER_54_279 ();
 sg13g2_decap_8 FILLER_54_292 ();
 sg13g2_decap_8 FILLER_54_299 ();
 sg13g2_fill_2 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_377 ();
 sg13g2_fill_2 FILLER_54_389 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_4 FILLER_55_42 ();
 sg13g2_fill_1 FILLER_55_46 ();
 sg13g2_fill_1 FILLER_55_89 ();
 sg13g2_fill_2 FILLER_55_108 ();
 sg13g2_fill_1 FILLER_55_110 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_4 FILLER_55_126 ();
 sg13g2_fill_2 FILLER_55_142 ();
 sg13g2_decap_4 FILLER_55_169 ();
 sg13g2_fill_2 FILLER_55_173 ();
 sg13g2_fill_1 FILLER_55_189 ();
 sg13g2_decap_4 FILLER_55_194 ();
 sg13g2_fill_1 FILLER_55_220 ();
 sg13g2_fill_2 FILLER_55_226 ();
 sg13g2_fill_1 FILLER_55_228 ();
 sg13g2_decap_4 FILLER_55_240 ();
 sg13g2_fill_2 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_289 ();
 sg13g2_decap_8 FILLER_55_300 ();
 sg13g2_decap_4 FILLER_55_307 ();
 sg13g2_fill_1 FILLER_55_311 ();
 sg13g2_fill_1 FILLER_55_320 ();
 sg13g2_fill_2 FILLER_55_340 ();
 sg13g2_decap_4 FILLER_55_355 ();
 sg13g2_fill_1 FILLER_55_359 ();
 sg13g2_decap_8 FILLER_55_365 ();
 sg13g2_decap_4 FILLER_55_372 ();
 sg13g2_fill_1 FILLER_55_376 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_fill_2 FILLER_56_49 ();
 sg13g2_fill_2 FILLER_56_55 ();
 sg13g2_fill_1 FILLER_56_57 ();
 sg13g2_fill_2 FILLER_56_80 ();
 sg13g2_fill_1 FILLER_56_87 ();
 sg13g2_fill_1 FILLER_56_93 ();
 sg13g2_fill_2 FILLER_56_106 ();
 sg13g2_fill_1 FILLER_56_108 ();
 sg13g2_fill_2 FILLER_56_143 ();
 sg13g2_fill_1 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_150 ();
 sg13g2_fill_2 FILLER_56_157 ();
 sg13g2_fill_1 FILLER_56_171 ();
 sg13g2_decap_4 FILLER_56_177 ();
 sg13g2_decap_4 FILLER_56_201 ();
 sg13g2_fill_2 FILLER_56_217 ();
 sg13g2_fill_1 FILLER_56_219 ();
 sg13g2_decap_4 FILLER_56_234 ();
 sg13g2_fill_2 FILLER_56_243 ();
 sg13g2_fill_1 FILLER_56_249 ();
 sg13g2_fill_1 FILLER_56_314 ();
 sg13g2_decap_4 FILLER_56_321 ();
 sg13g2_fill_1 FILLER_56_325 ();
 sg13g2_fill_2 FILLER_56_357 ();
 sg13g2_fill_1 FILLER_56_359 ();
 sg13g2_fill_1 FILLER_56_365 ();
 sg13g2_fill_2 FILLER_56_381 ();
 sg13g2_fill_1 FILLER_56_383 ();
 sg13g2_fill_2 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_4 FILLER_57_49 ();
 sg13g2_fill_2 FILLER_57_64 ();
 sg13g2_decap_4 FILLER_57_70 ();
 sg13g2_fill_1 FILLER_57_74 ();
 sg13g2_decap_8 FILLER_57_82 ();
 sg13g2_fill_1 FILLER_57_146 ();
 sg13g2_fill_2 FILLER_57_162 ();
 sg13g2_fill_1 FILLER_57_164 ();
 sg13g2_decap_4 FILLER_57_174 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_4 FILLER_57_217 ();
 sg13g2_fill_1 FILLER_57_221 ();
 sg13g2_decap_8 FILLER_57_234 ();
 sg13g2_decap_4 FILLER_57_241 ();
 sg13g2_fill_1 FILLER_57_245 ();
 sg13g2_fill_2 FILLER_57_254 ();
 sg13g2_fill_1 FILLER_57_282 ();
 sg13g2_fill_1 FILLER_57_314 ();
 sg13g2_fill_2 FILLER_57_350 ();
 sg13g2_fill_1 FILLER_57_352 ();
 sg13g2_fill_2 FILLER_57_365 ();
 sg13g2_fill_1 FILLER_57_367 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_fill_2 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_82 ();
 sg13g2_fill_2 FILLER_58_89 ();
 sg13g2_fill_1 FILLER_58_91 ();
 sg13g2_fill_2 FILLER_58_102 ();
 sg13g2_fill_1 FILLER_58_114 ();
 sg13g2_fill_2 FILLER_58_129 ();
 sg13g2_fill_1 FILLER_58_131 ();
 sg13g2_fill_1 FILLER_58_151 ();
 sg13g2_fill_1 FILLER_58_158 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_fill_1 FILLER_58_210 ();
 sg13g2_fill_1 FILLER_58_223 ();
 sg13g2_fill_1 FILLER_58_266 ();
 sg13g2_fill_2 FILLER_58_285 ();
 sg13g2_fill_1 FILLER_58_328 ();
 sg13g2_decap_4 FILLER_58_339 ();
 sg13g2_fill_2 FILLER_58_343 ();
 sg13g2_decap_4 FILLER_58_355 ();
 sg13g2_fill_1 FILLER_58_369 ();
 sg13g2_fill_1 FILLER_58_380 ();
 sg13g2_fill_2 FILLER_58_391 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_4 FILLER_59_28 ();
 sg13g2_fill_1 FILLER_59_63 ();
 sg13g2_fill_2 FILLER_59_90 ();
 sg13g2_fill_2 FILLER_59_113 ();
 sg13g2_fill_1 FILLER_59_115 ();
 sg13g2_fill_2 FILLER_59_151 ();
 sg13g2_decap_4 FILLER_59_195 ();
 sg13g2_fill_2 FILLER_59_264 ();
 sg13g2_decap_8 FILLER_59_270 ();
 sg13g2_decap_8 FILLER_59_277 ();
 sg13g2_decap_8 FILLER_59_284 ();
 sg13g2_fill_2 FILLER_59_291 ();
 sg13g2_fill_1 FILLER_59_293 ();
 sg13g2_fill_2 FILLER_59_298 ();
 sg13g2_decap_8 FILLER_59_343 ();
 sg13g2_decap_4 FILLER_59_350 ();
 sg13g2_fill_1 FILLER_59_354 ();
 sg13g2_fill_2 FILLER_59_360 ();
 sg13g2_decap_8 FILLER_59_367 ();
 sg13g2_fill_2 FILLER_59_374 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_4 FILLER_60_110 ();
 sg13g2_fill_2 FILLER_60_128 ();
 sg13g2_decap_8 FILLER_60_134 ();
 sg13g2_fill_2 FILLER_60_141 ();
 sg13g2_fill_1 FILLER_60_161 ();
 sg13g2_fill_2 FILLER_60_173 ();
 sg13g2_fill_1 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_187 ();
 sg13g2_fill_1 FILLER_60_194 ();
 sg13g2_decap_4 FILLER_60_211 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_fill_1 FILLER_60_243 ();
 sg13g2_fill_1 FILLER_60_252 ();
 sg13g2_fill_1 FILLER_60_262 ();
 sg13g2_decap_8 FILLER_60_269 ();
 sg13g2_decap_8 FILLER_60_276 ();
 sg13g2_fill_2 FILLER_60_283 ();
 sg13g2_fill_1 FILLER_60_285 ();
 sg13g2_decap_8 FILLER_60_291 ();
 sg13g2_fill_1 FILLER_60_305 ();
 sg13g2_fill_2 FILLER_60_316 ();
 sg13g2_fill_1 FILLER_60_318 ();
 sg13g2_fill_1 FILLER_60_323 ();
 sg13g2_fill_1 FILLER_60_339 ();
 sg13g2_decap_8 FILLER_60_345 ();
 sg13g2_fill_2 FILLER_60_352 ();
 sg13g2_fill_2 FILLER_60_359 ();
 sg13g2_fill_1 FILLER_60_361 ();
 sg13g2_decap_4 FILLER_60_368 ();
 sg13g2_fill_1 FILLER_60_372 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_2 FILLER_60_395 ();
 sg13g2_fill_1 FILLER_60_397 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_4 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_39 ();
 sg13g2_fill_1 FILLER_61_77 ();
 sg13g2_fill_2 FILLER_61_91 ();
 sg13g2_fill_1 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_138 ();
 sg13g2_fill_1 FILLER_61_149 ();
 sg13g2_fill_2 FILLER_61_160 ();
 sg13g2_fill_1 FILLER_61_162 ();
 sg13g2_fill_2 FILLER_61_173 ();
 sg13g2_fill_2 FILLER_61_181 ();
 sg13g2_decap_4 FILLER_61_188 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_217 ();
 sg13g2_decap_8 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_231 ();
 sg13g2_fill_2 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_240 ();
 sg13g2_fill_2 FILLER_61_246 ();
 sg13g2_fill_1 FILLER_61_248 ();
 sg13g2_fill_1 FILLER_61_260 ();
 sg13g2_decap_8 FILLER_61_299 ();
 sg13g2_decap_4 FILLER_61_306 ();
 sg13g2_fill_2 FILLER_61_333 ();
 sg13g2_fill_2 FILLER_61_367 ();
 sg13g2_fill_1 FILLER_61_369 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_fill_1 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_70 ();
 sg13g2_fill_2 FILLER_62_171 ();
 sg13g2_fill_1 FILLER_62_265 ();
 sg13g2_fill_1 FILLER_62_311 ();
 sg13g2_fill_2 FILLER_62_326 ();
 sg13g2_fill_1 FILLER_62_349 ();
 sg13g2_fill_1 FILLER_62_358 ();
 sg13g2_fill_2 FILLER_62_370 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_2 FILLER_62_388 ();
 sg13g2_fill_1 FILLER_62_390 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_4 FILLER_63_28 ();
 sg13g2_fill_1 FILLER_63_85 ();
 sg13g2_fill_1 FILLER_63_94 ();
 sg13g2_fill_2 FILLER_63_100 ();
 sg13g2_fill_1 FILLER_63_102 ();
 sg13g2_fill_2 FILLER_63_131 ();
 sg13g2_fill_1 FILLER_63_133 ();
 sg13g2_fill_2 FILLER_63_139 ();
 sg13g2_fill_2 FILLER_63_166 ();
 sg13g2_fill_1 FILLER_63_168 ();
 sg13g2_fill_2 FILLER_63_174 ();
 sg13g2_decap_4 FILLER_63_186 ();
 sg13g2_fill_1 FILLER_63_210 ();
 sg13g2_fill_2 FILLER_63_264 ();
 sg13g2_decap_4 FILLER_63_271 ();
 sg13g2_fill_2 FILLER_63_275 ();
 sg13g2_decap_4 FILLER_63_282 ();
 sg13g2_fill_1 FILLER_63_301 ();
 sg13g2_fill_2 FILLER_63_306 ();
 sg13g2_decap_8 FILLER_63_314 ();
 sg13g2_fill_1 FILLER_63_321 ();
 sg13g2_fill_2 FILLER_63_357 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_80 ();
 sg13g2_fill_2 FILLER_64_87 ();
 sg13g2_fill_2 FILLER_64_97 ();
 sg13g2_fill_2 FILLER_64_112 ();
 sg13g2_fill_2 FILLER_64_125 ();
 sg13g2_fill_1 FILLER_64_136 ();
 sg13g2_decap_4 FILLER_64_142 ();
 sg13g2_decap_8 FILLER_64_166 ();
 sg13g2_decap_8 FILLER_64_173 ();
 sg13g2_decap_8 FILLER_64_180 ();
 sg13g2_decap_8 FILLER_64_187 ();
 sg13g2_decap_8 FILLER_64_194 ();
 sg13g2_decap_4 FILLER_64_201 ();
 sg13g2_fill_1 FILLER_64_205 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_decap_4 FILLER_64_217 ();
 sg13g2_fill_1 FILLER_64_221 ();
 sg13g2_fill_1 FILLER_64_236 ();
 sg13g2_decap_8 FILLER_64_256 ();
 sg13g2_decap_8 FILLER_64_263 ();
 sg13g2_decap_4 FILLER_64_270 ();
 sg13g2_fill_1 FILLER_64_274 ();
 sg13g2_fill_1 FILLER_64_280 ();
 sg13g2_fill_2 FILLER_64_289 ();
 sg13g2_decap_8 FILLER_64_325 ();
 sg13g2_fill_2 FILLER_64_332 ();
 sg13g2_fill_1 FILLER_64_360 ();
 sg13g2_fill_2 FILLER_64_374 ();
 sg13g2_fill_1 FILLER_64_381 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_fill_2 FILLER_65_28 ();
 sg13g2_decap_4 FILLER_65_74 ();
 sg13g2_fill_1 FILLER_65_91 ();
 sg13g2_fill_2 FILLER_65_135 ();
 sg13g2_fill_1 FILLER_65_137 ();
 sg13g2_fill_2 FILLER_65_144 ();
 sg13g2_fill_1 FILLER_65_152 ();
 sg13g2_fill_2 FILLER_65_158 ();
 sg13g2_fill_2 FILLER_65_179 ();
 sg13g2_fill_2 FILLER_65_193 ();
 sg13g2_fill_1 FILLER_65_195 ();
 sg13g2_decap_4 FILLER_65_200 ();
 sg13g2_fill_1 FILLER_65_204 ();
 sg13g2_fill_1 FILLER_65_215 ();
 sg13g2_decap_8 FILLER_65_222 ();
 sg13g2_decap_4 FILLER_65_229 ();
 sg13g2_fill_1 FILLER_65_233 ();
 sg13g2_decap_8 FILLER_65_243 ();
 sg13g2_decap_4 FILLER_65_250 ();
 sg13g2_fill_1 FILLER_65_257 ();
 sg13g2_decap_4 FILLER_65_262 ();
 sg13g2_fill_2 FILLER_65_266 ();
 sg13g2_decap_8 FILLER_65_294 ();
 sg13g2_decap_4 FILLER_65_301 ();
 sg13g2_fill_1 FILLER_65_305 ();
 sg13g2_fill_1 FILLER_65_309 ();
 sg13g2_decap_8 FILLER_65_326 ();
 sg13g2_decap_4 FILLER_65_333 ();
 sg13g2_fill_1 FILLER_65_337 ();
 sg13g2_fill_1 FILLER_65_351 ();
 sg13g2_fill_1 FILLER_65_390 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_4 FILLER_66_21 ();
 sg13g2_fill_2 FILLER_66_25 ();
 sg13g2_fill_1 FILLER_66_94 ();
 sg13g2_fill_2 FILLER_66_101 ();
 sg13g2_fill_2 FILLER_66_111 ();
 sg13g2_fill_1 FILLER_66_113 ();
 sg13g2_fill_2 FILLER_66_134 ();
 sg13g2_fill_2 FILLER_66_157 ();
 sg13g2_fill_1 FILLER_66_159 ();
 sg13g2_fill_2 FILLER_66_193 ();
 sg13g2_fill_1 FILLER_66_195 ();
 sg13g2_fill_2 FILLER_66_216 ();
 sg13g2_decap_4 FILLER_66_224 ();
 sg13g2_fill_1 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_257 ();
 sg13g2_fill_2 FILLER_66_267 ();
 sg13g2_fill_2 FILLER_66_302 ();
 sg13g2_fill_1 FILLER_66_304 ();
 sg13g2_decap_4 FILLER_66_316 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_fill_2 FILLER_66_343 ();
 sg13g2_fill_2 FILLER_66_357 ();
 sg13g2_fill_2 FILLER_66_367 ();
 sg13g2_fill_1 FILLER_66_369 ();
 sg13g2_fill_1 FILLER_66_380 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_4 FILLER_67_35 ();
 sg13g2_fill_2 FILLER_67_87 ();
 sg13g2_fill_1 FILLER_67_102 ();
 sg13g2_fill_2 FILLER_67_109 ();
 sg13g2_fill_1 FILLER_67_111 ();
 sg13g2_fill_1 FILLER_67_118 ();
 sg13g2_fill_1 FILLER_67_129 ();
 sg13g2_fill_2 FILLER_67_135 ();
 sg13g2_fill_2 FILLER_67_142 ();
 sg13g2_fill_1 FILLER_67_166 ();
 sg13g2_fill_2 FILLER_67_202 ();
 sg13g2_fill_1 FILLER_67_204 ();
 sg13g2_decap_4 FILLER_67_219 ();
 sg13g2_fill_1 FILLER_67_254 ();
 sg13g2_fill_2 FILLER_67_281 ();
 sg13g2_fill_1 FILLER_67_283 ();
 sg13g2_fill_1 FILLER_67_292 ();
 sg13g2_fill_2 FILLER_67_319 ();
 sg13g2_fill_1 FILLER_67_321 ();
 sg13g2_fill_2 FILLER_67_328 ();
 sg13g2_decap_8 FILLER_67_370 ();
 sg13g2_decap_4 FILLER_67_377 ();
 sg13g2_fill_2 FILLER_67_381 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_fill_2 FILLER_68_49 ();
 sg13g2_fill_2 FILLER_68_62 ();
 sg13g2_fill_1 FILLER_68_64 ();
 sg13g2_fill_2 FILLER_68_74 ();
 sg13g2_fill_1 FILLER_68_89 ();
 sg13g2_fill_2 FILLER_68_124 ();
 sg13g2_fill_1 FILLER_68_126 ();
 sg13g2_fill_1 FILLER_68_146 ();
 sg13g2_fill_2 FILLER_68_176 ();
 sg13g2_fill_1 FILLER_68_184 ();
 sg13g2_fill_2 FILLER_68_191 ();
 sg13g2_decap_8 FILLER_68_215 ();
 sg13g2_fill_2 FILLER_68_222 ();
 sg13g2_fill_1 FILLER_68_239 ();
 sg13g2_fill_1 FILLER_68_256 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_2 FILLER_68_273 ();
 sg13g2_fill_1 FILLER_68_275 ();
 sg13g2_fill_1 FILLER_68_298 ();
 sg13g2_fill_1 FILLER_68_331 ();
 sg13g2_fill_2 FILLER_68_337 ();
 sg13g2_decap_4 FILLER_68_366 ();
 sg13g2_fill_2 FILLER_68_375 ();
 sg13g2_decap_4 FILLER_68_382 ();
 sg13g2_fill_2 FILLER_68_386 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_fill_1 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_75 ();
 sg13g2_decap_8 FILLER_69_82 ();
 sg13g2_decap_4 FILLER_69_89 ();
 sg13g2_fill_2 FILLER_69_93 ();
 sg13g2_fill_2 FILLER_69_140 ();
 sg13g2_fill_1 FILLER_69_178 ();
 sg13g2_fill_1 FILLER_69_197 ();
 sg13g2_decap_4 FILLER_69_219 ();
 sg13g2_fill_1 FILLER_69_242 ();
 sg13g2_fill_2 FILLER_69_248 ();
 sg13g2_decap_8 FILLER_69_253 ();
 sg13g2_fill_2 FILLER_69_260 ();
 sg13g2_fill_2 FILLER_69_265 ();
 sg13g2_fill_2 FILLER_69_276 ();
 sg13g2_fill_1 FILLER_69_299 ();
 sg13g2_fill_2 FILLER_69_357 ();
 sg13g2_fill_1 FILLER_69_359 ();
 sg13g2_fill_1 FILLER_69_365 ();
 sg13g2_fill_1 FILLER_69_379 ();
 sg13g2_fill_1 FILLER_69_393 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_fill_2 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_86 ();
 sg13g2_fill_1 FILLER_70_113 ();
 sg13g2_fill_1 FILLER_70_162 ();
 sg13g2_fill_2 FILLER_70_168 ();
 sg13g2_fill_1 FILLER_70_170 ();
 sg13g2_fill_2 FILLER_70_215 ();
 sg13g2_fill_1 FILLER_70_217 ();
 sg13g2_fill_1 FILLER_70_291 ();
 sg13g2_fill_2 FILLER_70_324 ();
 sg13g2_fill_1 FILLER_70_326 ();
 sg13g2_fill_2 FILLER_70_332 ();
 sg13g2_fill_1 FILLER_70_334 ();
 sg13g2_fill_2 FILLER_70_353 ();
 sg13g2_fill_1 FILLER_70_355 ();
 sg13g2_fill_2 FILLER_70_383 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_fill_2 FILLER_71_102 ();
 sg13g2_decap_4 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_128 ();
 sg13g2_fill_1 FILLER_71_135 ();
 sg13g2_fill_2 FILLER_71_144 ();
 sg13g2_fill_1 FILLER_71_146 ();
 sg13g2_decap_8 FILLER_71_156 ();
 sg13g2_fill_2 FILLER_71_172 ();
 sg13g2_fill_2 FILLER_71_183 ();
 sg13g2_fill_1 FILLER_71_185 ();
 sg13g2_fill_2 FILLER_71_202 ();
 sg13g2_fill_1 FILLER_71_254 ();
 sg13g2_fill_2 FILLER_71_269 ();
 sg13g2_decap_4 FILLER_71_342 ();
 sg13g2_fill_2 FILLER_71_367 ();
 sg13g2_fill_2 FILLER_71_381 ();
 sg13g2_fill_1 FILLER_71_383 ();
 sg13g2_fill_2 FILLER_71_406 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_fill_2 FILLER_72_112 ();
 sg13g2_fill_1 FILLER_72_114 ();
 sg13g2_fill_1 FILLER_72_123 ();
 sg13g2_decap_8 FILLER_72_129 ();
 sg13g2_fill_2 FILLER_72_142 ();
 sg13g2_decap_4 FILLER_72_149 ();
 sg13g2_decap_8 FILLER_72_162 ();
 sg13g2_decap_4 FILLER_72_169 ();
 sg13g2_fill_2 FILLER_72_173 ();
 sg13g2_fill_2 FILLER_72_183 ();
 sg13g2_fill_1 FILLER_72_185 ();
 sg13g2_fill_2 FILLER_72_197 ();
 sg13g2_fill_1 FILLER_72_199 ();
 sg13g2_decap_8 FILLER_72_212 ();
 sg13g2_fill_2 FILLER_72_219 ();
 sg13g2_fill_2 FILLER_72_247 ();
 sg13g2_fill_2 FILLER_72_275 ();
 sg13g2_fill_1 FILLER_72_277 ();
 sg13g2_fill_1 FILLER_72_336 ();
 sg13g2_fill_2 FILLER_72_342 ();
 sg13g2_fill_1 FILLER_72_352 ();
 sg13g2_decap_4 FILLER_72_400 ();
 sg13g2_fill_1 FILLER_72_404 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_fill_1 FILLER_73_119 ();
 sg13g2_fill_2 FILLER_73_135 ();
 sg13g2_fill_1 FILLER_73_137 ();
 sg13g2_fill_1 FILLER_73_147 ();
 sg13g2_fill_2 FILLER_73_152 ();
 sg13g2_decap_8 FILLER_73_162 ();
 sg13g2_decap_8 FILLER_73_169 ();
 sg13g2_decap_8 FILLER_73_176 ();
 sg13g2_decap_8 FILLER_73_183 ();
 sg13g2_decap_4 FILLER_73_190 ();
 sg13g2_fill_1 FILLER_73_194 ();
 sg13g2_fill_2 FILLER_73_229 ();
 sg13g2_fill_2 FILLER_73_235 ();
 sg13g2_fill_1 FILLER_73_237 ();
 sg13g2_fill_2 FILLER_73_331 ();
 sg13g2_fill_1 FILLER_73_333 ();
 sg13g2_fill_2 FILLER_73_338 ();
 sg13g2_fill_1 FILLER_73_340 ();
 sg13g2_fill_2 FILLER_73_346 ();
 sg13g2_fill_1 FILLER_73_360 ();
 sg13g2_fill_2 FILLER_73_388 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_fill_2 FILLER_74_105 ();
 sg13g2_fill_2 FILLER_74_143 ();
 sg13g2_fill_2 FILLER_74_156 ();
 sg13g2_fill_1 FILLER_74_158 ();
 sg13g2_decap_4 FILLER_74_171 ();
 sg13g2_decap_8 FILLER_74_185 ();
 sg13g2_decap_4 FILLER_74_192 ();
 sg13g2_decap_8 FILLER_74_199 ();
 sg13g2_fill_2 FILLER_74_206 ();
 sg13g2_fill_1 FILLER_74_216 ();
 sg13g2_fill_2 FILLER_74_222 ();
 sg13g2_fill_2 FILLER_74_233 ();
 sg13g2_fill_1 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_306 ();
 sg13g2_fill_2 FILLER_74_312 ();
 sg13g2_fill_1 FILLER_74_314 ();
 sg13g2_fill_1 FILLER_74_320 ();
 sg13g2_fill_2 FILLER_74_362 ();
 sg13g2_fill_1 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_fill_2 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_73 ();
 sg13g2_decap_8 FILLER_75_80 ();
 sg13g2_decap_8 FILLER_75_87 ();
 sg13g2_decap_8 FILLER_75_94 ();
 sg13g2_decap_4 FILLER_75_101 ();
 sg13g2_fill_1 FILLER_75_153 ();
 sg13g2_fill_2 FILLER_75_160 ();
 sg13g2_fill_1 FILLER_75_168 ();
 sg13g2_decap_4 FILLER_75_188 ();
 sg13g2_fill_2 FILLER_75_216 ();
 sg13g2_fill_1 FILLER_75_218 ();
 sg13g2_fill_1 FILLER_75_224 ();
 sg13g2_fill_1 FILLER_75_243 ();
 sg13g2_fill_2 FILLER_75_268 ();
 sg13g2_fill_1 FILLER_75_270 ();
 sg13g2_fill_2 FILLER_75_280 ();
 sg13g2_fill_2 FILLER_75_308 ();
 sg13g2_fill_1 FILLER_75_315 ();
 sg13g2_fill_2 FILLER_75_342 ();
 sg13g2_fill_1 FILLER_75_344 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_fill_2 FILLER_76_98 ();
 sg13g2_fill_1 FILLER_76_100 ();
 sg13g2_fill_2 FILLER_76_154 ();
 sg13g2_fill_1 FILLER_76_156 ();
 sg13g2_fill_2 FILLER_76_190 ();
 sg13g2_fill_1 FILLER_76_224 ();
 sg13g2_fill_2 FILLER_76_234 ();
 sg13g2_fill_1 FILLER_76_236 ();
 sg13g2_fill_2 FILLER_76_260 ();
 sg13g2_fill_1 FILLER_76_262 ();
 sg13g2_fill_1 FILLER_76_313 ();
 sg13g2_fill_1 FILLER_76_354 ();
 sg13g2_fill_2 FILLER_76_375 ();
 sg13g2_fill_1 FILLER_76_377 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_4 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_46 ();
 sg13g2_decap_8 FILLER_77_51 ();
 sg13g2_decap_8 FILLER_77_58 ();
 sg13g2_decap_8 FILLER_77_65 ();
 sg13g2_decap_8 FILLER_77_72 ();
 sg13g2_decap_8 FILLER_77_79 ();
 sg13g2_decap_8 FILLER_77_86 ();
 sg13g2_decap_8 FILLER_77_93 ();
 sg13g2_fill_1 FILLER_77_100 ();
 sg13g2_fill_1 FILLER_77_105 ();
 sg13g2_fill_2 FILLER_77_138 ();
 sg13g2_fill_2 FILLER_77_149 ();
 sg13g2_fill_1 FILLER_77_166 ();
 sg13g2_fill_1 FILLER_77_203 ();
 sg13g2_fill_1 FILLER_77_230 ();
 sg13g2_fill_1 FILLER_77_270 ();
 sg13g2_fill_2 FILLER_77_297 ();
 sg13g2_fill_2 FILLER_77_339 ();
 sg13g2_fill_1 FILLER_77_341 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_4 FILLER_78_42 ();
 sg13g2_fill_2 FILLER_78_46 ();
 sg13g2_decap_8 FILLER_78_51 ();
 sg13g2_decap_8 FILLER_78_58 ();
 sg13g2_decap_8 FILLER_78_65 ();
 sg13g2_decap_8 FILLER_78_72 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_fill_1 FILLER_78_105 ();
 sg13g2_decap_4 FILLER_78_207 ();
 sg13g2_fill_2 FILLER_78_219 ();
 sg13g2_fill_2 FILLER_78_235 ();
 sg13g2_fill_2 FILLER_78_251 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_fill_2 FILLER_79_105 ();
 sg13g2_decap_4 FILLER_79_174 ();
 sg13g2_fill_1 FILLER_79_178 ();
 sg13g2_decap_4 FILLER_79_404 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_8 FILLER_80_92 ();
 sg13g2_decap_8 FILLER_80_99 ();
 sg13g2_decap_8 FILLER_80_106 ();
 sg13g2_fill_2 FILLER_80_113 ();
 sg13g2_fill_1 FILLER_80_140 ();
 sg13g2_fill_2 FILLER_80_154 ();
 sg13g2_decap_8 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_179 ();
 sg13g2_decap_8 FILLER_80_186 ();
 sg13g2_decap_4 FILLER_80_193 ();
 sg13g2_fill_1 FILLER_80_197 ();
 sg13g2_decap_8 FILLER_80_202 ();
 sg13g2_decap_8 FILLER_80_209 ();
 sg13g2_fill_1 FILLER_80_216 ();
 sg13g2_fill_1 FILLER_80_262 ();
 sg13g2_fill_1 FILLER_80_332 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net151;
 assign uio_oe[6] = net152;
 assign uio_oe[7] = net153;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
endmodule

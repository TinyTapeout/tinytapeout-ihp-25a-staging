module tt_um_toivoh_demo_tt08 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire \dtop.detune_counter[10] ;
 wire \dtop.detune_counter[11] ;
 wire \dtop.detune_counter[12] ;
 wire \dtop.detune_counter[13] ;
 wire \dtop.detune_counter[14] ;
 wire \dtop.detune_counter[15] ;
 wire \dtop.detune_counter[16] ;
 wire \dtop.detune_counter[17] ;
 wire \dtop.detune_counter[4] ;
 wire \dtop.detune_counter[5] ;
 wire \dtop.detune_counter[6] ;
 wire \dtop.detune_counter[7] ;
 wire \dtop.detune_counter[8] ;
 wire \dtop.detune_counter[9] ;
 wire \dtop.enable ;
 wire \dtop.oct_counter[0] ;
 wire \dtop.oct_counter[1] ;
 wire \dtop.oct_counter[2] ;
 wire \dtop.oct_counter[3] ;
 wire \dtop.oct_counter[4] ;
 wire \dtop.oct_counter[5] ;
 wire \dtop.oct_counter[6] ;
 wire \dtop.out_sample[0] ;
 wire \dtop.out_sample[1] ;
 wire \dtop.out_sample[2] ;
 wire \dtop.out_sample[3] ;
 wire \dtop.out_sample[4] ;
 wire \dtop.out_sample[5] ;
 wire \dtop.out_sample[6] ;
 wire \dtop.player_inst.program_addr[0] ;
 wire \dtop.player_inst.program_addr[1] ;
 wire \dtop.player_inst.program_addr[2] ;
 wire \dtop.player_inst.program_addr[3] ;
 wire \dtop.player_inst.program_addr[4] ;
 wire \dtop.player_inst.program_addr[5] ;
 wire \dtop.player_inst.program_addr[6] ;
 wire \dtop.player_inst.synth.alu.acc[0] ;
 wire \dtop.player_inst.synth.alu.acc[10] ;
 wire \dtop.player_inst.synth.alu.acc[1] ;
 wire \dtop.player_inst.synth.alu.acc[2] ;
 wire \dtop.player_inst.synth.alu.acc[3] ;
 wire \dtop.player_inst.synth.alu.acc[4] ;
 wire \dtop.player_inst.synth.alu.acc[5] ;
 wire \dtop.player_inst.synth.alu.acc[6] ;
 wire \dtop.player_inst.synth.alu.acc[7] ;
 wire \dtop.player_inst.synth.alu.acc[8] ;
 wire \dtop.player_inst.synth.alu.acc[9] ;
 wire \dtop.player_inst.synth.alu.carry ;
 wire \dtop.player_inst.synth.alu.oct_en ;
 wire \dtop.player_inst.synth.alu.registers[0][0] ;
 wire \dtop.player_inst.synth.alu.registers[0][10] ;
 wire \dtop.player_inst.synth.alu.registers[0][1] ;
 wire \dtop.player_inst.synth.alu.registers[0][2] ;
 wire \dtop.player_inst.synth.alu.registers[0][3] ;
 wire \dtop.player_inst.synth.alu.registers[0][4] ;
 wire \dtop.player_inst.synth.alu.registers[0][5] ;
 wire \dtop.player_inst.synth.alu.registers[0][6] ;
 wire \dtop.player_inst.synth.alu.registers[0][7] ;
 wire \dtop.player_inst.synth.alu.registers[0][8] ;
 wire \dtop.player_inst.synth.alu.registers[0][9] ;
 wire \dtop.player_inst.synth.alu.registers[1][0] ;
 wire \dtop.player_inst.synth.alu.registers[1][10] ;
 wire \dtop.player_inst.synth.alu.registers[1][1] ;
 wire \dtop.player_inst.synth.alu.registers[1][2] ;
 wire \dtop.player_inst.synth.alu.registers[1][3] ;
 wire \dtop.player_inst.synth.alu.registers[1][4] ;
 wire \dtop.player_inst.synth.alu.registers[1][5] ;
 wire \dtop.player_inst.synth.alu.registers[1][6] ;
 wire \dtop.player_inst.synth.alu.registers[1][7] ;
 wire \dtop.player_inst.synth.alu.registers[1][8] ;
 wire \dtop.player_inst.synth.alu.registers[1][9] ;
 wire \dtop.player_inst.synth.alu.registers[2][0] ;
 wire \dtop.player_inst.synth.alu.registers[2][1] ;
 wire \dtop.player_inst.synth.alu.registers[2][2] ;
 wire \dtop.player_inst.synth.alu.registers[2][3] ;
 wire \dtop.player_inst.synth.alu.registers[2][4] ;
 wire \dtop.player_inst.synth.alu.registers[2][5] ;
 wire \dtop.player_inst.synth.alu.registers[2][6] ;
 wire \dtop.player_inst.synth.alu.registers[2][7] ;
 wire \dtop.player_inst.synth.alu.registers[3][0] ;
 wire \dtop.player_inst.synth.alu.registers[3][1] ;
 wire \dtop.player_inst.synth.alu.registers[3][2] ;
 wire \dtop.player_inst.synth.alu.registers[3][3] ;
 wire \dtop.player_inst.synth.alu.registers[3][4] ;
 wire \dtop.player_inst.synth.alu.registers[3][5] ;
 wire \dtop.player_inst.synth.alu.registers[3][6] ;
 wire \dtop.player_inst.synth.alu.registers[3][7] ;
 wire \dtop.player_inst.synth.alu.registers[4][0] ;
 wire \dtop.player_inst.synth.alu.registers[4][10] ;
 wire \dtop.player_inst.synth.alu.registers[4][1] ;
 wire \dtop.player_inst.synth.alu.registers[4][2] ;
 wire \dtop.player_inst.synth.alu.registers[4][3] ;
 wire \dtop.player_inst.synth.alu.registers[4][4] ;
 wire \dtop.player_inst.synth.alu.registers[4][5] ;
 wire \dtop.player_inst.synth.alu.registers[4][6] ;
 wire \dtop.player_inst.synth.alu.registers[4][7] ;
 wire \dtop.player_inst.synth.alu.registers[4][8] ;
 wire \dtop.player_inst.synth.alu.registers[4][9] ;
 wire \dtop.player_inst.synth.alu.registers[5][0] ;
 wire \dtop.player_inst.synth.alu.registers[5][1] ;
 wire \dtop.player_inst.synth.alu.registers[5][2] ;
 wire \dtop.player_inst.synth.alu.registers[5][3] ;
 wire \dtop.player_inst.synth.alu.registers[5][4] ;
 wire \dtop.player_inst.synth.alu.registers[5][5] ;
 wire \dtop.player_inst.synth.alu.registers[5][6] ;
 wire \dtop.vsync ;
 wire \dtop.vtop.color[4] ;
 wire \dtop.vtop.color[5] ;
 wire \dtop.vtop.color[6] ;
 wire \dtop.vtop.color[7] ;
 wire \dtop.vtop.dphases[0][0] ;
 wire \dtop.vtop.dphases[0][10] ;
 wire \dtop.vtop.dphases[0][1] ;
 wire \dtop.vtop.dphases[0][2] ;
 wire \dtop.vtop.dphases[0][3] ;
 wire \dtop.vtop.dphases[0][4] ;
 wire \dtop.vtop.dphases[0][5] ;
 wire \dtop.vtop.dphases[0][6] ;
 wire \dtop.vtop.dphases[0][7] ;
 wire \dtop.vtop.dphases[0][8] ;
 wire \dtop.vtop.dphases[0][9] ;
 wire \dtop.vtop.dphases[1][0] ;
 wire \dtop.vtop.dphases[1][10] ;
 wire \dtop.vtop.dphases[1][1] ;
 wire \dtop.vtop.dphases[1][2] ;
 wire \dtop.vtop.dphases[1][3] ;
 wire \dtop.vtop.dphases[1][4] ;
 wire \dtop.vtop.dphases[1][5] ;
 wire \dtop.vtop.dphases[1][6] ;
 wire \dtop.vtop.dphases[1][7] ;
 wire \dtop.vtop.dphases[1][8] ;
 wire \dtop.vtop.dphases[1][9] ;
 wire \dtop.vtop.dphases[2][0] ;
 wire \dtop.vtop.dphases[2][10] ;
 wire \dtop.vtop.dphases[2][1] ;
 wire \dtop.vtop.dphases[2][2] ;
 wire \dtop.vtop.dphases[2][3] ;
 wire \dtop.vtop.dphases[2][4] ;
 wire \dtop.vtop.dphases[2][5] ;
 wire \dtop.vtop.dphases[2][6] ;
 wire \dtop.vtop.dphases[2][7] ;
 wire \dtop.vtop.dphases[2][8] ;
 wire \dtop.vtop.dphases[2][9] ;
 wire \dtop.vtop.logo.addr[5] ;
 wire \dtop.vtop.logo.addr[6] ;
 wire \dtop.vtop.logo.addr[7] ;
 wire \dtop.vtop.logo.addr[8] ;
 wire \dtop.vtop.logo.addr[9] ;
 wire \dtop.vtop.pipeline.cosappr_acc[0] ;
 wire \dtop.vtop.pipeline.cosappr_acc[1] ;
 wire \dtop.vtop.pipeline.cosappr_acc[2] ;
 wire \dtop.vtop.pipeline.cosappr_acc[3] ;
 wire \dtop.vtop.pipeline.cosappr_acc[4] ;
 wire \dtop.vtop.pipeline.cosappr_acc[5] ;
 wire \dtop.vtop.pipeline.cosappr_acc[6] ;
 wire \dtop.vtop.pipeline.cosappr_acc[7] ;
 wire \dtop.vtop.pipeline.cosappr_acc[8] ;
 wire \dtop.vtop.pipeline.dz[0] ;
 wire \dtop.vtop.pipeline.dz[1] ;
 wire \dtop.vtop.pipeline.dz[2] ;
 wire \dtop.vtop.pipeline.dz[3] ;
 wire \dtop.vtop.pipeline.dz[4] ;
 wire \dtop.vtop.pipeline.dz[5] ;
 wire \dtop.vtop.pipeline.dz[6] ;
 wire \dtop.vtop.pipeline.dz[7] ;
 wire \dtop.vtop.pipeline.dz[8] ;
 wire \dtop.vtop.pipeline.neg_t[0] ;
 wire \dtop.vtop.pipeline.neg_t[1] ;
 wire \dtop.vtop.pipeline.neg_t[2] ;
 wire \dtop.vtop.pipeline.neg_t[3] ;
 wire \dtop.vtop.pipeline.neg_t[4] ;
 wire \dtop.vtop.pipeline.neg_t[5] ;
 wire \dtop.vtop.pipeline.neg_t[6] ;
 wire \dtop.vtop.pipeline.neg_t[7] ;
 wire \dtop.vtop.pipeline.neg_t[8] ;
 wire \dtop.vtop.pipeline.neg_t[9] ;
 wire \dtop.vtop.pipeline.next_nstep_counter[0] ;
 wire \dtop.vtop.pipeline.nstep[0] ;
 wire \dtop.vtop.pipeline.nstep[1] ;
 wire \dtop.vtop.pipeline.nstep_counter[0] ;
 wire \dtop.vtop.pipeline.nstep_counter[1] ;
 wire \dtop.vtop.pipeline.nstep_counter[2] ;
 wire \dtop.vtop.pipeline.nstep_counter[3] ;
 wire \dtop.vtop.pipeline.nstep_counter[4] ;
 wire \dtop.vtop.pipeline.nstep_zg[0] ;
 wire \dtop.vtop.pipeline.nstep_zg[1] ;
 wire \dtop.vtop.pipeline.phases[0][0] ;
 wire \dtop.vtop.pipeline.phases[0][10] ;
 wire \dtop.vtop.pipeline.phases[0][11] ;
 wire \dtop.vtop.pipeline.phases[0][12] ;
 wire \dtop.vtop.pipeline.phases[0][13] ;
 wire \dtop.vtop.pipeline.phases[0][14] ;
 wire \dtop.vtop.pipeline.phases[0][15] ;
 wire \dtop.vtop.pipeline.phases[0][1] ;
 wire \dtop.vtop.pipeline.phases[0][2] ;
 wire \dtop.vtop.pipeline.phases[0][3] ;
 wire \dtop.vtop.pipeline.phases[0][4] ;
 wire \dtop.vtop.pipeline.phases[0][5] ;
 wire \dtop.vtop.pipeline.phases[0][6] ;
 wire \dtop.vtop.pipeline.phases[0][7] ;
 wire \dtop.vtop.pipeline.phases[0][8] ;
 wire \dtop.vtop.pipeline.phases[0][9] ;
 wire \dtop.vtop.pipeline.phases[1][0] ;
 wire \dtop.vtop.pipeline.phases[1][10] ;
 wire \dtop.vtop.pipeline.phases[1][11] ;
 wire \dtop.vtop.pipeline.phases[1][12] ;
 wire \dtop.vtop.pipeline.phases[1][13] ;
 wire \dtop.vtop.pipeline.phases[1][14] ;
 wire \dtop.vtop.pipeline.phases[1][15] ;
 wire \dtop.vtop.pipeline.phases[1][1] ;
 wire \dtop.vtop.pipeline.phases[1][2] ;
 wire \dtop.vtop.pipeline.phases[1][3] ;
 wire \dtop.vtop.pipeline.phases[1][4] ;
 wire \dtop.vtop.pipeline.phases[1][5] ;
 wire \dtop.vtop.pipeline.phases[1][6] ;
 wire \dtop.vtop.pipeline.phases[1][7] ;
 wire \dtop.vtop.pipeline.phases[1][8] ;
 wire \dtop.vtop.pipeline.phases[1][9] ;
 wire \dtop.vtop.pipeline.phases[2][0] ;
 wire \dtop.vtop.pipeline.phases[2][10] ;
 wire \dtop.vtop.pipeline.phases[2][11] ;
 wire \dtop.vtop.pipeline.phases[2][12] ;
 wire \dtop.vtop.pipeline.phases[2][13] ;
 wire \dtop.vtop.pipeline.phases[2][14] ;
 wire \dtop.vtop.pipeline.phases[2][15] ;
 wire \dtop.vtop.pipeline.phases[2][1] ;
 wire \dtop.vtop.pipeline.phases[2][2] ;
 wire \dtop.vtop.pipeline.phases[2][3] ;
 wire \dtop.vtop.pipeline.phases[2][4] ;
 wire \dtop.vtop.pipeline.phases[2][5] ;
 wire \dtop.vtop.pipeline.phases[2][6] ;
 wire \dtop.vtop.pipeline.phases[2][7] ;
 wire \dtop.vtop.pipeline.phases[2][8] ;
 wire \dtop.vtop.pipeline.phases[2][9] ;
 wire \dtop.vtop.pipeline.wave_index[0] ;
 wire \dtop.vtop.pipeline.wave_index[1] ;
 wire \dtop.vtop.pipeline.z[0] ;
 wire \dtop.vtop.pipeline.z[10] ;
 wire \dtop.vtop.pipeline.z[11] ;
 wire \dtop.vtop.pipeline.z[12] ;
 wire \dtop.vtop.pipeline.z[13] ;
 wire \dtop.vtop.pipeline.z[14] ;
 wire \dtop.vtop.pipeline.z[1] ;
 wire \dtop.vtop.pipeline.z[2] ;
 wire \dtop.vtop.pipeline.z[3] ;
 wire \dtop.vtop.pipeline.z[4] ;
 wire \dtop.vtop.pipeline.z[5] ;
 wire \dtop.vtop.pipeline.z[6] ;
 wire \dtop.vtop.pipeline.z[7] ;
 wire \dtop.vtop.pipeline.z[8] ;
 wire \dtop.vtop.pipeline.z[9] ;
 wire \dtop.vtop.pipeline.zg[0] ;
 wire \dtop.vtop.pipeline.zg[1] ;
 wire \dtop.vtop.pipeline.zg[2] ;
 wire \dtop.vtop.pipeline.zg[3] ;
 wire \dtop.vtop.pipeline.zg[4] ;
 wire \dtop.vtop.pipeline.zg[5] ;
 wire \dtop.vtop.pipeline.zg[6] ;
 wire \dtop.vtop.pipeline.zg[7] ;
 wire \dtop.vtop.pipeline.zg[8] ;
 wire \dtop.vtop.pipeline.zg[9] ;
 wire \dtop.vtop.pipeline.zg_acc[0] ;
 wire \dtop.vtop.pipeline.zg_acc[1] ;
 wire \dtop.vtop.pipeline.zg_acc[2] ;
 wire \dtop.vtop.pipeline.zg_acc[3] ;
 wire \dtop.vtop.pipeline.zg_acc[4] ;
 wire \dtop.vtop.pipeline.zg_acc[5] ;
 wire \dtop.vtop.pipeline.zg_acc[6] ;
 wire \dtop.vtop.pipeline.zg_acc[7] ;
 wire \dtop.vtop.pipeline.zg_acc[8] ;
 wire \dtop.vtop.pipeline.zg_acc[9] ;
 wire \dtop.vtop.pipeline.zg_valid ;
 wire \dtop.vtop.rs.saturated ;
 wire \dtop.vtop.rs.scan_y.phase[0] ;
 wire \dtop.vtop.rs.scan_y.phase[1] ;
 wire \dtop.vtop.rs.x_scan.phase[0] ;
 wire \dtop.vtop.rs.x_scan.phase[1] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_leaf_0_clk;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;

 sg13g2_inv_4 _3442_ (.A(net654),
    .Y(_2630_));
 sg13g2_inv_4 _3443_ (.A(net652),
    .Y(_2631_));
 sg13g2_inv_4 _3444_ (.A(net649),
    .Y(_2632_));
 sg13g2_inv_4 _3445_ (.A(\dtop.player_inst.synth.alu.acc[3] ),
    .Y(_2633_));
 sg13g2_inv_4 _3446_ (.A(\dtop.player_inst.synth.alu.acc[2] ),
    .Y(_2634_));
 sg13g2_inv_4 _3447_ (.A(\dtop.player_inst.synth.alu.acc[1] ),
    .Y(_2635_));
 sg13g2_inv_4 _3448_ (.A(net650),
    .Y(_2636_));
 sg13g2_inv_4 _3449_ (.A(\dtop.player_inst.synth.alu.acc[7] ),
    .Y(_2637_));
 sg13g2_inv_2 _3450_ (.Y(_2638_),
    .A(net1164));
 sg13g2_inv_1 _3451_ (.Y(_2639_),
    .A(\dtop.player_inst.synth.alu.acc[9] ));
 sg13g2_inv_2 _3452_ (.Y(_2640_),
    .A(\dtop.player_inst.synth.alu.acc[8] ));
 sg13g2_inv_1 _3453_ (.Y(_2641_),
    .A(net651));
 sg13g2_inv_1 _3454_ (.Y(_2642_),
    .A(net600));
 sg13g2_inv_1 _3455_ (.Y(_2643_),
    .A(\dtop.vtop.pipeline.z[12] ));
 sg13g2_inv_1 _3456_ (.Y(_2644_),
    .A(\dtop.vtop.pipeline.z[11] ));
 sg13g2_inv_1 _3457_ (.Y(_2645_),
    .A(\dtop.vtop.pipeline.z[10] ));
 sg13g2_inv_1 _3458_ (.Y(_2646_),
    .A(\dtop.vtop.pipeline.z[9] ));
 sg13g2_inv_1 _3459_ (.Y(_2647_),
    .A(\dtop.vtop.pipeline.z[8] ));
 sg13g2_inv_1 _3460_ (.Y(_2648_),
    .A(net562));
 sg13g2_inv_1 _3461_ (.Y(_2649_),
    .A(net491));
 sg13g2_inv_1 _3462_ (.Y(_2650_),
    .A(net490));
 sg13g2_inv_1 _3463_ (.Y(_2651_),
    .A(\dtop.vtop.pipeline.dz[8] ));
 sg13g2_inv_1 _3464_ (.Y(_2652_),
    .A(\dtop.vtop.pipeline.neg_t[6] ));
 sg13g2_inv_1 _3465_ (.Y(_2653_),
    .A(\dtop.oct_counter[2] ));
 sg13g2_inv_2 _3466_ (.Y(_2654_),
    .A(\dtop.player_inst.program_addr[6] ));
 sg13g2_inv_1 _3467_ (.Y(_2655_),
    .A(net1204));
 sg13g2_inv_4 _3468_ (.A(net1207),
    .Y(_2656_));
 sg13g2_inv_2 _3469_ (.Y(_2657_),
    .A(net1199));
 sg13g2_inv_2 _3470_ (.Y(_2658_),
    .A(\dtop.detune_counter[14] ));
 sg13g2_inv_4 _3471_ (.A(\dtop.detune_counter[12] ),
    .Y(_2659_));
 sg13g2_inv_1 _3472_ (.Y(_2660_),
    .A(net1230));
 sg13g2_inv_2 _3473_ (.Y(_2661_),
    .A(net1232));
 sg13g2_inv_2 _3474_ (.Y(_2662_),
    .A(\dtop.detune_counter[9] ));
 sg13g2_inv_2 _3475_ (.Y(_2663_),
    .A(\dtop.vtop.logo.addr[9] ));
 sg13g2_inv_1 _3476_ (.Y(_2664_),
    .A(net1166));
 sg13g2_inv_2 _3477_ (.Y(_2665_),
    .A(net1167));
 sg13g2_inv_1 _3478_ (.Y(_2666_),
    .A(net1168));
 sg13g2_inv_1 _3479_ (.Y(_2667_),
    .A(net1170));
 sg13g2_inv_4 _3480_ (.A(\dtop.player_inst.program_addr[0] ),
    .Y(_2668_));
 sg13g2_inv_4 _3481_ (.A(net1219),
    .Y(_2669_));
 sg13g2_inv_1 _3482_ (.Y(_2670_),
    .A(net1211));
 sg13g2_inv_2 _3483_ (.Y(_2671_),
    .A(net1215));
 sg13g2_inv_1 _3484_ (.Y(_2672_),
    .A(net575));
 sg13g2_inv_1 _3485_ (.Y(_2673_),
    .A(\dtop.detune_counter[4] ));
 sg13g2_inv_1 _3486_ (.Y(_2674_),
    .A(\dtop.detune_counter[17] ));
 sg13g2_inv_2 _3487_ (.Y(_2675_),
    .A(\dtop.vtop.pipeline.zg[9] ));
 sg13g2_inv_2 _3488_ (.Y(_2676_),
    .A(net641));
 sg13g2_inv_2 _3489_ (.Y(_2677_),
    .A(net571));
 sg13g2_inv_1 _3490_ (.Y(_2678_),
    .A(net533));
 sg13g2_inv_1 _3491_ (.Y(_2679_),
    .A(net478));
 sg13g2_inv_2 _3492_ (.Y(_2680_),
    .A(net1194));
 sg13g2_inv_1 _3493_ (.Y(_2681_),
    .A(_0061_));
 sg13g2_inv_1 _3494_ (.Y(_2682_),
    .A(\dtop.vtop.rs.x_scan.phase[1] ));
 sg13g2_inv_4 _3495_ (.A(net570),
    .Y(_2683_));
 sg13g2_inv_2 _3496_ (.Y(_2684_),
    .A(_0078_));
 sg13g2_inv_1 _3497_ (.Y(_2685_),
    .A(_0088_));
 sg13g2_inv_2 _3498_ (.Y(_2686_),
    .A(net607));
 sg13g2_inv_1 _3499_ (.Y(_2687_),
    .A(net516));
 sg13g2_inv_1 _3500_ (.Y(_2688_),
    .A(\dtop.vtop.pipeline.phases[2][15] ));
 sg13g2_inv_1 _3501_ (.Y(_2689_),
    .A(\dtop.vtop.pipeline.phases[1][15] ));
 sg13g2_inv_1 _3502_ (.Y(_2690_),
    .A(\dtop.vtop.dphases[1][0] ));
 sg13g2_inv_2 _3503_ (.Y(_2691_),
    .A(net1188));
 sg13g2_inv_1 _3504_ (.Y(_2692_),
    .A(\dtop.vtop.dphases[1][1] ));
 sg13g2_inv_1 _3505_ (.Y(_2693_),
    .A(\dtop.vtop.dphases[1][2] ));
 sg13g2_inv_1 _3506_ (.Y(_2694_),
    .A(\dtop.vtop.dphases[1][3] ));
 sg13g2_inv_1 _3507_ (.Y(_2695_),
    .A(\dtop.vtop.dphases[1][4] ));
 sg13g2_inv_1 _3508_ (.Y(_2696_),
    .A(\dtop.vtop.dphases[1][5] ));
 sg13g2_inv_1 _3509_ (.Y(_2697_),
    .A(_0025_));
 sg13g2_inv_1 _3510_ (.Y(_2698_),
    .A(\dtop.vtop.dphases[1][9] ));
 sg13g2_inv_1 _3511_ (.Y(_2699_),
    .A(net444));
 sg13g2_inv_1 _3512_ (.Y(_2700_),
    .A(net473));
 sg13g2_inv_1 _3513_ (.Y(_2701_),
    .A(net469));
 sg13g2_inv_1 _3514_ (.Y(_2702_),
    .A(net531));
 sg13g2_nor2_2 _3515_ (.A(net1202),
    .B(net1199),
    .Y(_2703_));
 sg13g2_or2_2 _3516_ (.X(_2704_),
    .B(net1198),
    .A(net1202));
 sg13g2_nor2_1 _3517_ (.A(_2656_),
    .B(_2704_),
    .Y(_2705_));
 sg13g2_nand2_2 _3518_ (.Y(_2706_),
    .A(net1205),
    .B(_2703_));
 sg13g2_nor2b_1 _3519_ (.A(net1214),
    .B_N(net1209),
    .Y(_2707_));
 sg13g2_nand2b_1 _3520_ (.Y(_2708_),
    .B(net1209),
    .A_N(net1212));
 sg13g2_nand3b_1 _3521_ (.B(net1210),
    .C(net1218),
    .Y(_2709_),
    .A_N(net1213));
 sg13g2_and2_1 _3522_ (.A(net1221),
    .B(net1216),
    .X(_2710_));
 sg13g2_nand2_1 _3523_ (.Y(_2711_),
    .A(net1221),
    .B(net1216));
 sg13g2_nor2_2 _3524_ (.A(net1158),
    .B(net1157),
    .Y(_2712_));
 sg13g2_and2_2 _3525_ (.A(net1139),
    .B(net1136),
    .X(_2713_));
 sg13g2_nand2_2 _3526_ (.Y(_2714_),
    .A(net1139),
    .B(net1136));
 sg13g2_and3_1 _3527_ (.X(_2715_),
    .A(net1201),
    .B(net1206),
    .C(net1198));
 sg13g2_nand3_1 _3528_ (.B(net1206),
    .C(net1198),
    .A(net1201),
    .Y(_2716_));
 sg13g2_nor2b_2 _3529_ (.A(net1209),
    .B_N(net1212),
    .Y(_2717_));
 sg13g2_nand2b_1 _3530_ (.Y(_2718_),
    .B(net1212),
    .A_N(net1209));
 sg13g2_nor2_2 _3531_ (.A(net1153),
    .B(net1151),
    .Y(_2719_));
 sg13g2_nor2_2 _3532_ (.A(net1156),
    .B(net1151),
    .Y(_2720_));
 sg13g2_nor3_2 _3533_ (.A(net1156),
    .B(_2716_),
    .C(net1152),
    .Y(_2721_));
 sg13g2_nor2_2 _3534_ (.A(net1202),
    .B(net1205),
    .Y(_2722_));
 sg13g2_or2_2 _3535_ (.X(_2723_),
    .B(net1205),
    .A(net1201));
 sg13g2_nor3_2 _3536_ (.A(net1201),
    .B(net1206),
    .C(net1198),
    .Y(_2724_));
 sg13g2_or3_2 _3537_ (.A(net1201),
    .B(net1206),
    .C(net1198),
    .X(_2725_));
 sg13g2_nor2_2 _3538_ (.A(net1221),
    .B(net1217),
    .Y(_2726_));
 sg13g2_or2_2 _3539_ (.X(_2727_),
    .B(net1217),
    .A(net1221));
 sg13g2_nor2_2 _3540_ (.A(net1152),
    .B(_2727_),
    .Y(_2728_));
 sg13g2_a21oi_2 _3541_ (.B1(_2721_),
    .Y(_2729_),
    .A2(_2728_),
    .A1(net1149));
 sg13g2_nor2_2 _3542_ (.A(_2657_),
    .B(_2723_),
    .Y(_2730_));
 sg13g2_nand2_1 _3543_ (.Y(_2731_),
    .A(net1199),
    .B(_2722_));
 sg13g2_nor2_1 _3544_ (.A(net1209),
    .B(net1212),
    .Y(_2732_));
 sg13g2_or2_2 _3545_ (.X(_2733_),
    .B(net1213),
    .A(net1209));
 sg13g2_nor2_2 _3546_ (.A(net1156),
    .B(_2733_),
    .Y(_2734_));
 sg13g2_nand2_1 _3547_ (.Y(_2735_),
    .A(net1135),
    .B(_2734_));
 sg13g2_nand3_1 _3548_ (.B(_2729_),
    .C(_2735_),
    .A(_2714_),
    .Y(_2736_));
 sg13g2_nand2b_2 _3549_ (.Y(_2737_),
    .B(net1201),
    .A_N(net1206));
 sg13g2_nor2_1 _3550_ (.A(\dtop.player_inst.program_addr[6] ),
    .B(_2737_),
    .Y(_2738_));
 sg13g2_nand2b_2 _3551_ (.Y(_2739_),
    .B(_2654_),
    .A_N(_2737_));
 sg13g2_nor3_2 _3552_ (.A(net1216),
    .B(net1210),
    .C(net1213),
    .Y(_2740_));
 sg13g2_and2_1 _3553_ (.A(net1222),
    .B(_2740_),
    .X(_2741_));
 sg13g2_nand2_1 _3554_ (.Y(_2742_),
    .A(net1222),
    .B(_2740_));
 sg13g2_nor2b_2 _3555_ (.A(net1221),
    .B_N(net1216),
    .Y(_2743_));
 sg13g2_nand2b_1 _3556_ (.Y(_2744_),
    .B(net1219),
    .A_N(net1224));
 sg13g2_nor2_2 _3557_ (.A(_2733_),
    .B(net1146),
    .Y(_2745_));
 sg13g2_o21ai_1 _3558_ (.B1(net1133),
    .Y(_2746_),
    .A1(_2741_),
    .A2(_2745_));
 sg13g2_and2_2 _3559_ (.A(net1209),
    .B(net1212),
    .X(_2747_));
 sg13g2_nand2_1 _3560_ (.Y(_2748_),
    .A(net1210),
    .B(net1213));
 sg13g2_nor2_2 _3561_ (.A(net1217),
    .B(_2748_),
    .Y(_2749_));
 sg13g2_nand3b_1 _3562_ (.B(net1210),
    .C(net1213),
    .Y(_2750_),
    .A_N(net1216));
 sg13g2_nand2b_2 _3563_ (.Y(_2751_),
    .B(net1222),
    .A_N(net1216));
 sg13g2_nor2_2 _3564_ (.A(_2668_),
    .B(_2750_),
    .Y(_2752_));
 sg13g2_nand2_1 _3565_ (.Y(_2753_),
    .A(net1133),
    .B(_2752_));
 sg13g2_nor3_2 _3566_ (.A(\dtop.player_inst.program_addr[6] ),
    .B(net1160),
    .C(_2737_),
    .Y(_2754_));
 sg13g2_nor4_2 _3567_ (.A(\dtop.player_inst.program_addr[6] ),
    .B(net1157),
    .C(net1152),
    .Y(_2755_),
    .D(_2737_));
 sg13g2_nor2_1 _3568_ (.A(_2754_),
    .B(_2755_),
    .Y(_2756_));
 sg13g2_nor2_1 _3569_ (.A(net1157),
    .B(net1145),
    .Y(_2757_));
 sg13g2_nand4_1 _3570_ (.B(net1218),
    .C(net1210),
    .A(net1223),
    .Y(_2758_),
    .D(net1213));
 sg13g2_nor3_2 _3571_ (.A(net1202),
    .B(_2656_),
    .C(_2657_),
    .Y(_2759_));
 sg13g2_nand3b_1 _3572_ (.B(net1205),
    .C(net1198),
    .Y(_2760_),
    .A_N(net1201));
 sg13g2_nand2_1 _3573_ (.Y(_2761_),
    .A(net1131),
    .B(net1130));
 sg13g2_nor2_2 _3574_ (.A(net1147),
    .B(net1145),
    .Y(_2762_));
 sg13g2_nor4_2 _3575_ (.A(\dtop.player_inst.program_addr[6] ),
    .B(_2737_),
    .C(net1147),
    .Y(_2763_),
    .D(net1145));
 sg13g2_nor4_2 _3576_ (.A(net1221),
    .B(net1216),
    .C(net1209),
    .Y(_2764_),
    .D(net1212));
 sg13g2_or4_2 _3577_ (.A(net1223),
    .B(net1218),
    .C(net1210),
    .D(net1213),
    .X(_2765_));
 sg13g2_nor2_1 _3578_ (.A(net1152),
    .B(net1146),
    .Y(_2766_));
 sg13g2_nand2_2 _3579_ (.Y(_2767_),
    .A(_2717_),
    .B(_2743_));
 sg13g2_nand3_1 _3580_ (.B(net1133),
    .C(_2743_),
    .A(net1212),
    .Y(_2768_));
 sg13g2_o21ai_1 _3581_ (.B1(_2761_),
    .Y(_2769_),
    .A1(_2739_),
    .A2(_2765_));
 sg13g2_nand4_1 _3582_ (.B(_2753_),
    .C(_2756_),
    .A(_2746_),
    .Y(_2770_),
    .D(_2768_));
 sg13g2_nor2_1 _3583_ (.A(_2769_),
    .B(_2770_),
    .Y(_2771_));
 sg13g2_nor2_2 _3584_ (.A(net1158),
    .B(_2751_),
    .Y(_2772_));
 sg13g2_or2_2 _3585_ (.X(_2773_),
    .B(_2751_),
    .A(net1158));
 sg13g2_nor2_2 _3586_ (.A(net1223),
    .B(_2750_),
    .Y(_2774_));
 sg13g2_nand2_1 _3587_ (.Y(_2775_),
    .A(_2726_),
    .B(_2747_));
 sg13g2_o21ai_1 _3588_ (.B1(_2709_),
    .Y(_2776_),
    .A1(net1223),
    .A2(_2750_));
 sg13g2_o21ai_1 _3589_ (.B1(net1134),
    .Y(_2777_),
    .A1(_2772_),
    .A2(_2776_));
 sg13g2_nand2_2 _3590_ (.Y(_2778_),
    .A(_2707_),
    .B(_2743_));
 sg13g2_nor2_2 _3591_ (.A(_2725_),
    .B(_2778_),
    .Y(_2779_));
 sg13g2_nor2_2 _3592_ (.A(net1148),
    .B(_2773_),
    .Y(_2780_));
 sg13g2_nor2_1 _3593_ (.A(net1158),
    .B(_2727_),
    .Y(_2781_));
 sg13g2_nor3_2 _3594_ (.A(net1159),
    .B(net1153),
    .C(_2727_),
    .Y(_2782_));
 sg13g2_nor3_2 _3595_ (.A(net1158),
    .B(net1156),
    .C(net1153),
    .Y(_2783_));
 sg13g2_or4_1 _3596_ (.A(_2779_),
    .B(_2780_),
    .C(_2782_),
    .D(_2783_),
    .X(_2784_));
 sg13g2_a22oi_1 _3597_ (.Y(_2785_),
    .B1(_2732_),
    .B2(_2710_),
    .A2(_2726_),
    .A1(_2717_));
 sg13g2_nor4_2 _3598_ (.A(_2656_),
    .B(_2704_),
    .C(net1152),
    .Y(_2786_),
    .D(_2727_));
 sg13g2_a21oi_1 _3599_ (.A1(_2706_),
    .A2(_2739_),
    .Y(_2787_),
    .B1(_2785_));
 sg13g2_nand3_1 _3600_ (.B(_2722_),
    .C(_2764_),
    .A(net1198),
    .Y(_2788_));
 sg13g2_nand2_1 _3601_ (.Y(_2789_),
    .A(net1150),
    .B(_2749_));
 sg13g2_nor3_2 _3602_ (.A(net1158),
    .B(net1148),
    .C(_2727_),
    .Y(_2790_));
 sg13g2_a21oi_1 _3603_ (.A1(_2712_),
    .A2(net1150),
    .Y(_2791_),
    .B1(_2790_));
 sg13g2_nand2_1 _3604_ (.Y(_2792_),
    .A(net1154),
    .B(_2747_));
 sg13g2_nor2_2 _3605_ (.A(net1151),
    .B(_2751_),
    .Y(_2793_));
 sg13g2_or2_2 _3606_ (.X(_2794_),
    .B(_2751_),
    .A(net1151));
 sg13g2_a21oi_1 _3607_ (.A1(_2758_),
    .A2(_2794_),
    .Y(_2795_),
    .B1(net1148));
 sg13g2_nor2b_1 _3608_ (.A(_2795_),
    .B_N(_2792_),
    .Y(_2796_));
 sg13g2_nand4_1 _3609_ (.B(_2789_),
    .C(_2791_),
    .A(_2788_),
    .Y(_2797_),
    .D(_2796_));
 sg13g2_nor3_1 _3610_ (.A(_2784_),
    .B(_2787_),
    .C(_2797_),
    .Y(_2798_));
 sg13g2_nand3_1 _3611_ (.B(_2777_),
    .C(_2798_),
    .A(_2771_),
    .Y(_2799_));
 sg13g2_nor3_2 _3612_ (.A(net1156),
    .B(net1148),
    .C(_2733_),
    .Y(_2800_));
 sg13g2_nand4_1 _3613_ (.B(_2722_),
    .C(_2732_),
    .A(net1198),
    .Y(_2801_),
    .D(_2743_));
 sg13g2_o21ai_1 _3614_ (.B1(_2801_),
    .Y(_2802_),
    .A1(_2706_),
    .A2(_2778_));
 sg13g2_or2_1 _3615_ (.X(_2803_),
    .B(_2802_),
    .A(_2800_));
 sg13g2_nand4_1 _3616_ (.B(_2703_),
    .C(_2707_),
    .A(net1205),
    .Y(_2804_),
    .D(_2726_));
 sg13g2_nand3_1 _3617_ (.B(net1150),
    .C(_2740_),
    .A(net1222),
    .Y(_2805_));
 sg13g2_nand2_1 _3618_ (.Y(_2806_),
    .A(_2804_),
    .B(_2805_));
 sg13g2_nor2_2 _3619_ (.A(_2654_),
    .B(_2737_),
    .Y(_2807_));
 sg13g2_nand3b_1 _3620_ (.B(net1201),
    .C(\dtop.player_inst.program_addr[6] ),
    .Y(_2808_),
    .A_N(net1206));
 sg13g2_or2_1 _3621_ (.X(_2809_),
    .B(_2808_),
    .A(_2765_));
 sg13g2_nor3_2 _3622_ (.A(_2657_),
    .B(_2723_),
    .C(_2758_),
    .Y(_2810_));
 sg13g2_nor3_2 _3623_ (.A(_2733_),
    .B(net1146),
    .C(_2808_),
    .Y(_2811_));
 sg13g2_nand4_1 _3624_ (.B(net1217),
    .C(_2703_),
    .A(net1205),
    .Y(_2812_),
    .D(_2747_));
 sg13g2_nor4_2 _3625_ (.A(_2656_),
    .B(_2704_),
    .C(net1151),
    .Y(_2813_),
    .D(_2751_));
 sg13g2_nand2_1 _3626_ (.Y(_2814_),
    .A(net1137),
    .B(_2745_));
 sg13g2_a22oi_1 _3627_ (.Y(_2815_),
    .B1(_2757_),
    .B2(net1133),
    .A2(_2740_),
    .A1(net1155));
 sg13g2_nor3_2 _3628_ (.A(net1153),
    .B(_2733_),
    .C(net1146),
    .Y(_2816_));
 sg13g2_a221oi_1 _3629_ (.B2(net1132),
    .C1(_2816_),
    .B1(_2757_),
    .A1(net1155),
    .Y(_2817_),
    .A2(_2740_));
 sg13g2_nand2b_1 _3630_ (.Y(_2818_),
    .B(_2815_),
    .A_N(_2816_));
 sg13g2_nor3_1 _3631_ (.A(_2657_),
    .B(net1151),
    .C(_2723_),
    .Y(_2819_));
 sg13g2_a22oi_1 _3632_ (.Y(_2820_),
    .B1(_2774_),
    .B2(net1139),
    .A2(net1135),
    .A1(_2728_));
 sg13g2_a21oi_1 _3633_ (.A1(_2750_),
    .A2(_2794_),
    .Y(_2821_),
    .B1(net1143));
 sg13g2_nor3_2 _3634_ (.A(net1152),
    .B(net1146),
    .C(net1143),
    .Y(_2822_));
 sg13g2_nand2_2 _3635_ (.Y(_2823_),
    .A(net1138),
    .B(_2764_));
 sg13g2_xnor2_1 _3636_ (.Y(_2824_),
    .A(net1221),
    .B(net1216));
 sg13g2_nor3_2 _3637_ (.A(net1159),
    .B(net1143),
    .C(_2824_),
    .Y(_2825_));
 sg13g2_nor3_1 _3638_ (.A(net1157),
    .B(net1151),
    .C(net1143),
    .Y(_2826_));
 sg13g2_nor3_1 _3639_ (.A(net1159),
    .B(_2727_),
    .C(net1144),
    .Y(_2827_));
 sg13g2_nor2_1 _3640_ (.A(_2826_),
    .B(_2827_),
    .Y(_2828_));
 sg13g2_nand2_1 _3641_ (.Y(_2829_),
    .A(_2823_),
    .B(_2828_));
 sg13g2_nor4_2 _3642_ (.A(_2821_),
    .B(_2822_),
    .C(_2825_),
    .Y(_2830_),
    .D(_2829_));
 sg13g2_nand4_1 _3643_ (.B(_2722_),
    .C(_2743_),
    .A(net1199),
    .Y(_2831_),
    .D(_2747_));
 sg13g2_nor2_2 _3644_ (.A(_2733_),
    .B(net1143),
    .Y(_2832_));
 sg13g2_a221oi_1 _3645_ (.B2(_2807_),
    .C1(_2806_),
    .B1(_2764_),
    .A1(net1138),
    .Y(_2833_),
    .A2(_2745_));
 sg13g2_o21ai_1 _3646_ (.B1(net1134),
    .Y(_2834_),
    .A1(_2720_),
    .A2(_2781_));
 sg13g2_nand3_1 _3647_ (.B(_2717_),
    .C(_2726_),
    .A(net1154),
    .Y(_2835_));
 sg13g2_nor2_2 _3648_ (.A(_2716_),
    .B(_2767_),
    .Y(_2836_));
 sg13g2_a221oi_1 _3649_ (.B2(_2762_),
    .C1(_2832_),
    .B1(net1134),
    .A1(_2668_),
    .Y(_2837_),
    .A2(_2719_));
 sg13g2_nand4_1 _3650_ (.B(_2833_),
    .C(_2834_),
    .A(_2812_),
    .Y(_2838_),
    .D(_2837_));
 sg13g2_nor3_1 _3651_ (.A(_2810_),
    .B(_2811_),
    .C(_2813_),
    .Y(_2839_));
 sg13g2_nand2_1 _3652_ (.Y(_2840_),
    .A(_2820_),
    .B(_2839_));
 sg13g2_nor4_1 _3653_ (.A(_2803_),
    .B(_2818_),
    .C(_2838_),
    .D(_2840_),
    .Y(_2841_));
 sg13g2_and2_1 _3654_ (.A(_2830_),
    .B(_2841_),
    .X(_2842_));
 sg13g2_nor2b_1 _3655_ (.A(_2799_),
    .B_N(_2842_),
    .Y(_2843_));
 sg13g2_nand2b_1 _3656_ (.Y(_2844_),
    .B(_2843_),
    .A_N(net1100));
 sg13g2_nor3_1 _3657_ (.A(net1153),
    .B(net1146),
    .C(net1145),
    .Y(_2845_));
 sg13g2_nand2_1 _3658_ (.Y(_2846_),
    .A(net1227),
    .B(_0057_));
 sg13g2_nor2_2 _3659_ (.A(net1229),
    .B(_2846_),
    .Y(_2847_));
 sg13g2_or2_2 _3660_ (.X(_2848_),
    .B(_2846_),
    .A(net1228));
 sg13g2_a21o_1 _3661_ (.A2(_2774_),
    .A1(net1150),
    .B1(_2786_),
    .X(_2849_));
 sg13g2_or4_1 _3662_ (.A(net1139),
    .B(_2811_),
    .C(_2845_),
    .D(_2847_),
    .X(_2850_));
 sg13g2_nor4_1 _3663_ (.A(_2779_),
    .B(_2780_),
    .C(_2849_),
    .D(_2850_),
    .Y(_2851_));
 sg13g2_nor2_1 _3664_ (.A(_2706_),
    .B(_2750_),
    .Y(_2852_));
 sg13g2_nor3_2 _3665_ (.A(net1156),
    .B(_2733_),
    .C(_2808_),
    .Y(_2853_));
 sg13g2_nand2_2 _3666_ (.Y(_2854_),
    .A(_2734_),
    .B(_2807_));
 sg13g2_a221oi_1 _3667_ (.B2(_2741_),
    .C1(_2853_),
    .B1(_2807_),
    .A1(net1138),
    .Y(_2855_),
    .A2(_2749_));
 sg13g2_nor3_2 _3668_ (.A(net1158),
    .B(_2716_),
    .C(_2751_),
    .Y(_2856_));
 sg13g2_nor3_2 _3669_ (.A(net1158),
    .B(net1153),
    .C(net1146),
    .Y(_2857_));
 sg13g2_nor2_1 _3670_ (.A(_2856_),
    .B(_2857_),
    .Y(_2858_));
 sg13g2_nor2_1 _3671_ (.A(net1160),
    .B(net1153),
    .Y(_2859_));
 sg13g2_a21oi_1 _3672_ (.A1(_2785_),
    .A2(_2794_),
    .Y(_2860_),
    .B1(_2739_));
 sg13g2_a21oi_1 _3673_ (.A1(net1132),
    .A2(_2745_),
    .Y(_2861_),
    .B1(_2860_));
 sg13g2_a22oi_1 _3674_ (.Y(_2862_),
    .B1(net1131),
    .B2(net1154),
    .A2(_2752_),
    .A1(net1149));
 sg13g2_nor2_1 _3675_ (.A(net1148),
    .B(_2765_),
    .Y(_2863_));
 sg13g2_nand2_1 _3676_ (.Y(_2864_),
    .A(net1149),
    .B(_2764_));
 sg13g2_o21ai_1 _3677_ (.B1(_2864_),
    .Y(_2865_),
    .A1(_2706_),
    .A2(_2709_));
 sg13g2_o21ai_1 _3678_ (.B1(_2809_),
    .Y(_2866_),
    .A1(_2706_),
    .A2(_2758_));
 sg13g2_nand3_1 _3679_ (.B(_2743_),
    .C(_2747_),
    .A(net1150),
    .Y(_2867_));
 sg13g2_nor2_2 _3680_ (.A(_2725_),
    .B(_2767_),
    .Y(_2868_));
 sg13g2_nor3_1 _3681_ (.A(net1162),
    .B(net1148),
    .C(net1147),
    .Y(_2869_));
 sg13g2_nor4_1 _3682_ (.A(_2795_),
    .B(_2865_),
    .C(_2866_),
    .D(_2869_),
    .Y(_2870_));
 sg13g2_nand3_1 _3683_ (.B(_2717_),
    .C(net1150),
    .A(_2710_),
    .Y(_2871_));
 sg13g2_nand4_1 _3684_ (.B(net1221),
    .C(_2703_),
    .A(net1205),
    .Y(_2872_),
    .D(_2740_));
 sg13g2_and2_1 _3685_ (.A(_2871_),
    .B(_2872_),
    .X(_2873_));
 sg13g2_nand2_1 _3686_ (.Y(_2874_),
    .A(net1154),
    .B(_2749_));
 sg13g2_and4_1 _3687_ (.A(_2862_),
    .B(_2870_),
    .C(_2873_),
    .D(_2874_),
    .X(_2875_));
 sg13g2_nand3b_1 _3688_ (.B(net1227),
    .C(net1228),
    .Y(_2876_),
    .A_N(\dtop.detune_counter[17] ));
 sg13g2_nor2_1 _3689_ (.A(_2659_),
    .B(_2661_),
    .Y(_2877_));
 sg13g2_nand2_2 _3690_ (.Y(_2878_),
    .A(\dtop.detune_counter[12] ),
    .B(net1231));
 sg13g2_nand4_1 _3691_ (.B(\dtop.detune_counter[12] ),
    .C(net1230),
    .A(\dtop.detune_counter[14] ),
    .Y(_2879_),
    .D(net1231));
 sg13g2_nand3b_1 _3692_ (.B(_2879_),
    .C(\dtop.detune_counter[14] ),
    .Y(_2880_),
    .A_N(\dtop.detune_counter[10] ));
 sg13g2_nor2b_2 _3693_ (.A(_2876_),
    .B_N(_2880_),
    .Y(_2881_));
 sg13g2_nand2b_2 _3694_ (.Y(_2882_),
    .B(_2880_),
    .A_N(_2876_));
 sg13g2_nand2_1 _3695_ (.Y(_2883_),
    .A(_2845_),
    .B(net1120));
 sg13g2_or2_2 _3696_ (.X(_2884_),
    .B(_2878_),
    .A(_0087_));
 sg13g2_or4_1 _3697_ (.A(_2706_),
    .B(net1147),
    .C(net1145),
    .D(_2884_),
    .X(_2885_));
 sg13g2_a22oi_1 _3698_ (.Y(_2886_),
    .B1(_2734_),
    .B2(net1137),
    .A2(net1149),
    .A1(_2712_));
 sg13g2_nand2_1 _3699_ (.Y(_2887_),
    .A(net1139),
    .B(_2766_));
 sg13g2_or2_1 _3700_ (.X(_2888_),
    .B(_2887_),
    .A(_2848_));
 sg13g2_and2_2 _3701_ (.A(\dtop.detune_counter[10] ),
    .B(\dtop.detune_counter[9] ),
    .X(_2889_));
 sg13g2_xnor2_1 _3702_ (.Y(_2890_),
    .A(_0061_),
    .B(_2889_));
 sg13g2_nor3_2 _3703_ (.A(net1229),
    .B(net1227),
    .C(_0057_),
    .Y(_2891_));
 sg13g2_or3_2 _3704_ (.A(net1228),
    .B(\dtop.detune_counter[16] ),
    .C(_0057_),
    .X(_2892_));
 sg13g2_nor2_1 _3705_ (.A(net1160),
    .B(_2892_),
    .Y(_2893_));
 sg13g2_nor3_1 _3706_ (.A(net1147),
    .B(net1145),
    .C(net1143),
    .Y(_2894_));
 sg13g2_or3_1 _3707_ (.A(net1146),
    .B(net1145),
    .C(net1143),
    .X(_2895_));
 sg13g2_nor4_1 _3708_ (.A(net1134),
    .B(_2790_),
    .C(_2832_),
    .D(_2894_),
    .Y(_2896_));
 sg13g2_and2_1 _3709_ (.A(net1137),
    .B(_2720_),
    .X(_2897_));
 sg13g2_nor2_1 _3710_ (.A(net1148),
    .B(_2785_),
    .Y(_2898_));
 sg13g2_a221oi_1 _3711_ (.B2(_2728_),
    .C1(_2800_),
    .B1(net1149),
    .A1(net1138),
    .Y(_2899_),
    .A2(_2720_));
 sg13g2_and2_1 _3712_ (.A(_2817_),
    .B(_2899_),
    .X(_2900_));
 sg13g2_nand2_1 _3713_ (.Y(_2901_),
    .A(net1149),
    .B(_2745_));
 sg13g2_a22oi_1 _3714_ (.Y(_2902_),
    .B1(_2772_),
    .B2(net1138),
    .A2(_2745_),
    .A1(_2724_));
 sg13g2_nand3b_1 _3715_ (.B(_2814_),
    .C(_2902_),
    .Y(_2903_),
    .A_N(_2813_));
 sg13g2_nor3_1 _3716_ (.A(_2719_),
    .B(_2806_),
    .C(_2903_),
    .Y(_2904_));
 sg13g2_nand3_1 _3717_ (.B(_2900_),
    .C(_2904_),
    .A(_2830_),
    .Y(_2905_));
 sg13g2_nor2_2 _3718_ (.A(_2876_),
    .B(_2879_),
    .Y(_2906_));
 sg13g2_or2_2 _3719_ (.X(_2907_),
    .B(_2879_),
    .A(_2876_));
 sg13g2_nor2b_1 _3720_ (.A(net1227),
    .B_N(net1229),
    .Y(_2908_));
 sg13g2_and2_2 _3721_ (.A(\dtop.detune_counter[17] ),
    .B(_2908_),
    .X(_2909_));
 sg13g2_nand3b_1 _3722_ (.B(\dtop.detune_counter[17] ),
    .C(net1228),
    .Y(_2910_),
    .A_N(net1227));
 sg13g2_and2_1 _3723_ (.A(_2892_),
    .B(net1142),
    .X(_2911_));
 sg13g2_nand2_1 _3724_ (.Y(_2912_),
    .A(_2892_),
    .B(net1141));
 sg13g2_nor2_1 _3725_ (.A(_2906_),
    .B(_2912_),
    .Y(_2913_));
 sg13g2_nand2_2 _3726_ (.Y(_2914_),
    .A(_2907_),
    .B(_2911_));
 sg13g2_nor4_2 _3727_ (.A(net1228),
    .B(\dtop.detune_counter[16] ),
    .C(_2674_),
    .Y(_2915_),
    .D(_2879_));
 sg13g2_or4_2 _3728_ (.A(net1228),
    .B(net1227),
    .C(_2674_),
    .D(_2879_),
    .X(_2916_));
 sg13g2_nand2_1 _3729_ (.Y(_2917_),
    .A(_2907_),
    .B(_2916_));
 sg13g2_nor3_2 _3730_ (.A(_2906_),
    .B(_2911_),
    .C(_2915_),
    .Y(_2918_));
 sg13g2_nand2_1 _3731_ (.Y(_2919_),
    .A(_0072_),
    .B(_2909_));
 sg13g2_nand2_1 _3732_ (.Y(_2920_),
    .A(_0072_),
    .B(_2889_));
 sg13g2_o21ai_1 _3733_ (.B1(net1142),
    .Y(_2921_),
    .A1(_2918_),
    .A2(_2920_));
 sg13g2_nand3_1 _3734_ (.B(_2919_),
    .C(_2921_),
    .A(_2849_),
    .Y(_2922_));
 sg13g2_nand4_1 _3735_ (.B(_2855_),
    .C(_2883_),
    .A(_2771_),
    .Y(_2923_),
    .D(_2886_));
 sg13g2_a22oi_1 _3736_ (.Y(_2924_),
    .B1(_2890_),
    .B2(_2893_),
    .A2(_2811_),
    .A1(net1182));
 sg13g2_and4_1 _3737_ (.A(_2861_),
    .B(_2885_),
    .C(_2888_),
    .D(_2924_),
    .X(_2925_));
 sg13g2_nor2b_1 _3738_ (.A(_2859_),
    .B_N(_2896_),
    .Y(_2926_));
 sg13g2_nand4_1 _3739_ (.B(_2922_),
    .C(_2925_),
    .A(_2875_),
    .Y(_2927_),
    .D(_2926_));
 sg13g2_nor4_1 _3740_ (.A(_2851_),
    .B(_2905_),
    .C(_2923_),
    .D(_2927_),
    .Y(_2928_));
 sg13g2_nor2b_2 _3741_ (.A(_2928_),
    .B_N(net1192),
    .Y(_2929_));
 sg13g2_inv_1 _3742_ (.Y(_2930_),
    .A(_2929_));
 sg13g2_and2_1 _3743_ (.A(net1251),
    .B(_2929_),
    .X(_2931_));
 sg13g2_nand2_1 _3744_ (.Y(_2932_),
    .A(_2844_),
    .B(_2931_));
 sg13g2_nand2_1 _3745_ (.Y(_2933_),
    .A(net596),
    .B(net1251));
 sg13g2_nor4_2 _3746_ (.A(_2657_),
    .B(_2668_),
    .C(_2723_),
    .Y(_2934_),
    .D(_2750_));
 sg13g2_a221oi_1 _3747_ (.B2(net1136),
    .C1(_2853_),
    .B1(net1130),
    .A1(net1135),
    .Y(_2935_),
    .A2(_2752_));
 sg13g2_or2_1 _3748_ (.X(_2936_),
    .B(_2822_),
    .A(_2763_));
 sg13g2_nor2_1 _3749_ (.A(_2755_),
    .B(_2810_),
    .Y(_2937_));
 sg13g2_nor4_2 _3750_ (.A(_2755_),
    .B(_2763_),
    .C(_2810_),
    .Y(_2938_),
    .D(_2822_));
 sg13g2_a22oi_1 _3751_ (.Y(_2939_),
    .B1(_2781_),
    .B2(net1135),
    .A2(_2764_),
    .A1(net1132));
 sg13g2_and2_1 _3752_ (.A(_2938_),
    .B(_2939_),
    .X(_2940_));
 sg13g2_nand2_1 _3753_ (.Y(_2941_),
    .A(_2938_),
    .B(_2939_));
 sg13g2_o21ai_1 _3754_ (.B1(_2887_),
    .Y(_2942_),
    .A1(_2742_),
    .A2(_2808_));
 sg13g2_nand3_1 _3755_ (.B(_2872_),
    .C(_2895_),
    .A(_2871_),
    .Y(_2943_));
 sg13g2_a21oi_1 _3756_ (.A1(_2775_),
    .A2(_2794_),
    .Y(_2944_),
    .B1(_2739_));
 sg13g2_nand3_1 _3757_ (.B(net1154),
    .C(_2732_),
    .A(_2710_),
    .Y(_2945_));
 sg13g2_nand2_1 _3758_ (.Y(_2946_),
    .A(_2867_),
    .B(_2945_));
 sg13g2_or4_1 _3759_ (.A(_2868_),
    .B(_2943_),
    .C(_2944_),
    .D(_2946_),
    .X(_2947_));
 sg13g2_nand2_1 _3760_ (.Y(_2948_),
    .A(net1155),
    .B(_2793_));
 sg13g2_nor3_1 _3761_ (.A(net1152),
    .B(_2727_),
    .C(net1144),
    .Y(_2949_));
 sg13g2_a21oi_1 _3762_ (.A1(net1156),
    .A2(_2819_),
    .Y(_2950_),
    .B1(_2949_));
 sg13g2_a22oi_1 _3763_ (.Y(_2951_),
    .B1(_2749_),
    .B2(net1130),
    .A2(_2740_),
    .A1(net1134));
 sg13g2_nand2b_1 _3764_ (.Y(_2952_),
    .B(net1222),
    .A_N(_2951_));
 sg13g2_o21ai_1 _3765_ (.B1(net1137),
    .Y(_2953_),
    .A1(_2764_),
    .A2(_2772_));
 sg13g2_a21oi_1 _3766_ (.A1(_2765_),
    .A2(_2773_),
    .Y(_2954_),
    .B1(_2706_));
 sg13g2_a21oi_2 _3767_ (.B1(_2782_),
    .Y(_2955_),
    .A2(_2793_),
    .A1(net1149));
 sg13g2_o21ai_1 _3768_ (.B1(net1155),
    .Y(_2956_),
    .A1(net1131),
    .A2(_2793_));
 sg13g2_o21ai_1 _3769_ (.B1(net1137),
    .Y(_2957_),
    .A1(_2749_),
    .A2(_2762_));
 sg13g2_nand4_1 _3770_ (.B(_2901_),
    .C(_2940_),
    .A(_2864_),
    .Y(_2958_),
    .D(_2955_));
 sg13g2_nand3_1 _3771_ (.B(_2952_),
    .C(_2953_),
    .A(_2950_),
    .Y(_2959_));
 sg13g2_nor2_1 _3772_ (.A(_2947_),
    .B(_2959_),
    .Y(_2960_));
 sg13g2_nand4_1 _3773_ (.B(_2935_),
    .C(_2956_),
    .A(_2858_),
    .Y(_2961_),
    .D(_2957_));
 sg13g2_nor4_1 _3774_ (.A(_2897_),
    .B(_2942_),
    .C(_2958_),
    .D(_2961_),
    .Y(_0374_));
 sg13g2_nand2_1 _3775_ (.Y(_0375_),
    .A(_2960_),
    .B(_0374_));
 sg13g2_a22oi_1 _3776_ (.Y(_0376_),
    .B1(net1134),
    .B2(_2740_),
    .A2(_2719_),
    .A1(_2669_));
 sg13g2_nand4_1 _3777_ (.B(_2804_),
    .C(_2805_),
    .A(_2788_),
    .Y(_0377_),
    .D(_2835_));
 sg13g2_or3_1 _3778_ (.A(net1099),
    .B(net1054),
    .C(_0377_),
    .X(_0378_));
 sg13g2_a21oi_1 _3779_ (.A1(net1137),
    .A2(net1131),
    .Y(_0379_),
    .B1(_2779_));
 sg13g2_o21ai_1 _3780_ (.B1(_0379_),
    .Y(_0380_),
    .A1(net1153),
    .A2(_2775_));
 sg13g2_o21ai_1 _3781_ (.B1(_2809_),
    .Y(_0381_),
    .A1(_2731_),
    .A2(_2773_));
 sg13g2_a221oi_1 _3782_ (.B2(_2720_),
    .C1(_0381_),
    .B1(_2759_),
    .A1(net1132),
    .Y(_0382_),
    .A2(net1131));
 sg13g2_nor2_1 _3783_ (.A(_2754_),
    .B(_2832_),
    .Y(_0383_));
 sg13g2_o21ai_1 _3784_ (.B1(_2726_),
    .Y(_0384_),
    .A1(_2754_),
    .A2(_2832_));
 sg13g2_a22oi_1 _3785_ (.Y(_0385_),
    .B1(_2752_),
    .B2(net1155),
    .A2(_2741_),
    .A1(net1133));
 sg13g2_nand4_1 _3786_ (.B(_0382_),
    .C(_0384_),
    .A(_2886_),
    .Y(_0386_),
    .D(_0385_));
 sg13g2_or2_1 _3787_ (.X(_0387_),
    .B(_0386_),
    .A(_0380_));
 sg13g2_a22oi_1 _3788_ (.Y(_0388_),
    .B1(net1130),
    .B2(_2793_),
    .A2(_2752_),
    .A1(net1132));
 sg13g2_a22oi_1 _3789_ (.Y(_0389_),
    .B1(_2766_),
    .B2(net1132),
    .A2(_2762_),
    .A1(net1134));
 sg13g2_o21ai_1 _3790_ (.B1(_2831_),
    .Y(_0390_),
    .A1(_2739_),
    .A2(_2767_));
 sg13g2_a22oi_1 _3791_ (.Y(_0391_),
    .B1(net1131),
    .B2(net1130),
    .A2(net1134),
    .A1(_2720_));
 sg13g2_a221oi_1 _3792_ (.B2(net1139),
    .C1(_2790_),
    .B1(_2745_),
    .A1(net1136),
    .Y(_0392_),
    .A2(net1154));
 sg13g2_nand4_1 _3793_ (.B(_0389_),
    .C(_0391_),
    .A(_0388_),
    .Y(_0393_),
    .D(_0392_));
 sg13g2_a21oi_2 _3794_ (.B1(net1148),
    .Y(_0394_),
    .A2(_2773_),
    .A1(_2758_));
 sg13g2_nor2_1 _3795_ (.A(net1144),
    .B(_2775_),
    .Y(_0395_));
 sg13g2_or4_1 _3796_ (.A(_2803_),
    .B(_2811_),
    .C(_0393_),
    .D(_0395_),
    .X(_0396_));
 sg13g2_nor4_1 _3797_ (.A(_2836_),
    .B(_0387_),
    .C(_0394_),
    .D(_0396_),
    .Y(_0397_));
 sg13g2_nor2b_1 _3798_ (.A(_0378_),
    .B_N(_0397_),
    .Y(_0398_));
 sg13g2_or2_1 _3799_ (.X(_0399_),
    .B(_0398_),
    .A(_0375_));
 sg13g2_xnor2_1 _3800_ (.Y(_0400_),
    .A(net1165),
    .B(\dtop.player_inst.synth.alu.acc[9] ));
 sg13g2_a22oi_1 _3801_ (.Y(_0401_),
    .B1(_0400_),
    .B2(_0380_),
    .A2(_0399_),
    .A1(net1165));
 sg13g2_o21ai_1 _3802_ (.B1(net1248),
    .Y(_0402_),
    .A1(net1099),
    .A2(_2811_));
 sg13g2_nor2b_1 _3803_ (.A(_0070_),
    .B_N(net1141),
    .Y(_0403_));
 sg13g2_nor4_2 _3804_ (.A(_0070_),
    .B(_2906_),
    .C(_2909_),
    .Y(_0404_),
    .D(_2915_));
 sg13g2_nand3_1 _3805_ (.B(_2916_),
    .C(_0403_),
    .A(_2907_),
    .Y(_0405_));
 sg13g2_and4_1 _3806_ (.A(net1232),
    .B(_2907_),
    .C(_2916_),
    .D(_0403_),
    .X(_0406_));
 sg13g2_nand4_1 _3807_ (.B(_2907_),
    .C(_2916_),
    .A(net1232),
    .Y(_0407_),
    .D(_0403_));
 sg13g2_nand2_1 _3808_ (.Y(_0408_),
    .A(_2848_),
    .B(_0406_));
 sg13g2_o21ai_1 _3809_ (.B1(_0402_),
    .Y(_0409_),
    .A1(_2939_),
    .A2(_0408_));
 sg13g2_inv_2 _3810_ (.Y(_0410_),
    .A(_0409_));
 sg13g2_nand3_1 _3811_ (.B(_2812_),
    .C(_2945_),
    .A(_2801_),
    .Y(_0411_));
 sg13g2_nor3_1 _3812_ (.A(_2825_),
    .B(_2894_),
    .C(_0411_),
    .Y(_0412_));
 sg13g2_o21ai_1 _3813_ (.B1(net1130),
    .Y(_0413_),
    .A1(net1136),
    .A2(_2774_));
 sg13g2_inv_1 _3814_ (.Y(_0414_),
    .A(_0413_));
 sg13g2_and4_1 _3815_ (.A(_2777_),
    .B(_2861_),
    .C(_0412_),
    .D(_0413_),
    .X(_0415_));
 sg13g2_nor2_1 _3816_ (.A(_2811_),
    .B(_2832_),
    .Y(_0416_));
 sg13g2_o21ai_1 _3817_ (.B1(net1132),
    .Y(_0417_),
    .A1(_2741_),
    .A2(_2774_));
 sg13g2_nand3_1 _3818_ (.B(_0416_),
    .C(_0417_),
    .A(_2855_),
    .Y(_0418_));
 sg13g2_nor3_1 _3819_ (.A(net1217),
    .B(net1159),
    .C(net1143),
    .Y(_0419_));
 sg13g2_nor2_1 _3820_ (.A(_2826_),
    .B(_0419_),
    .Y(_0420_));
 sg13g2_a221oi_1 _3821_ (.B2(_2707_),
    .C1(_2934_),
    .B1(net1133),
    .A1(net1212),
    .Y(_0421_),
    .A2(net1154));
 sg13g2_nand4_1 _3822_ (.B(_2950_),
    .C(_0420_),
    .A(_2817_),
    .Y(_0422_),
    .D(_0421_));
 sg13g2_nand4_1 _3823_ (.B(_2735_),
    .C(_2809_),
    .A(_2704_),
    .Y(_0423_),
    .D(_2951_));
 sg13g2_nor4_2 _3824_ (.A(_2859_),
    .B(_0418_),
    .C(_0422_),
    .Y(_0424_),
    .D(_0423_));
 sg13g2_and2_1 _3825_ (.A(_0415_),
    .B(_0424_),
    .X(_0425_));
 sg13g2_nor3_1 _3826_ (.A(net1156),
    .B(_2733_),
    .C(net1144),
    .Y(_0426_));
 sg13g2_a221oi_1 _3827_ (.B2(net1150),
    .C1(_2786_),
    .B1(_2776_),
    .A1(net1138),
    .Y(_0427_),
    .A2(_2734_));
 sg13g2_a21o_1 _3828_ (.A2(_2785_),
    .A1(_2742_),
    .B1(_2731_),
    .X(_0428_));
 sg13g2_nand2_1 _3829_ (.Y(_0429_),
    .A(net1217),
    .B(_2719_));
 sg13g2_nor4_1 _3830_ (.A(_2657_),
    .B(net1151),
    .C(_2723_),
    .D(_2824_),
    .Y(_0430_));
 sg13g2_or3_2 _3831_ (.A(_2856_),
    .B(_2857_),
    .C(_0430_),
    .X(_0431_));
 sg13g2_or2_1 _3832_ (.X(_0432_),
    .B(_2949_),
    .A(_2934_));
 sg13g2_a221oi_1 _3833_ (.B2(_2703_),
    .C1(_2790_),
    .B1(_2745_),
    .A1(net1136),
    .Y(_0433_),
    .A2(net1154));
 sg13g2_nand2_1 _3834_ (.Y(_0434_),
    .A(_2938_),
    .B(_0433_));
 sg13g2_nand3_1 _3835_ (.B(_2948_),
    .C(_0388_),
    .A(_2834_),
    .Y(_0435_));
 sg13g2_nor3_1 _3836_ (.A(_2769_),
    .B(_0434_),
    .C(_0435_),
    .Y(_0436_));
 sg13g2_or4_1 _3837_ (.A(_2954_),
    .B(_0377_),
    .C(_0390_),
    .D(_0431_),
    .X(_0437_));
 sg13g2_nor4_1 _3838_ (.A(_2754_),
    .B(_2782_),
    .C(_2826_),
    .D(_2827_),
    .Y(_0438_));
 sg13g2_nor4_1 _3839_ (.A(_2813_),
    .B(_2934_),
    .C(_2949_),
    .D(_0426_),
    .Y(_0439_));
 sg13g2_nand4_1 _3840_ (.B(_2899_),
    .C(_0438_),
    .A(_2817_),
    .Y(_0440_),
    .D(_0439_));
 sg13g2_a221oi_1 _3841_ (.B2(net1150),
    .C1(_2845_),
    .B1(_2772_),
    .A1(net1139),
    .Y(_0441_),
    .A2(_2766_));
 sg13g2_nand4_1 _3842_ (.B(_0428_),
    .C(_0429_),
    .A(_0427_),
    .Y(_0442_),
    .D(_0441_));
 sg13g2_nor4_1 _3843_ (.A(_0418_),
    .B(_0437_),
    .C(_0440_),
    .D(_0442_),
    .Y(_0443_));
 sg13g2_nand4_1 _3844_ (.B(_0415_),
    .C(_0436_),
    .A(_2875_),
    .Y(_0444_),
    .D(_0443_));
 sg13g2_a21o_2 _3845_ (.A2(_0444_),
    .A1(_2823_),
    .B1(_0425_),
    .X(_0445_));
 sg13g2_a22oi_1 _3846_ (.Y(_0446_),
    .B1(net1131),
    .B2(net1137),
    .A2(net1133),
    .A1(_2734_));
 sg13g2_nand3_1 _3847_ (.B(_2815_),
    .C(_0446_),
    .A(_2746_),
    .Y(_0447_));
 sg13g2_a21oi_1 _3848_ (.A1(_2792_),
    .A2(_0383_),
    .Y(_0448_),
    .B1(_2710_));
 sg13g2_nand3_1 _3849_ (.B(_0420_),
    .C(_0427_),
    .A(_2777_),
    .Y(_0449_));
 sg13g2_nor3_2 _3850_ (.A(_0447_),
    .B(_0448_),
    .C(_0449_),
    .Y(_0450_));
 sg13g2_nor2b_1 _3851_ (.A(_2780_),
    .B_N(_0450_),
    .Y(_0451_));
 sg13g2_nand2_1 _3852_ (.Y(_0452_),
    .A(_0445_),
    .B(_0451_));
 sg13g2_nand4_1 _3853_ (.B(_2805_),
    .C(_2902_),
    .A(_2804_),
    .Y(_0453_),
    .D(_0376_));
 sg13g2_nor2_2 _3854_ (.A(_2941_),
    .B(_0393_),
    .Y(_0454_));
 sg13g2_inv_2 _3855_ (.Y(_0455_),
    .A(net1072));
 sg13g2_o21ai_1 _3856_ (.B1(_2809_),
    .Y(_0456_),
    .A1(net1144),
    .A2(_2778_));
 sg13g2_nor3_1 _3857_ (.A(_2811_),
    .B(_2816_),
    .C(_0456_),
    .Y(_0457_));
 sg13g2_or2_1 _3858_ (.X(_0458_),
    .B(_2728_),
    .A(net1136));
 sg13g2_a221oi_1 _3859_ (.B2(net1132),
    .C1(_2813_),
    .B1(_0458_),
    .A1(_2734_),
    .Y(_0459_),
    .A2(_2759_));
 sg13g2_nand3_1 _3860_ (.B(_0457_),
    .C(_0459_),
    .A(_2862_),
    .Y(_0460_));
 sg13g2_nor3_1 _3861_ (.A(_0453_),
    .B(_0455_),
    .C(_0460_),
    .Y(_0461_));
 sg13g2_nand3_1 _3862_ (.B(_0451_),
    .C(_0461_),
    .A(_0445_),
    .Y(_0462_));
 sg13g2_nand3_1 _3863_ (.B(net1139),
    .C(_2743_),
    .A(net1210),
    .Y(_0463_));
 sg13g2_nor3_2 _3864_ (.A(_2670_),
    .B(_2706_),
    .C(net1147),
    .Y(_0464_));
 sg13g2_and4_1 _3865_ (.A(_2862_),
    .B(_0457_),
    .C(_0459_),
    .D(_0463_),
    .X(_0465_));
 sg13g2_nand2_1 _3866_ (.Y(_0466_),
    .A(_0450_),
    .B(_0465_));
 sg13g2_a221oi_1 _3867_ (.B2(_2728_),
    .C1(_2863_),
    .B1(net1130),
    .A1(net1137),
    .Y(_0467_),
    .A2(_2752_));
 sg13g2_nand2b_1 _3868_ (.Y(_0468_),
    .B(_0467_),
    .A_N(_0431_));
 sg13g2_nor4_2 _3869_ (.A(_2897_),
    .B(_2942_),
    .C(_2947_),
    .Y(_0469_),
    .D(_0468_));
 sg13g2_nand2_1 _3870_ (.Y(_0470_),
    .A(_2820_),
    .B(_2955_));
 sg13g2_nor4_2 _3871_ (.A(_2836_),
    .B(_2898_),
    .C(_0394_),
    .Y(_0471_),
    .D(_0470_));
 sg13g2_nor2_1 _3872_ (.A(_2731_),
    .B(_2767_),
    .Y(_0472_));
 sg13g2_nor3_1 _3873_ (.A(_2721_),
    .B(_2934_),
    .C(_0472_),
    .Y(_0473_));
 sg13g2_nand3_1 _3874_ (.B(_2801_),
    .C(_2854_),
    .A(_2714_),
    .Y(_0474_));
 sg13g2_nor2_1 _3875_ (.A(_0414_),
    .B(_0474_),
    .Y(_0475_));
 sg13g2_nand4_1 _3876_ (.B(_0471_),
    .C(_0473_),
    .A(_0469_),
    .Y(_0476_),
    .D(_0475_));
 sg13g2_nor4_2 _3877_ (.A(_0453_),
    .B(net1062),
    .C(_0466_),
    .Y(_0477_),
    .D(_0476_));
 sg13g2_nand2_2 _3878_ (.Y(_0478_),
    .A(_0445_),
    .B(_0477_));
 sg13g2_nand2b_1 _3879_ (.Y(_0479_),
    .B(_0478_),
    .A_N(_0462_));
 sg13g2_nor2_1 _3880_ (.A(net1098),
    .B(_0470_),
    .Y(_0480_));
 sg13g2_nand3_1 _3881_ (.B(_0465_),
    .C(_0480_),
    .A(_0450_),
    .Y(_0481_));
 sg13g2_a21o_2 _3882_ (.A2(net1131),
    .A1(net1149),
    .B1(_2800_),
    .X(_0482_));
 sg13g2_nor3_2 _3883_ (.A(_2721_),
    .B(_0481_),
    .C(_0482_),
    .Y(_0483_));
 sg13g2_or3_1 _3884_ (.A(_2721_),
    .B(_0481_),
    .C(_0482_),
    .X(_0484_));
 sg13g2_nand2_1 _3885_ (.Y(_0485_),
    .A(_0478_),
    .B(_0483_));
 sg13g2_nand2_2 _3886_ (.Y(_0486_),
    .A(_0450_),
    .B(_0471_));
 sg13g2_nand3_1 _3887_ (.B(_2729_),
    .C(_0480_),
    .A(_2714_),
    .Y(_0487_));
 sg13g2_nor4_2 _3888_ (.A(_0479_),
    .B(_0485_),
    .C(_0486_),
    .Y(_0488_),
    .D(_0487_));
 sg13g2_a221oi_1 _3889_ (.B2(_0445_),
    .C1(_0484_),
    .B1(_0477_),
    .A1(_0450_),
    .Y(_0489_),
    .A2(_0471_));
 sg13g2_nor2_1 _3890_ (.A(_0452_),
    .B(_0487_),
    .Y(_0490_));
 sg13g2_nor2_1 _3891_ (.A(_0037_),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_nand3_1 _3892_ (.B(_0489_),
    .C(_0491_),
    .A(_0479_),
    .Y(_0492_));
 sg13g2_nor2_1 _3893_ (.A(_2772_),
    .B(_0481_),
    .Y(_0493_));
 sg13g2_and2_1 _3894_ (.A(_0462_),
    .B(_0493_),
    .X(_0494_));
 sg13g2_nand2_1 _3895_ (.Y(_0495_),
    .A(_0462_),
    .B(_0493_));
 sg13g2_a221oi_1 _3896_ (.B2(\dtop.player_inst.synth.alu.registers[0][10] ),
    .C1(_0494_),
    .B1(_0488_),
    .A1(\dtop.player_inst.synth.alu.registers[1][10] ),
    .Y(_0496_),
    .A2(_0464_));
 sg13g2_nand4_1 _3897_ (.B(_2940_),
    .C(net1118),
    .A(_2848_),
    .Y(_0497_),
    .D(_0425_));
 sg13g2_nor2_2 _3898_ (.A(net1232),
    .B(_0405_),
    .Y(_0498_));
 sg13g2_nand2_1 _3899_ (.Y(_0499_),
    .A(_2661_),
    .B(_0404_));
 sg13g2_nand3_1 _3900_ (.B(_0390_),
    .C(_0498_),
    .A(_2848_),
    .Y(_0500_));
 sg13g2_and3_2 _3901_ (.X(_0501_),
    .A(_0445_),
    .B(_0497_),
    .C(_0500_));
 sg13g2_nand3_1 _3902_ (.B(_0497_),
    .C(_0500_),
    .A(_0445_),
    .Y(_0502_));
 sg13g2_a21oi_1 _3903_ (.A1(_0436_),
    .A2(_0444_),
    .Y(_0503_),
    .B1(_0425_));
 sg13g2_nand3_1 _3904_ (.B(_0415_),
    .C(_0424_),
    .A(_2848_),
    .Y(_0504_));
 sg13g2_nor3_1 _3905_ (.A(net1232),
    .B(_0390_),
    .C(_0405_),
    .Y(_0505_));
 sg13g2_a21oi_1 _3906_ (.A1(_2937_),
    .A2(_0405_),
    .Y(_0506_),
    .B1(_0505_));
 sg13g2_o21ai_1 _3907_ (.B1(_0506_),
    .Y(_0507_),
    .A1(_2938_),
    .A2(_0407_));
 sg13g2_nand2b_1 _3908_ (.Y(_0508_),
    .B(_0507_),
    .A_N(_0504_));
 sg13g2_nand2b_2 _3909_ (.Y(_0509_),
    .B(_0508_),
    .A_N(_0503_));
 sg13g2_or3_1 _3910_ (.A(_2954_),
    .B(_0390_),
    .C(_0434_),
    .X(_0510_));
 sg13g2_a21o_1 _3911_ (.A2(_0424_),
    .A1(_0415_),
    .B1(_0510_),
    .X(_0511_));
 sg13g2_nand2_2 _3912_ (.Y(_0512_),
    .A(net1232),
    .B(net1142));
 sg13g2_nor2_2 _3913_ (.A(_0404_),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_nand2b_1 _3914_ (.Y(_0514_),
    .B(_0405_),
    .A_N(_0512_));
 sg13g2_o21ai_1 _3915_ (.B1(_2938_),
    .Y(_0515_),
    .A1(_0505_),
    .A2(_0513_));
 sg13g2_nand3_1 _3916_ (.B(_0388_),
    .C(_0389_),
    .A(_2938_),
    .Y(_0516_));
 sg13g2_and2_2 _3917_ (.A(_0405_),
    .B(_0512_),
    .X(_0517_));
 sg13g2_nand2_1 _3918_ (.Y(_0518_),
    .A(_0405_),
    .B(_0512_));
 sg13g2_nand2_1 _3919_ (.Y(_0519_),
    .A(_2936_),
    .B(net1118));
 sg13g2_nand3b_1 _3920_ (.B(_0516_),
    .C(_0517_),
    .Y(_0520_),
    .A_N(_2936_));
 sg13g2_nand3_1 _3921_ (.B(_0519_),
    .C(_0520_),
    .A(_0515_),
    .Y(_0521_));
 sg13g2_o21ai_1 _3922_ (.B1(_0511_),
    .Y(_0522_),
    .A1(_0504_),
    .A2(_0521_));
 sg13g2_mux2_1 _3923_ (.A0(\dtop.player_inst.synth.alu.registers[4][3] ),
    .A1(\dtop.detune_counter[10] ),
    .S(net1074),
    .X(_0523_));
 sg13g2_nor2_1 _3924_ (.A(_2661_),
    .B(net1062),
    .Y(_0524_));
 sg13g2_a21oi_1 _3925_ (.A1(\dtop.player_inst.synth.alu.registers[4][4] ),
    .A2(net1062),
    .Y(_0525_),
    .B1(_0524_));
 sg13g2_nor2_1 _3926_ (.A(net1053),
    .B(_0523_),
    .Y(_0526_));
 sg13g2_a21oi_1 _3927_ (.A1(net1052),
    .A2(_0525_),
    .Y(_0527_),
    .B1(_0526_));
 sg13g2_nor2b_1 _3928_ (.A(_0454_),
    .B_N(_0044_),
    .Y(_0528_));
 sg13g2_a21oi_1 _3929_ (.A1(_0087_),
    .A2(net1074),
    .Y(_0529_),
    .B1(_0528_));
 sg13g2_nand2_1 _3930_ (.Y(_0530_),
    .A(net1052),
    .B(_0529_));
 sg13g2_nor2_1 _3931_ (.A(_2659_),
    .B(net1062),
    .Y(_0531_));
 sg13g2_a21oi_1 _3932_ (.A1(\dtop.player_inst.synth.alu.registers[4][5] ),
    .A2(net1062),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_o21ai_1 _3933_ (.B1(_0530_),
    .Y(_0533_),
    .A1(net1052),
    .A2(_0532_));
 sg13g2_mux2_1 _3934_ (.A0(_0533_),
    .A1(_0527_),
    .S(net1035),
    .X(_0534_));
 sg13g2_nor2_2 _3935_ (.A(net1036),
    .B(net1053),
    .Y(_0535_));
 sg13g2_mux2_1 _3936_ (.A0(_0047_),
    .A1(_0058_),
    .S(net1074),
    .X(_0536_));
 sg13g2_nor2b_2 _3937_ (.A(net1036),
    .B_N(net1053),
    .Y(_0537_));
 sg13g2_mux2_1 _3938_ (.A0(_0048_),
    .A1(_0057_),
    .S(net1074),
    .X(_0538_));
 sg13g2_mux2_1 _3939_ (.A0(_0046_),
    .A1(_0000_),
    .S(net1074),
    .X(_0539_));
 sg13g2_nor2_1 _3940_ (.A(_0045_),
    .B(_0454_),
    .Y(_0540_));
 sg13g2_a21oi_1 _3941_ (.A1(_2681_),
    .A2(net1074),
    .Y(_0541_),
    .B1(_0540_));
 sg13g2_mux2_1 _3942_ (.A0(_0541_),
    .A1(_0539_),
    .S(_0522_),
    .X(_0542_));
 sg13g2_a22oi_1 _3943_ (.Y(_0543_),
    .B1(_0537_),
    .B2(_0538_),
    .A2(_0536_),
    .A1(_0535_));
 sg13g2_a21oi_1 _3944_ (.A1(net1036),
    .A2(_0542_),
    .Y(_0544_),
    .B1(net1038));
 sg13g2_a22oi_1 _3945_ (.Y(_0545_),
    .B1(_0543_),
    .B2(_0544_),
    .A2(_0534_),
    .A1(net1037));
 sg13g2_a22oi_1 _3946_ (.Y(_0546_),
    .B1(_0545_),
    .B2(_0494_),
    .A2(_0496_),
    .A1(_0492_));
 sg13g2_xnor2_1 _3947_ (.Y(_0547_),
    .A(_0409_),
    .B(_0546_));
 sg13g2_nor2_1 _3948_ (.A(_0401_),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_xor2_1 _3949_ (.B(_0547_),
    .A(_0401_),
    .X(_0549_));
 sg13g2_xor2_1 _3950_ (.B(\dtop.player_inst.synth.alu.acc[8] ),
    .A(net1165),
    .X(_0550_));
 sg13g2_a22oi_1 _3951_ (.Y(_0551_),
    .B1(_0380_),
    .B2(_0550_),
    .A2(net1100),
    .A1(\dtop.player_inst.synth.alu.acc[1] ));
 sg13g2_a22oi_1 _3952_ (.Y(_0552_),
    .B1(_0398_),
    .B2(net1165),
    .A2(net1054),
    .A1(\dtop.player_inst.synth.alu.acc[9] ));
 sg13g2_nand2_1 _3953_ (.Y(_0553_),
    .A(_0551_),
    .B(_0552_));
 sg13g2_nor2_2 _3954_ (.A(_0483_),
    .B(_0486_),
    .Y(_0554_));
 sg13g2_nor2_1 _3955_ (.A(_0489_),
    .B(_0554_),
    .Y(_0555_));
 sg13g2_nor2_1 _3956_ (.A(\dtop.detune_counter[14] ),
    .B(net1230),
    .Y(_0556_));
 sg13g2_or2_2 _3957_ (.X(_0557_),
    .B(_0556_),
    .A(net1141));
 sg13g2_nor2_1 _3958_ (.A(\dtop.detune_counter[12] ),
    .B(net1231),
    .Y(_0558_));
 sg13g2_nor2_1 _3959_ (.A(\dtop.detune_counter[10] ),
    .B(\dtop.detune_counter[9] ),
    .Y(_0559_));
 sg13g2_or2_1 _3960_ (.X(_0560_),
    .B(\dtop.detune_counter[9] ),
    .A(\dtop.detune_counter[10] ));
 sg13g2_nor2_1 _3961_ (.A(net1234),
    .B(_0560_),
    .Y(_0561_));
 sg13g2_o21ai_1 _3962_ (.B1(_0561_),
    .Y(_0562_),
    .A1(net1141),
    .A2(_0558_));
 sg13g2_nand2_1 _3963_ (.Y(_0563_),
    .A(_0557_),
    .B(_0562_));
 sg13g2_inv_1 _3964_ (.Y(_0564_),
    .A(_0563_));
 sg13g2_nor3_2 _3965_ (.A(_0489_),
    .B(_0554_),
    .C(_0563_),
    .Y(_0565_));
 sg13g2_o21ai_1 _3966_ (.B1(_0518_),
    .Y(_0566_),
    .A1(_2848_),
    .A2(_0407_));
 sg13g2_a21oi_1 _3967_ (.A1(_0070_),
    .A2(_0556_),
    .Y(_0567_),
    .B1(net1141));
 sg13g2_a21oi_2 _3968_ (.B1(_0567_),
    .Y(_0568_),
    .A2(net1119),
    .A1(_2658_));
 sg13g2_and2_1 _3969_ (.A(_0489_),
    .B(_0568_),
    .X(_0569_));
 sg13g2_nand2_1 _3970_ (.Y(_0570_),
    .A(net1119),
    .B(net1118));
 sg13g2_nand4_1 _3971_ (.B(_2907_),
    .C(_2912_),
    .A(_2889_),
    .Y(_0571_),
    .D(_2916_));
 sg13g2_or2_1 _3972_ (.X(_0572_),
    .B(net1237),
    .A(net1234));
 sg13g2_a21oi_1 _3973_ (.A1(_0407_),
    .A2(_0572_),
    .Y(_0573_),
    .B1(_0571_));
 sg13g2_nor4_1 _3974_ (.A(net1233),
    .B(_0075_),
    .C(_2684_),
    .D(_2909_),
    .Y(_0574_));
 sg13g2_o21ai_1 _3975_ (.B1(_0570_),
    .Y(_0575_),
    .A1(_0573_),
    .A2(_0574_));
 sg13g2_or4_1 _3976_ (.A(_2891_),
    .B(_2906_),
    .C(_2915_),
    .D(_0512_),
    .X(_0576_));
 sg13g2_inv_1 _3977_ (.Y(_0577_),
    .A(_0576_));
 sg13g2_nor4_2 _3978_ (.A(net1233),
    .B(_0075_),
    .C(_0078_),
    .Y(_0578_),
    .D(_2909_));
 sg13g2_o21ai_1 _3979_ (.B1(_0075_),
    .Y(_0579_),
    .A1(net1233),
    .A2(_0078_));
 sg13g2_a21oi_1 _3980_ (.A1(net1233),
    .A2(_0078_),
    .Y(_0580_),
    .B1(_0579_));
 sg13g2_a22oi_1 _3981_ (.Y(_0581_),
    .B1(_0580_),
    .B2(net1141),
    .A2(_0578_),
    .A1(_0577_));
 sg13g2_nor3_1 _3982_ (.A(_0518_),
    .B(_0571_),
    .C(_0572_),
    .Y(_0582_));
 sg13g2_a21oi_2 _3983_ (.B1(_0582_),
    .Y(_0583_),
    .A2(_0581_),
    .A1(_0575_));
 sg13g2_a21o_1 _3984_ (.A2(_0581_),
    .A1(_0575_),
    .B1(_0582_),
    .X(_0584_));
 sg13g2_a21o_1 _3985_ (.A2(_0078_),
    .A1(net1233),
    .B1(_0075_),
    .X(_0585_));
 sg13g2_nand3_1 _3986_ (.B(_0579_),
    .C(_0585_),
    .A(net1141),
    .Y(_0586_));
 sg13g2_a22oi_1 _3987_ (.Y(_0587_),
    .B1(_0576_),
    .B2(_0578_),
    .A2(_0574_),
    .A1(_2918_));
 sg13g2_a21o_1 _3988_ (.A2(_0587_),
    .A1(_0586_),
    .B1(_0573_),
    .X(_0588_));
 sg13g2_nand4_1 _3989_ (.B(_2889_),
    .C(_2918_),
    .A(_2684_),
    .Y(_0589_),
    .D(net1118));
 sg13g2_and2_1 _3990_ (.A(_0588_),
    .B(_0589_),
    .X(_0590_));
 sg13g2_nand2_2 _3991_ (.Y(_0591_),
    .A(_0588_),
    .B(_0589_));
 sg13g2_nor2_1 _3992_ (.A(_0584_),
    .B(_0591_),
    .Y(_0592_));
 sg13g2_nand2_1 _3993_ (.Y(_0593_),
    .A(_0583_),
    .B(_0590_));
 sg13g2_a21oi_1 _3994_ (.A1(_0512_),
    .A2(_0588_),
    .Y(_0594_),
    .B1(net1118));
 sg13g2_a22oi_1 _3995_ (.Y(_0595_),
    .B1(_0593_),
    .B2(_0594_),
    .A2(_0583_),
    .A1(_0404_));
 sg13g2_nor3_2 _3996_ (.A(net1228),
    .B(net1227),
    .C(\dtop.detune_counter[17] ),
    .Y(_0596_));
 sg13g2_and2_1 _3997_ (.A(_2658_),
    .B(_0596_),
    .X(_0597_));
 sg13g2_nand2_2 _3998_ (.Y(_0598_),
    .A(_2658_),
    .B(_0596_));
 sg13g2_nor2_2 _3999_ (.A(_2889_),
    .B(_0559_),
    .Y(_0599_));
 sg13g2_nand2b_1 _4000_ (.Y(_0600_),
    .B(net1237),
    .A_N(net1234));
 sg13g2_nand2b_2 _4001_ (.Y(_0601_),
    .B(net1235),
    .A_N(net1237));
 sg13g2_mux2_1 _4002_ (.A0(_0600_),
    .A1(_0601_),
    .S(_0599_),
    .X(_0602_));
 sg13g2_a21oi_2 _4003_ (.B1(net1236),
    .Y(_0603_),
    .A2(_0599_),
    .A1(net1234));
 sg13g2_o21ai_1 _4004_ (.B1(_0597_),
    .Y(_0604_),
    .A1(_0407_),
    .A2(_0602_));
 sg13g2_a21o_1 _4005_ (.A2(_0603_),
    .A1(_0407_),
    .B1(_0604_),
    .X(_0605_));
 sg13g2_nand2_1 _4006_ (.Y(_0606_),
    .A(\dtop.detune_counter[10] ),
    .B(_2662_));
 sg13g2_a21oi_1 _4007_ (.A1(net1237),
    .A2(_0606_),
    .Y(_0607_),
    .B1(net1234));
 sg13g2_a22oi_1 _4008_ (.Y(_0608_),
    .B1(_0560_),
    .B2(net1234),
    .A2(net1237),
    .A1(_2662_));
 sg13g2_inv_1 _4009_ (.Y(_0609_),
    .A(_0608_));
 sg13g2_a21oi_1 _4010_ (.A1(_2878_),
    .A2(_0609_),
    .Y(_0610_),
    .B1(net1118));
 sg13g2_o21ai_1 _4011_ (.B1(_0610_),
    .Y(_0611_),
    .A1(_2878_),
    .A2(_0607_));
 sg13g2_nand2_1 _4012_ (.Y(_0612_),
    .A(_2877_),
    .B(_0601_));
 sg13g2_mux2_1 _4013_ (.A0(_0600_),
    .A1(_0601_),
    .S(_0560_),
    .X(_0613_));
 sg13g2_nand2_1 _4014_ (.Y(_0614_),
    .A(_2878_),
    .B(_0613_));
 sg13g2_nand3_1 _4015_ (.B(_0612_),
    .C(_0614_),
    .A(net1118),
    .Y(_0615_));
 sg13g2_nand3_1 _4016_ (.B(_0611_),
    .C(_0615_),
    .A(_0598_),
    .Y(_0616_));
 sg13g2_and3_1 _4017_ (.X(_0617_),
    .A(_0554_),
    .B(_0605_),
    .C(_0616_));
 sg13g2_a221oi_1 _4018_ (.B2(_0595_),
    .C1(_0617_),
    .B1(_0569_),
    .A1(_0565_),
    .Y(_0618_),
    .A2(_0566_));
 sg13g2_xnor2_1 _4019_ (.Y(_0619_),
    .A(_2914_),
    .B(_0618_));
 sg13g2_xnor2_1 _4020_ (.Y(_0620_),
    .A(_2913_),
    .B(_0618_));
 sg13g2_nand2b_1 _4021_ (.Y(_0621_),
    .B(_2917_),
    .A_N(_0606_));
 sg13g2_nor2_1 _4022_ (.A(_0593_),
    .B(_0621_),
    .Y(_0622_));
 sg13g2_nor2_1 _4023_ (.A(_0583_),
    .B(_0591_),
    .Y(_0623_));
 sg13g2_a221oi_1 _4024_ (.B2(_2917_),
    .C1(_0514_),
    .B1(_0623_),
    .A1(_0592_),
    .Y(_0624_),
    .A2(_0621_));
 sg13g2_a21oi_1 _4025_ (.A1(_0584_),
    .A2(_0591_),
    .Y(_0625_),
    .B1(_0499_));
 sg13g2_o21ai_1 _4026_ (.B1(_0498_),
    .Y(_0626_),
    .A1(_0583_),
    .A2(_0590_));
 sg13g2_a21oi_1 _4027_ (.A1(_0407_),
    .A2(_0626_),
    .Y(_0627_),
    .B1(_0592_));
 sg13g2_or3_1 _4028_ (.A(_0517_),
    .B(_0624_),
    .C(_0627_),
    .X(_0628_));
 sg13g2_nand2_1 _4029_ (.Y(_0629_),
    .A(_0583_),
    .B(_0591_));
 sg13g2_nand3_1 _4030_ (.B(_0583_),
    .C(_0591_),
    .A(_0517_),
    .Y(_0630_));
 sg13g2_and3_1 _4031_ (.X(_0631_),
    .A(_0489_),
    .B(_0568_),
    .C(_0630_));
 sg13g2_a21oi_1 _4032_ (.A1(_0512_),
    .A2(_0608_),
    .Y(_0632_),
    .B1(_2877_));
 sg13g2_o21ai_1 _4033_ (.B1(_0632_),
    .Y(_0633_),
    .A1(_0498_),
    .A2(_0613_));
 sg13g2_a21oi_1 _4034_ (.A1(_2909_),
    .A2(_0607_),
    .Y(_0634_),
    .B1(_2878_));
 sg13g2_nand2_1 _4035_ (.Y(_0635_),
    .A(_0601_),
    .B(_0634_));
 sg13g2_a21oi_1 _4036_ (.A1(_0633_),
    .A2(_0635_),
    .Y(_0636_),
    .B1(_0597_));
 sg13g2_nor2_1 _4037_ (.A(_0498_),
    .B(_0602_),
    .Y(_0637_));
 sg13g2_a21o_1 _4038_ (.A2(_0603_),
    .A1(_0512_),
    .B1(_0598_),
    .X(_0638_));
 sg13g2_nor2_1 _4039_ (.A(_0637_),
    .B(_0638_),
    .Y(_0639_));
 sg13g2_nor4_1 _4040_ (.A(_0483_),
    .B(_0486_),
    .C(_0636_),
    .D(_0639_),
    .Y(_0640_));
 sg13g2_o21ai_1 _4041_ (.B1(_0404_),
    .Y(_0641_),
    .A1(_2661_),
    .A2(_2848_));
 sg13g2_a221oi_1 _4042_ (.B2(_0565_),
    .C1(_0640_),
    .B1(_0641_),
    .A1(_0628_),
    .Y(_0642_),
    .A2(_0631_));
 sg13g2_nor3_1 _4043_ (.A(net1119),
    .B(_0618_),
    .C(_0642_),
    .Y(_0643_));
 sg13g2_or3_2 _4044_ (.A(net1119),
    .B(_0618_),
    .C(_0642_),
    .X(_0644_));
 sg13g2_o21ai_1 _4045_ (.B1(_0642_),
    .Y(_0645_),
    .A1(net1119),
    .A2(_0618_));
 sg13g2_nand2_1 _4046_ (.Y(_0646_),
    .A(_0644_),
    .B(_0645_));
 sg13g2_a21oi_1 _4047_ (.A1(_0644_),
    .A2(_0645_),
    .Y(_0647_),
    .B1(_0619_));
 sg13g2_a21o_1 _4048_ (.A2(_0645_),
    .A1(_0644_),
    .B1(_0619_),
    .X(_0648_));
 sg13g2_o21ai_1 _4049_ (.B1(_0590_),
    .Y(_0649_),
    .A1(net1119),
    .A2(_0621_));
 sg13g2_nand3b_1 _4050_ (.B(_0649_),
    .C(_0513_),
    .Y(_0650_),
    .A_N(_0623_));
 sg13g2_nor3_1 _4051_ (.A(_2914_),
    .B(_0583_),
    .C(_0591_),
    .Y(_0651_));
 sg13g2_a221oi_1 _4052_ (.B2(net1118),
    .C1(_0625_),
    .B1(_0629_),
    .A1(_0517_),
    .Y(_0652_),
    .A2(_0593_));
 sg13g2_o21ai_1 _4053_ (.B1(_0650_),
    .Y(_0653_),
    .A1(_0651_),
    .A2(_0652_));
 sg13g2_a21oi_1 _4054_ (.A1(_0514_),
    .A2(_0607_),
    .Y(_0654_),
    .B1(_0612_));
 sg13g2_nor2_2 _4055_ (.A(net1232),
    .B(_2914_),
    .Y(_0655_));
 sg13g2_nor2_1 _4056_ (.A(_0513_),
    .B(_0655_),
    .Y(_0656_));
 sg13g2_a21oi_1 _4057_ (.A1(_0608_),
    .A2(_0656_),
    .Y(_0657_),
    .B1(_0614_));
 sg13g2_o21ai_1 _4058_ (.B1(_0598_),
    .Y(_0658_),
    .A1(_0654_),
    .A2(_0657_));
 sg13g2_o21ai_1 _4059_ (.B1(net1236),
    .Y(_0659_),
    .A1(net1234),
    .A2(_0599_));
 sg13g2_nand2_1 _4060_ (.Y(_0660_),
    .A(_0603_),
    .B(_0656_));
 sg13g2_nand3_1 _4061_ (.B(_0602_),
    .C(_0660_),
    .A(_0597_),
    .Y(_0661_));
 sg13g2_and2_1 _4062_ (.A(_0658_),
    .B(_0661_),
    .X(_0662_));
 sg13g2_a22oi_1 _4063_ (.Y(_0663_),
    .B1(_0662_),
    .B2(_0485_),
    .A2(_0653_),
    .A1(_0569_));
 sg13g2_nand2_1 _4064_ (.Y(_0664_),
    .A(_0405_),
    .B(_0655_));
 sg13g2_nand3_1 _4065_ (.B(_0565_),
    .C(_0664_),
    .A(_0408_),
    .Y(_0665_));
 sg13g2_o21ai_1 _4066_ (.B1(_0665_),
    .Y(_0666_),
    .A1(_0555_),
    .A2(_0663_));
 sg13g2_xnor2_1 _4067_ (.Y(_0667_),
    .A(_0644_),
    .B(_0666_));
 sg13g2_nand2_2 _4068_ (.Y(_0668_),
    .A(_2729_),
    .B(_0478_));
 sg13g2_nand2_1 _4069_ (.Y(_0669_),
    .A(_0517_),
    .B(_0565_));
 sg13g2_o21ai_1 _4070_ (.B1(_0598_),
    .Y(_0670_),
    .A1(_0632_),
    .A2(_0634_));
 sg13g2_nand3_1 _4071_ (.B(_0638_),
    .C(_0670_),
    .A(_0554_),
    .Y(_0671_));
 sg13g2_a21oi_1 _4072_ (.A1(_0499_),
    .A2(_0591_),
    .Y(_0672_),
    .B1(_0583_));
 sg13g2_o21ai_1 _4073_ (.B1(_0569_),
    .Y(_0673_),
    .A1(_0622_),
    .A2(_0672_));
 sg13g2_and3_1 _4074_ (.X(_0674_),
    .A(_0669_),
    .B(_0671_),
    .C(_0673_));
 sg13g2_a21o_1 _4075_ (.A2(_0666_),
    .A1(_0643_),
    .B1(_0674_),
    .X(_0675_));
 sg13g2_nand3_1 _4076_ (.B(_0666_),
    .C(_0674_),
    .A(_0643_),
    .Y(_0676_));
 sg13g2_and2_2 _4077_ (.A(_0675_),
    .B(_0676_),
    .X(_0677_));
 sg13g2_nand2_1 _4078_ (.Y(_0678_),
    .A(_0668_),
    .B(_0677_));
 sg13g2_a21oi_1 _4079_ (.A1(_0648_),
    .A2(_0667_),
    .Y(_0679_),
    .B1(_0678_));
 sg13g2_nand2_1 _4080_ (.Y(_0680_),
    .A(\dtop.player_inst.synth.alu.registers[1][9] ),
    .B(net1117));
 sg13g2_nand2_1 _4081_ (.Y(_0681_),
    .A(net1053),
    .B(_0541_));
 sg13g2_o21ai_1 _4082_ (.B1(_0681_),
    .Y(_0682_),
    .A1(net1053),
    .A2(_0529_));
 sg13g2_and2_1 _4083_ (.A(_0509_),
    .B(_0682_),
    .X(_0683_));
 sg13g2_a221oi_1 _4084_ (.B2(_0535_),
    .C1(_0683_),
    .B1(_0539_),
    .A1(_0536_),
    .Y(_0684_),
    .A2(_0537_));
 sg13g2_mux2_1 _4085_ (.A0(_0525_),
    .A1(_0532_),
    .S(net1052),
    .X(_0685_));
 sg13g2_nor2_1 _4086_ (.A(\dtop.player_inst.synth.alu.registers[4][2] ),
    .B(net1073),
    .Y(_0686_));
 sg13g2_a21oi_1 _4087_ (.A1(_2662_),
    .A2(net1073),
    .Y(_0687_),
    .B1(_0686_));
 sg13g2_mux2_1 _4088_ (.A0(_0687_),
    .A1(_0523_),
    .S(net1053),
    .X(_0688_));
 sg13g2_nor2_1 _4089_ (.A(net1035),
    .B(_0685_),
    .Y(_0689_));
 sg13g2_a21oi_1 _4090_ (.A1(net1035),
    .A2(_0688_),
    .Y(_0690_),
    .B1(_0689_));
 sg13g2_a21oi_1 _4091_ (.A1(net1037),
    .A2(_0690_),
    .Y(_0691_),
    .B1(net998));
 sg13g2_o21ai_1 _4092_ (.B1(_0691_),
    .Y(_0692_),
    .A1(net1037),
    .A2(_0684_));
 sg13g2_a22oi_1 _4093_ (.Y(_0693_),
    .B1(_0488_),
    .B2(\dtop.player_inst.synth.alu.registers[0][9] ),
    .A2(_2713_),
    .A1(\dtop.detune_counter[6] ));
 sg13g2_nand3_1 _4094_ (.B(_0692_),
    .C(_0693_),
    .A(_0680_),
    .Y(_0694_));
 sg13g2_nor2_1 _4095_ (.A(_0679_),
    .B(_0694_),
    .Y(_0695_));
 sg13g2_xnor2_1 _4096_ (.Y(_0696_),
    .A(_0409_),
    .B(_0695_));
 sg13g2_nor2_1 _4097_ (.A(_0553_),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_nand2_1 _4098_ (.Y(_0698_),
    .A(_0553_),
    .B(_0696_));
 sg13g2_nand2_1 _4099_ (.Y(_0699_),
    .A(\dtop.player_inst.synth.alu.acc[9] ),
    .B(net1000));
 sg13g2_nand2_1 _4100_ (.Y(_0700_),
    .A(\dtop.player_inst.synth.alu.acc[2] ),
    .B(net1100));
 sg13g2_xor2_1 _4101_ (.B(net1165),
    .A(\dtop.player_inst.synth.alu.acc[7] ),
    .X(_0701_));
 sg13g2_a22oi_1 _4102_ (.Y(_0702_),
    .B1(net1075),
    .B2(_0701_),
    .A2(_0375_),
    .A1(\dtop.player_inst.synth.alu.acc[8] ));
 sg13g2_nand3_1 _4103_ (.B(_0700_),
    .C(_0702_),
    .A(_0699_),
    .Y(_0703_));
 sg13g2_mux2_1 _4104_ (.A0(_0646_),
    .A1(_0648_),
    .S(_0667_),
    .X(_0704_));
 sg13g2_nand3_1 _4105_ (.B(_0677_),
    .C(_0704_),
    .A(_0668_),
    .Y(_0705_));
 sg13g2_mux2_1 _4106_ (.A0(\dtop.player_inst.synth.alu.registers[4][1] ),
    .A1(net1235),
    .S(net1073),
    .X(_0706_));
 sg13g2_inv_1 _4107_ (.Y(_0707_),
    .A(_0706_));
 sg13g2_nand2_1 _4108_ (.Y(_0708_),
    .A(net1052),
    .B(_0687_));
 sg13g2_o21ai_1 _4109_ (.B1(_0708_),
    .Y(_0709_),
    .A1(net1052),
    .A2(_0707_));
 sg13g2_mux2_1 _4110_ (.A0(_0527_),
    .A1(_0709_),
    .S(net1035),
    .X(_0710_));
 sg13g2_a21oi_1 _4111_ (.A1(net1036),
    .A2(_0533_),
    .Y(_0711_),
    .B1(net1037));
 sg13g2_o21ai_1 _4112_ (.B1(_0711_),
    .Y(_0712_),
    .A1(net1035),
    .A2(_0542_));
 sg13g2_o21ai_1 _4113_ (.B1(_0712_),
    .Y(_0713_),
    .A1(_0501_),
    .A2(_0710_));
 sg13g2_a22oi_1 _4114_ (.Y(_0714_),
    .B1(_0464_),
    .B2(\dtop.player_inst.synth.alu.registers[1][8] ),
    .A2(_2713_),
    .A1(\dtop.detune_counter[5] ));
 sg13g2_o21ai_1 _4115_ (.B1(_0714_),
    .Y(_0715_),
    .A1(net998),
    .A2(_0713_));
 sg13g2_a21oi_1 _4116_ (.A1(\dtop.player_inst.synth.alu.registers[0][8] ),
    .A2(_0488_),
    .Y(_0716_),
    .B1(_0715_));
 sg13g2_nand2_1 _4117_ (.Y(_0717_),
    .A(_0705_),
    .B(_0716_));
 sg13g2_xnor2_1 _4118_ (.Y(_0718_),
    .A(_0410_),
    .B(_0717_));
 sg13g2_nand2_1 _4119_ (.Y(_0719_),
    .A(_0703_),
    .B(_0718_));
 sg13g2_xor2_1 _4120_ (.B(_0718_),
    .A(_0703_),
    .X(_0720_));
 sg13g2_nand2_1 _4121_ (.Y(_0721_),
    .A(\dtop.player_inst.synth.alu.acc[8] ),
    .B(net1000));
 sg13g2_xor2_1 _4122_ (.B(net1165),
    .A(\dtop.player_inst.synth.alu.acc[6] ),
    .X(_0722_));
 sg13g2_and2_1 _4123_ (.A(net1075),
    .B(_0722_),
    .X(_0723_));
 sg13g2_a221oi_1 _4124_ (.B2(\dtop.player_inst.synth.alu.acc[7] ),
    .C1(_0723_),
    .B1(_0375_),
    .A1(\dtop.player_inst.synth.alu.acc[3] ),
    .Y(_0724_),
    .A2(net1100));
 sg13g2_nor2_1 _4125_ (.A(net1035),
    .B(_0688_),
    .Y(_0725_));
 sg13g2_nand2b_1 _4126_ (.Y(_0726_),
    .B(net1072),
    .A_N(net1236));
 sg13g2_o21ai_1 _4127_ (.B1(_0726_),
    .Y(_0727_),
    .A1(\dtop.player_inst.synth.alu.registers[4][0] ),
    .A2(net1073));
 sg13g2_mux2_1 _4128_ (.A0(_0727_),
    .A1(_0707_),
    .S(net1051),
    .X(_0728_));
 sg13g2_a21oi_1 _4129_ (.A1(net1034),
    .A2(_0728_),
    .Y(_0729_),
    .B1(_0725_));
 sg13g2_nand2b_1 _4130_ (.Y(_0730_),
    .B(_0682_),
    .A_N(net1035));
 sg13g2_a21oi_1 _4131_ (.A1(net1035),
    .A2(_0685_),
    .Y(_0731_),
    .B1(net1037));
 sg13g2_a221oi_1 _4132_ (.B2(_0731_),
    .C1(net999),
    .B1(_0730_),
    .A1(net1037),
    .Y(_0732_),
    .A2(_0729_));
 sg13g2_nand2_1 _4133_ (.Y(_0733_),
    .A(_0619_),
    .B(_0642_));
 sg13g2_nand2_1 _4134_ (.Y(_0734_),
    .A(_0667_),
    .B(_0733_));
 sg13g2_o21ai_1 _4135_ (.B1(_0734_),
    .Y(_0735_),
    .A1(_0620_),
    .A2(_0667_));
 sg13g2_o21ai_1 _4136_ (.B1(_0668_),
    .Y(_0736_),
    .A1(_0646_),
    .A2(_0674_));
 sg13g2_a21o_1 _4137_ (.A2(_0735_),
    .A1(_0677_),
    .B1(_0736_),
    .X(_0737_));
 sg13g2_a22oi_1 _4138_ (.Y(_0738_),
    .B1(net1116),
    .B2(\dtop.player_inst.synth.alu.registers[3][7] ),
    .A2(_2713_),
    .A1(\dtop.detune_counter[4] ));
 sg13g2_a22oi_1 _4139_ (.Y(_0739_),
    .B1(_0464_),
    .B2(\dtop.player_inst.synth.alu.registers[1][7] ),
    .A2(net1121),
    .A1(\dtop.player_inst.synth.alu.registers[2][7] ));
 sg13g2_nand3_1 _4140_ (.B(_0738_),
    .C(_0739_),
    .A(net998),
    .Y(_0740_));
 sg13g2_a21oi_1 _4141_ (.A1(\dtop.player_inst.synth.alu.registers[0][7] ),
    .A2(net994),
    .Y(_0741_),
    .B1(_0740_));
 sg13g2_a21oi_2 _4142_ (.B1(_0732_),
    .Y(_0742_),
    .A2(_0741_),
    .A1(_0737_));
 sg13g2_xnor2_1 _4143_ (.Y(_0743_),
    .A(_0409_),
    .B(_0742_));
 sg13g2_and3_1 _4144_ (.X(_0744_),
    .A(_0721_),
    .B(_0724_),
    .C(_0743_));
 sg13g2_a21oi_1 _4145_ (.A1(_0721_),
    .A2(_0724_),
    .Y(_0745_),
    .B1(_0743_));
 sg13g2_nor3_1 _4146_ (.A(net1099),
    .B(_2811_),
    .C(_0399_),
    .Y(_0746_));
 sg13g2_or2_1 _4147_ (.X(_0747_),
    .B(_0386_),
    .A(_0378_));
 sg13g2_nor2_1 _4148_ (.A(_0746_),
    .B(_0747_),
    .Y(_0748_));
 sg13g2_or3_1 _4149_ (.A(net1100),
    .B(_0387_),
    .C(net1000),
    .X(_0749_));
 sg13g2_inv_1 _4150_ (.Y(_0750_),
    .A(_0749_));
 sg13g2_o21ai_1 _4151_ (.B1(_0748_),
    .Y(_0751_),
    .A1(\dtop.player_inst.synth.alu.acc[7] ),
    .A2(_0750_));
 sg13g2_nand2_1 _4152_ (.Y(_0752_),
    .A(\dtop.player_inst.synth.alu.acc[4] ),
    .B(net1099));
 sg13g2_xor2_1 _4153_ (.B(net1164),
    .A(\dtop.player_inst.synth.alu.acc[5] ),
    .X(_0753_));
 sg13g2_a22oi_1 _4154_ (.Y(_0754_),
    .B1(net1075),
    .B2(_0753_),
    .A2(net1054),
    .A1(\dtop.player_inst.synth.alu.acc[6] ));
 sg13g2_nand3_1 _4155_ (.B(_0752_),
    .C(_0754_),
    .A(_0751_),
    .Y(_0755_));
 sg13g2_nand2b_1 _4156_ (.Y(_0756_),
    .B(net1072),
    .A_N(_0080_));
 sg13g2_nor2b_1 _4157_ (.A(net1051),
    .B_N(_0756_),
    .Y(_0757_));
 sg13g2_a21oi_1 _4158_ (.A1(net1051),
    .A2(_0727_),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_mux2_1 _4159_ (.A0(_0709_),
    .A1(_0758_),
    .S(net1034),
    .X(_0759_));
 sg13g2_nand2_1 _4160_ (.Y(_0760_),
    .A(net1037),
    .B(_0759_));
 sg13g2_a21oi_1 _4161_ (.A1(_0501_),
    .A2(_0534_),
    .Y(_0761_),
    .B1(net999));
 sg13g2_nand3_1 _4162_ (.B(_0645_),
    .C(_0666_),
    .A(_0644_),
    .Y(_0762_));
 sg13g2_a21oi_1 _4163_ (.A1(_0677_),
    .A2(_0762_),
    .Y(_0763_),
    .B1(_0620_));
 sg13g2_a22oi_1 _4164_ (.Y(_0764_),
    .B1(_0647_),
    .B2(_0677_),
    .A2(_0478_),
    .A1(_2729_));
 sg13g2_nand2b_1 _4165_ (.Y(_0765_),
    .B(_0764_),
    .A_N(_0763_));
 sg13g2_nor2_2 _4166_ (.A(net1226),
    .B(_2714_),
    .Y(_0766_));
 sg13g2_nand2_1 _4167_ (.Y(_0767_),
    .A(\dtop.vtop.logo.addr[9] ),
    .B(_0766_));
 sg13g2_a22oi_1 _4168_ (.Y(_0768_),
    .B1(net1117),
    .B2(\dtop.player_inst.synth.alu.registers[1][6] ),
    .A2(net1121),
    .A1(\dtop.player_inst.synth.alu.registers[2][6] ));
 sg13g2_a22oi_1 _4169_ (.Y(_0769_),
    .B1(_0460_),
    .B2(\dtop.player_inst.synth.alu.registers[5][6] ),
    .A2(net1098),
    .A1(\dtop.oct_counter[6] ));
 sg13g2_nand4_1 _4170_ (.B(_0767_),
    .C(_0768_),
    .A(net999),
    .Y(_0770_),
    .D(_0769_));
 sg13g2_a221oi_1 _4171_ (.B2(\dtop.player_inst.synth.alu.registers[0][6] ),
    .C1(_0770_),
    .B1(net994),
    .A1(\dtop.player_inst.synth.alu.registers[3][6] ),
    .Y(_0771_),
    .A2(net1116));
 sg13g2_a22oi_1 _4172_ (.Y(_0772_),
    .B1(_0765_),
    .B2(_0771_),
    .A2(_0761_),
    .A1(_0760_));
 sg13g2_xnor2_1 _4173_ (.Y(_0773_),
    .A(_0410_),
    .B(_0772_));
 sg13g2_nand2_1 _4174_ (.Y(_0774_),
    .A(_0755_),
    .B(_0773_));
 sg13g2_xor2_1 _4175_ (.B(_0773_),
    .A(_0755_),
    .X(_0775_));
 sg13g2_o21ai_1 _4176_ (.B1(_0748_),
    .Y(_0776_),
    .A1(\dtop.player_inst.synth.alu.acc[6] ),
    .A2(_0750_));
 sg13g2_xor2_1 _4177_ (.B(net1164),
    .A(\dtop.player_inst.synth.alu.acc[4] ),
    .X(_0777_));
 sg13g2_or2_1 _4178_ (.X(_0778_),
    .B(net1054),
    .A(net1099));
 sg13g2_a22oi_1 _4179_ (.Y(_0779_),
    .B1(_0778_),
    .B2(\dtop.player_inst.synth.alu.acc[5] ),
    .A2(_0777_),
    .A1(net1075));
 sg13g2_nand2_1 _4180_ (.Y(_0780_),
    .A(_0776_),
    .B(_0779_));
 sg13g2_nor2_1 _4181_ (.A(_0619_),
    .B(_0646_),
    .Y(_0781_));
 sg13g2_nand2b_1 _4182_ (.Y(_0782_),
    .B(_0733_),
    .A_N(_0667_));
 sg13g2_or2_1 _4183_ (.X(_0783_),
    .B(_0782_),
    .A(_0781_));
 sg13g2_a21oi_1 _4184_ (.A1(_0762_),
    .A2(_0783_),
    .Y(_0784_),
    .B1(_0678_));
 sg13g2_nand2b_1 _4185_ (.Y(_0785_),
    .B(net1072),
    .A_N(_0051_));
 sg13g2_mux2_1 _4186_ (.A0(_0785_),
    .A1(_0756_),
    .S(net1051),
    .X(_0786_));
 sg13g2_mux2_1 _4187_ (.A0(_0728_),
    .A1(_0786_),
    .S(net1034),
    .X(_0787_));
 sg13g2_a21o_1 _4188_ (.A2(_0787_),
    .A1(net1037),
    .B1(net998),
    .X(_0788_));
 sg13g2_a21oi_1 _4189_ (.A1(_0501_),
    .A2(_0690_),
    .Y(_0789_),
    .B1(_0788_));
 sg13g2_nand2_1 _4190_ (.Y(_0790_),
    .A(\dtop.player_inst.synth.alu.registers[0][5] ),
    .B(net994));
 sg13g2_nor2_1 _4191_ (.A(_2664_),
    .B(\dtop.vtop.rs.saturated ),
    .Y(_0791_));
 sg13g2_a22oi_1 _4192_ (.Y(_0792_),
    .B1(net1117),
    .B2(\dtop.player_inst.synth.alu.registers[1][5] ),
    .A2(net1121),
    .A1(\dtop.player_inst.synth.alu.registers[2][5] ));
 sg13g2_a22oi_1 _4193_ (.Y(_0793_),
    .B1(net1116),
    .B2(\dtop.player_inst.synth.alu.registers[3][5] ),
    .A2(net1098),
    .A1(\dtop.oct_counter[5] ));
 sg13g2_a22oi_1 _4194_ (.Y(_0794_),
    .B1(_0766_),
    .B2(net1166),
    .A2(_0460_),
    .A1(\dtop.player_inst.synth.alu.registers[5][5] ));
 sg13g2_nand4_1 _4195_ (.B(_0792_),
    .C(_0793_),
    .A(_0790_),
    .Y(_0795_),
    .D(_0794_));
 sg13g2_nor3_2 _4196_ (.A(_0784_),
    .B(_0789_),
    .C(_0795_),
    .Y(_0796_));
 sg13g2_xnor2_1 _4197_ (.Y(_0797_),
    .A(_0409_),
    .B(_0796_));
 sg13g2_nand2_1 _4198_ (.Y(_0798_),
    .A(_0780_),
    .B(_0797_));
 sg13g2_or2_1 _4199_ (.X(_0799_),
    .B(_0797_),
    .A(_0780_));
 sg13g2_nand2_1 _4200_ (.Y(_0800_),
    .A(\dtop.player_inst.synth.alu.acc[5] ),
    .B(net1000));
 sg13g2_nand2_1 _4201_ (.Y(_0801_),
    .A(\dtop.player_inst.synth.alu.acc[4] ),
    .B(net1054));
 sg13g2_nand2_1 _4202_ (.Y(_0802_),
    .A(\dtop.player_inst.synth.alu.acc[6] ),
    .B(net1099));
 sg13g2_xor2_1 _4203_ (.B(net1164),
    .A(\dtop.player_inst.synth.alu.acc[3] ),
    .X(_0803_));
 sg13g2_a22oi_1 _4204_ (.Y(_0804_),
    .B1(_0803_),
    .B2(net1075),
    .A2(_0386_),
    .A1(_0037_));
 sg13g2_nand4_1 _4205_ (.B(_0801_),
    .C(_0802_),
    .A(_0800_),
    .Y(_0805_),
    .D(_0804_));
 sg13g2_nand2_1 _4206_ (.Y(_0806_),
    .A(_0620_),
    .B(_0667_));
 sg13g2_nand3_1 _4207_ (.B(_0782_),
    .C(_0806_),
    .A(_0677_),
    .Y(_0807_));
 sg13g2_and2_1 _4208_ (.A(\dtop.player_inst.synth.alu.registers[1][4] ),
    .B(net1117),
    .X(_0808_));
 sg13g2_a22oi_1 _4209_ (.Y(_0809_),
    .B1(net1116),
    .B2(\dtop.player_inst.synth.alu.registers[3][4] ),
    .A2(net1098),
    .A1(\dtop.oct_counter[4] ));
 sg13g2_a22oi_1 _4210_ (.Y(_0810_),
    .B1(_0766_),
    .B2(\dtop.vtop.logo.addr[7] ),
    .A2(_0460_),
    .A1(\dtop.player_inst.synth.alu.registers[5][4] ));
 sg13g2_a221oi_1 _4211_ (.B2(\dtop.player_inst.synth.alu.registers[0][4] ),
    .C1(_0808_),
    .B1(net994),
    .A1(\dtop.player_inst.synth.alu.registers[2][4] ),
    .Y(_0811_),
    .A2(net1121));
 sg13g2_nor2_1 _4212_ (.A(_0083_),
    .B(net1062),
    .Y(_0812_));
 sg13g2_nand2b_1 _4213_ (.Y(_0813_),
    .B(net1072),
    .A_N(_0083_));
 sg13g2_mux2_1 _4214_ (.A0(_0813_),
    .A1(_0785_),
    .S(net1051),
    .X(_0814_));
 sg13g2_nand2_1 _4215_ (.Y(_0815_),
    .A(net1033),
    .B(_0814_));
 sg13g2_o21ai_1 _4216_ (.B1(_0815_),
    .Y(_0816_),
    .A1(net1033),
    .A2(_0758_));
 sg13g2_a21oi_1 _4217_ (.A1(net1038),
    .A2(_0816_),
    .Y(_0817_),
    .B1(net998));
 sg13g2_o21ai_1 _4218_ (.B1(_0817_),
    .Y(_0818_),
    .A1(net1038),
    .A2(_0710_));
 sg13g2_nand4_1 _4219_ (.B(_0810_),
    .C(_0811_),
    .A(_0809_),
    .Y(_0819_),
    .D(_0818_));
 sg13g2_a21oi_2 _4220_ (.B1(_0819_),
    .Y(_0820_),
    .A2(_0807_),
    .A1(_0668_));
 sg13g2_xnor2_1 _4221_ (.Y(_0821_),
    .A(_0409_),
    .B(_0820_));
 sg13g2_and2_1 _4222_ (.A(_0805_),
    .B(_0821_),
    .X(_0822_));
 sg13g2_nor2_1 _4223_ (.A(\dtop.player_inst.synth.alu.acc[3] ),
    .B(_0749_),
    .Y(_0823_));
 sg13g2_a21oi_1 _4224_ (.A1(_2637_),
    .A2(_0749_),
    .Y(_0824_),
    .B1(_0823_));
 sg13g2_xor2_1 _4225_ (.B(net1164),
    .A(\dtop.player_inst.synth.alu.acc[2] ),
    .X(_0825_));
 sg13g2_a22oi_1 _4226_ (.Y(_0826_),
    .B1(_0825_),
    .B2(net1075),
    .A2(_0386_),
    .A1(\dtop.player_inst.synth.alu.acc[9] ));
 sg13g2_a22oi_1 _4227_ (.Y(_0827_),
    .B1(_0778_),
    .B2(_0824_),
    .A2(net1000),
    .A1(\dtop.player_inst.synth.alu.acc[4] ));
 sg13g2_and2_2 _4228_ (.A(_0826_),
    .B(_0827_),
    .X(_0828_));
 sg13g2_a21oi_1 _4229_ (.A1(_0675_),
    .A2(_0676_),
    .Y(_0829_),
    .B1(_0647_));
 sg13g2_a221oi_1 _4230_ (.B2(_0704_),
    .C1(_0829_),
    .B1(_0677_),
    .A1(_2729_),
    .Y(_0830_),
    .A2(_0478_));
 sg13g2_nor3_1 _4231_ (.A(_2663_),
    .B(net1226),
    .C(net1062),
    .Y(_0831_));
 sg13g2_nand3b_1 _4232_ (.B(net1072),
    .C(\dtop.vtop.logo.addr[9] ),
    .Y(_0832_),
    .A_N(\dtop.vtop.rs.saturated ));
 sg13g2_mux2_1 _4233_ (.A0(_0831_),
    .A1(_0812_),
    .S(net1051),
    .X(_0833_));
 sg13g2_o21ai_1 _4234_ (.B1(net1038),
    .Y(_0834_),
    .A1(net1033),
    .A2(_0786_));
 sg13g2_a21oi_1 _4235_ (.A1(net1034),
    .A2(_0833_),
    .Y(_0835_),
    .B1(_0834_));
 sg13g2_nor2_1 _4236_ (.A(net998),
    .B(_0835_),
    .Y(_0836_));
 sg13g2_o21ai_1 _4237_ (.B1(_0836_),
    .Y(_0837_),
    .A1(net1038),
    .A2(_0729_));
 sg13g2_nand2_1 _4238_ (.Y(_0838_),
    .A(net1169),
    .B(_0766_));
 sg13g2_a22oi_1 _4239_ (.Y(_0839_),
    .B1(net1116),
    .B2(\dtop.player_inst.synth.alu.registers[3][3] ),
    .A2(net1117),
    .A1(\dtop.player_inst.synth.alu.registers[1][3] ));
 sg13g2_a22oi_1 _4240_ (.Y(_0840_),
    .B1(_0460_),
    .B2(\dtop.player_inst.synth.alu.registers[5][3] ),
    .A2(net1121),
    .A1(\dtop.player_inst.synth.alu.registers[2][3] ));
 sg13g2_nand3_1 _4241_ (.B(_0839_),
    .C(_0840_),
    .A(_0838_),
    .Y(_0841_));
 sg13g2_a221oi_1 _4242_ (.B2(\dtop.player_inst.synth.alu.registers[0][3] ),
    .C1(_0841_),
    .B1(net994),
    .A1(\dtop.oct_counter[3] ),
    .Y(_0842_),
    .A2(net1098));
 sg13g2_nand2_2 _4243_ (.Y(_0843_),
    .A(_0837_),
    .B(_0842_));
 sg13g2_o21ai_1 _4244_ (.B1(_0410_),
    .Y(_0844_),
    .A1(_0830_),
    .A2(_0843_));
 sg13g2_or3_1 _4245_ (.A(_0410_),
    .B(_0830_),
    .C(_0843_),
    .X(_0845_));
 sg13g2_a21o_1 _4246_ (.A2(_0845_),
    .A1(_0844_),
    .B1(_0828_),
    .X(_0846_));
 sg13g2_nand3_1 _4247_ (.B(_0747_),
    .C(_0749_),
    .A(\dtop.player_inst.synth.alu.acc[8] ),
    .Y(_0847_));
 sg13g2_xor2_1 _4248_ (.B(net1164),
    .A(\dtop.player_inst.synth.alu.acc[1] ),
    .X(_0848_));
 sg13g2_nand2_1 _4249_ (.Y(_0849_),
    .A(\dtop.player_inst.synth.alu.acc[3] ),
    .B(net1000));
 sg13g2_nand2_1 _4250_ (.Y(_0850_),
    .A(_0847_),
    .B(_0849_));
 sg13g2_a221oi_1 _4251_ (.B2(_0848_),
    .C1(_0850_),
    .B1(net1075),
    .A1(\dtop.player_inst.synth.alu.acc[2] ),
    .Y(_0851_),
    .A2(net1054));
 sg13g2_nand2_1 _4252_ (.Y(_0852_),
    .A(net1072),
    .B(_0791_));
 sg13g2_mux2_1 _4253_ (.A0(_0852_),
    .A1(_0832_),
    .S(net1051),
    .X(_0853_));
 sg13g2_nand2b_1 _4254_ (.Y(_0854_),
    .B(_0814_),
    .A_N(net1033));
 sg13g2_a21oi_1 _4255_ (.A1(net1033),
    .A2(_0853_),
    .Y(_0855_),
    .B1(_0501_));
 sg13g2_a22oi_1 _4256_ (.Y(_0856_),
    .B1(_0854_),
    .B2(_0855_),
    .A2(_0759_),
    .A1(_0501_));
 sg13g2_nand2_1 _4257_ (.Y(_0857_),
    .A(\dtop.player_inst.synth.alu.registers[5][2] ),
    .B(_0460_));
 sg13g2_a22oi_1 _4258_ (.Y(_0858_),
    .B1(net1116),
    .B2(\dtop.player_inst.synth.alu.registers[3][2] ),
    .A2(net1117),
    .A1(\dtop.player_inst.synth.alu.registers[1][2] ));
 sg13g2_a22oi_1 _4259_ (.Y(_0859_),
    .B1(_0766_),
    .B2(net1175),
    .A2(net1121),
    .A1(\dtop.player_inst.synth.alu.registers[2][2] ));
 sg13g2_nand3_1 _4260_ (.B(_0858_),
    .C(_0859_),
    .A(_0857_),
    .Y(_0860_));
 sg13g2_a221oi_1 _4261_ (.B2(\dtop.player_inst.synth.alu.registers[0][2] ),
    .C1(_0860_),
    .B1(net994),
    .A1(net1179),
    .Y(_0861_),
    .A2(net1098));
 sg13g2_o21ai_1 _4262_ (.B1(_0861_),
    .Y(_0862_),
    .A1(net998),
    .A2(_0856_));
 sg13g2_xnor2_1 _4263_ (.Y(_0863_),
    .A(_0410_),
    .B(_0862_));
 sg13g2_nor2b_1 _4264_ (.A(_0851_),
    .B_N(_0863_),
    .Y(_0864_));
 sg13g2_nand2_1 _4265_ (.Y(_0865_),
    .A(\dtop.player_inst.synth.alu.acc[9] ),
    .B(net1099));
 sg13g2_xor2_1 _4266_ (.B(net1164),
    .A(\dtop.player_inst.synth.alu.acc[0] ),
    .X(_0866_));
 sg13g2_a22oi_1 _4267_ (.Y(_0867_),
    .B1(_0866_),
    .B2(net1075),
    .A2(_0386_),
    .A1(\dtop.player_inst.synth.alu.acc[7] ));
 sg13g2_nand2_1 _4268_ (.Y(_0868_),
    .A(_0865_),
    .B(_0867_));
 sg13g2_a221oi_1 _4269_ (.B2(\dtop.player_inst.synth.alu.acc[2] ),
    .C1(_0868_),
    .B1(net1000),
    .A1(\dtop.player_inst.synth.alu.acc[1] ),
    .Y(_0869_),
    .A2(net1054));
 sg13g2_nand2b_1 _4270_ (.Y(_0870_),
    .B(_0833_),
    .A_N(net1033));
 sg13g2_and2_2 _4271_ (.A(net1034),
    .B(net1052),
    .X(_0871_));
 sg13g2_nand4_1 _4272_ (.B(net1033),
    .C(net1051),
    .A(net1072),
    .Y(_0872_),
    .D(_0791_));
 sg13g2_nand3_1 _4273_ (.B(_0870_),
    .C(_0872_),
    .A(net1038),
    .Y(_0873_));
 sg13g2_a21oi_1 _4274_ (.A1(_0501_),
    .A2(_0787_),
    .Y(_0874_),
    .B1(net998));
 sg13g2_nand2_1 _4275_ (.Y(_0875_),
    .A(\dtop.player_inst.synth.alu.registers[5][1] ),
    .B(_0460_));
 sg13g2_a22oi_1 _4276_ (.Y(_0876_),
    .B1(_0766_),
    .B2(net1176),
    .A2(net1116),
    .A1(\dtop.player_inst.synth.alu.registers[3][1] ));
 sg13g2_a22oi_1 _4277_ (.Y(_0877_),
    .B1(net1117),
    .B2(\dtop.player_inst.synth.alu.registers[1][1] ),
    .A2(net1121),
    .A1(\dtop.player_inst.synth.alu.registers[2][1] ));
 sg13g2_nor2b_1 _4278_ (.A(\dtop.player_inst.synth.alu.acc[0] ),
    .B_N(\dtop.player_inst.synth.alu.carry ),
    .Y(_0878_));
 sg13g2_nand2_1 _4279_ (.Y(_0879_),
    .A(_2636_),
    .B(\dtop.player_inst.synth.alu.carry ));
 sg13g2_a21oi_1 _4280_ (.A1(_2820_),
    .A2(_2955_),
    .Y(_0880_),
    .B1(_2699_));
 sg13g2_a22oi_1 _4281_ (.Y(_0881_),
    .B1(_0878_),
    .B2(_0880_),
    .A2(net1098),
    .A1(net1180));
 sg13g2_nand4_1 _4282_ (.B(_0876_),
    .C(_0877_),
    .A(_0875_),
    .Y(_0882_),
    .D(_0881_));
 sg13g2_a221oi_1 _4283_ (.B2(_0874_),
    .C1(_0882_),
    .B1(_0873_),
    .A1(\dtop.player_inst.synth.alu.registers[0][1] ),
    .Y(_0883_),
    .A2(net994));
 sg13g2_xnor2_1 _4284_ (.Y(_0884_),
    .A(_0409_),
    .B(_0883_));
 sg13g2_nor2b_1 _4285_ (.A(_0869_),
    .B_N(_0884_),
    .Y(_0885_));
 sg13g2_nor3_1 _4286_ (.A(_2665_),
    .B(net1226),
    .C(net1062),
    .Y(_0886_));
 sg13g2_o21ai_1 _4287_ (.B1(net1038),
    .Y(_0887_),
    .A1(net1033),
    .A2(_0853_));
 sg13g2_a21oi_1 _4288_ (.A1(_0871_),
    .A2(_0886_),
    .Y(_0888_),
    .B1(_0887_));
 sg13g2_a21o_1 _4289_ (.A2(_0816_),
    .A1(_0501_),
    .B1(_0888_),
    .X(_0889_));
 sg13g2_and2_1 _4290_ (.A(\dtop.player_inst.synth.alu.registers[3][0] ),
    .B(net1116),
    .X(_0890_));
 sg13g2_a221oi_1 _4291_ (.B2(\dtop.oct_counter[5] ),
    .C1(_0890_),
    .B1(_0766_),
    .A1(\dtop.player_inst.synth.alu.registers[2][0] ),
    .Y(_0891_),
    .A2(net1121));
 sg13g2_a22oi_1 _4292_ (.Y(_0892_),
    .B1(net1117),
    .B2(\dtop.player_inst.synth.alu.registers[1][0] ),
    .A2(_0460_),
    .A1(\dtop.player_inst.synth.alu.registers[5][0] ));
 sg13g2_a22oi_1 _4293_ (.Y(_0893_),
    .B1(_0879_),
    .B2(_0880_),
    .A2(net1098),
    .A1(net1183));
 sg13g2_nand3_1 _4294_ (.B(_0892_),
    .C(_0893_),
    .A(_0891_),
    .Y(_0894_));
 sg13g2_a21oi_1 _4295_ (.A1(\dtop.player_inst.synth.alu.registers[0][0] ),
    .A2(net994),
    .Y(_0895_),
    .B1(_0894_));
 sg13g2_o21ai_1 _4296_ (.B1(_0895_),
    .Y(_0896_),
    .A1(net999),
    .A2(_0889_));
 sg13g2_a221oi_1 _4297_ (.B2(\dtop.player_inst.synth.alu.acc[6] ),
    .C1(_0377_),
    .B1(_0386_),
    .A1(net1164),
    .Y(_0897_),
    .A2(net1099));
 sg13g2_a22oi_1 _4298_ (.Y(_0898_),
    .B1(net1000),
    .B2(\dtop.player_inst.synth.alu.acc[1] ),
    .A2(net1054),
    .A1(\dtop.player_inst.synth.alu.acc[0] ));
 sg13g2_nand2_2 _4299_ (.Y(_0899_),
    .A(_0897_),
    .B(_0898_));
 sg13g2_mux2_1 _4300_ (.A0(_0409_),
    .A1(_0899_),
    .S(_0896_),
    .X(_0900_));
 sg13g2_xnor2_1 _4301_ (.Y(_0901_),
    .A(_0869_),
    .B(_0884_));
 sg13g2_a21oi_1 _4302_ (.A1(_0900_),
    .A2(_0901_),
    .Y(_0902_),
    .B1(_0885_));
 sg13g2_xor2_1 _4303_ (.B(_0863_),
    .A(_0851_),
    .X(_0903_));
 sg13g2_nor2_1 _4304_ (.A(_0902_),
    .B(_0903_),
    .Y(_0904_));
 sg13g2_nor2_1 _4305_ (.A(_0864_),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_and3_1 _4306_ (.X(_0906_),
    .A(_0828_),
    .B(_0844_),
    .C(_0845_));
 sg13g2_nand3_1 _4307_ (.B(_0844_),
    .C(_0845_),
    .A(_0828_),
    .Y(_0907_));
 sg13g2_nand2_1 _4308_ (.Y(_0908_),
    .A(_0846_),
    .B(_0907_));
 sg13g2_o21ai_1 _4309_ (.B1(_0846_),
    .Y(_0909_),
    .A1(_0905_),
    .A2(_0906_));
 sg13g2_xor2_1 _4310_ (.B(_0821_),
    .A(_0805_),
    .X(_0910_));
 sg13g2_a21o_1 _4311_ (.A2(_0910_),
    .A1(_0909_),
    .B1(_0822_),
    .X(_0911_));
 sg13g2_nand2_1 _4312_ (.Y(_0912_),
    .A(_0799_),
    .B(_0911_));
 sg13g2_a221oi_1 _4313_ (.B2(_0910_),
    .C1(_0822_),
    .B1(_0909_),
    .A1(_0780_),
    .Y(_0913_),
    .A2(_0797_));
 sg13g2_nand3b_1 _4314_ (.B(_0775_),
    .C(_0799_),
    .Y(_0914_),
    .A_N(_0913_));
 sg13g2_nand2_1 _4315_ (.Y(_0915_),
    .A(_0774_),
    .B(_0914_));
 sg13g2_a21oi_1 _4316_ (.A1(_0774_),
    .A2(_0914_),
    .Y(_0916_),
    .B1(_0744_));
 sg13g2_o21ai_1 _4317_ (.B1(_0720_),
    .Y(_0917_),
    .A1(_0745_),
    .A2(_0916_));
 sg13g2_and2_1 _4318_ (.A(_0719_),
    .B(_0917_),
    .X(_0918_));
 sg13g2_o21ai_1 _4319_ (.B1(_0698_),
    .Y(_0919_),
    .A1(_0697_),
    .A2(_0918_));
 sg13g2_nand2_1 _4320_ (.Y(_0920_),
    .A(_0549_),
    .B(_0919_));
 sg13g2_nor2_1 _4321_ (.A(_2932_),
    .B(_0548_),
    .Y(_0921_));
 sg13g2_a22oi_1 _4322_ (.Y(_0089_),
    .B1(_0920_),
    .B2(_0921_),
    .A2(_2933_),
    .A1(_2932_));
 sg13g2_nor2_1 _4323_ (.A(net557),
    .B(_2854_),
    .Y(_0922_));
 sg13g2_nor3_1 _4324_ (.A(net557),
    .B(net617),
    .C(_2854_),
    .Y(_0923_));
 sg13g2_nor4_2 _4325_ (.A(net557),
    .B(_0056_),
    .C(net604),
    .Y(_0924_),
    .D(_2854_));
 sg13g2_nor2b_2 _4326_ (.A(net1178),
    .B_N(_0924_),
    .Y(_0925_));
 sg13g2_nor2b_1 _4327_ (.A(_0054_),
    .B_N(_0925_),
    .Y(_0926_));
 sg13g2_and3_1 _4328_ (.X(_0927_),
    .A(net1177),
    .B(_2672_),
    .C(_0926_));
 sg13g2_and2_1 _4329_ (.A(net1176),
    .B(_0927_),
    .X(_0928_));
 sg13g2_and3_1 _4330_ (.X(_0929_),
    .A(net1169),
    .B(net1175),
    .C(_0928_));
 sg13g2_nor2_2 _4331_ (.A(net1168),
    .B(net1173),
    .Y(_0930_));
 sg13g2_nor3_1 _4332_ (.A(\dtop.vtop.logo.addr[9] ),
    .B(net1166),
    .C(net1167),
    .Y(_0931_));
 sg13g2_nand3_1 _4333_ (.B(_0930_),
    .C(_0931_),
    .A(net1177),
    .Y(_0932_));
 sg13g2_nor2_1 _4334_ (.A(\dtop.oct_counter[4] ),
    .B(\dtop.oct_counter[3] ),
    .Y(_0933_));
 sg13g2_nand4_1 _4335_ (.B(net1226),
    .C(_0925_),
    .A(net1176),
    .Y(_0934_),
    .D(_0933_));
 sg13g2_o21ai_1 _4336_ (.B1(net1243),
    .Y(_0935_),
    .A1(_0932_),
    .A2(_0934_));
 sg13g2_nand3_1 _4337_ (.B(net580),
    .C(_0929_),
    .A(net616),
    .Y(_0936_));
 sg13g2_nor2_1 _4338_ (.A(net615),
    .B(_0936_),
    .Y(_0937_));
 sg13g2_xnor2_1 _4339_ (.Y(_0938_),
    .A(net1226),
    .B(_0937_));
 sg13g2_nor2_1 _4340_ (.A(_0935_),
    .B(_0938_),
    .Y(_0138_));
 sg13g2_nor4_2 _4341_ (.A(net4),
    .B(net1226),
    .C(net1050),
    .Y(_0939_),
    .D(_0938_));
 sg13g2_nor2_1 _4342_ (.A(net5),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_o21ai_1 _4343_ (.B1(\dtop.detune_counter[4] ),
    .Y(_0941_),
    .A1(net5),
    .A2(_0939_));
 sg13g2_nor2_1 _4344_ (.A(_0051_),
    .B(_0941_),
    .Y(_0942_));
 sg13g2_and2_1 _4345_ (.A(net577),
    .B(_0942_),
    .X(_0943_));
 sg13g2_and3_1 _4346_ (.X(_0944_),
    .A(net1235),
    .B(net1236),
    .C(_0943_));
 sg13g2_and2_1 _4347_ (.A(_2889_),
    .B(_0944_),
    .X(_0945_));
 sg13g2_nand2_2 _4348_ (.Y(_0946_),
    .A(net1231),
    .B(_0945_));
 sg13g2_nor2_1 _4349_ (.A(_2659_),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_nor4_1 _4350_ (.A(_2658_),
    .B(_2659_),
    .C(_2660_),
    .D(_0946_),
    .Y(_0948_));
 sg13g2_nor2b_1 _4351_ (.A(_2879_),
    .B_N(_0945_),
    .Y(_0949_));
 sg13g2_nand2_1 _4352_ (.Y(_0950_),
    .A(net1229),
    .B(_0949_));
 sg13g2_a22oi_1 _4353_ (.Y(_0951_),
    .B1(_0950_),
    .B2(net1227),
    .A2(_0949_),
    .A1(_2908_));
 sg13g2_nor2_1 _4354_ (.A(net621),
    .B(_0950_),
    .Y(_0952_));
 sg13g2_xnor2_1 _4355_ (.Y(_0953_),
    .A(_0057_),
    .B(_0952_));
 sg13g2_inv_1 _4356_ (.Y(_0954_),
    .A(net622));
 sg13g2_nand2b_1 _4357_ (.Y(_0955_),
    .B(_0953_),
    .A_N(_0951_));
 sg13g2_a21oi_1 _4358_ (.A1(net1247),
    .A2(_0955_),
    .Y(_0956_),
    .B1(net5));
 sg13g2_xnor2_1 _4359_ (.Y(_0957_),
    .A(net637),
    .B(_0940_));
 sg13g2_nor2_1 _4360_ (.A(net953),
    .B(_0957_),
    .Y(_0090_));
 sg13g2_xor2_1 _4361_ (.B(_0941_),
    .A(net573),
    .X(_0958_));
 sg13g2_nor2_1 _4362_ (.A(net953),
    .B(_0958_),
    .Y(_0091_));
 sg13g2_nor2_1 _4363_ (.A(net577),
    .B(_0942_),
    .Y(_0959_));
 sg13g2_nor3_1 _4364_ (.A(_0943_),
    .B(net953),
    .C(_0959_),
    .Y(_0092_));
 sg13g2_nor3_1 _4365_ (.A(_0051_),
    .B(net633),
    .C(_0941_),
    .Y(_0960_));
 sg13g2_xnor2_1 _4366_ (.Y(_0961_),
    .A(net1236),
    .B(_0960_));
 sg13g2_nor2_1 _4367_ (.A(net953),
    .B(net634),
    .Y(_0093_));
 sg13g2_a21oi_1 _4368_ (.A1(net1236),
    .A2(_0943_),
    .Y(_0962_),
    .B1(net1235));
 sg13g2_nor3_1 _4369_ (.A(_0944_),
    .B(net952),
    .C(net591),
    .Y(_0094_));
 sg13g2_nand3_1 _4370_ (.B(_2684_),
    .C(_0943_),
    .A(net1236),
    .Y(_0963_));
 sg13g2_xnor2_1 _4371_ (.Y(_0964_),
    .A(_2662_),
    .B(_0963_));
 sg13g2_nor2_1 _4372_ (.A(net953),
    .B(_0964_),
    .Y(_0095_));
 sg13g2_a21oi_1 _4373_ (.A1(\dtop.detune_counter[9] ),
    .A2(_0944_),
    .Y(_0965_),
    .B1(net628));
 sg13g2_nor3_1 _4374_ (.A(_0945_),
    .B(net952),
    .C(net629),
    .Y(_0096_));
 sg13g2_nand3b_1 _4375_ (.B(_0944_),
    .C(net647),
    .Y(_0966_),
    .A_N(net1233));
 sg13g2_xnor2_1 _4376_ (.Y(_0967_),
    .A(_2661_),
    .B(_0966_));
 sg13g2_nor2_1 _4377_ (.A(net952),
    .B(_0967_),
    .Y(_0097_));
 sg13g2_xnor2_1 _4378_ (.Y(_0968_),
    .A(net644),
    .B(_0946_));
 sg13g2_nor2_1 _4379_ (.A(net952),
    .B(_0968_),
    .Y(_0098_));
 sg13g2_nor3_2 _4380_ (.A(_2659_),
    .B(_2660_),
    .C(_0946_),
    .Y(_0969_));
 sg13g2_nor2_1 _4381_ (.A(net1230),
    .B(_0947_),
    .Y(_0970_));
 sg13g2_nor3_1 _4382_ (.A(net952),
    .B(_0969_),
    .C(_0970_),
    .Y(_0099_));
 sg13g2_nor2_1 _4383_ (.A(net569),
    .B(_0969_),
    .Y(_0971_));
 sg13g2_nor3_1 _4384_ (.A(_0948_),
    .B(net952),
    .C(_0971_),
    .Y(_0100_));
 sg13g2_nand2_1 _4385_ (.Y(_0972_),
    .A(_2681_),
    .B(_0969_));
 sg13g2_xor2_1 _4386_ (.B(_0972_),
    .A(net1229),
    .X(_0973_));
 sg13g2_nor2_1 _4387_ (.A(net952),
    .B(_0973_),
    .Y(_0101_));
 sg13g2_nor2_1 _4388_ (.A(_0951_),
    .B(net953),
    .Y(_0102_));
 sg13g2_nor2_1 _4389_ (.A(_0954_),
    .B(net952),
    .Y(_0103_));
 sg13g2_nor2_1 _4390_ (.A(net1183),
    .B(net1181),
    .Y(_0974_));
 sg13g2_and3_1 _4391_ (.X(_0975_),
    .A(net1178),
    .B(_2730_),
    .C(_0974_));
 sg13g2_nand4_1 _4392_ (.B(net1200),
    .C(_2722_),
    .A(net1178),
    .Y(_0976_),
    .D(_0974_));
 sg13g2_nor2_1 _4393_ (.A(net1220),
    .B(net1123),
    .Y(_0977_));
 sg13g2_nand2b_1 _4394_ (.Y(_0978_),
    .B(\dtop.vtop.pipeline.wave_index[1] ),
    .A_N(\dtop.vtop.pipeline.wave_index[0] ));
 sg13g2_nor2_1 _4395_ (.A(net1114),
    .B(_0978_),
    .Y(_0979_));
 sg13g2_a21o_1 _4396_ (.A2(net1111),
    .A1(_0001_),
    .B1(_0979_),
    .X(_0980_));
 sg13g2_nand3b_1 _4397_ (.B(_0057_),
    .C(net1228),
    .Y(_0981_),
    .A_N(\dtop.detune_counter[16] ));
 sg13g2_nand3b_1 _4398_ (.B(_2660_),
    .C(_2659_),
    .Y(_0982_),
    .A_N(_2876_));
 sg13g2_a21o_2 _4399_ (.A2(_0982_),
    .A1(_0981_),
    .B1(\dtop.detune_counter[17] ),
    .X(_0983_));
 sg13g2_and3_1 _4400_ (.X(_0984_),
    .A(\dtop.vtop.pipeline.wave_index[0] ),
    .B(\dtop.vtop.pipeline.wave_index[1] ),
    .C(_0983_));
 sg13g2_a21oi_1 _4401_ (.A1(\dtop.vtop.pipeline.wave_index[0] ),
    .A2(\dtop.vtop.pipeline.wave_index[1] ),
    .Y(_0985_),
    .B1(_0003_));
 sg13g2_or3_1 _4402_ (.A(net1114),
    .B(_0984_),
    .C(_0985_),
    .X(_0986_));
 sg13g2_o21ai_1 _4403_ (.B1(_0986_),
    .Y(_0987_),
    .A1(_2669_),
    .A2(net1125));
 sg13g2_inv_1 _4404_ (.Y(_0988_),
    .A(_0987_));
 sg13g2_mux2_1 _4405_ (.A0(_0001_),
    .A1(_0004_),
    .S(net1123),
    .X(_0989_));
 sg13g2_mux2_2 _4406_ (.A0(_2685_),
    .A1(_2686_),
    .S(net1122),
    .X(_0990_));
 sg13g2_mux2_2 _4407_ (.A0(_0088_),
    .A1(_0003_),
    .S(net1124),
    .X(_0991_));
 sg13g2_and2_1 _4408_ (.A(net1108),
    .B(net1104),
    .X(_0992_));
 sg13g2_nand2_1 _4409_ (.Y(_0993_),
    .A(net1106),
    .B(net1104));
 sg13g2_nor2_2 _4410_ (.A(net1108),
    .B(net1103),
    .Y(_0994_));
 sg13g2_o21ai_1 _4411_ (.B1(net1103),
    .Y(_0995_),
    .A1(\dtop.vtop.pipeline.phases[2][15] ),
    .A2(net1107));
 sg13g2_a22oi_1 _4412_ (.Y(_0996_),
    .B1(_0994_),
    .B2(\dtop.vtop.pipeline.zg_acc[8] ),
    .A2(net1107),
    .A1(\dtop.vtop.pipeline.phases[1][15] ));
 sg13g2_a22oi_1 _4413_ (.Y(_0997_),
    .B1(_0995_),
    .B2(_0996_),
    .A2(net1097),
    .A1(_0002_));
 sg13g2_mux4_1 _4414_ (.S0(_0991_),
    .A0(_2687_),
    .A1(_2688_),
    .A2(_2689_),
    .A3(_0002_),
    .S1(net1107),
    .X(_0998_));
 sg13g2_nor2_1 _4415_ (.A(_2658_),
    .B(_0981_),
    .Y(_0999_));
 sg13g2_nor3_1 _4416_ (.A(_2659_),
    .B(net1230),
    .C(_2876_),
    .Y(_1000_));
 sg13g2_a221oi_1 _4417_ (.B2(net1230),
    .C1(_1000_),
    .B1(_0999_),
    .A1(_2658_),
    .Y(_1001_),
    .A2(_2847_));
 sg13g2_a21oi_1 _4418_ (.A1(\dtop.detune_counter[13] ),
    .A2(_0999_),
    .Y(_1002_),
    .B1(net1124));
 sg13g2_or2_1 _4419_ (.X(_1003_),
    .B(_1002_),
    .A(_1001_));
 sg13g2_nand2_1 _4420_ (.Y(_1004_),
    .A(_0997_),
    .B(_1003_));
 sg13g2_and2_1 _4421_ (.A(_0035_),
    .B(net1097),
    .X(_1005_));
 sg13g2_nand2_1 _4422_ (.Y(_1006_),
    .A(_0035_),
    .B(net1097));
 sg13g2_nor3_1 _4423_ (.A(_0036_),
    .B(net1107),
    .C(net1103),
    .Y(_1007_));
 sg13g2_or2_1 _4424_ (.X(_1008_),
    .B(net1107),
    .A(\dtop.vtop.pipeline.phases[2][14] ));
 sg13g2_a21o_1 _4425_ (.A2(net1107),
    .A1(\dtop.vtop.pipeline.phases[1][14] ),
    .B1(net1103),
    .X(_1009_));
 sg13g2_nor2_2 _4426_ (.A(net1106),
    .B(_0990_),
    .Y(_1010_));
 sg13g2_nand2b_2 _4427_ (.Y(_1011_),
    .B(net1104),
    .A_N(net1105));
 sg13g2_a221oi_1 _4428_ (.B2(_1008_),
    .C1(_1007_),
    .B1(net1103),
    .A1(\dtop.vtop.pipeline.phases[1][14] ),
    .Y(_1012_),
    .A2(net1107));
 sg13g2_a21o_1 _4429_ (.A2(_1009_),
    .A1(_1008_),
    .B1(_1007_),
    .X(_1013_));
 sg13g2_nand2_1 _4430_ (.Y(_1014_),
    .A(_1006_),
    .B(_1013_));
 sg13g2_nor2_1 _4431_ (.A(_0998_),
    .B(_1003_),
    .Y(_1015_));
 sg13g2_or2_1 _4432_ (.X(_1016_),
    .B(_1003_),
    .A(_0998_));
 sg13g2_a21oi_2 _4433_ (.B1(_1016_),
    .Y(_1017_),
    .A2(_1013_),
    .A1(_1006_));
 sg13g2_o21ai_1 _4434_ (.B1(_1015_),
    .Y(_1018_),
    .A1(_1005_),
    .A2(_1012_));
 sg13g2_nor3_2 _4435_ (.A(_1005_),
    .B(_1012_),
    .C(_1015_),
    .Y(_1019_));
 sg13g2_nand3_1 _4436_ (.B(_1013_),
    .C(_1016_),
    .A(_1006_),
    .Y(_1020_));
 sg13g2_nand2_1 _4437_ (.Y(_1021_),
    .A(net1061),
    .B(net1060));
 sg13g2_and2_1 _4438_ (.A(net1105),
    .B(_0990_),
    .X(_1022_));
 sg13g2_a22oi_1 _4439_ (.Y(_1023_),
    .B1(_1022_),
    .B2(\dtop.vtop.pipeline.phases[1][12] ),
    .A2(net1093),
    .A1(\dtop.vtop.pipeline.phases[2][12] ));
 sg13g2_a21oi_2 _4440_ (.B1(net1097),
    .Y(_1024_),
    .A2(net1094),
    .A1(\dtop.vtop.pipeline.zg_acc[5] ));
 sg13g2_a22oi_1 _4441_ (.Y(_1025_),
    .B1(_1023_),
    .B2(_1024_),
    .A2(net1096),
    .A1(_0032_));
 sg13g2_xor2_1 _4442_ (.B(_1025_),
    .A(net1046),
    .X(_1026_));
 sg13g2_xnor2_1 _4443_ (.Y(_1027_),
    .A(net1046),
    .B(_1025_));
 sg13g2_nor3_1 _4444_ (.A(_0034_),
    .B(net1108),
    .C(net1103),
    .Y(_1028_));
 sg13g2_or2_1 _4445_ (.X(_1029_),
    .B(net1108),
    .A(\dtop.vtop.pipeline.phases[2][13] ));
 sg13g2_a221oi_1 _4446_ (.B2(_1029_),
    .C1(_1028_),
    .B1(_0991_),
    .A1(\dtop.vtop.pipeline.phases[1][13] ),
    .Y(_1030_),
    .A2(net1107));
 sg13g2_a21o_2 _4447_ (.A2(_0992_),
    .A1(_0033_),
    .B1(_1030_),
    .X(_1031_));
 sg13g2_xnor2_1 _4448_ (.Y(_1032_),
    .A(net1046),
    .B(_1031_));
 sg13g2_xor2_1 _4449_ (.B(_1031_),
    .A(net1046),
    .X(_1033_));
 sg13g2_nor2_2 _4450_ (.A(net1032),
    .B(_1032_),
    .Y(_1034_));
 sg13g2_nand2_2 _4451_ (.Y(_1035_),
    .A(_1027_),
    .B(_1033_));
 sg13g2_o21ai_1 _4452_ (.B1(net1106),
    .Y(_1036_),
    .A1(\dtop.vtop.pipeline.phases[1][10] ),
    .A2(net1104));
 sg13g2_a22oi_1 _4453_ (.Y(_1037_),
    .B1(net1093),
    .B2(\dtop.vtop.pipeline.phases[2][10] ),
    .A2(net1094),
    .A1(\dtop.vtop.pipeline.zg_acc[3] ));
 sg13g2_a22oi_1 _4454_ (.Y(_1038_),
    .B1(_1036_),
    .B2(_1037_),
    .A2(net1096),
    .A1(_0029_));
 sg13g2_xor2_1 _4455_ (.B(_1038_),
    .A(net1046),
    .X(_1039_));
 sg13g2_xnor2_1 _4456_ (.Y(_1040_),
    .A(net1046),
    .B(_1038_));
 sg13g2_a22oi_1 _4457_ (.Y(_1041_),
    .B1(_1010_),
    .B2(\dtop.vtop.pipeline.phases[2][11] ),
    .A2(net1094),
    .A1(\dtop.vtop.pipeline.zg_acc[4] ));
 sg13g2_o21ai_1 _4458_ (.B1(net1108),
    .Y(_1042_),
    .A1(\dtop.vtop.pipeline.phases[1][11] ),
    .A2(net1103));
 sg13g2_a22oi_1 _4459_ (.Y(_1043_),
    .B1(_1041_),
    .B2(_1042_),
    .A2(net1097),
    .A1(_0031_));
 sg13g2_xor2_1 _4460_ (.B(_1043_),
    .A(net1046),
    .X(_1044_));
 sg13g2_xnor2_1 _4461_ (.Y(_1045_),
    .A(net1046),
    .B(_1043_));
 sg13g2_nand2_2 _4462_ (.Y(_1046_),
    .A(net1028),
    .B(net1022));
 sg13g2_o21ai_1 _4463_ (.B1(net1106),
    .Y(_1047_),
    .A1(\dtop.vtop.pipeline.phases[1][9] ),
    .A2(net1104));
 sg13g2_a22oi_1 _4464_ (.Y(_1048_),
    .B1(_1010_),
    .B2(\dtop.vtop.pipeline.phases[2][9] ),
    .A2(net1094),
    .A1(\dtop.vtop.pipeline.zg_acc[2] ));
 sg13g2_a22oi_1 _4465_ (.Y(_1049_),
    .B1(_1047_),
    .B2(_1048_),
    .A2(net1097),
    .A1(_0027_));
 sg13g2_nand2_1 _4466_ (.Y(_1050_),
    .A(_1021_),
    .B(_1049_));
 sg13g2_or2_1 _4467_ (.X(_1051_),
    .B(_1049_),
    .A(_1021_));
 sg13g2_nand3_1 _4468_ (.B(net1060),
    .C(_1049_),
    .A(net1061),
    .Y(_1052_));
 sg13g2_a21o_1 _4469_ (.A2(net1060),
    .A1(net1061),
    .B1(_1049_),
    .X(_1053_));
 sg13g2_nand2_1 _4470_ (.Y(_1054_),
    .A(_1052_),
    .B(_1053_));
 sg13g2_and2_1 _4471_ (.A(_1052_),
    .B(_1053_),
    .X(_1055_));
 sg13g2_and2_1 _4472_ (.A(_0022_),
    .B(net1097),
    .X(_1056_));
 sg13g2_o21ai_1 _4473_ (.B1(net1103),
    .Y(_1057_),
    .A1(\dtop.vtop.pipeline.phases[2][7] ),
    .A2(net1108));
 sg13g2_a22oi_1 _4474_ (.Y(_1058_),
    .B1(net1094),
    .B2(\dtop.vtop.pipeline.zg_acc[0] ),
    .A2(net1108),
    .A1(\dtop.vtop.pipeline.phases[1][7] ));
 sg13g2_a21oi_2 _4475_ (.B1(_1056_),
    .Y(_1059_),
    .A2(_1058_),
    .A1(_1057_));
 sg13g2_a21o_2 _4476_ (.A2(_1058_),
    .A1(_1057_),
    .B1(_1056_),
    .X(_1060_));
 sg13g2_o21ai_1 _4477_ (.B1(_1059_),
    .Y(_1061_),
    .A1(_1017_),
    .A2(_1019_));
 sg13g2_nand3_1 _4478_ (.B(net1060),
    .C(_1060_),
    .A(net1061),
    .Y(_1062_));
 sg13g2_nand3_1 _4479_ (.B(net1060),
    .C(_1059_),
    .A(net1061),
    .Y(_1063_));
 sg13g2_o21ai_1 _4480_ (.B1(_1060_),
    .Y(_1064_),
    .A1(_1017_),
    .A2(_1019_));
 sg13g2_nand2_2 _4481_ (.Y(_1065_),
    .A(_1063_),
    .B(_1064_));
 sg13g2_nand2_2 _4482_ (.Y(_1066_),
    .A(_1061_),
    .B(_1062_));
 sg13g2_a221oi_1 _4483_ (.B2(\dtop.vtop.pipeline.phases[1][6] ),
    .C1(net1095),
    .B1(_1022_),
    .A1(\dtop.vtop.pipeline.phases[2][6] ),
    .Y(_1067_),
    .A2(net1093));
 sg13g2_a21oi_2 _4484_ (.B1(_1067_),
    .Y(_1068_),
    .A2(net1095),
    .A1(_0020_));
 sg13g2_a21o_2 _4485_ (.A2(net1096),
    .A1(_0020_),
    .B1(_1067_),
    .X(_1069_));
 sg13g2_nand3_1 _4486_ (.B(net1060),
    .C(_1068_),
    .A(net1061),
    .Y(_1070_));
 sg13g2_o21ai_1 _4487_ (.B1(_1069_),
    .Y(_1071_),
    .A1(_1017_),
    .A2(_1019_));
 sg13g2_o21ai_1 _4488_ (.B1(_1068_),
    .Y(_1072_),
    .A1(_1017_),
    .A2(_1019_));
 sg13g2_nand3_1 _4489_ (.B(_1020_),
    .C(_1069_),
    .A(_1018_),
    .Y(_1073_));
 sg13g2_nand2_1 _4490_ (.Y(_1074_),
    .A(_1072_),
    .B(_1073_));
 sg13g2_nand2_2 _4491_ (.Y(_1075_),
    .A(_1070_),
    .B(_1071_));
 sg13g2_nand4_1 _4492_ (.B(_1064_),
    .C(_1070_),
    .A(_1063_),
    .Y(_1076_),
    .D(_1071_));
 sg13g2_and2_1 _4493_ (.A(net1017),
    .B(_1076_),
    .X(_1077_));
 sg13g2_a22oi_1 _4494_ (.Y(_1078_),
    .B1(_1070_),
    .B2(_1071_),
    .A2(_1064_),
    .A1(_1063_));
 sg13g2_nand4_1 _4495_ (.B(_1062_),
    .C(_1072_),
    .A(_1061_),
    .Y(_1079_),
    .D(_1073_));
 sg13g2_a22oi_1 _4496_ (.Y(_1080_),
    .B1(_1070_),
    .B2(_1071_),
    .A2(_1062_),
    .A1(_1061_));
 sg13g2_a22oi_1 _4497_ (.Y(_1081_),
    .B1(_1072_),
    .B2(_1073_),
    .A2(_1064_),
    .A1(_1063_));
 sg13g2_xnor2_1 _4498_ (.Y(_1082_),
    .A(_1059_),
    .B(_1068_));
 sg13g2_xnor2_1 _4499_ (.Y(_1083_),
    .A(_1060_),
    .B(_1068_));
 sg13g2_nor2_1 _4500_ (.A(net1013),
    .B(_1082_),
    .Y(_1084_));
 sg13g2_a22oi_1 _4501_ (.Y(_1085_),
    .B1(_1010_),
    .B2(\dtop.vtop.pipeline.phases[2][8] ),
    .A2(net1094),
    .A1(_2697_));
 sg13g2_o21ai_1 _4502_ (.B1(net1106),
    .Y(_1086_),
    .A1(\dtop.vtop.pipeline.phases[1][8] ),
    .A2(net1104));
 sg13g2_a22oi_1 _4503_ (.Y(_1087_),
    .B1(_1085_),
    .B2(_1086_),
    .A2(net1097),
    .A1(_0024_));
 sg13g2_o21ai_1 _4504_ (.B1(_1087_),
    .Y(_1088_),
    .A1(_1017_),
    .A2(_1019_));
 sg13g2_or3_1 _4505_ (.A(_1017_),
    .B(_1019_),
    .C(_1087_),
    .X(_1089_));
 sg13g2_nand3_1 _4506_ (.B(net1060),
    .C(_1087_),
    .A(net1061),
    .Y(_1090_));
 sg13g2_a21o_2 _4507_ (.A2(net1060),
    .A1(net1061),
    .B1(_1087_),
    .X(_1091_));
 sg13g2_nand2_1 _4508_ (.Y(_1092_),
    .A(_1090_),
    .B(_1091_));
 sg13g2_nand2_2 _4509_ (.Y(_1093_),
    .A(_1088_),
    .B(_1089_));
 sg13g2_a22oi_1 _4510_ (.Y(_1094_),
    .B1(_1088_),
    .B2(_1089_),
    .A2(_1064_),
    .A1(_1063_));
 sg13g2_nand2b_1 _4511_ (.Y(_1095_),
    .B(net1009),
    .A_N(_1080_));
 sg13g2_nand2_1 _4512_ (.Y(_1096_),
    .A(_1082_),
    .B(net1009));
 sg13g2_nand2_1 _4513_ (.Y(_1097_),
    .A(_1079_),
    .B(net1012));
 sg13g2_xnor2_1 _4514_ (.Y(_1098_),
    .A(_1083_),
    .B(net1011));
 sg13g2_inv_1 _4515_ (.Y(_1099_),
    .A(_1098_));
 sg13g2_a21oi_1 _4516_ (.A1(net1013),
    .A2(_1098_),
    .Y(_1100_),
    .B1(_1084_));
 sg13g2_or2_1 _4517_ (.X(_1101_),
    .B(_1100_),
    .A(_1046_));
 sg13g2_nor2_1 _4518_ (.A(net1030),
    .B(_1080_),
    .Y(_1102_));
 sg13g2_nand2_1 _4519_ (.Y(_1103_),
    .A(net1028),
    .B(_1082_));
 sg13g2_nand4_1 _4520_ (.B(_1064_),
    .C(_1090_),
    .A(_1063_),
    .Y(_1104_),
    .D(_1091_));
 sg13g2_nor2_1 _4521_ (.A(_1078_),
    .B(net1011),
    .Y(_1105_));
 sg13g2_nor2_1 _4522_ (.A(net1018),
    .B(net1011),
    .Y(_1106_));
 sg13g2_nand4_1 _4523_ (.B(_1053_),
    .C(_1090_),
    .A(_1052_),
    .Y(_1107_),
    .D(_1091_));
 sg13g2_nor2_2 _4524_ (.A(_1078_),
    .B(net1007),
    .Y(_1108_));
 sg13g2_or2_1 _4525_ (.X(_1109_),
    .B(_1108_),
    .A(_1103_));
 sg13g2_a21oi_1 _4526_ (.A1(net1031),
    .A2(_1083_),
    .Y(_1110_),
    .B1(net1022));
 sg13g2_nor2_2 _4527_ (.A(net1030),
    .B(net1023),
    .Y(_1111_));
 sg13g2_nor2_2 _4528_ (.A(net1026),
    .B(net1022),
    .Y(_1112_));
 sg13g2_nor2_1 _4529_ (.A(net1025),
    .B(net1020),
    .Y(_1113_));
 sg13g2_nand2_1 _4530_ (.Y(_1114_),
    .A(net1031),
    .B(net1024));
 sg13g2_mux2_1 _4531_ (.A0(_1075_),
    .A1(_1082_),
    .S(net1011),
    .X(_1115_));
 sg13g2_mux2_1 _4532_ (.A0(_1083_),
    .A1(_1115_),
    .S(net1018),
    .X(_1116_));
 sg13g2_a22oi_1 _4533_ (.Y(_1117_),
    .B1(_1113_),
    .B2(_1116_),
    .A2(_1110_),
    .A1(_1109_));
 sg13g2_a21o_1 _4534_ (.A2(_1117_),
    .A1(_1101_),
    .B1(_1035_),
    .X(_1118_));
 sg13g2_mux2_1 _4535_ (.A0(_1098_),
    .A1(_1115_),
    .S(net1018),
    .X(_1119_));
 sg13g2_nand2b_1 _4536_ (.Y(_1120_),
    .B(net1012),
    .A_N(_1081_));
 sg13g2_a21oi_2 _4537_ (.B1(_1083_),
    .Y(_1121_),
    .A2(_1091_),
    .A1(_1090_));
 sg13g2_a21oi_2 _4538_ (.B1(_1121_),
    .Y(_1122_),
    .A2(net1010),
    .A1(_1074_));
 sg13g2_nor2_1 _4539_ (.A(_1066_),
    .B(net1009),
    .Y(_1123_));
 sg13g2_nand4_1 _4540_ (.B(_1062_),
    .C(_1088_),
    .A(_1061_),
    .Y(_1124_),
    .D(_1089_));
 sg13g2_and2_1 _4541_ (.A(net1013),
    .B(_1104_),
    .X(_1125_));
 sg13g2_xnor2_1 _4542_ (.Y(_1126_),
    .A(_1059_),
    .B(_1087_));
 sg13g2_xnor2_1 _4543_ (.Y(_1127_),
    .A(_1060_),
    .B(_1087_));
 sg13g2_nand2_2 _4544_ (.Y(_1128_),
    .A(net1013),
    .B(_1127_));
 sg13g2_xnor2_1 _4545_ (.Y(_1129_),
    .A(_1122_),
    .B(_1128_));
 sg13g2_nand2_2 _4546_ (.Y(_1130_),
    .A(net1032),
    .B(_1033_));
 sg13g2_mux4_1 _4547_ (.S0(net1020),
    .A0(_1099_),
    .A1(_1116_),
    .A2(_1129_),
    .A3(_1119_),
    .S1(net1031),
    .X(_1131_));
 sg13g2_or2_1 _4548_ (.X(_1132_),
    .B(_1131_),
    .A(_1130_));
 sg13g2_a21oi_1 _4549_ (.A1(_1066_),
    .A2(net1011),
    .Y(_1133_),
    .B1(net1015));
 sg13g2_o21ai_1 _4550_ (.B1(net1019),
    .Y(_1134_),
    .A1(_1065_),
    .A2(net1010));
 sg13g2_xnor2_1 _4551_ (.Y(_1135_),
    .A(_1122_),
    .B(_1133_));
 sg13g2_a21oi_1 _4552_ (.A1(net1014),
    .A2(_1115_),
    .Y(_1136_),
    .B1(_1084_));
 sg13g2_nand2_1 _4553_ (.Y(_1137_),
    .A(net1019),
    .B(_1065_));
 sg13g2_nor3_1 _4554_ (.A(net1031),
    .B(net1013),
    .C(_1124_),
    .Y(_1138_));
 sg13g2_xnor2_1 _4555_ (.Y(_1139_),
    .A(_1075_),
    .B(_1138_));
 sg13g2_nand2_2 _4556_ (.Y(_1140_),
    .A(_1027_),
    .B(_1032_));
 sg13g2_a221oi_1 _4557_ (.B2(net1020),
    .C1(_1140_),
    .B1(_1139_),
    .A1(_1113_),
    .Y(_1141_),
    .A2(_1136_));
 sg13g2_o21ai_1 _4558_ (.B1(_1141_),
    .Y(_1142_),
    .A1(_1046_),
    .A2(_1135_));
 sg13g2_nor2_1 _4559_ (.A(net1018),
    .B(_1094_),
    .Y(_1143_));
 sg13g2_or2_1 _4560_ (.X(_1144_),
    .B(_1094_),
    .A(net1017));
 sg13g2_nand3_1 _4561_ (.B(_1127_),
    .C(_1144_),
    .A(net1028),
    .Y(_1145_));
 sg13g2_and2_1 _4562_ (.A(net1030),
    .B(net1007),
    .X(_1146_));
 sg13g2_nand2_1 _4563_ (.Y(_1147_),
    .A(net1030),
    .B(net1018));
 sg13g2_a21oi_2 _4564_ (.B1(net1028),
    .Y(_1148_),
    .A2(_1066_),
    .A1(net1014));
 sg13g2_a21oi_2 _4565_ (.B1(net1026),
    .Y(_1149_),
    .A2(_1124_),
    .A1(net1014));
 sg13g2_nand2_1 _4566_ (.Y(_1150_),
    .A(net1007),
    .B(_1148_));
 sg13g2_nor4_2 _4567_ (.A(_1027_),
    .B(_1033_),
    .C(net1021),
    .Y(_1151_),
    .D(_1149_));
 sg13g2_nand3_1 _4568_ (.B(_1137_),
    .C(_1144_),
    .A(net1027),
    .Y(_1152_));
 sg13g2_nand3_1 _4569_ (.B(_1032_),
    .C(net1021),
    .A(net1032),
    .Y(_1153_));
 sg13g2_a21oi_1 _4570_ (.A1(_1134_),
    .A2(_1148_),
    .Y(_1154_),
    .B1(_1153_));
 sg13g2_a22oi_1 _4571_ (.Y(_1155_),
    .B1(_1152_),
    .B2(_1154_),
    .A2(_1151_),
    .A1(_1145_));
 sg13g2_nand4_1 _4572_ (.B(_1132_),
    .C(_1142_),
    .A(_1118_),
    .Y(_1156_),
    .D(_1155_));
 sg13g2_xnor2_1 _4573_ (.Y(_1157_),
    .A(net1047),
    .B(_1156_));
 sg13g2_xor2_1 _4574_ (.B(_1156_),
    .A(net1047),
    .X(_1158_));
 sg13g2_a22oi_1 _4575_ (.Y(_1159_),
    .B1(_1090_),
    .B2(_1091_),
    .A2(_1053_),
    .A1(_1052_));
 sg13g2_nand2_2 _4576_ (.Y(_1160_),
    .A(net1016),
    .B(_1104_));
 sg13g2_and2_1 _4577_ (.A(net1016),
    .B(_1104_),
    .X(_1161_));
 sg13g2_nor2_1 _4578_ (.A(net1030),
    .B(net1018),
    .Y(_1162_));
 sg13g2_nand2_1 _4579_ (.Y(_1163_),
    .A(net1027),
    .B(net1013));
 sg13g2_a221oi_1 _4580_ (.B2(_1147_),
    .C1(_1082_),
    .B1(_1163_),
    .A1(net1007),
    .Y(_1164_),
    .A2(_1160_));
 sg13g2_nand2_1 _4581_ (.Y(_1165_),
    .A(_1080_),
    .B(net1012));
 sg13g2_and2_1 _4582_ (.A(_1095_),
    .B(_1165_),
    .X(_1166_));
 sg13g2_nor2_1 _4583_ (.A(_1164_),
    .B(_1166_),
    .Y(_1167_));
 sg13g2_a21o_1 _4584_ (.A2(_1166_),
    .A1(_1164_),
    .B1(net1020),
    .X(_1168_));
 sg13g2_nand2_1 _4585_ (.Y(_1169_),
    .A(_1081_),
    .B(net1009));
 sg13g2_xnor2_1 _4586_ (.Y(_1170_),
    .A(_1081_),
    .B(net1012));
 sg13g2_a221oi_1 _4587_ (.B2(_1103_),
    .C1(net1022),
    .B1(_1170_),
    .A1(net1027),
    .Y(_1171_),
    .A2(_1121_));
 sg13g2_nor2b_1 _4588_ (.A(_1171_),
    .B_N(_1034_),
    .Y(_1172_));
 sg13g2_o21ai_1 _4589_ (.B1(_1172_),
    .Y(_1173_),
    .A1(_1167_),
    .A2(_1168_));
 sg13g2_mux2_1 _4590_ (.A0(_1079_),
    .A1(_1082_),
    .S(net1010),
    .X(_1174_));
 sg13g2_a21o_1 _4591_ (.A2(_1104_),
    .A1(_1082_),
    .B1(net1014),
    .X(_1175_));
 sg13g2_a221oi_1 _4592_ (.B2(_1175_),
    .C1(_1114_),
    .B1(_1174_),
    .A1(_1084_),
    .Y(_1176_),
    .A2(net1009));
 sg13g2_nor2_1 _4593_ (.A(_1079_),
    .B(net1009),
    .Y(_1177_));
 sg13g2_nand2_1 _4594_ (.Y(_1178_),
    .A(_1078_),
    .B(net1011));
 sg13g2_a221oi_1 _4595_ (.B2(net1012),
    .C1(_1094_),
    .B1(_1078_),
    .A1(_1050_),
    .Y(_1179_),
    .A2(_1051_));
 sg13g2_a221oi_1 _4596_ (.B2(_1178_),
    .C1(_1046_),
    .B1(_1143_),
    .A1(_1096_),
    .Y(_1180_),
    .A2(_1133_));
 sg13g2_nand2_1 _4597_ (.Y(_1181_),
    .A(net1021),
    .B(_1083_));
 sg13g2_a21oi_1 _4598_ (.A1(_1102_),
    .A2(_1159_),
    .Y(_1182_),
    .B1(_1181_));
 sg13g2_or4_1 _4599_ (.A(net1032),
    .B(_1176_),
    .C(_1180_),
    .D(_1182_),
    .X(_1183_));
 sg13g2_o21ai_1 _4600_ (.B1(net1026),
    .Y(_1184_),
    .A1(net1013),
    .A2(_1124_));
 sg13g2_nand2_1 _4601_ (.Y(_1185_),
    .A(net1023),
    .B(_1184_));
 sg13g2_o21ai_1 _4602_ (.B1(net1022),
    .Y(_1186_),
    .A1(_1106_),
    .A2(_1184_));
 sg13g2_nand2_1 _4603_ (.Y(_1187_),
    .A(net1016),
    .B(_1124_));
 sg13g2_nand3_1 _4604_ (.B(_1112_),
    .C(_1187_),
    .A(net1007),
    .Y(_1188_));
 sg13g2_nand3_1 _4605_ (.B(_1111_),
    .C(_1127_),
    .A(net1008),
    .Y(_1189_));
 sg13g2_nand4_1 _4606_ (.B(_1186_),
    .C(_1188_),
    .A(net1032),
    .Y(_1190_),
    .D(_1189_));
 sg13g2_nand3_1 _4607_ (.B(_1183_),
    .C(_1190_),
    .A(_1032_),
    .Y(_1191_));
 sg13g2_nand4_1 _4608_ (.B(net1017),
    .C(_1076_),
    .A(net1027),
    .Y(_1192_),
    .D(_1127_));
 sg13g2_o21ai_1 _4609_ (.B1(_1192_),
    .Y(_1193_),
    .A1(_1163_),
    .A2(_1170_));
 sg13g2_nor2_1 _4610_ (.A(net1017),
    .B(_1081_),
    .Y(_1194_));
 sg13g2_a221oi_1 _4611_ (.B2(_1095_),
    .C1(net1027),
    .B1(_1194_),
    .A1(_1077_),
    .Y(_1195_),
    .A2(_1127_));
 sg13g2_nor2_1 _4612_ (.A(net1023),
    .B(_1130_),
    .Y(_1196_));
 sg13g2_nor4_1 _4613_ (.A(net1024),
    .B(_1130_),
    .C(_1193_),
    .D(_1195_),
    .Y(_1197_));
 sg13g2_a221oi_1 _4614_ (.B2(_1074_),
    .C1(net1014),
    .B1(_1094_),
    .A1(_1080_),
    .Y(_1198_),
    .A2(net1011));
 sg13g2_a21oi_1 _4615_ (.A1(_1165_),
    .A2(_1169_),
    .Y(_1199_),
    .B1(net1017));
 sg13g2_o21ai_1 _4616_ (.B1(net1027),
    .Y(_1200_),
    .A1(_1198_),
    .A2(_1199_));
 sg13g2_nor2_1 _4617_ (.A(net1020),
    .B(_1130_),
    .Y(_1201_));
 sg13g2_a221oi_1 _4618_ (.B2(_1194_),
    .C1(net1027),
    .B1(_1165_),
    .A1(_1120_),
    .Y(_1202_),
    .A2(_1161_));
 sg13g2_nor2b_1 _4619_ (.A(_1202_),
    .B_N(_1201_),
    .Y(_1203_));
 sg13g2_a21oi_1 _4620_ (.A1(_1200_),
    .A2(_1203_),
    .Y(_1204_),
    .B1(_1197_));
 sg13g2_nand3_1 _4621_ (.B(_1191_),
    .C(_1204_),
    .A(_1173_),
    .Y(_1205_));
 sg13g2_xor2_1 _4622_ (.B(_1205_),
    .A(net1048),
    .X(_1206_));
 sg13g2_nand2_1 _4623_ (.Y(_1207_),
    .A(net1049),
    .B(_1206_));
 sg13g2_nand2_1 _4624_ (.Y(_1208_),
    .A(_0987_),
    .B(_1157_));
 sg13g2_nand3_1 _4625_ (.B(_1207_),
    .C(_1208_),
    .A(net1070),
    .Y(_1209_));
 sg13g2_nand4_1 _4626_ (.B(net1162),
    .C(net1208),
    .A(_2669_),
    .Y(_1210_),
    .D(net1111));
 sg13g2_nand2_1 _4627_ (.Y(_1211_),
    .A(net315),
    .B(net1088));
 sg13g2_o21ai_1 _4628_ (.B1(_1211_),
    .Y(_0104_),
    .A1(_1209_),
    .A2(net1088));
 sg13g2_and2_1 _4629_ (.A(net1030),
    .B(_1121_),
    .X(_1212_));
 sg13g2_nand2b_1 _4630_ (.Y(_1213_),
    .B(_1127_),
    .A_N(_1080_));
 sg13g2_nor3_1 _4631_ (.A(net1014),
    .B(_1080_),
    .C(_1126_),
    .Y(_1214_));
 sg13g2_xnor2_1 _4632_ (.Y(_1215_),
    .A(net1016),
    .B(_1213_));
 sg13g2_xnor2_1 _4633_ (.Y(_1216_),
    .A(_1212_),
    .B(_1215_));
 sg13g2_a21oi_2 _4634_ (.B1(net1031),
    .Y(_1217_),
    .A2(_1104_),
    .A1(net1015));
 sg13g2_a221oi_1 _4635_ (.B2(net1009),
    .C1(net1016),
    .B1(_1075_),
    .A1(_1061_),
    .Y(_1218_),
    .A2(_1062_));
 sg13g2_a221oi_1 _4636_ (.B2(_1217_),
    .C1(_1218_),
    .B1(_1187_),
    .A1(_1077_),
    .Y(_1219_),
    .A2(_1097_));
 sg13g2_o21ai_1 _4637_ (.B1(_1027_),
    .Y(_1220_),
    .A1(net1021),
    .A2(_1219_));
 sg13g2_a21o_1 _4638_ (.A2(_1216_),
    .A1(net1021),
    .B1(_1220_),
    .X(_1221_));
 sg13g2_a21oi_1 _4639_ (.A1(net1016),
    .A2(_1126_),
    .Y(_1222_),
    .B1(net1031));
 sg13g2_o21ai_1 _4640_ (.B1(_1222_),
    .Y(_1223_),
    .A1(_1198_),
    .A2(_1213_));
 sg13g2_a221oi_1 _4641_ (.B2(net1014),
    .C1(net1027),
    .B1(_1213_),
    .A1(_1079_),
    .Y(_1224_),
    .A2(_1159_));
 sg13g2_nand3b_1 _4642_ (.B(net1024),
    .C(_1223_),
    .Y(_1225_),
    .A_N(_1224_));
 sg13g2_o21ai_1 _4643_ (.B1(_1111_),
    .Y(_1226_),
    .A1(_1179_),
    .A2(_1214_));
 sg13g2_nand3_1 _4644_ (.B(_1128_),
    .C(_1134_),
    .A(_1112_),
    .Y(_1227_));
 sg13g2_and3_1 _4645_ (.X(_1228_),
    .A(net1032),
    .B(_1226_),
    .C(_1227_));
 sg13g2_a21oi_1 _4646_ (.A1(_1225_),
    .A2(_1228_),
    .Y(_1229_),
    .B1(_1032_));
 sg13g2_o21ai_1 _4647_ (.B1(net1016),
    .Y(_1230_),
    .A1(_1076_),
    .A2(net1012));
 sg13g2_o21ai_1 _4648_ (.B1(net1007),
    .Y(_1231_),
    .A1(_1123_),
    .A2(_1230_));
 sg13g2_or2_1 _4649_ (.X(_1232_),
    .B(_1231_),
    .A(_1046_));
 sg13g2_nor3_1 _4650_ (.A(_1105_),
    .B(_1138_),
    .C(_1177_),
    .Y(_1233_));
 sg13g2_nand2b_1 _4651_ (.Y(_1234_),
    .B(_1230_),
    .A_N(_1108_));
 sg13g2_a221oi_1 _4652_ (.B2(_1113_),
    .C1(net1032),
    .B1(_1234_),
    .A1(net1020),
    .Y(_1235_),
    .A2(_1233_));
 sg13g2_a221oi_1 _4653_ (.B2(_1147_),
    .C1(net1022),
    .B1(_1184_),
    .A1(_1124_),
    .Y(_1236_),
    .A2(_1162_));
 sg13g2_nor2_1 _4654_ (.A(_1046_),
    .B(net1007),
    .Y(_1237_));
 sg13g2_nor2_1 _4655_ (.A(_1236_),
    .B(_1237_),
    .Y(_1238_));
 sg13g2_a22oi_1 _4656_ (.Y(_1239_),
    .B1(_1238_),
    .B2(net1032),
    .A2(_1235_),
    .A1(_1232_));
 sg13g2_a22oi_1 _4657_ (.Y(_1240_),
    .B1(_1239_),
    .B2(_1032_),
    .A2(_1229_),
    .A1(_1221_));
 sg13g2_xnor2_1 _4658_ (.Y(_1241_),
    .A(net1047),
    .B(_1240_));
 sg13g2_xor2_1 _4659_ (.B(_1240_),
    .A(net1047),
    .X(_1242_));
 sg13g2_nand2_1 _4660_ (.Y(_1243_),
    .A(net1049),
    .B(_1241_));
 sg13g2_o21ai_1 _4661_ (.B1(_1243_),
    .Y(_1244_),
    .A1(net1049),
    .A2(_1206_));
 sg13g2_nor2_1 _4662_ (.A(net1071),
    .B(_0987_),
    .Y(_1245_));
 sg13g2_a22oi_1 _4663_ (.Y(_1246_),
    .B1(_1245_),
    .B2(_1158_),
    .A2(_1244_),
    .A1(net1070));
 sg13g2_nand2_1 _4664_ (.Y(_1247_),
    .A(net309),
    .B(net1088));
 sg13g2_o21ai_1 _4665_ (.B1(_1247_),
    .Y(_0105_),
    .A1(net1088),
    .A2(_1246_));
 sg13g2_nor2b_1 _4666_ (.A(_1046_),
    .B_N(_1231_),
    .Y(_1248_));
 sg13g2_o21ai_1 _4667_ (.B1(_1146_),
    .Y(_1249_),
    .A1(_1177_),
    .A2(_1230_));
 sg13g2_a21oi_1 _4668_ (.A1(_1076_),
    .A2(net1012),
    .Y(_1250_),
    .B1(net1016));
 sg13g2_nand3b_1 _4669_ (.B(_1160_),
    .C(_1112_),
    .Y(_1251_),
    .A_N(_1250_));
 sg13g2_o21ai_1 _4670_ (.B1(_1111_),
    .Y(_1252_),
    .A1(_1161_),
    .A2(_1250_));
 sg13g2_nand3_1 _4671_ (.B(_1251_),
    .C(_1252_),
    .A(_1249_),
    .Y(_1253_));
 sg13g2_o21ai_1 _4672_ (.B1(_1034_),
    .Y(_1254_),
    .A1(_1248_),
    .A2(_1253_));
 sg13g2_nor2_1 _4673_ (.A(net1025),
    .B(_1230_),
    .Y(_1255_));
 sg13g2_a21oi_2 _4674_ (.B1(net1013),
    .Y(_1256_),
    .A2(net1009),
    .A1(_1079_));
 sg13g2_o21ai_1 _4675_ (.B1(net1018),
    .Y(_1257_),
    .A1(_1078_),
    .A2(net1011));
 sg13g2_o21ai_1 _4676_ (.B1(net1020),
    .Y(_1258_),
    .A1(_1108_),
    .A2(_1256_));
 sg13g2_o21ai_1 _4677_ (.B1(_1258_),
    .Y(_1259_),
    .A1(_1186_),
    .A2(_1255_));
 sg13g2_nand2b_1 _4678_ (.Y(_1260_),
    .B(_1259_),
    .A_N(_1140_));
 sg13g2_nor3_1 _4679_ (.A(net1026),
    .B(_1159_),
    .C(_1250_),
    .Y(_1261_));
 sg13g2_o21ai_1 _4680_ (.B1(_1201_),
    .Y(_1262_),
    .A1(_1125_),
    .A2(_1184_));
 sg13g2_or2_1 _4681_ (.X(_1263_),
    .B(_1262_),
    .A(_1261_));
 sg13g2_o21ai_1 _4682_ (.B1(net1025),
    .Y(_1264_),
    .A1(_1106_),
    .A2(_1161_));
 sg13g2_o21ai_1 _4683_ (.B1(_1264_),
    .Y(_1265_),
    .A1(_1150_),
    .A2(_1159_));
 sg13g2_a21oi_1 _4684_ (.A1(_1124_),
    .A2(_1162_),
    .Y(_1266_),
    .B1(_1153_));
 sg13g2_a22oi_1 _4685_ (.Y(_1267_),
    .B1(_1266_),
    .B2(_1147_),
    .A2(_1265_),
    .A1(_1196_));
 sg13g2_nand4_1 _4686_ (.B(_1260_),
    .C(_1263_),
    .A(_1254_),
    .Y(_1268_),
    .D(_1267_));
 sg13g2_xnor2_1 _4687_ (.Y(_1269_),
    .A(net1047),
    .B(_1268_));
 sg13g2_xor2_1 _4688_ (.B(_1268_),
    .A(net1047),
    .X(_1270_));
 sg13g2_mux2_1 _4689_ (.A0(_1241_),
    .A1(_1270_),
    .S(net1049),
    .X(_1271_));
 sg13g2_mux4_1 _4690_ (.S0(net1049),
    .A0(_1157_),
    .A1(_1206_),
    .A2(_1242_),
    .A3(_1269_),
    .S1(net1070),
    .X(_1272_));
 sg13g2_nand2_1 _4691_ (.Y(_1273_),
    .A(net311),
    .B(net1089));
 sg13g2_o21ai_1 _4692_ (.B1(_1273_),
    .Y(_0106_),
    .A1(net1089),
    .A2(_1272_));
 sg13g2_a21oi_1 _4693_ (.A1(_1078_),
    .A2(_1159_),
    .Y(_1274_),
    .B1(net1025));
 sg13g2_a22oi_1 _4694_ (.Y(_1275_),
    .B1(_1274_),
    .B2(net1008),
    .A2(_1160_),
    .A1(net1025));
 sg13g2_o21ai_1 _4695_ (.B1(net1023),
    .Y(_1276_),
    .A1(net1030),
    .A2(_1230_));
 sg13g2_mux2_1 _4696_ (.A0(_1276_),
    .A1(net1023),
    .S(_1275_),
    .X(_1277_));
 sg13g2_and2_1 _4697_ (.A(_1034_),
    .B(_1277_),
    .X(_1278_));
 sg13g2_o21ai_1 _4698_ (.B1(net1022),
    .Y(_1279_),
    .A1(net1025),
    .A2(_1159_));
 sg13g2_a21oi_1 _4699_ (.A1(_1187_),
    .A2(_1217_),
    .Y(_1280_),
    .B1(_1279_));
 sg13g2_nor2_1 _4700_ (.A(net1023),
    .B(_1149_),
    .Y(_1281_));
 sg13g2_a221oi_1 _4701_ (.B2(net1025),
    .C1(net1022),
    .B1(_1160_),
    .A1(net1007),
    .Y(_1282_),
    .A2(_1148_));
 sg13g2_nor2_1 _4702_ (.A(_1130_),
    .B(_1281_),
    .Y(_1283_));
 sg13g2_nor3_1 _4703_ (.A(_1130_),
    .B(_1280_),
    .C(_1282_),
    .Y(_1284_));
 sg13g2_nor3_2 _4704_ (.A(_1123_),
    .B(_1153_),
    .C(_1163_),
    .Y(_1285_));
 sg13g2_nand2_1 _4705_ (.Y(_1286_),
    .A(net1030),
    .B(_1257_));
 sg13g2_a22oi_1 _4706_ (.Y(_1287_),
    .B1(_1256_),
    .B2(_1111_),
    .A2(_1184_),
    .A1(net1023));
 sg13g2_a21oi_1 _4707_ (.A1(_1286_),
    .A2(_1287_),
    .Y(_1288_),
    .B1(_1140_));
 sg13g2_nor4_2 _4708_ (.A(_1278_),
    .B(_1284_),
    .C(_1285_),
    .Y(_1289_),
    .D(_1288_));
 sg13g2_xor2_1 _4709_ (.B(_1289_),
    .A(net1047),
    .X(_1290_));
 sg13g2_xnor2_1 _4710_ (.Y(_1291_),
    .A(net1047),
    .B(_1289_));
 sg13g2_nor2_1 _4711_ (.A(net1049),
    .B(_1269_),
    .Y(_1292_));
 sg13g2_nor2_1 _4712_ (.A(_0987_),
    .B(_1290_),
    .Y(_1293_));
 sg13g2_mux4_1 _4713_ (.S0(net1049),
    .A0(_1206_),
    .A1(_1242_),
    .A2(_1269_),
    .A3(_1290_),
    .S1(net1070),
    .X(_1294_));
 sg13g2_nand2_1 _4714_ (.Y(_1295_),
    .A(net322),
    .B(net1089));
 sg13g2_o21ai_1 _4715_ (.B1(_1295_),
    .Y(_0107_),
    .A1(net1090),
    .A2(_1294_));
 sg13g2_and2_1 _4716_ (.A(_1111_),
    .B(_1257_),
    .X(_1296_));
 sg13g2_nor2_1 _4717_ (.A(_1140_),
    .B(_1296_),
    .Y(_1297_));
 sg13g2_or2_1 _4718_ (.X(_1298_),
    .B(_1297_),
    .A(_1283_));
 sg13g2_nor2_1 _4719_ (.A(_1274_),
    .B(_1276_),
    .Y(_1299_));
 sg13g2_a21oi_1 _4720_ (.A1(net1008),
    .A2(_1112_),
    .Y(_1300_),
    .B1(_1299_));
 sg13g2_a22oi_1 _4721_ (.Y(_1301_),
    .B1(_1300_),
    .B2(_1034_),
    .A2(_1298_),
    .A1(_1185_));
 sg13g2_xnor2_1 _4722_ (.Y(_1302_),
    .A(net1048),
    .B(_1301_));
 sg13g2_mux2_1 _4723_ (.A0(_1291_),
    .A1(_1302_),
    .S(_0988_),
    .X(_1303_));
 sg13g2_mux2_2 _4724_ (.A0(_1271_),
    .A1(_1303_),
    .S(net1070),
    .X(_1304_));
 sg13g2_mux2_1 _4725_ (.A0(_1304_),
    .A1(net407),
    .S(net1090),
    .X(_0108_));
 sg13g2_a21o_1 _4726_ (.A2(_1230_),
    .A1(net1025),
    .B1(net1020),
    .X(_1305_));
 sg13g2_a221oi_1 _4727_ (.B2(_1034_),
    .C1(_1283_),
    .B1(_1305_),
    .A1(_1027_),
    .Y(_1306_),
    .A2(_1296_));
 sg13g2_xor2_1 _4728_ (.B(_1306_),
    .A(net1048),
    .X(_1307_));
 sg13g2_nand2_1 _4729_ (.Y(_1308_),
    .A(_0988_),
    .B(_1307_));
 sg13g2_o21ai_1 _4730_ (.B1(_1308_),
    .Y(_1309_),
    .A1(net1049),
    .A2(_1302_));
 sg13g2_nor3_1 _4731_ (.A(net1070),
    .B(_1292_),
    .C(_1293_),
    .Y(_1310_));
 sg13g2_a21oi_2 _4732_ (.B1(_1310_),
    .Y(_1311_),
    .A2(_1309_),
    .A1(net1070));
 sg13g2_mux2_1 _4733_ (.A0(_1311_),
    .A1(net421),
    .S(net1089),
    .X(_0109_));
 sg13g2_o21ai_1 _4734_ (.B1(_1033_),
    .Y(_1312_),
    .A1(_1027_),
    .A2(_1281_));
 sg13g2_xnor2_1 _4735_ (.Y(_1313_),
    .A(net1048),
    .B(_1312_));
 sg13g2_nand2_1 _4736_ (.Y(_1314_),
    .A(_0987_),
    .B(_1307_));
 sg13g2_o21ai_1 _4737_ (.B1(_1314_),
    .Y(_1315_),
    .A1(_0987_),
    .A2(_1313_));
 sg13g2_inv_1 _4738_ (.Y(_1316_),
    .A(_1315_));
 sg13g2_nand2_1 _4739_ (.Y(_1317_),
    .A(net1071),
    .B(_1315_));
 sg13g2_o21ai_1 _4740_ (.B1(_1317_),
    .Y(_1318_),
    .A1(net1070),
    .A2(_1303_));
 sg13g2_nand2_1 _4741_ (.Y(_1319_),
    .A(net312),
    .B(net1089));
 sg13g2_o21ai_1 _4742_ (.B1(_1319_),
    .Y(_0110_),
    .A1(net1089),
    .A2(_1318_));
 sg13g2_nand2_1 _4743_ (.Y(_1320_),
    .A(_0987_),
    .B(_1313_));
 sg13g2_o21ai_1 _4744_ (.B1(_1320_),
    .Y(_1321_),
    .A1(_0987_),
    .A2(_0998_));
 sg13g2_nand2_1 _4745_ (.Y(_1322_),
    .A(net1071),
    .B(_1321_));
 sg13g2_o21ai_1 _4746_ (.B1(_1322_),
    .Y(_1323_),
    .A1(net1071),
    .A2(_1309_));
 sg13g2_mux2_1 _4747_ (.A0(_1323_),
    .A1(net413),
    .S(net1088),
    .X(_0111_));
 sg13g2_nand2_1 _4748_ (.Y(_1324_),
    .A(net1071),
    .B(_0998_));
 sg13g2_o21ai_1 _4749_ (.B1(_1324_),
    .Y(_1325_),
    .A1(net1071),
    .A2(_1316_));
 sg13g2_inv_1 _4750_ (.Y(_1326_),
    .A(_1325_));
 sg13g2_nand2_1 _4751_ (.Y(_1327_),
    .A(net310),
    .B(net1088));
 sg13g2_o21ai_1 _4752_ (.B1(_1327_),
    .Y(_0112_),
    .A1(net1090),
    .A2(_1325_));
 sg13g2_nand2_1 _4753_ (.Y(_1328_),
    .A(net316),
    .B(net1088));
 sg13g2_o21ai_1 _4754_ (.B1(_1324_),
    .Y(_1329_),
    .A1(net1071),
    .A2(_1321_));
 sg13g2_o21ai_1 _4755_ (.B1(_1328_),
    .Y(_0113_),
    .A1(net1088),
    .A2(_1329_));
 sg13g2_nand2_1 _4756_ (.Y(_1330_),
    .A(net308),
    .B(net1089));
 sg13g2_o21ai_1 _4757_ (.B1(_1330_),
    .Y(_0114_),
    .A1(net1089),
    .A2(_1329_));
 sg13g2_nand3_1 _4758_ (.B(net1162),
    .C(net1114),
    .A(net1220),
    .Y(_1331_));
 sg13g2_nand4_1 _4759_ (.B(net1162),
    .C(net1208),
    .A(net1220),
    .Y(_1332_),
    .D(net1111));
 sg13g2_nand2_1 _4760_ (.Y(_1333_),
    .A(net329),
    .B(net1085));
 sg13g2_o21ai_1 _4761_ (.B1(_1333_),
    .Y(_0115_),
    .A1(_1209_),
    .A2(net1085));
 sg13g2_nand2_1 _4762_ (.Y(_1334_),
    .A(net366),
    .B(net1086));
 sg13g2_o21ai_1 _4763_ (.B1(_1334_),
    .Y(_0116_),
    .A1(_1246_),
    .A2(net1085));
 sg13g2_nand2_1 _4764_ (.Y(_1335_),
    .A(net367),
    .B(net1087));
 sg13g2_o21ai_1 _4765_ (.B1(_1335_),
    .Y(_0117_),
    .A1(_1272_),
    .A2(net1087));
 sg13g2_nand2_1 _4766_ (.Y(_1336_),
    .A(net385),
    .B(net1087));
 sg13g2_o21ai_1 _4767_ (.B1(_1336_),
    .Y(_0118_),
    .A1(_1294_),
    .A2(net1087));
 sg13g2_mux2_1 _4768_ (.A0(_1304_),
    .A1(net460),
    .S(net1086),
    .X(_0119_));
 sg13g2_mux2_1 _4769_ (.A0(_1311_),
    .A1(net476),
    .S(net1086),
    .X(_0120_));
 sg13g2_nand2_1 _4770_ (.Y(_1337_),
    .A(net320),
    .B(net1086));
 sg13g2_o21ai_1 _4771_ (.B1(_1337_),
    .Y(_0121_),
    .A1(_1318_),
    .A2(net1086));
 sg13g2_mux2_1 _4772_ (.A0(_1323_),
    .A1(net493),
    .S(net1085),
    .X(_0122_));
 sg13g2_nand2_1 _4773_ (.Y(_1338_),
    .A(net334),
    .B(net1085));
 sg13g2_o21ai_1 _4774_ (.B1(_1338_),
    .Y(_0123_),
    .A1(_1325_),
    .A2(net1085));
 sg13g2_nand2_1 _4775_ (.Y(_1339_),
    .A(net341),
    .B(net1085));
 sg13g2_o21ai_1 _4776_ (.B1(_1339_),
    .Y(_0124_),
    .A1(_1329_),
    .A2(net1085));
 sg13g2_nand2_1 _4777_ (.Y(_1340_),
    .A(net463),
    .B(net1087));
 sg13g2_o21ai_1 _4778_ (.B1(_1340_),
    .Y(_0125_),
    .A1(_0998_),
    .A2(net1087));
 sg13g2_nand4_1 _4779_ (.B(net1215),
    .C(net1208),
    .A(_2669_),
    .Y(_1341_),
    .D(net1111));
 sg13g2_nand2_1 _4780_ (.Y(_1342_),
    .A(net370),
    .B(net1083));
 sg13g2_o21ai_1 _4781_ (.B1(_1342_),
    .Y(_0126_),
    .A1(_1209_),
    .A2(net1082));
 sg13g2_nand2_1 _4782_ (.Y(_1343_),
    .A(net388),
    .B(net1082));
 sg13g2_o21ai_1 _4783_ (.B1(_1343_),
    .Y(_0127_),
    .A1(_1246_),
    .A2(net1082));
 sg13g2_nand2_1 _4784_ (.Y(_1344_),
    .A(net335),
    .B(net1083));
 sg13g2_o21ai_1 _4785_ (.B1(_1344_),
    .Y(_0128_),
    .A1(_1272_),
    .A2(net1083));
 sg13g2_nand2_1 _4786_ (.Y(_1345_),
    .A(net453),
    .B(net1083));
 sg13g2_o21ai_1 _4787_ (.B1(_1345_),
    .Y(_0129_),
    .A1(_1294_),
    .A2(net1084));
 sg13g2_mux2_1 _4788_ (.A0(_1304_),
    .A1(net488),
    .S(net1084),
    .X(_0130_));
 sg13g2_mux2_1 _4789_ (.A0(_1311_),
    .A1(net487),
    .S(net1083),
    .X(_0131_));
 sg13g2_nand2_1 _4790_ (.Y(_1346_),
    .A(net323),
    .B(net1083));
 sg13g2_o21ai_1 _4791_ (.B1(_1346_),
    .Y(_0132_),
    .A1(_1318_),
    .A2(net1083));
 sg13g2_mux2_1 _4792_ (.A0(_1323_),
    .A1(net458),
    .S(net1082),
    .X(_0133_));
 sg13g2_nand2_1 _4793_ (.Y(_1347_),
    .A(net343),
    .B(net1082));
 sg13g2_o21ai_1 _4794_ (.B1(_1347_),
    .Y(_0134_),
    .A1(_1325_),
    .A2(net1082));
 sg13g2_nand2_1 _4795_ (.Y(_1348_),
    .A(net358),
    .B(net1082));
 sg13g2_o21ai_1 _4796_ (.B1(_1348_),
    .Y(_0135_),
    .A1(_1329_),
    .A2(net1082));
 sg13g2_nand2_1 _4797_ (.Y(_1349_),
    .A(net321),
    .B(net1084));
 sg13g2_o21ai_1 _4798_ (.B1(_1349_),
    .Y(_0136_),
    .A1(_1329_),
    .A2(net1084));
 sg13g2_nand2_1 _4799_ (.Y(_1350_),
    .A(_0537_),
    .B(_0564_));
 sg13g2_nor2_1 _4800_ (.A(net1119),
    .B(_0518_),
    .Y(_1351_));
 sg13g2_nand2_1 _4801_ (.Y(_1352_),
    .A(_2914_),
    .B(_0517_));
 sg13g2_nand2b_1 _4802_ (.Y(_1353_),
    .B(net1036),
    .A_N(net1053));
 sg13g2_a21oi_1 _4803_ (.A1(net1119),
    .A2(_0622_),
    .Y(_1354_),
    .B1(_0623_));
 sg13g2_nor2_1 _4804_ (.A(_0513_),
    .B(_0651_),
    .Y(_1355_));
 sg13g2_nor2_1 _4805_ (.A(_1354_),
    .B(_1355_),
    .Y(_1356_));
 sg13g2_nand2b_1 _4806_ (.Y(_1357_),
    .B(_1356_),
    .A_N(_1353_));
 sg13g2_nor2_1 _4807_ (.A(_0568_),
    .B(_1353_),
    .Y(_1358_));
 sg13g2_o21ai_1 _4808_ (.B1(net1120),
    .Y(_1359_),
    .A1(net1234),
    .A2(net2));
 sg13g2_a21oi_1 _4809_ (.A1(net1142),
    .A2(_1359_),
    .Y(_1360_),
    .B1(net1036));
 sg13g2_nor3_2 _4810_ (.A(_0537_),
    .B(_1358_),
    .C(_1360_),
    .Y(_1361_));
 sg13g2_a21oi_1 _4811_ (.A1(_0603_),
    .A2(_0655_),
    .Y(_1362_),
    .B1(_0598_));
 sg13g2_nand2_1 _4812_ (.Y(_1363_),
    .A(_0608_),
    .B(_0655_));
 sg13g2_a21oi_1 _4813_ (.A1(_0598_),
    .A2(_1363_),
    .Y(_1364_),
    .B1(_1362_));
 sg13g2_and2_1 _4814_ (.A(net1),
    .B(net1120),
    .X(_1365_));
 sg13g2_o21ai_1 _4815_ (.B1(_1364_),
    .Y(_1366_),
    .A1(net3),
    .A2(_2882_));
 sg13g2_or2_1 _4816_ (.X(_1367_),
    .B(_1366_),
    .A(_1365_));
 sg13g2_nand2_1 _4817_ (.Y(_1368_),
    .A(_0871_),
    .B(_1367_));
 sg13g2_nand2_1 _4818_ (.Y(_1369_),
    .A(_2684_),
    .B(_0535_));
 sg13g2_nand4_1 _4819_ (.B(_1361_),
    .C(_1368_),
    .A(_1357_),
    .Y(_1370_),
    .D(_1369_));
 sg13g2_o21ai_1 _4820_ (.B1(_1370_),
    .Y(_1371_),
    .A1(_1350_),
    .A2(_1352_));
 sg13g2_or2_1 _4821_ (.X(_1372_),
    .B(_1356_),
    .A(_1353_));
 sg13g2_nand2_1 _4822_ (.Y(_1373_),
    .A(_0659_),
    .B(_1362_));
 sg13g2_nand2_1 _4823_ (.Y(_1374_),
    .A(_0609_),
    .B(_0613_));
 sg13g2_nand2_1 _4824_ (.Y(_1375_),
    .A(_1363_),
    .B(_1374_));
 sg13g2_nor2_1 _4825_ (.A(_2878_),
    .B(_0600_),
    .Y(_1376_));
 sg13g2_xor2_1 _4826_ (.B(_1376_),
    .A(_1375_),
    .X(_1377_));
 sg13g2_o21ai_1 _4827_ (.B1(_1373_),
    .Y(_1378_),
    .A1(_0597_),
    .A2(_1377_));
 sg13g2_nor3_1 _4828_ (.A(net1),
    .B(net3),
    .C(_2882_),
    .Y(_1379_));
 sg13g2_nand3b_1 _4829_ (.B(_1378_),
    .C(_1379_),
    .Y(_1380_),
    .A_N(_1364_));
 sg13g2_nand3_1 _4830_ (.B(_1367_),
    .C(_1380_),
    .A(_0871_),
    .Y(_1381_));
 sg13g2_nand2b_1 _4831_ (.Y(_1382_),
    .B(_0535_),
    .A_N(_0079_));
 sg13g2_nand4_1 _4832_ (.B(_1372_),
    .C(_1381_),
    .A(_1361_),
    .Y(_1383_),
    .D(_1382_));
 sg13g2_a21oi_1 _4833_ (.A1(_1364_),
    .A2(_1379_),
    .Y(_1384_),
    .B1(_1378_));
 sg13g2_o21ai_1 _4834_ (.B1(_0871_),
    .Y(_1385_),
    .A1(_1365_),
    .A2(_1384_));
 sg13g2_a22oi_1 _4835_ (.Y(_1386_),
    .B1(_1361_),
    .B2(_1385_),
    .A2(_0564_),
    .A1(_0537_));
 sg13g2_o21ai_1 _4836_ (.B1(_1383_),
    .Y(_1387_),
    .A1(_1350_),
    .A2(_1351_));
 sg13g2_nand3_1 _4837_ (.B(_2935_),
    .C(_0469_),
    .A(net1001),
    .Y(_1388_));
 sg13g2_nor2_2 _4838_ (.A(_2844_),
    .B(_1388_),
    .Y(_1389_));
 sg13g2_nor4_1 _4839_ (.A(_0851_),
    .B(_0862_),
    .C(_1371_),
    .D(_1387_),
    .Y(_1390_));
 sg13g2_nor2b_1 _4840_ (.A(_0896_),
    .B_N(_0899_),
    .Y(_1391_));
 sg13g2_or3_1 _4841_ (.A(_0828_),
    .B(_0830_),
    .C(_0843_),
    .X(_1392_));
 sg13g2_and2_1 _4842_ (.A(_0805_),
    .B(_0820_),
    .X(_1393_));
 sg13g2_o21ai_1 _4843_ (.B1(_1371_),
    .Y(_1394_),
    .A1(_1387_),
    .A2(_1393_));
 sg13g2_a21o_1 _4844_ (.A2(_1392_),
    .A1(_1387_),
    .B1(_1394_),
    .X(_1395_));
 sg13g2_nand2_1 _4845_ (.Y(_1396_),
    .A(_1386_),
    .B(_1395_));
 sg13g2_nand3b_1 _4846_ (.B(_0883_),
    .C(_1387_),
    .Y(_1397_),
    .A_N(_0869_));
 sg13g2_nor2_1 _4847_ (.A(_1386_),
    .B(_1390_),
    .Y(_1398_));
 sg13g2_o21ai_1 _4848_ (.B1(_1371_),
    .Y(_1399_),
    .A1(_1387_),
    .A2(_1391_));
 sg13g2_nand3_1 _4849_ (.B(_1398_),
    .C(_1399_),
    .A(_1397_),
    .Y(_1400_));
 sg13g2_nand3_1 _4850_ (.B(_1396_),
    .C(_1400_),
    .A(_1389_),
    .Y(_1401_));
 sg13g2_o21ai_1 _4851_ (.B1(_1401_),
    .Y(_0137_),
    .A1(_2699_),
    .A2(_1389_));
 sg13g2_nand3_1 _4852_ (.B(net1181),
    .C(_0063_),
    .A(net1179),
    .Y(_1402_));
 sg13g2_o21ai_1 _4853_ (.B1(_2682_),
    .Y(_1403_),
    .A1(net1200),
    .A2(_1402_));
 sg13g2_nor3_1 _4854_ (.A(net1203),
    .B(_2962_),
    .C(net1157),
    .Y(_1404_));
 sg13g2_o21ai_1 _4855_ (.B1(_2656_),
    .Y(_1405_),
    .A1(net1200),
    .A2(\dtop.vtop.rs.x_scan.phase[0] ));
 sg13g2_nand3_1 _4856_ (.B(_1404_),
    .C(_1405_),
    .A(_1403_),
    .Y(_1406_));
 sg13g2_o21ai_1 _4857_ (.B1(\dtop.vtop.rs.x_scan.phase[0] ),
    .Y(_1407_),
    .A1(net1200),
    .A2(_2682_));
 sg13g2_nor2_1 _4858_ (.A(net1179),
    .B(net1181),
    .Y(_1408_));
 sg13g2_nand2b_1 _4859_ (.Y(_1409_),
    .B(_1408_),
    .A_N(_0063_));
 sg13g2_a221oi_1 _4860_ (.B2(\dtop.vtop.rs.x_scan.phase[1] ),
    .C1(_1406_),
    .B1(_1409_),
    .A1(net1205),
    .Y(_1410_),
    .A2(_1407_));
 sg13g2_nor2_2 _4861_ (.A(_2682_),
    .B(net653),
    .Y(_1411_));
 sg13g2_and2_1 _4862_ (.A(net1214),
    .B(_0056_),
    .X(_1412_));
 sg13g2_nand3_1 _4863_ (.B(_1411_),
    .C(_1412_),
    .A(_1410_),
    .Y(_1413_));
 sg13g2_nand2_1 _4864_ (.Y(_1414_),
    .A(net1250),
    .B(_1413_));
 sg13g2_nor2_1 _4865_ (.A(net390),
    .B(_1414_),
    .Y(_1415_));
 sg13g2_o21ai_1 _4866_ (.B1(_1414_),
    .Y(_1416_),
    .A1(_2683_),
    .A2(\dtop.vtop.rs.scan_y.phase[0] ));
 sg13g2_nor2b_1 _4867_ (.A(_1415_),
    .B_N(_1416_),
    .Y(_0139_));
 sg13g2_nor3_1 _4868_ (.A(net1226),
    .B(_0085_),
    .C(_0084_),
    .Y(_1417_));
 sg13g2_nand2_1 _4869_ (.Y(_1418_),
    .A(\dtop.vtop.rs.scan_y.phase[1] ),
    .B(\dtop.vtop.rs.scan_y.phase[0] ));
 sg13g2_nor2_1 _4870_ (.A(_0054_),
    .B(_0052_),
    .Y(_1419_));
 sg13g2_nand3_1 _4871_ (.B(_1418_),
    .C(_1419_),
    .A(_1417_),
    .Y(_1420_));
 sg13g2_and2_1 _4872_ (.A(\dtop.oct_counter[5] ),
    .B(_0052_),
    .X(_1421_));
 sg13g2_nand4_1 _4873_ (.B(_0085_),
    .C(_0084_),
    .A(net1226),
    .Y(_1422_),
    .D(_1421_));
 sg13g2_o21ai_1 _4874_ (.B1(_1420_),
    .Y(_1423_),
    .A1(_1418_),
    .A2(_1422_));
 sg13g2_xnor2_1 _4875_ (.Y(_1424_),
    .A(_0053_),
    .B(\dtop.vtop.rs.scan_y.phase[0] ));
 sg13g2_or2_2 _4876_ (.X(_1425_),
    .B(\dtop.vtop.rs.scan_y.phase[0] ),
    .A(\dtop.vtop.rs.scan_y.phase[1] ));
 sg13g2_nand2_1 _4877_ (.Y(_1426_),
    .A(net1174),
    .B(_1425_));
 sg13g2_a21oi_1 _4878_ (.A1(net1168),
    .A2(_1425_),
    .Y(_1427_),
    .B1(net1177));
 sg13g2_nand2_1 _4879_ (.Y(_1428_),
    .A(_2666_),
    .B(net1171));
 sg13g2_o21ai_1 _4880_ (.B1(_2666_),
    .Y(_1429_),
    .A1(net1174),
    .A2(_0054_));
 sg13g2_a21oi_1 _4881_ (.A1(net1177),
    .A2(_1429_),
    .Y(_1430_),
    .B1(_1427_));
 sg13g2_and4_1 _4882_ (.A(net1176),
    .B(_1424_),
    .C(_1426_),
    .D(_1430_),
    .X(_1431_));
 sg13g2_and3_1 _4883_ (.X(_1432_),
    .A(_0925_),
    .B(_1423_),
    .C(_1431_));
 sg13g2_nand2_1 _4884_ (.Y(_1433_),
    .A(\dtop.vtop.rs.scan_y.phase[0] ),
    .B(_1432_));
 sg13g2_o21ai_1 _4885_ (.B1(net1243),
    .Y(_1434_),
    .A1(\dtop.vtop.rs.scan_y.phase[0] ),
    .A2(_1432_));
 sg13g2_nor2b_1 _4886_ (.A(_1434_),
    .B_N(_1433_),
    .Y(_0140_));
 sg13g2_o21ai_1 _4887_ (.B1(net1243),
    .Y(_1435_),
    .A1(_2683_),
    .A2(_1433_));
 sg13g2_a21oi_1 _4888_ (.A1(_2683_),
    .A2(_1433_),
    .Y(_0141_),
    .B1(_1435_));
 sg13g2_nor2_1 _4889_ (.A(net1214),
    .B(_0056_),
    .Y(_1436_));
 sg13g2_mux2_1 _4890_ (.A0(_1436_),
    .A1(_1412_),
    .S(_1411_),
    .X(_1437_));
 sg13g2_a21oi_1 _4891_ (.A1(_1410_),
    .A2(_1437_),
    .Y(_1438_),
    .B1(net581));
 sg13g2_nand3_1 _4892_ (.B(_1410_),
    .C(_1436_),
    .A(\dtop.vtop.rs.x_scan.phase[0] ),
    .Y(_1439_));
 sg13g2_nand2_1 _4893_ (.Y(_1440_),
    .A(net1250),
    .B(_1439_));
 sg13g2_nor2_1 _4894_ (.A(net582),
    .B(_1440_),
    .Y(_0142_));
 sg13g2_o21ai_1 _4895_ (.B1(net1250),
    .Y(_1441_),
    .A1(net584),
    .A2(_1439_));
 sg13g2_a21o_1 _4896_ (.A2(_1439_),
    .A1(net584),
    .B1(_1441_),
    .X(_0143_));
 sg13g2_o21ai_1 _4897_ (.B1(net1250),
    .Y(_1442_),
    .A1(_2962_),
    .A2(_2854_));
 sg13g2_nand2_2 _4898_ (.Y(_1443_),
    .A(net1192),
    .B(net1224));
 sg13g2_xnor2_1 _4899_ (.Y(_1444_),
    .A(net1191),
    .B(net1225));
 sg13g2_nor2_1 _4900_ (.A(_1442_),
    .B(_1444_),
    .Y(_0144_));
 sg13g2_xnor2_1 _4901_ (.Y(_1445_),
    .A(_2669_),
    .B(_1443_));
 sg13g2_nor2_1 _4902_ (.A(_1442_),
    .B(_1445_),
    .Y(_0145_));
 sg13g2_nor2_1 _4903_ (.A(_0088_),
    .B(_1443_),
    .Y(_1446_));
 sg13g2_xnor2_1 _4904_ (.Y(_1447_),
    .A(net1214),
    .B(_1446_));
 sg13g2_nor2_1 _4905_ (.A(_1442_),
    .B(_1447_),
    .Y(_0146_));
 sg13g2_nor3_1 _4906_ (.A(_0088_),
    .B(_0001_),
    .C(_1443_),
    .Y(_1448_));
 sg13g2_xnor2_1 _4907_ (.Y(_1449_),
    .A(net1211),
    .B(_1448_));
 sg13g2_nor2_1 _4908_ (.A(_1442_),
    .B(net627),
    .Y(_0147_));
 sg13g2_nor4_2 _4909_ (.A(_2656_),
    .B(_0088_),
    .C(net1145),
    .Y(_1450_),
    .D(_1443_));
 sg13g2_a21oi_1 _4910_ (.A1(_2747_),
    .A2(_1446_),
    .Y(_1451_),
    .B1(net1206));
 sg13g2_nor3_1 _4911_ (.A(_1442_),
    .B(_1450_),
    .C(_1451_),
    .Y(_0148_));
 sg13g2_nand2_1 _4912_ (.Y(_1452_),
    .A(net1204),
    .B(_1450_));
 sg13g2_xnor2_1 _4913_ (.Y(_1453_),
    .A(net1203),
    .B(_1450_));
 sg13g2_nor2_1 _4914_ (.A(_1442_),
    .B(_1453_),
    .Y(_0149_));
 sg13g2_xnor2_1 _4915_ (.Y(_1454_),
    .A(_2654_),
    .B(_1452_));
 sg13g2_nor2_1 _4916_ (.A(_1442_),
    .B(_1454_),
    .Y(_0150_));
 sg13g2_nor2_1 _4917_ (.A(\dtop.vtop.pipeline.z[14] ),
    .B(_2675_),
    .Y(_1455_));
 sg13g2_nand2b_1 _4918_ (.Y(_1456_),
    .B(\dtop.vtop.pipeline.zg[9] ),
    .A_N(\dtop.vtop.pipeline.z[14] ));
 sg13g2_nand2b_1 _4919_ (.Y(_1457_),
    .B(\dtop.vtop.pipeline.zg[2] ),
    .A_N(\dtop.vtop.pipeline.z[7] ));
 sg13g2_nor2b_1 _4920_ (.A(\dtop.vtop.pipeline.z[6] ),
    .B_N(\dtop.vtop.pipeline.zg[1] ),
    .Y(_1458_));
 sg13g2_nor2b_1 _4921_ (.A(\dtop.vtop.pipeline.z[5] ),
    .B_N(\dtop.vtop.pipeline.zg[0] ),
    .Y(_1459_));
 sg13g2_nand2b_1 _4922_ (.Y(_1460_),
    .B(\dtop.vtop.pipeline.z[6] ),
    .A_N(\dtop.vtop.pipeline.zg[1] ));
 sg13g2_o21ai_1 _4923_ (.B1(_1460_),
    .Y(_1461_),
    .A1(_1458_),
    .A2(_1459_));
 sg13g2_nor2b_1 _4924_ (.A(\dtop.vtop.pipeline.zg[2] ),
    .B_N(\dtop.vtop.pipeline.z[7] ),
    .Y(_1462_));
 sg13g2_a221oi_1 _4925_ (.B2(_1461_),
    .C1(_1462_),
    .B1(_1457_),
    .A1(\dtop.vtop.pipeline.z[8] ),
    .Y(_1463_),
    .A2(_2679_));
 sg13g2_nand2_1 _4926_ (.Y(_1464_),
    .A(_2647_),
    .B(\dtop.vtop.pipeline.zg[3] ));
 sg13g2_o21ai_1 _4927_ (.B1(_1464_),
    .Y(_1465_),
    .A1(\dtop.vtop.pipeline.z[9] ),
    .A2(_2678_));
 sg13g2_a22oi_1 _4928_ (.Y(_1466_),
    .B1(_2678_),
    .B2(\dtop.vtop.pipeline.z[9] ),
    .A2(_2677_),
    .A1(\dtop.vtop.pipeline.z[10] ));
 sg13g2_o21ai_1 _4929_ (.B1(_1466_),
    .Y(_1467_),
    .A1(_1463_),
    .A2(_1465_));
 sg13g2_a22oi_1 _4930_ (.Y(_1468_),
    .B1(\dtop.vtop.pipeline.zg[5] ),
    .B2(_2645_),
    .A2(\dtop.vtop.pipeline.zg[6] ),
    .A1(_2644_));
 sg13g2_nand2b_1 _4931_ (.Y(_1469_),
    .B(\dtop.vtop.pipeline.z[12] ),
    .A_N(\dtop.vtop.pipeline.zg[7] ));
 sg13g2_o21ai_1 _4932_ (.B1(_1469_),
    .Y(_1470_),
    .A1(_2644_),
    .A2(\dtop.vtop.pipeline.zg[6] ));
 sg13g2_a21o_1 _4933_ (.A2(_1468_),
    .A1(_1467_),
    .B1(_1470_),
    .X(_1471_));
 sg13g2_a22oi_1 _4934_ (.Y(_1472_),
    .B1(\dtop.vtop.pipeline.zg[7] ),
    .B2(_2643_),
    .A2(\dtop.vtop.pipeline.zg[8] ),
    .A1(_2642_));
 sg13g2_a22oi_1 _4935_ (.Y(_1473_),
    .B1(_2676_),
    .B2(\dtop.vtop.pipeline.z[13] ),
    .A2(_2675_),
    .A1(\dtop.vtop.pipeline.z[14] ));
 sg13g2_inv_1 _4936_ (.Y(_1474_),
    .A(_1473_));
 sg13g2_a21oi_1 _4937_ (.A1(_1471_),
    .A2(_1472_),
    .Y(_1475_),
    .B1(_1474_));
 sg13g2_a21o_1 _4938_ (.A2(_1472_),
    .A1(_1471_),
    .B1(_1474_),
    .X(_1476_));
 sg13g2_nand2_1 _4939_ (.Y(_1477_),
    .A(_1456_),
    .B(_1476_));
 sg13g2_inv_2 _4940_ (.Y(_1478_),
    .A(net1042));
 sg13g2_nand3_1 _4941_ (.B(_0983_),
    .C(_1478_),
    .A(net639),
    .Y(_1479_));
 sg13g2_nor3_1 _4942_ (.A(\dtop.detune_counter[12] ),
    .B(_2660_),
    .C(_2876_),
    .Y(_1480_));
 sg13g2_a221oi_1 _4943_ (.B2(_2660_),
    .C1(_1480_),
    .B1(_0999_),
    .A1(_2681_),
    .Y(_1481_),
    .A2(_2847_));
 sg13g2_nor2_1 _4944_ (.A(\dtop.vtop.pipeline.wave_index[0] ),
    .B(_1481_),
    .Y(_1482_));
 sg13g2_nand2b_1 _4945_ (.Y(_1483_),
    .B(\dtop.vtop.pipeline.wave_index[1] ),
    .A_N(_1481_));
 sg13g2_and2_1 _4946_ (.A(_0978_),
    .B(_1483_),
    .X(_1484_));
 sg13g2_nor2_1 _4947_ (.A(_1482_),
    .B(_1484_),
    .Y(_1485_));
 sg13g2_inv_1 _4948_ (.Y(_1486_),
    .A(net1059));
 sg13g2_nand2_1 _4949_ (.Y(_1487_),
    .A(_1479_),
    .B(net1059));
 sg13g2_nand3_1 _4950_ (.B(_1479_),
    .C(net1059),
    .A(net1129),
    .Y(_1488_));
 sg13g2_mux2_1 _4951_ (.A0(net1189),
    .A1(net1197),
    .S(_1488_),
    .X(_0151_));
 sg13g2_mux2_1 _4952_ (.A0(net1186),
    .A1(net1195),
    .S(_1488_),
    .X(_0152_));
 sg13g2_nor2_1 _4953_ (.A(_0062_),
    .B(_1478_),
    .Y(_1489_));
 sg13g2_o21ai_1 _4954_ (.B1(net1044),
    .Y(_1490_),
    .A1(\dtop.vtop.pipeline.nstep_zg[0] ),
    .A2(net1193));
 sg13g2_mux2_1 _4955_ (.A0(_0060_),
    .A1(_0059_),
    .S(net1044),
    .X(_1491_));
 sg13g2_nand2_1 _4956_ (.Y(_1492_),
    .A(_1490_),
    .B(_1491_));
 sg13g2_xor2_1 _4957_ (.B(_1491_),
    .A(_1490_),
    .X(_1493_));
 sg13g2_o21ai_1 _4958_ (.B1(net1128),
    .Y(_1494_),
    .A1(net558),
    .A2(net996));
 sg13g2_a21oi_1 _4959_ (.A1(net996),
    .A2(_1493_),
    .Y(_0153_),
    .B1(_1494_));
 sg13g2_nand3_1 _4960_ (.B(_2680_),
    .C(net1044),
    .A(net1196),
    .Y(_1495_));
 sg13g2_mux2_1 _4961_ (.A0(_0039_),
    .A1(_0082_),
    .S(net1044),
    .X(_1496_));
 sg13g2_xnor2_1 _4962_ (.Y(_1497_),
    .A(_1495_),
    .B(_1496_));
 sg13g2_xor2_1 _4963_ (.B(_1497_),
    .A(_1492_),
    .X(_1498_));
 sg13g2_inv_1 _4964_ (.Y(_1499_),
    .A(_1498_));
 sg13g2_o21ai_1 _4965_ (.B1(net1128),
    .Y(_1500_),
    .A1(net560),
    .A2(net996));
 sg13g2_a21oi_1 _4966_ (.A1(net996),
    .A2(_1499_),
    .Y(_0154_),
    .B1(_1500_));
 sg13g2_nand2_1 _4967_ (.Y(_1501_),
    .A(_1496_),
    .B(_1498_));
 sg13g2_nor3_1 _4968_ (.A(net1196),
    .B(_2680_),
    .C(_1478_),
    .Y(_1502_));
 sg13g2_mux2_1 _4969_ (.A0(_0069_),
    .A1(_0081_),
    .S(net1044),
    .X(_1503_));
 sg13g2_xor2_1 _4970_ (.B(_1503_),
    .A(_1502_),
    .X(_1504_));
 sg13g2_xnor2_1 _4971_ (.Y(_1505_),
    .A(_1501_),
    .B(_1504_));
 sg13g2_inv_1 _4972_ (.Y(_1506_),
    .A(_1505_));
 sg13g2_o21ai_1 _4973_ (.B1(net1128),
    .Y(_1507_),
    .A1(net549),
    .A2(net996));
 sg13g2_a21oi_1 _4974_ (.A1(net996),
    .A2(_1505_),
    .Y(_0155_),
    .B1(_1507_));
 sg13g2_o21ai_1 _4975_ (.B1(_1506_),
    .Y(_1508_),
    .A1(_1502_),
    .A2(_1503_));
 sg13g2_nand2b_1 _4976_ (.Y(_1509_),
    .B(net1044),
    .A_N(_0040_));
 sg13g2_o21ai_1 _4977_ (.B1(_1509_),
    .Y(_1510_),
    .A1(_0068_),
    .A2(net1045));
 sg13g2_nand3_1 _4978_ (.B(net1193),
    .C(net1045),
    .A(net1196),
    .Y(_1511_));
 sg13g2_xor2_1 _4979_ (.B(_1511_),
    .A(_1510_),
    .X(_1512_));
 sg13g2_xnor2_1 _4980_ (.Y(_1513_),
    .A(_1508_),
    .B(_1512_));
 sg13g2_o21ai_1 _4981_ (.B1(net1128),
    .Y(_1514_),
    .A1(net585),
    .A2(net996));
 sg13g2_a21oi_1 _4982_ (.A1(net996),
    .A2(_1513_),
    .Y(_0156_),
    .B1(_1514_));
 sg13g2_mux2_1 _4983_ (.A0(\dtop.vtop.pipeline.dz[4] ),
    .A1(\dtop.vtop.pipeline.neg_t[4] ),
    .S(net1045),
    .X(_1515_));
 sg13g2_nor3_2 _4984_ (.A(_1510_),
    .B(_1513_),
    .C(_1515_),
    .Y(_1516_));
 sg13g2_o21ai_1 _4985_ (.B1(_1515_),
    .Y(_1517_),
    .A1(_1510_),
    .A2(_1513_));
 sg13g2_nand2b_1 _4986_ (.Y(_1518_),
    .B(_1517_),
    .A_N(_1516_));
 sg13g2_inv_1 _4987_ (.Y(_1519_),
    .A(_1518_));
 sg13g2_o21ai_1 _4988_ (.B1(net1128),
    .Y(_1520_),
    .A1(net518),
    .A2(net997));
 sg13g2_a21oi_1 _4989_ (.A1(net997),
    .A2(_1519_),
    .Y(_0157_),
    .B1(net519));
 sg13g2_mux2_1 _4990_ (.A0(\dtop.vtop.pipeline.dz[5] ),
    .A1(\dtop.vtop.pipeline.neg_t[5] ),
    .S(net1045),
    .X(_1521_));
 sg13g2_nor2b_1 _4991_ (.A(_1521_),
    .B_N(_1516_),
    .Y(_1522_));
 sg13g2_xnor2_1 _4992_ (.Y(_1523_),
    .A(_1516_),
    .B(_1521_));
 sg13g2_o21ai_1 _4993_ (.B1(net1129),
    .Y(_1524_),
    .A1(net564),
    .A2(net995));
 sg13g2_a21oi_1 _4994_ (.A1(net995),
    .A2(_1523_),
    .Y(_0158_),
    .B1(_1524_));
 sg13g2_mux2_1 _4995_ (.A0(_0066_),
    .A1(_0074_),
    .S(net1045),
    .X(_1525_));
 sg13g2_nand2_1 _4996_ (.Y(_1526_),
    .A(_1522_),
    .B(_1525_));
 sg13g2_xor2_1 _4997_ (.B(_1525_),
    .A(_1522_),
    .X(_1527_));
 sg13g2_o21ai_1 _4998_ (.B1(net1129),
    .Y(_1528_),
    .A1(net512),
    .A2(net995));
 sg13g2_a21oi_1 _4999_ (.A1(net995),
    .A2(_1527_),
    .Y(_0159_),
    .B1(_1528_));
 sg13g2_mux2_1 _5000_ (.A0(\dtop.vtop.pipeline.dz[7] ),
    .A1(\dtop.vtop.pipeline.neg_t[7] ),
    .S(net1041),
    .X(_1529_));
 sg13g2_or2_1 _5001_ (.X(_1530_),
    .B(_1529_),
    .A(_1526_));
 sg13g2_xor2_1 _5002_ (.B(_1529_),
    .A(_1526_),
    .X(_1531_));
 sg13g2_o21ai_1 _5003_ (.B1(net1129),
    .Y(_1532_),
    .A1(net588),
    .A2(net997));
 sg13g2_a21oi_1 _5004_ (.A1(net997),
    .A2(_1531_),
    .Y(_0160_),
    .B1(_1532_));
 sg13g2_mux2_1 _5005_ (.A0(_0064_),
    .A1(_0071_),
    .S(net1041),
    .X(_1533_));
 sg13g2_nor2b_1 _5006_ (.A(_1530_),
    .B_N(_1533_),
    .Y(_1534_));
 sg13g2_xor2_1 _5007_ (.B(_1533_),
    .A(_1530_),
    .X(_1535_));
 sg13g2_inv_1 _5008_ (.Y(_1536_),
    .A(_1535_));
 sg13g2_o21ai_1 _5009_ (.B1(net1129),
    .Y(_1537_),
    .A1(net517),
    .A2(net995));
 sg13g2_a21oi_1 _5010_ (.A1(net995),
    .A2(_1536_),
    .Y(_0161_),
    .B1(_1537_));
 sg13g2_nor2b_1 _5011_ (.A(net995),
    .B_N(net566),
    .Y(_1538_));
 sg13g2_xnor2_1 _5012_ (.Y(_1539_),
    .A(_0041_),
    .B(_1534_));
 sg13g2_a21oi_1 _5013_ (.A1(net995),
    .A2(_1539_),
    .Y(_1540_),
    .B1(_1538_));
 sg13g2_nor2_1 _5014_ (.A(net1114),
    .B(net567),
    .Y(_0162_));
 sg13g2_nand2_1 _5015_ (.Y(_1541_),
    .A(net1180),
    .B(net1178));
 sg13g2_nand2b_1 _5016_ (.Y(_1542_),
    .B(net1180),
    .A_N(net1182));
 sg13g2_a22oi_1 _5017_ (.Y(_1543_),
    .B1(_1542_),
    .B2(_2653_),
    .A2(_1541_),
    .A1(net1182));
 sg13g2_xnor2_1 _5018_ (.Y(_1544_),
    .A(net1204),
    .B(_1543_));
 sg13g2_nand2_1 _5019_ (.Y(_1545_),
    .A(net1179),
    .B(net1207));
 sg13g2_xnor2_1 _5020_ (.Y(_1546_),
    .A(net1179),
    .B(net1207));
 sg13g2_xor2_1 _5021_ (.B(_0063_),
    .A(net1180),
    .X(_1547_));
 sg13g2_or3_2 _5022_ (.A(net1162),
    .B(_1543_),
    .C(_1547_),
    .X(_1548_));
 sg13g2_nand2_1 _5023_ (.Y(_1549_),
    .A(net1180),
    .B(net1211));
 sg13g2_a21o_2 _5024_ (.A2(_1549_),
    .A1(_1548_),
    .B1(_1546_),
    .X(_1550_));
 sg13g2_and2_1 _5025_ (.A(_1545_),
    .B(_1550_),
    .X(_1551_));
 sg13g2_nand2b_1 _5026_ (.Y(_1552_),
    .B(_1544_),
    .A_N(_1551_));
 sg13g2_o21ai_1 _5027_ (.B1(_1552_),
    .Y(_1553_),
    .A1(_2655_),
    .A2(_1543_));
 sg13g2_nand2_1 _5028_ (.Y(_1554_),
    .A(net1182),
    .B(net1181));
 sg13g2_nand2b_1 _5029_ (.Y(_1555_),
    .B(net1179),
    .A_N(net1182));
 sg13g2_nor2_1 _5030_ (.A(net1178),
    .B(_1542_),
    .Y(_1556_));
 sg13g2_a21oi_1 _5031_ (.A1(_1554_),
    .A2(_1555_),
    .Y(_1557_),
    .B1(_1556_));
 sg13g2_xnor2_1 _5032_ (.Y(_1558_),
    .A(_2654_),
    .B(_1557_));
 sg13g2_nand2b_1 _5033_ (.Y(_1559_),
    .B(_1553_),
    .A_N(_1558_));
 sg13g2_o21ai_1 _5034_ (.B1(_1559_),
    .Y(_1560_),
    .A1(_0050_),
    .A2(_1557_));
 sg13g2_xnor2_1 _5035_ (.Y(_1561_),
    .A(_2653_),
    .B(_1542_));
 sg13g2_nand2_1 _5036_ (.Y(_1562_),
    .A(_1560_),
    .B(_1561_));
 sg13g2_o21ai_1 _5037_ (.B1(net1180),
    .Y(_1563_),
    .A1(net1182),
    .A2(net1178));
 sg13g2_nand3_1 _5038_ (.B(_1561_),
    .C(_1563_),
    .A(_1560_),
    .Y(_1564_));
 sg13g2_nor2_1 _5039_ (.A(net1178),
    .B(_1554_),
    .Y(_1565_));
 sg13g2_nor2_1 _5040_ (.A(_1408_),
    .B(_1565_),
    .Y(_1566_));
 sg13g2_xor2_1 _5041_ (.B(_1566_),
    .A(_1564_),
    .X(_1567_));
 sg13g2_nor3_2 _5042_ (.A(\dtop.vtop.rs.x_scan.phase[1] ),
    .B(\dtop.vtop.rs.x_scan.phase[0] ),
    .C(_1567_),
    .Y(_1568_));
 sg13g2_inv_1 _5043_ (.Y(_1569_),
    .A(_1568_));
 sg13g2_xor2_1 _5044_ (.B(_1561_),
    .A(_1560_),
    .X(_1570_));
 sg13g2_xnor2_1 _5045_ (.Y(_1571_),
    .A(_1560_),
    .B(_1561_));
 sg13g2_nor2_1 _5046_ (.A(_0065_),
    .B(net988),
    .Y(_1572_));
 sg13g2_xnor2_1 _5047_ (.Y(_1573_),
    .A(_1553_),
    .B(_1558_));
 sg13g2_xor2_1 _5048_ (.B(_1558_),
    .A(_1553_),
    .X(_1574_));
 sg13g2_xnor2_1 _5049_ (.Y(_1575_),
    .A(\dtop.vtop.pipeline.dz[6] ),
    .B(_1573_));
 sg13g2_a21oi_1 _5050_ (.A1(_0065_),
    .A2(net988),
    .Y(_1576_),
    .B1(_1575_));
 sg13g2_nand2b_1 _5051_ (.Y(_1577_),
    .B(_1576_),
    .A_N(_1572_));
 sg13g2_xnor2_1 _5052_ (.Y(_1578_),
    .A(_1544_),
    .B(_1551_));
 sg13g2_xor2_1 _5053_ (.B(_1551_),
    .A(_1544_),
    .X(_1579_));
 sg13g2_xnor2_1 _5054_ (.Y(_1580_),
    .A(\dtop.vtop.pipeline.dz[5] ),
    .B(_1578_));
 sg13g2_nand3_1 _5055_ (.B(_1548_),
    .C(_1549_),
    .A(_1546_),
    .Y(_1581_));
 sg13g2_and2_1 _5056_ (.A(_1550_),
    .B(_1581_),
    .X(_1582_));
 sg13g2_nand2_2 _5057_ (.Y(_1583_),
    .A(_1550_),
    .B(_1581_));
 sg13g2_xnor2_1 _5058_ (.Y(_1584_),
    .A(\dtop.vtop.pipeline.dz[4] ),
    .B(_1582_));
 sg13g2_nor3_1 _5059_ (.A(_1577_),
    .B(_1580_),
    .C(_1584_),
    .Y(_1585_));
 sg13g2_xnor2_1 _5060_ (.Y(_1586_),
    .A(_1562_),
    .B(_1563_));
 sg13g2_inv_1 _5061_ (.Y(_1587_),
    .A(_1586_));
 sg13g2_xnor2_1 _5062_ (.Y(_1588_),
    .A(_0064_),
    .B(_1586_));
 sg13g2_o21ai_1 _5063_ (.B1(_1547_),
    .Y(_1589_),
    .A1(net1162),
    .A2(_1543_));
 sg13g2_nand2_2 _5064_ (.Y(_1590_),
    .A(_1548_),
    .B(_1589_));
 sg13g2_and2_1 _5065_ (.A(_0068_),
    .B(_1590_),
    .X(_1591_));
 sg13g2_xnor2_1 _5066_ (.Y(_1592_),
    .A(_2671_),
    .B(_1543_));
 sg13g2_xor2_1 _5067_ (.B(_1592_),
    .A(\dtop.vtop.pipeline.dz[2] ),
    .X(_1593_));
 sg13g2_nor2_1 _5068_ (.A(_0068_),
    .B(_1590_),
    .Y(_1594_));
 sg13g2_nor3_1 _5069_ (.A(_1591_),
    .B(_1593_),
    .C(_1594_),
    .Y(_1595_));
 sg13g2_nor2_1 _5070_ (.A(\dtop.vtop.pipeline.dz[1] ),
    .B(net1219),
    .Y(_1596_));
 sg13g2_a22oi_1 _5071_ (.Y(_1597_),
    .B1(net1219),
    .B2(\dtop.vtop.pipeline.dz[1] ),
    .A2(net1225),
    .A1(\dtop.vtop.pipeline.dz[0] ));
 sg13g2_nor2b_1 _5072_ (.A(_1596_),
    .B_N(_1597_),
    .Y(_1598_));
 sg13g2_or2_1 _5073_ (.X(_1599_),
    .B(net1225),
    .A(\dtop.vtop.pipeline.dz[0] ));
 sg13g2_nand4_1 _5074_ (.B(_1595_),
    .C(_1598_),
    .A(_1588_),
    .Y(_1600_),
    .D(_1599_));
 sg13g2_nor4_2 _5075_ (.A(_1577_),
    .B(_1580_),
    .C(_1584_),
    .Y(_1601_),
    .D(_1600_));
 sg13g2_o21ai_1 _5076_ (.B1(_1595_),
    .Y(_1602_),
    .A1(_1596_),
    .A2(_1598_));
 sg13g2_a22oi_1 _5077_ (.Y(_1603_),
    .B1(_1592_),
    .B2(_0069_),
    .A2(_1590_),
    .A1(_0068_));
 sg13g2_o21ai_1 _5078_ (.B1(_1602_),
    .Y(_1604_),
    .A1(_1594_),
    .A2(_1603_));
 sg13g2_a22oi_1 _5079_ (.Y(_1605_),
    .B1(_1574_),
    .B2(_0066_),
    .A2(net988),
    .A1(_0065_));
 sg13g2_nor3_1 _5080_ (.A(\dtop.vtop.pipeline.dz[4] ),
    .B(_1580_),
    .C(net1069),
    .Y(_1606_));
 sg13g2_a21oi_1 _5081_ (.A1(_0067_),
    .A2(_1579_),
    .Y(_1607_),
    .B1(_1606_));
 sg13g2_nor2_1 _5082_ (.A(_1577_),
    .B(_1607_),
    .Y(_1608_));
 sg13g2_a21oi_1 _5083_ (.A1(_1585_),
    .A2(_1604_),
    .Y(_1609_),
    .B1(_1608_));
 sg13g2_o21ai_1 _5084_ (.B1(_1609_),
    .Y(_1610_),
    .A1(_1572_),
    .A2(_1605_));
 sg13g2_a22oi_1 _5085_ (.Y(_1611_),
    .B1(_1588_),
    .B2(_1610_),
    .A2(_1587_),
    .A1(_2651_));
 sg13g2_o21ai_1 _5086_ (.B1(_1568_),
    .Y(_1612_),
    .A1(_1601_),
    .A2(_1611_));
 sg13g2_or4_2 _5087_ (.A(_2641_),
    .B(_0062_),
    .C(net1042),
    .D(_1612_),
    .X(_1613_));
 sg13g2_a21oi_1 _5088_ (.A1(net554),
    .A2(net957),
    .Y(_1614_),
    .B1(net1113));
 sg13g2_o21ai_1 _5089_ (.B1(_1614_),
    .Y(_0163_),
    .A1(_1493_),
    .A2(_1613_));
 sg13g2_a21oi_1 _5090_ (.A1(net542),
    .A2(_1613_),
    .Y(_1615_),
    .B1(net1113));
 sg13g2_o21ai_1 _5091_ (.B1(_1615_),
    .Y(_0164_),
    .A1(_1499_),
    .A2(net957));
 sg13g2_a21oi_1 _5092_ (.A1(net522),
    .A2(net957),
    .Y(_1616_),
    .B1(net1113));
 sg13g2_o21ai_1 _5093_ (.B1(_1616_),
    .Y(_0165_),
    .A1(_1505_),
    .A2(net957));
 sg13g2_a21oi_1 _5094_ (.A1(net454),
    .A2(net957),
    .Y(_1617_),
    .B1(net1113));
 sg13g2_o21ai_1 _5095_ (.B1(_1617_),
    .Y(_0166_),
    .A1(_1513_),
    .A2(net957));
 sg13g2_a21oi_1 _5096_ (.A1(net578),
    .A2(net957),
    .Y(_1618_),
    .B1(net1113));
 sg13g2_o21ai_1 _5097_ (.B1(_1618_),
    .Y(_0167_),
    .A1(_1519_),
    .A2(net957));
 sg13g2_a21oi_1 _5098_ (.A1(net543),
    .A2(net958),
    .Y(_1619_),
    .B1(net1114));
 sg13g2_o21ai_1 _5099_ (.B1(_1619_),
    .Y(_0168_),
    .A1(_1523_),
    .A2(net958));
 sg13g2_a21oi_1 _5100_ (.A1(net544),
    .A2(net958),
    .Y(_1620_),
    .B1(net1115));
 sg13g2_o21ai_1 _5101_ (.B1(_1620_),
    .Y(_0169_),
    .A1(_1527_),
    .A2(net958));
 sg13g2_a21oi_1 _5102_ (.A1(net536),
    .A2(net958),
    .Y(_1621_),
    .B1(net1113));
 sg13g2_o21ai_1 _5103_ (.B1(_1621_),
    .Y(_0170_),
    .A1(_1531_),
    .A2(net958));
 sg13g2_a21oi_1 _5104_ (.A1(net556),
    .A2(net958),
    .Y(_1622_),
    .B1(net1113));
 sg13g2_o21ai_1 _5105_ (.B1(_1622_),
    .Y(_0171_),
    .A1(_1536_),
    .A2(net958));
 sg13g2_a21oi_1 _5106_ (.A1(_1478_),
    .A2(_1612_),
    .Y(_1623_),
    .B1(_2641_));
 sg13g2_a21o_2 _5107_ (.A2(_1612_),
    .A1(_1478_),
    .B1(_2641_),
    .X(_1624_));
 sg13g2_nor2b_1 _5108_ (.A(net1196),
    .B_N(\dtop.vtop.pipeline.dz[0] ),
    .Y(_1625_));
 sg13g2_nand2_1 _5109_ (.Y(_1626_),
    .A(_2680_),
    .B(_1625_));
 sg13g2_nand3_1 _5110_ (.B(_1456_),
    .C(_1476_),
    .A(_0059_),
    .Y(_1627_));
 sg13g2_o21ai_1 _5111_ (.B1(_1626_),
    .Y(_1628_),
    .A1(_1455_),
    .A2(_1475_));
 sg13g2_and2_1 _5112_ (.A(_1627_),
    .B(_1628_),
    .X(_1629_));
 sg13g2_a21oi_1 _5113_ (.A1(net956),
    .A2(_1629_),
    .Y(_1630_),
    .B1(net387));
 sg13g2_nand3_1 _5114_ (.B(_1627_),
    .C(_1628_),
    .A(net387),
    .Y(_1631_));
 sg13g2_o21ai_1 _5115_ (.B1(net1127),
    .Y(_1632_),
    .A1(_1624_),
    .A2(_1631_));
 sg13g2_nor2_1 _5116_ (.A(_1630_),
    .B(_1632_),
    .Y(_0172_));
 sg13g2_mux2_1 _5117_ (.A0(_0039_),
    .A1(_0060_),
    .S(net1196),
    .X(_1633_));
 sg13g2_nand2b_1 _5118_ (.Y(_1634_),
    .B(_2680_),
    .A_N(_1633_));
 sg13g2_nor3_2 _5119_ (.A(_0082_),
    .B(_1455_),
    .C(_1475_),
    .Y(_1635_));
 sg13g2_a21oi_1 _5120_ (.A1(_1456_),
    .A2(_1476_),
    .Y(_1636_),
    .B1(_1634_));
 sg13g2_nor2_1 _5121_ (.A(_1635_),
    .B(_1636_),
    .Y(_1637_));
 sg13g2_o21ai_1 _5122_ (.B1(\dtop.vtop.pipeline.z[1] ),
    .Y(_1638_),
    .A1(_1635_),
    .A2(_1636_));
 sg13g2_nor3_1 _5123_ (.A(\dtop.vtop.pipeline.z[1] ),
    .B(_1635_),
    .C(_1636_),
    .Y(_1639_));
 sg13g2_xor2_1 _5124_ (.B(_1637_),
    .A(net568),
    .X(_1640_));
 sg13g2_xnor2_1 _5125_ (.Y(_1641_),
    .A(_1631_),
    .B(_1640_));
 sg13g2_o21ai_1 _5126_ (.B1(net1127),
    .Y(_1642_),
    .A1(net568),
    .A2(net956));
 sg13g2_a21oi_1 _5127_ (.A1(net956),
    .A2(_1641_),
    .Y(_0173_),
    .B1(_1642_));
 sg13g2_mux2_1 _5128_ (.A0(_0069_),
    .A1(_0039_),
    .S(\dtop.vtop.pipeline.nstep_zg[0] ),
    .X(_1643_));
 sg13g2_nor2_1 _5129_ (.A(net1194),
    .B(_1643_),
    .Y(_1644_));
 sg13g2_a21oi_1 _5130_ (.A1(net1193),
    .A2(_1625_),
    .Y(_1645_),
    .B1(_1644_));
 sg13g2_mux2_1 _5131_ (.A0(_0081_),
    .A1(_1645_),
    .S(net1043),
    .X(_1646_));
 sg13g2_nor2_1 _5132_ (.A(_2650_),
    .B(_1646_),
    .Y(_1647_));
 sg13g2_xnor2_1 _5133_ (.Y(_1648_),
    .A(\dtop.vtop.pipeline.z[2] ),
    .B(_1646_));
 sg13g2_o21ai_1 _5134_ (.B1(_1638_),
    .Y(_1649_),
    .A1(_1631_),
    .A2(_1639_));
 sg13g2_xor2_1 _5135_ (.B(_1649_),
    .A(_1648_),
    .X(_1650_));
 sg13g2_o21ai_1 _5136_ (.B1(net1126),
    .Y(_1651_),
    .A1(_1624_),
    .A2(_1650_));
 sg13g2_a21oi_1 _5137_ (.A1(_2650_),
    .A2(_1624_),
    .Y(_0174_),
    .B1(_1651_));
 sg13g2_a21oi_1 _5138_ (.A1(_1648_),
    .A2(_1649_),
    .Y(_1652_),
    .B1(_1647_));
 sg13g2_nand2_1 _5139_ (.Y(_1653_),
    .A(net1193),
    .B(_1633_));
 sg13g2_nor2b_1 _5140_ (.A(net1196),
    .B_N(_0068_),
    .Y(_1654_));
 sg13g2_a21oi_1 _5141_ (.A1(\dtop.vtop.pipeline.nstep_zg[0] ),
    .A2(_0069_),
    .Y(_1655_),
    .B1(_1654_));
 sg13g2_o21ai_1 _5142_ (.B1(_1653_),
    .Y(_1656_),
    .A1(net1194),
    .A2(_1655_));
 sg13g2_mux2_1 _5143_ (.A0(_0040_),
    .A1(_1656_),
    .S(net1043),
    .X(_1657_));
 sg13g2_inv_1 _5144_ (.Y(_1658_),
    .A(_1657_));
 sg13g2_nand2_1 _5145_ (.Y(_1659_),
    .A(\dtop.vtop.pipeline.z[3] ),
    .B(_1658_));
 sg13g2_xor2_1 _5146_ (.B(_1657_),
    .A(net561),
    .X(_1660_));
 sg13g2_xnor2_1 _5147_ (.Y(_1661_),
    .A(_1652_),
    .B(_1660_));
 sg13g2_o21ai_1 _5148_ (.B1(net1126),
    .Y(_1662_),
    .A1(net561),
    .A2(net956));
 sg13g2_a21oi_1 _5149_ (.A1(net956),
    .A2(_1661_),
    .Y(_0175_),
    .B1(_1662_));
 sg13g2_o21ai_1 _5150_ (.B1(_1659_),
    .Y(_1663_),
    .A1(_1652_),
    .A2(_1660_));
 sg13g2_mux2_1 _5151_ (.A0(_0042_),
    .A1(_0068_),
    .S(net1196),
    .X(_1664_));
 sg13g2_mux2_1 _5152_ (.A0(_1643_),
    .A1(_1664_),
    .S(_2680_),
    .X(_1665_));
 sg13g2_mux2_1 _5153_ (.A0(_0077_),
    .A1(_1665_),
    .S(net1043),
    .X(_1666_));
 sg13g2_nor2_1 _5154_ (.A(_2649_),
    .B(_1666_),
    .Y(_1667_));
 sg13g2_xnor2_1 _5155_ (.Y(_1668_),
    .A(_2649_),
    .B(_1666_));
 sg13g2_inv_1 _5156_ (.Y(_1669_),
    .A(_1668_));
 sg13g2_xnor2_1 _5157_ (.Y(_1670_),
    .A(_1663_),
    .B(_1668_));
 sg13g2_o21ai_1 _5158_ (.B1(net1126),
    .Y(_1671_),
    .A1(_1624_),
    .A2(_1670_));
 sg13g2_a21oi_1 _5159_ (.A1(_2649_),
    .A2(_1624_),
    .Y(_0176_),
    .B1(_1671_));
 sg13g2_a21oi_1 _5160_ (.A1(_1663_),
    .A2(_1669_),
    .Y(_1672_),
    .B1(_1667_));
 sg13g2_mux2_1 _5161_ (.A0(_0067_),
    .A1(_0042_),
    .S(net1196),
    .X(_1673_));
 sg13g2_nand2_1 _5162_ (.Y(_1674_),
    .A(net1194),
    .B(_1655_));
 sg13g2_o21ai_1 _5163_ (.B1(_1674_),
    .Y(_1675_),
    .A1(net1193),
    .A2(_1673_));
 sg13g2_nor2_1 _5164_ (.A(_0076_),
    .B(net1041),
    .Y(_1676_));
 sg13g2_a21oi_1 _5165_ (.A1(net1042),
    .A2(_1675_),
    .Y(_1677_),
    .B1(_1676_));
 sg13g2_inv_1 _5166_ (.Y(_1678_),
    .A(_1677_));
 sg13g2_nor2_1 _5167_ (.A(\dtop.vtop.pipeline.z[5] ),
    .B(_1678_),
    .Y(_1679_));
 sg13g2_xor2_1 _5168_ (.B(_1677_),
    .A(net592),
    .X(_1680_));
 sg13g2_xnor2_1 _5169_ (.Y(_1681_),
    .A(_1672_),
    .B(_1680_));
 sg13g2_o21ai_1 _5170_ (.B1(net1126),
    .Y(_1682_),
    .A1(net592),
    .A2(net956));
 sg13g2_a21oi_1 _5171_ (.A1(_1623_),
    .A2(_1681_),
    .Y(_0177_),
    .B1(_1682_));
 sg13g2_mux2_1 _5172_ (.A0(_0066_),
    .A1(_0067_),
    .S(net1197),
    .X(_1683_));
 sg13g2_mux2_1 _5173_ (.A0(_1664_),
    .A1(_1683_),
    .S(_2680_),
    .X(_1684_));
 sg13g2_mux2_1 _5174_ (.A0(_0074_),
    .A1(_1684_),
    .S(net1042),
    .X(_1685_));
 sg13g2_nor2_1 _5175_ (.A(_2648_),
    .B(_1685_),
    .Y(_1686_));
 sg13g2_xnor2_1 _5176_ (.Y(_1687_),
    .A(_2648_),
    .B(_1685_));
 sg13g2_a221oi_1 _5177_ (.B2(\dtop.vtop.pipeline.z[5] ),
    .C1(_1667_),
    .B1(_1678_),
    .A1(_1663_),
    .Y(_1688_),
    .A2(_1669_));
 sg13g2_nor3_2 _5178_ (.A(_1679_),
    .B(_1687_),
    .C(_1688_),
    .Y(_1689_));
 sg13g2_o21ai_1 _5179_ (.B1(_1687_),
    .Y(_1690_),
    .A1(_1679_),
    .A2(_1688_));
 sg13g2_nor2b_1 _5180_ (.A(_1689_),
    .B_N(_1690_),
    .Y(_1691_));
 sg13g2_o21ai_1 _5181_ (.B1(net1126),
    .Y(_1692_),
    .A1(_1624_),
    .A2(_1691_));
 sg13g2_a21oi_1 _5182_ (.A1(_2648_),
    .A2(_1624_),
    .Y(_0178_),
    .B1(_1692_));
 sg13g2_nor2_1 _5183_ (.A(_1686_),
    .B(_1689_),
    .Y(_1693_));
 sg13g2_and2_1 _5184_ (.A(net1193),
    .B(_1673_),
    .X(_1694_));
 sg13g2_mux2_1 _5185_ (.A0(_0065_),
    .A1(_0066_),
    .S(net1197),
    .X(_1695_));
 sg13g2_a21oi_1 _5186_ (.A1(_2680_),
    .A2(_1695_),
    .Y(_1696_),
    .B1(_1694_));
 sg13g2_nor2_1 _5187_ (.A(_0043_),
    .B(net1041),
    .Y(_1697_));
 sg13g2_a21oi_1 _5188_ (.A1(net1042),
    .A2(_1696_),
    .Y(_1698_),
    .B1(_1697_));
 sg13g2_inv_1 _5189_ (.Y(_1699_),
    .A(_1698_));
 sg13g2_nand2_1 _5190_ (.Y(_1700_),
    .A(\dtop.vtop.pipeline.z[7] ),
    .B(_1699_));
 sg13g2_xor2_1 _5191_ (.B(_1698_),
    .A(\dtop.vtop.pipeline.z[7] ),
    .X(_1701_));
 sg13g2_inv_1 _5192_ (.Y(_1702_),
    .A(_1701_));
 sg13g2_o21ai_1 _5193_ (.B1(_1702_),
    .Y(_1703_),
    .A1(_1686_),
    .A2(_1689_));
 sg13g2_xnor2_1 _5194_ (.Y(_1704_),
    .A(_1693_),
    .B(_1701_));
 sg13g2_o21ai_1 _5195_ (.B1(net1127),
    .Y(_1705_),
    .A1(net597),
    .A2(net954));
 sg13g2_a21oi_1 _5196_ (.A1(net954),
    .A2(_1704_),
    .Y(_0179_),
    .B1(_1705_));
 sg13g2_nor2b_1 _5197_ (.A(net1197),
    .B_N(_0064_),
    .Y(_1706_));
 sg13g2_a21oi_1 _5198_ (.A1(net1197),
    .A2(_0065_),
    .Y(_1707_),
    .B1(_1706_));
 sg13g2_nor2_1 _5199_ (.A(net1195),
    .B(_1707_),
    .Y(_1708_));
 sg13g2_a21oi_1 _5200_ (.A1(net1193),
    .A2(_1683_),
    .Y(_1709_),
    .B1(_1708_));
 sg13g2_nor2_1 _5201_ (.A(_0071_),
    .B(net1041),
    .Y(_1710_));
 sg13g2_a21oi_1 _5202_ (.A1(net1041),
    .A2(_1709_),
    .Y(_1711_),
    .B1(_1710_));
 sg13g2_xnor2_1 _5203_ (.Y(_1712_),
    .A(_2647_),
    .B(_1711_));
 sg13g2_a21o_1 _5204_ (.A2(_1703_),
    .A1(_1700_),
    .B1(_1712_),
    .X(_1713_));
 sg13g2_nand3_1 _5205_ (.B(_1703_),
    .C(_1712_),
    .A(_1700_),
    .Y(_1714_));
 sg13g2_nand2_1 _5206_ (.Y(_1715_),
    .A(_1713_),
    .B(_1714_));
 sg13g2_o21ai_1 _5207_ (.B1(net1127),
    .Y(_1716_),
    .A1(net547),
    .A2(net954));
 sg13g2_a21oi_1 _5208_ (.A1(net954),
    .A2(_1715_),
    .Y(_0180_),
    .B1(_1716_));
 sg13g2_o21ai_1 _5209_ (.B1(_1713_),
    .Y(_1717_),
    .A1(_2647_),
    .A2(_1711_));
 sg13g2_a21oi_1 _5210_ (.A1(\dtop.vtop.pipeline.dz[8] ),
    .A2(net1197),
    .Y(_1718_),
    .B1(net1195));
 sg13g2_a21oi_1 _5211_ (.A1(net1195),
    .A2(_1695_),
    .Y(_1719_),
    .B1(_1718_));
 sg13g2_nor2_1 _5212_ (.A(_0041_),
    .B(net1041),
    .Y(_1720_));
 sg13g2_a21oi_1 _5213_ (.A1(net1041),
    .A2(_1719_),
    .Y(_1721_),
    .B1(_1720_));
 sg13g2_nor2_1 _5214_ (.A(_2646_),
    .B(_1721_),
    .Y(_1722_));
 sg13g2_nand2_1 _5215_ (.Y(_1723_),
    .A(_2646_),
    .B(_1721_));
 sg13g2_nor2b_1 _5216_ (.A(_1722_),
    .B_N(_1723_),
    .Y(_1724_));
 sg13g2_xnor2_1 _5217_ (.Y(_1725_),
    .A(_1717_),
    .B(_1724_));
 sg13g2_o21ai_1 _5218_ (.B1(net1127),
    .Y(_1726_),
    .A1(net572),
    .A2(net954));
 sg13g2_a21oi_1 _5219_ (.A1(net954),
    .A2(_1725_),
    .Y(_0181_),
    .B1(_1726_));
 sg13g2_a21oi_1 _5220_ (.A1(net1193),
    .A2(_1707_),
    .Y(_1727_),
    .B1(_1478_));
 sg13g2_xnor2_1 _5221_ (.Y(_1728_),
    .A(\dtop.vtop.pipeline.z[10] ),
    .B(_1727_));
 sg13g2_and2_1 _5222_ (.A(_1717_),
    .B(_1723_),
    .X(_1729_));
 sg13g2_nor2_1 _5223_ (.A(_1722_),
    .B(_1729_),
    .Y(_1730_));
 sg13g2_o21ai_1 _5224_ (.B1(_1728_),
    .Y(_1731_),
    .A1(_1722_),
    .A2(_1729_));
 sg13g2_xor2_1 _5225_ (.B(_1730_),
    .A(_1728_),
    .X(_1732_));
 sg13g2_o21ai_1 _5226_ (.B1(net1127),
    .Y(_1733_),
    .A1(net574),
    .A2(net954));
 sg13g2_a21oi_1 _5227_ (.A1(net954),
    .A2(_1732_),
    .Y(_0182_),
    .B1(_1733_));
 sg13g2_nand3_1 _5228_ (.B(net1197),
    .C(net1195),
    .A(\dtop.vtop.pipeline.dz[8] ),
    .Y(_1734_));
 sg13g2_nand3_1 _5229_ (.B(net1042),
    .C(_1734_),
    .A(_2644_),
    .Y(_1735_));
 sg13g2_a21oi_1 _5230_ (.A1(net1042),
    .A2(_1734_),
    .Y(_1736_),
    .B1(_2644_));
 sg13g2_a21o_1 _5231_ (.A2(_1734_),
    .A1(net1042),
    .B1(_2644_),
    .X(_1737_));
 sg13g2_and2_1 _5232_ (.A(_1735_),
    .B(_1737_),
    .X(_1738_));
 sg13g2_o21ai_1 _5233_ (.B1(_1731_),
    .Y(_1739_),
    .A1(_2645_),
    .A2(_1727_));
 sg13g2_xnor2_1 _5234_ (.Y(_1740_),
    .A(_1738_),
    .B(_1739_));
 sg13g2_o21ai_1 _5235_ (.B1(net1127),
    .Y(_1741_),
    .A1(net546),
    .A2(net955));
 sg13g2_a21oi_1 _5236_ (.A1(net955),
    .A2(_1740_),
    .Y(_0183_),
    .B1(_1741_));
 sg13g2_nor2_1 _5237_ (.A(\dtop.vtop.pipeline.z[12] ),
    .B(net1043),
    .Y(_1742_));
 sg13g2_nor2_1 _5238_ (.A(_2643_),
    .B(_1478_),
    .Y(_1743_));
 sg13g2_nand2_1 _5239_ (.Y(_1744_),
    .A(\dtop.vtop.pipeline.z[12] ),
    .B(net1043));
 sg13g2_nor2_1 _5240_ (.A(_1742_),
    .B(_1743_),
    .Y(_1745_));
 sg13g2_a21oi_2 _5241_ (.B1(_1736_),
    .Y(_1746_),
    .A2(_1739_),
    .A1(_1735_));
 sg13g2_xnor2_1 _5242_ (.Y(_1747_),
    .A(_1745_),
    .B(_1746_));
 sg13g2_o21ai_1 _5243_ (.B1(net1126),
    .Y(_1748_),
    .A1(net583),
    .A2(net955));
 sg13g2_a21oi_1 _5244_ (.A1(net955),
    .A2(_1747_),
    .Y(_0184_),
    .B1(_1748_));
 sg13g2_mux2_1 _5245_ (.A0(_1743_),
    .A1(_1742_),
    .S(_1746_),
    .X(_1749_));
 sg13g2_nand2_1 _5246_ (.Y(_1750_),
    .A(net955),
    .B(_1749_));
 sg13g2_o21ai_1 _5247_ (.B1(net1126),
    .Y(_1751_),
    .A1(_2642_),
    .A2(_1750_));
 sg13g2_a21oi_1 _5248_ (.A1(_2642_),
    .A2(_1750_),
    .Y(_0185_),
    .B1(_1751_));
 sg13g2_o21ai_1 _5249_ (.B1(\dtop.vtop.pipeline.z[13] ),
    .Y(_1752_),
    .A1(_1744_),
    .A2(_1746_));
 sg13g2_o21ai_1 _5250_ (.B1(_1752_),
    .Y(_1753_),
    .A1(\dtop.vtop.pipeline.z[13] ),
    .A2(_1478_));
 sg13g2_nor2_1 _5251_ (.A(_1750_),
    .B(_1753_),
    .Y(_1754_));
 sg13g2_o21ai_1 _5252_ (.B1(net1126),
    .Y(_1755_),
    .A1(net499),
    .A2(_1754_));
 sg13g2_a21oi_1 _5253_ (.A1(net499),
    .A2(_1754_),
    .Y(_0186_),
    .B1(_1755_));
 sg13g2_nand2b_1 _5254_ (.Y(_1756_),
    .B(net610),
    .A_N(\dtop.vtop.pipeline.wave_index[1] ));
 sg13g2_o21ai_1 _5255_ (.B1(_1331_),
    .Y(_1757_),
    .A1(net1114),
    .A2(_1756_));
 sg13g2_a221oi_1 _5256_ (.B2(\dtop.vtop.pipeline.phases[1][0] ),
    .C1(net1095),
    .B1(net1092),
    .A1(\dtop.vtop.pipeline.phases[2][0] ),
    .Y(_1758_),
    .A2(net1093));
 sg13g2_a21oi_1 _5257_ (.A1(_0007_),
    .A2(net1095),
    .Y(_1759_),
    .B1(_1758_));
 sg13g2_xnor2_1 _5258_ (.Y(_1760_),
    .A(net1105),
    .B(net1104));
 sg13g2_nor3_1 _5259_ (.A(\dtop.vtop.dphases[2][0] ),
    .B(net1105),
    .C(_0990_),
    .Y(_1761_));
 sg13g2_a221oi_1 _5260_ (.B2(_0009_),
    .C1(_1761_),
    .B1(net1081),
    .A1(_2690_),
    .Y(_1762_),
    .A2(net1091));
 sg13g2_and2_1 _5261_ (.A(net1161),
    .B(_1762_),
    .X(_1763_));
 sg13g2_a21oi_1 _5262_ (.A1(_0008_),
    .A2(_1763_),
    .Y(_1764_),
    .B1(_1759_));
 sg13g2_nand3_1 _5263_ (.B(_1759_),
    .C(_1763_),
    .A(_0008_),
    .Y(_1765_));
 sg13g2_nand2_1 _5264_ (.Y(_1766_),
    .A(net1122),
    .B(_1765_));
 sg13g2_nor2_1 _5265_ (.A(_1764_),
    .B(_1766_),
    .Y(_1767_));
 sg13g2_mux2_1 _5266_ (.A0(net405),
    .A1(_1767_),
    .S(net1067),
    .X(_0187_));
 sg13g2_nand2_1 _5267_ (.Y(_1768_),
    .A(\dtop.vtop.pipeline.phases[1][1] ),
    .B(net1106));
 sg13g2_nor2_1 _5268_ (.A(\dtop.vtop.pipeline.phases[2][1] ),
    .B(net1105),
    .Y(_1769_));
 sg13g2_a221oi_1 _5269_ (.B2(_0990_),
    .C1(_1769_),
    .B1(_1768_),
    .A1(_0010_),
    .Y(_1770_),
    .A2(net1096));
 sg13g2_nor3_1 _5270_ (.A(\dtop.vtop.dphases[2][1] ),
    .B(net1105),
    .C(_0990_),
    .Y(_1771_));
 sg13g2_a221oi_1 _5271_ (.B2(_0011_),
    .C1(_1771_),
    .B1(net1081),
    .A1(_2692_),
    .Y(_1772_),
    .A2(net1091));
 sg13g2_mux2_1 _5272_ (.A0(_1762_),
    .A1(_1772_),
    .S(net1161),
    .X(_1773_));
 sg13g2_nand3_1 _5273_ (.B(_1770_),
    .C(_1773_),
    .A(_0008_),
    .Y(_1774_));
 sg13g2_a21oi_1 _5274_ (.A1(_0008_),
    .A2(_1773_),
    .Y(_1775_),
    .B1(_1770_));
 sg13g2_a21o_1 _5275_ (.A2(_1773_),
    .A1(_0008_),
    .B1(_1770_),
    .X(_1776_));
 sg13g2_nand2_1 _5276_ (.Y(_1777_),
    .A(_1774_),
    .B(_1776_));
 sg13g2_xnor2_1 _5277_ (.Y(_1778_),
    .A(_1765_),
    .B(_1777_));
 sg13g2_nand2_2 _5278_ (.Y(_1779_),
    .A(net1211),
    .B(_2891_));
 sg13g2_xnor2_1 _5279_ (.Y(_1780_),
    .A(net1231),
    .B(net1220));
 sg13g2_nor2_1 _5280_ (.A(_1779_),
    .B(_1780_),
    .Y(_1781_));
 sg13g2_a21oi_1 _5281_ (.A1(_0088_),
    .A2(_1779_),
    .Y(_1782_),
    .B1(net1123));
 sg13g2_nor2b_2 _5282_ (.A(_1781_),
    .B_N(_1782_),
    .Y(_1783_));
 sg13g2_nand2b_2 _5283_ (.Y(_1784_),
    .B(_1782_),
    .A_N(_1781_));
 sg13g2_a21oi_2 _5284_ (.B1(net1112),
    .Y(_1785_),
    .A2(_1589_),
    .A1(_1548_));
 sg13g2_a21o_1 _5285_ (.A2(_1589_),
    .A1(_1548_),
    .B1(net1112),
    .X(_1786_));
 sg13g2_nor2_1 _5286_ (.A(_1783_),
    .B(_1785_),
    .Y(_1787_));
 sg13g2_xnor2_1 _5287_ (.Y(_1788_),
    .A(\dtop.detune_counter[12] ),
    .B(net1215));
 sg13g2_xnor2_1 _5288_ (.Y(_1789_),
    .A(_1780_),
    .B(_1788_));
 sg13g2_nand2_1 _5289_ (.Y(_1790_),
    .A(_0001_),
    .B(_1779_));
 sg13g2_o21ai_1 _5290_ (.B1(_1790_),
    .Y(_1791_),
    .A1(_1779_),
    .A2(_1789_));
 sg13g2_o21ai_1 _5291_ (.B1(_1791_),
    .Y(_1792_),
    .A1(_1783_),
    .A2(_1785_));
 sg13g2_and3_1 _5292_ (.X(_1793_),
    .A(_2891_),
    .B(_1780_),
    .C(_1788_));
 sg13g2_nor3_2 _5293_ (.A(net1208),
    .B(net1123),
    .C(_1793_),
    .Y(_1794_));
 sg13g2_or3_1 _5294_ (.A(net1208),
    .B(net1123),
    .C(_1793_),
    .X(_1795_));
 sg13g2_nand4_1 _5295_ (.B(_1783_),
    .C(_1791_),
    .A(net1110),
    .Y(_1796_),
    .D(net1101));
 sg13g2_o21ai_1 _5296_ (.B1(_1796_),
    .Y(_1797_),
    .A1(net1109),
    .A2(_1778_));
 sg13g2_mux2_1 _5297_ (.A0(net401),
    .A1(_1797_),
    .S(net1067),
    .X(_0188_));
 sg13g2_o21ai_1 _5298_ (.B1(_1774_),
    .Y(_1798_),
    .A1(_1765_),
    .A2(_1775_));
 sg13g2_a221oi_1 _5299_ (.B2(\dtop.vtop.pipeline.phases[1][2] ),
    .C1(net1095),
    .B1(net1092),
    .A1(\dtop.vtop.pipeline.phases[2][2] ),
    .Y(_1799_),
    .A2(net1093));
 sg13g2_a21oi_2 _5300_ (.B1(_1799_),
    .Y(_1800_),
    .A2(net1095),
    .A1(_0012_));
 sg13g2_nor3_1 _5301_ (.A(\dtop.vtop.dphases[2][2] ),
    .B(net1106),
    .C(_0990_),
    .Y(_1801_));
 sg13g2_a221oi_1 _5302_ (.B2(_0013_),
    .C1(_1801_),
    .B1(_1760_),
    .A1(_2693_),
    .Y(_1802_),
    .A2(net1091));
 sg13g2_mux2_1 _5303_ (.A0(_1772_),
    .A1(_1802_),
    .S(net1161),
    .X(_1803_));
 sg13g2_mux2_1 _5304_ (.A0(_1803_),
    .A1(_1763_),
    .S(net1184),
    .X(_1804_));
 sg13g2_and2_1 _5305_ (.A(_1800_),
    .B(_1804_),
    .X(_1805_));
 sg13g2_xor2_1 _5306_ (.B(_1804_),
    .A(_1800_),
    .X(_1806_));
 sg13g2_xnor2_1 _5307_ (.Y(_1807_),
    .A(_1798_),
    .B(_1806_));
 sg13g2_o21ai_1 _5308_ (.B1(_1796_),
    .Y(_1808_),
    .A1(net1109),
    .A2(_1807_));
 sg13g2_mux2_1 _5309_ (.A0(net416),
    .A1(_1808_),
    .S(net1067),
    .X(_0189_));
 sg13g2_a21oi_2 _5310_ (.B1(_1805_),
    .Y(_1809_),
    .A2(_1806_),
    .A1(_1798_));
 sg13g2_nand2_1 _5311_ (.Y(_1810_),
    .A(\dtop.vtop.pipeline.phases[1][3] ),
    .B(net1105));
 sg13g2_nor2_1 _5312_ (.A(\dtop.vtop.pipeline.phases[2][3] ),
    .B(net1105),
    .Y(_1811_));
 sg13g2_a221oi_1 _5313_ (.B2(_0990_),
    .C1(_1811_),
    .B1(_1810_),
    .A1(_0014_),
    .Y(_1812_),
    .A2(net1096));
 sg13g2_a22oi_1 _5314_ (.Y(_1813_),
    .B1(_1760_),
    .B2(_0015_),
    .A2(net1091),
    .A1(_2694_));
 sg13g2_o21ai_1 _5315_ (.B1(_1813_),
    .Y(_1814_),
    .A1(\dtop.vtop.dphases[2][3] ),
    .A2(_1011_));
 sg13g2_nand2_1 _5316_ (.Y(_1815_),
    .A(net1188),
    .B(_1802_));
 sg13g2_o21ai_1 _5317_ (.B1(_1815_),
    .Y(_1816_),
    .A1(net1188),
    .A2(_1814_));
 sg13g2_mux2_1 _5318_ (.A0(_1816_),
    .A1(_1773_),
    .S(net1184),
    .X(_1817_));
 sg13g2_nand2_1 _5319_ (.Y(_1818_),
    .A(_1812_),
    .B(_1817_));
 sg13g2_xnor2_1 _5320_ (.Y(_1819_),
    .A(_1812_),
    .B(_1817_));
 sg13g2_o21ai_1 _5321_ (.B1(net1122),
    .Y(_1820_),
    .A1(_1809_),
    .A2(_1819_));
 sg13g2_a21o_1 _5322_ (.A2(_1819_),
    .A1(_1809_),
    .B1(_1820_),
    .X(_1821_));
 sg13g2_o21ai_1 _5323_ (.B1(_1821_),
    .Y(_1822_),
    .A1(_1784_),
    .A2(_1794_));
 sg13g2_mux2_1 _5324_ (.A0(net428),
    .A1(_1822_),
    .S(net1067),
    .X(_0190_));
 sg13g2_a21oi_2 _5325_ (.B1(_1785_),
    .Y(_1823_),
    .A2(_1791_),
    .A1(net1110));
 sg13g2_a21o_2 _5326_ (.A2(_1791_),
    .A1(net1110),
    .B1(_1785_),
    .X(_1824_));
 sg13g2_nor2_1 _5327_ (.A(_1783_),
    .B(_1824_),
    .Y(_1825_));
 sg13g2_o21ai_1 _5328_ (.B1(net1066),
    .Y(_1826_),
    .A1(_2673_),
    .A2(_1823_));
 sg13g2_nand3_1 _5329_ (.B(net1101),
    .C(_1826_),
    .A(net1110),
    .Y(_1827_));
 sg13g2_o21ai_1 _5330_ (.B1(_1818_),
    .Y(_1828_),
    .A1(_1809_),
    .A2(_1819_));
 sg13g2_a221oi_1 _5331_ (.B2(\dtop.vtop.pipeline.phases[1][4] ),
    .C1(net1095),
    .B1(net1092),
    .A1(\dtop.vtop.pipeline.phases[2][4] ),
    .Y(_1829_),
    .A2(net1093));
 sg13g2_a21oi_2 _5332_ (.B1(_1829_),
    .Y(_1830_),
    .A2(net1095),
    .A1(_0016_));
 sg13g2_a22oi_1 _5333_ (.Y(_1831_),
    .B1(_1760_),
    .B2(_0017_),
    .A2(net1092),
    .A1(_2695_));
 sg13g2_o21ai_1 _5334_ (.B1(_1831_),
    .Y(_1832_),
    .A1(\dtop.vtop.dphases[2][4] ),
    .A2(_1011_));
 sg13g2_nand2b_1 _5335_ (.Y(_1833_),
    .B(net1161),
    .A_N(_1832_));
 sg13g2_o21ai_1 _5336_ (.B1(_1833_),
    .Y(_1834_),
    .A1(net1161),
    .A2(_1814_));
 sg13g2_mux2_1 _5337_ (.A0(_1834_),
    .A1(_1803_),
    .S(net1184),
    .X(_1835_));
 sg13g2_and2_1 _5338_ (.A(_1830_),
    .B(_1835_),
    .X(_1836_));
 sg13g2_xor2_1 _5339_ (.B(_1835_),
    .A(_1830_),
    .X(_1837_));
 sg13g2_xnor2_1 _5340_ (.Y(_1838_),
    .A(_1828_),
    .B(_1837_));
 sg13g2_o21ai_1 _5341_ (.B1(_1827_),
    .Y(_1839_),
    .A1(net1110),
    .A2(_1838_));
 sg13g2_mux2_1 _5342_ (.A0(net402),
    .A1(_1839_),
    .S(net1067),
    .X(_0191_));
 sg13g2_a21o_1 _5343_ (.A2(_1837_),
    .A1(_1828_),
    .B1(_1836_),
    .X(_1840_));
 sg13g2_a22oi_1 _5344_ (.Y(_1841_),
    .B1(net1092),
    .B2(\dtop.vtop.pipeline.phases[1][5] ),
    .A2(net1093),
    .A1(\dtop.vtop.pipeline.phases[2][5] ));
 sg13g2_o21ai_1 _5345_ (.B1(_1841_),
    .Y(_1842_),
    .A1(_0018_),
    .A2(_0993_));
 sg13g2_a22oi_1 _5346_ (.Y(_1843_),
    .B1(net1081),
    .B2(_0019_),
    .A2(net1092),
    .A1(_2696_));
 sg13g2_o21ai_1 _5347_ (.B1(_1843_),
    .Y(_1844_),
    .A1(\dtop.vtop.dphases[2][5] ),
    .A2(_1011_));
 sg13g2_nand2b_1 _5348_ (.Y(_1845_),
    .B(net1161),
    .A_N(_1844_));
 sg13g2_o21ai_1 _5349_ (.B1(_1845_),
    .Y(_1846_),
    .A1(net1161),
    .A2(_1832_));
 sg13g2_mux2_1 _5350_ (.A0(_1846_),
    .A1(_1816_),
    .S(net1184),
    .X(_1847_));
 sg13g2_and2_1 _5351_ (.A(_1842_),
    .B(_1847_),
    .X(_1848_));
 sg13g2_or2_1 _5352_ (.X(_1849_),
    .B(_1847_),
    .A(_1842_));
 sg13g2_nand2b_1 _5353_ (.Y(_1850_),
    .B(_1849_),
    .A_N(_1848_));
 sg13g2_inv_1 _5354_ (.Y(_1851_),
    .A(_1850_));
 sg13g2_o21ai_1 _5355_ (.B1(net1122),
    .Y(_1852_),
    .A1(_1840_),
    .A2(_1851_));
 sg13g2_a21oi_1 _5356_ (.A1(_1840_),
    .A2(_1851_),
    .Y(_1853_),
    .B1(_1852_));
 sg13g2_nand2_1 _5357_ (.Y(_1854_),
    .A(_2658_),
    .B(net1230));
 sg13g2_or3_1 _5358_ (.A(net1208),
    .B(_0556_),
    .C(_0981_),
    .X(_1855_));
 sg13g2_o21ai_1 _5359_ (.B1(net1208),
    .Y(_1856_),
    .A1(_0981_),
    .A2(_1854_));
 sg13g2_nand3_1 _5360_ (.B(_1855_),
    .C(_1856_),
    .A(net1112),
    .Y(_1857_));
 sg13g2_nand2b_1 _5361_ (.Y(_1858_),
    .B(net1080),
    .A_N(_0054_));
 sg13g2_nand3_1 _5362_ (.B(_1784_),
    .C(_1786_),
    .A(_0051_),
    .Y(_1859_));
 sg13g2_o21ai_1 _5363_ (.B1(\dtop.detune_counter[4] ),
    .Y(_1860_),
    .A1(_1783_),
    .A2(_1785_));
 sg13g2_nand2_1 _5364_ (.Y(_1861_),
    .A(_1859_),
    .B(_1860_));
 sg13g2_a21oi_1 _5365_ (.A1(_1859_),
    .A2(_1860_),
    .Y(_1862_),
    .B1(_1823_));
 sg13g2_o21ai_1 _5366_ (.B1(net1101),
    .Y(_1863_),
    .A1(_1825_),
    .A2(_1862_));
 sg13g2_nand2_2 _5367_ (.Y(_1864_),
    .A(_1792_),
    .B(_1794_));
 sg13g2_nand2_1 _5368_ (.Y(_1865_),
    .A(_1863_),
    .B(_1864_));
 sg13g2_nand3b_1 _5369_ (.B(_1863_),
    .C(_1864_),
    .Y(_1866_),
    .A_N(_1858_));
 sg13g2_a21oi_1 _5370_ (.A1(_1858_),
    .A2(_1865_),
    .Y(_1867_),
    .B1(net1122));
 sg13g2_a21o_1 _5371_ (.A2(_1867_),
    .A1(_1866_),
    .B1(_1853_),
    .X(_1868_));
 sg13g2_mux2_1 _5372_ (.A0(net399),
    .A1(_1868_),
    .S(net1067),
    .X(_0192_));
 sg13g2_a21o_1 _5373_ (.A2(_1849_),
    .A1(_1840_),
    .B1(_1848_),
    .X(_1869_));
 sg13g2_nand2b_1 _5374_ (.Y(_1870_),
    .B(net1092),
    .A_N(\dtop.vtop.dphases[1][6] ));
 sg13g2_o21ai_1 _5375_ (.B1(_1870_),
    .Y(_1871_),
    .A1(\dtop.vtop.dphases[2][6] ),
    .A2(_1011_));
 sg13g2_a21oi_1 _5376_ (.A1(_0021_),
    .A2(net1081),
    .Y(_1872_),
    .B1(_1871_));
 sg13g2_nor2_1 _5377_ (.A(net1187),
    .B(_1872_),
    .Y(_1873_));
 sg13g2_a21oi_1 _5378_ (.A1(net1187),
    .A2(_1844_),
    .Y(_1874_),
    .B1(_1873_));
 sg13g2_mux2_1 _5379_ (.A0(_1874_),
    .A1(_1834_),
    .S(net1184),
    .X(_1875_));
 sg13g2_and2_1 _5380_ (.A(_1068_),
    .B(_1875_),
    .X(_1876_));
 sg13g2_xnor2_1 _5381_ (.Y(_1877_),
    .A(_1069_),
    .B(_1875_));
 sg13g2_xor2_1 _5382_ (.B(_1877_),
    .A(_1869_),
    .X(_1878_));
 sg13g2_and2_1 _5383_ (.A(_2672_),
    .B(net1080),
    .X(_1879_));
 sg13g2_a21oi_1 _5384_ (.A1(_1784_),
    .A2(_1786_),
    .Y(_1880_),
    .B1(\dtop.detune_counter[5] ));
 sg13g2_nor3_1 _5385_ (.A(_0080_),
    .B(_1783_),
    .C(_1785_),
    .Y(_1881_));
 sg13g2_nor3_1 _5386_ (.A(_1823_),
    .B(_1880_),
    .C(_1881_),
    .Y(_1882_));
 sg13g2_nor3_1 _5387_ (.A(\dtop.detune_counter[4] ),
    .B(_1783_),
    .C(_1824_),
    .Y(_1883_));
 sg13g2_o21ai_1 _5388_ (.B1(net1101),
    .Y(_1884_),
    .A1(_1882_),
    .A2(_1883_));
 sg13g2_and3_1 _5389_ (.X(_1885_),
    .A(_1864_),
    .B(_1879_),
    .C(_1884_));
 sg13g2_nand3_1 _5390_ (.B(_1879_),
    .C(_1884_),
    .A(_1864_),
    .Y(_1886_));
 sg13g2_a21oi_1 _5391_ (.A1(_1864_),
    .A2(_1884_),
    .Y(_1887_),
    .B1(_1879_));
 sg13g2_nor2_1 _5392_ (.A(_1885_),
    .B(_1887_),
    .Y(_1888_));
 sg13g2_xnor2_1 _5393_ (.Y(_1889_),
    .A(_1866_),
    .B(_1888_));
 sg13g2_mux2_1 _5394_ (.A0(_1878_),
    .A1(_1889_),
    .S(net1109),
    .X(_1890_));
 sg13g2_mux2_1 _5395_ (.A0(net433),
    .A1(_1890_),
    .S(net1067),
    .X(_0193_));
 sg13g2_a22oi_1 _5396_ (.Y(_1891_),
    .B1(net1091),
    .B2(\dtop.vtop.dphases[1][7] ),
    .A2(net1093),
    .A1(\dtop.vtop.dphases[2][7] ));
 sg13g2_mux2_1 _5397_ (.A0(_1891_),
    .A1(_0023_),
    .S(net1081),
    .X(_1892_));
 sg13g2_nand2_1 _5398_ (.Y(_1893_),
    .A(net1187),
    .B(_1872_));
 sg13g2_o21ai_1 _5399_ (.B1(_1893_),
    .Y(_1894_),
    .A1(net1187),
    .A2(_1892_));
 sg13g2_mux2_1 _5400_ (.A0(_1894_),
    .A1(_1846_),
    .S(net1184),
    .X(_1895_));
 sg13g2_nand2_1 _5401_ (.Y(_1896_),
    .A(_1059_),
    .B(_1895_));
 sg13g2_xnor2_1 _5402_ (.Y(_1897_),
    .A(_1059_),
    .B(_1895_));
 sg13g2_a21oi_2 _5403_ (.B1(_1876_),
    .Y(_1898_),
    .A2(_1877_),
    .A1(_1869_));
 sg13g2_xnor2_1 _5404_ (.Y(_1899_),
    .A(_1897_),
    .B(_1898_));
 sg13g2_o21ai_1 _5405_ (.B1(_1886_),
    .Y(_1900_),
    .A1(_1866_),
    .A2(_1887_));
 sg13g2_nand2_1 _5406_ (.Y(_1901_),
    .A(net1177),
    .B(net1080));
 sg13g2_mux2_1 _5407_ (.A0(\dtop.detune_counter[6] ),
    .A1(_0079_),
    .S(net1066),
    .X(_1902_));
 sg13g2_mux2_1 _5408_ (.A0(_1861_),
    .A1(_1902_),
    .S(_1824_),
    .X(_1903_));
 sg13g2_mux2_1 _5409_ (.A0(net1066),
    .A1(_1903_),
    .S(net1102),
    .X(_1904_));
 sg13g2_nor2_1 _5410_ (.A(_1901_),
    .B(_1904_),
    .Y(_1905_));
 sg13g2_xor2_1 _5411_ (.B(_1904_),
    .A(_1901_),
    .X(_1906_));
 sg13g2_o21ai_1 _5412_ (.B1(net1110),
    .Y(_1907_),
    .A1(_1900_),
    .A2(_1906_));
 sg13g2_a21o_1 _5413_ (.A2(_1906_),
    .A1(_1900_),
    .B1(_1907_),
    .X(_1908_));
 sg13g2_o21ai_1 _5414_ (.B1(_1908_),
    .Y(_1909_),
    .A1(net1109),
    .A2(_1899_));
 sg13g2_mux2_1 _5415_ (.A0(net389),
    .A1(_1909_),
    .S(net1068),
    .X(_0194_));
 sg13g2_o21ai_1 _5416_ (.B1(_1896_),
    .Y(_1910_),
    .A1(_1897_),
    .A2(_1898_));
 sg13g2_nand2b_1 _5417_ (.Y(_1911_),
    .B(net1091),
    .A_N(\dtop.vtop.dphases[1][8] ));
 sg13g2_o21ai_1 _5418_ (.B1(_1911_),
    .Y(_1912_),
    .A1(\dtop.vtop.dphases[2][8] ),
    .A2(_1011_));
 sg13g2_a21oi_1 _5419_ (.A1(_0026_),
    .A2(net1081),
    .Y(_1913_),
    .B1(_1912_));
 sg13g2_nor2_1 _5420_ (.A(net1187),
    .B(_1913_),
    .Y(_1914_));
 sg13g2_a21oi_1 _5421_ (.A1(net1187),
    .A2(_1892_),
    .Y(_1915_),
    .B1(_1914_));
 sg13g2_mux2_1 _5422_ (.A0(_1915_),
    .A1(_1874_),
    .S(net1185),
    .X(_1916_));
 sg13g2_and2_1 _5423_ (.A(_1087_),
    .B(_1916_),
    .X(_1917_));
 sg13g2_xor2_1 _5424_ (.B(_1916_),
    .A(_1087_),
    .X(_1918_));
 sg13g2_o21ai_1 _5425_ (.B1(net1122),
    .Y(_1919_),
    .A1(_1910_),
    .A2(_1918_));
 sg13g2_a21o_1 _5426_ (.A2(_1918_),
    .A1(_1910_),
    .B1(_1919_),
    .X(_1920_));
 sg13g2_a21oi_1 _5427_ (.A1(_1900_),
    .A2(_1906_),
    .Y(_1921_),
    .B1(_1905_));
 sg13g2_nand2_1 _5428_ (.Y(_1922_),
    .A(net1176),
    .B(net1080));
 sg13g2_nand2b_1 _5429_ (.Y(_1923_),
    .B(_1794_),
    .A_N(_1826_));
 sg13g2_nor2_1 _5430_ (.A(net1236),
    .B(net1064),
    .Y(_1924_));
 sg13g2_a21oi_1 _5431_ (.A1(_2684_),
    .A2(net1064),
    .Y(_1925_),
    .B1(_1924_));
 sg13g2_o21ai_1 _5432_ (.B1(_1823_),
    .Y(_1926_),
    .A1(_1880_),
    .A2(_1881_));
 sg13g2_o21ai_1 _5433_ (.B1(_1926_),
    .Y(_1927_),
    .A1(_1823_),
    .A2(_1925_));
 sg13g2_o21ai_1 _5434_ (.B1(_1923_),
    .Y(_1928_),
    .A1(_1794_),
    .A2(_1927_));
 sg13g2_or2_1 _5435_ (.X(_1929_),
    .B(_1928_),
    .A(_1922_));
 sg13g2_xnor2_1 _5436_ (.Y(_1930_),
    .A(_1922_),
    .B(_1928_));
 sg13g2_xnor2_1 _5437_ (.Y(_1931_),
    .A(_1921_),
    .B(_1930_));
 sg13g2_o21ai_1 _5438_ (.B1(_1920_),
    .Y(_1932_),
    .A1(net1122),
    .A2(_1931_));
 sg13g2_mux2_1 _5439_ (.A0(net436),
    .A1(_1932_),
    .S(net1068),
    .X(_0195_));
 sg13g2_o21ai_1 _5440_ (.B1(_1929_),
    .Y(_1933_),
    .A1(_1921_),
    .A2(_1930_));
 sg13g2_nand2_1 _5441_ (.Y(_1934_),
    .A(net1174),
    .B(net1080));
 sg13g2_mux2_1 _5442_ (.A0(net1235),
    .A1(_0075_),
    .S(net1064),
    .X(_1935_));
 sg13g2_mux4_1 _5443_ (.S0(_1824_),
    .A0(net1066),
    .A1(_1861_),
    .A2(_1902_),
    .A3(_1935_),
    .S1(net1101),
    .X(_1936_));
 sg13g2_nor2_1 _5444_ (.A(_1934_),
    .B(_1936_),
    .Y(_1937_));
 sg13g2_xor2_1 _5445_ (.B(_1936_),
    .A(_1934_),
    .X(_1938_));
 sg13g2_xnor2_1 _5446_ (.Y(_1939_),
    .A(_1933_),
    .B(_1938_));
 sg13g2_a21oi_1 _5447_ (.A1(_1910_),
    .A2(_1918_),
    .Y(_1940_),
    .B1(_1917_));
 sg13g2_a22oi_1 _5448_ (.Y(_1941_),
    .B1(net1081),
    .B2(_0028_),
    .A2(net1091),
    .A1(_2698_));
 sg13g2_o21ai_1 _5449_ (.B1(_1941_),
    .Y(_1942_),
    .A1(\dtop.vtop.dphases[2][9] ),
    .A2(_1011_));
 sg13g2_nand2_1 _5450_ (.Y(_1943_),
    .A(net1187),
    .B(_1913_));
 sg13g2_o21ai_1 _5451_ (.B1(_1943_),
    .Y(_1944_),
    .A1(net1187),
    .A2(_1942_));
 sg13g2_mux2_1 _5452_ (.A0(_1944_),
    .A1(_1894_),
    .S(net1185),
    .X(_1945_));
 sg13g2_or2_1 _5453_ (.X(_1946_),
    .B(_1945_),
    .A(_1049_));
 sg13g2_inv_1 _5454_ (.Y(_1947_),
    .A(_1946_));
 sg13g2_nand2_1 _5455_ (.Y(_1948_),
    .A(_1049_),
    .B(_1945_));
 sg13g2_nand2_1 _5456_ (.Y(_1949_),
    .A(_1946_),
    .B(_1948_));
 sg13g2_xor2_1 _5457_ (.B(_1949_),
    .A(_1940_),
    .X(_1950_));
 sg13g2_nor2_1 _5458_ (.A(net1110),
    .B(_1950_),
    .Y(_1951_));
 sg13g2_a21oi_2 _5459_ (.B1(_1951_),
    .Y(_1952_),
    .A2(_1939_),
    .A1(net1109));
 sg13g2_mux2_1 _5460_ (.A0(net468),
    .A1(_1952_),
    .S(_1757_),
    .X(_0196_));
 sg13g2_nand2b_1 _5461_ (.Y(_1953_),
    .B(net1091),
    .A_N(\dtop.vtop.dphases[1][10] ));
 sg13g2_o21ai_1 _5462_ (.B1(_1953_),
    .Y(_1954_),
    .A1(\dtop.vtop.dphases[2][10] ),
    .A2(_1011_));
 sg13g2_a21oi_2 _5463_ (.B1(_1954_),
    .Y(_1955_),
    .A2(net1081),
    .A1(_0030_));
 sg13g2_inv_1 _5464_ (.Y(_1956_),
    .A(_1955_));
 sg13g2_nor2_1 _5465_ (.A(net1161),
    .B(_1942_),
    .Y(_1957_));
 sg13g2_a21oi_1 _5466_ (.A1(_2691_),
    .A2(_1955_),
    .Y(_1958_),
    .B1(_1957_));
 sg13g2_nand2_1 _5467_ (.Y(_1959_),
    .A(net1185),
    .B(_1915_));
 sg13g2_o21ai_1 _5468_ (.B1(_1959_),
    .Y(_1960_),
    .A1(net1185),
    .A2(_1958_));
 sg13g2_xnor2_1 _5469_ (.Y(_1961_),
    .A(_1038_),
    .B(_1960_));
 sg13g2_o21ai_1 _5470_ (.B1(_1948_),
    .Y(_1962_),
    .A1(_1940_),
    .A2(_1947_));
 sg13g2_nor2b_1 _5471_ (.A(_1961_),
    .B_N(_1962_),
    .Y(_1963_));
 sg13g2_xor2_1 _5472_ (.B(_1962_),
    .A(_1961_),
    .X(_1964_));
 sg13g2_a21oi_1 _5473_ (.A1(_1933_),
    .A2(_1938_),
    .Y(_1965_),
    .B1(_1937_));
 sg13g2_nand2_1 _5474_ (.Y(_1966_),
    .A(net1169),
    .B(net1080));
 sg13g2_o21ai_1 _5475_ (.B1(_1794_),
    .Y(_1967_),
    .A1(_1882_),
    .A2(_1883_));
 sg13g2_nand2_1 _5476_ (.Y(_1968_),
    .A(net1233),
    .B(net1064));
 sg13g2_o21ai_1 _5477_ (.B1(_1968_),
    .Y(_1969_),
    .A1(_2662_),
    .A2(net1064));
 sg13g2_mux2_1 _5478_ (.A0(_1925_),
    .A1(_1969_),
    .S(_1824_),
    .X(_1970_));
 sg13g2_nand2_1 _5479_ (.Y(_1971_),
    .A(net1101),
    .B(_1970_));
 sg13g2_and2_1 _5480_ (.A(_1967_),
    .B(_1971_),
    .X(_1972_));
 sg13g2_nand2b_1 _5481_ (.Y(_1973_),
    .B(_1972_),
    .A_N(_1966_));
 sg13g2_xnor2_1 _5482_ (.Y(_1974_),
    .A(_1966_),
    .B(_1972_));
 sg13g2_inv_1 _5483_ (.Y(_1975_),
    .A(_1974_));
 sg13g2_xnor2_1 _5484_ (.Y(_1976_),
    .A(_1965_),
    .B(_1974_));
 sg13g2_nand2_1 _5485_ (.Y(_1977_),
    .A(net1109),
    .B(_1976_));
 sg13g2_o21ai_1 _5486_ (.B1(_1977_),
    .Y(_1978_),
    .A1(net1109),
    .A2(_1964_));
 sg13g2_mux2_1 _5487_ (.A0(net403),
    .A1(_1978_),
    .S(net1068),
    .X(_0197_));
 sg13g2_a21oi_1 _5488_ (.A1(_1038_),
    .A2(_1960_),
    .Y(_1979_),
    .B1(_1963_));
 sg13g2_nor2_1 _5489_ (.A(net1185),
    .B(_1955_),
    .Y(_1980_));
 sg13g2_mux2_1 _5490_ (.A0(_1955_),
    .A1(_1944_),
    .S(net1184),
    .X(_1981_));
 sg13g2_and2_1 _5491_ (.A(_1043_),
    .B(_1981_),
    .X(_1982_));
 sg13g2_inv_1 _5492_ (.Y(_1983_),
    .A(_1982_));
 sg13g2_nor2_1 _5493_ (.A(_1043_),
    .B(_1981_),
    .Y(_1984_));
 sg13g2_or2_1 _5494_ (.X(_1985_),
    .B(_1984_),
    .A(_1982_));
 sg13g2_a21oi_1 _5495_ (.A1(_1979_),
    .A2(_1985_),
    .Y(_1986_),
    .B1(net1109));
 sg13g2_o21ai_1 _5496_ (.B1(_1986_),
    .Y(_1987_),
    .A1(_1979_),
    .A2(_1985_));
 sg13g2_o21ai_1 _5497_ (.B1(_1973_),
    .Y(_1988_),
    .A1(_1965_),
    .A2(_1975_));
 sg13g2_nand2_1 _5498_ (.Y(_1989_),
    .A(net1167),
    .B(net1080));
 sg13g2_mux2_1 _5499_ (.A0(\dtop.detune_counter[10] ),
    .A1(_0072_),
    .S(net1064),
    .X(_1990_));
 sg13g2_mux2_1 _5500_ (.A0(_1935_),
    .A1(_1990_),
    .S(_1824_),
    .X(_1991_));
 sg13g2_mux2_1 _5501_ (.A0(_1903_),
    .A1(_1991_),
    .S(net1101),
    .X(_1992_));
 sg13g2_nor2_1 _5502_ (.A(_1989_),
    .B(_1992_),
    .Y(_1993_));
 sg13g2_nand2_1 _5503_ (.Y(_1994_),
    .A(_1989_),
    .B(_1992_));
 sg13g2_nand2b_1 _5504_ (.Y(_1995_),
    .B(_1994_),
    .A_N(_1993_));
 sg13g2_xor2_1 _5505_ (.B(_1995_),
    .A(_1988_),
    .X(_1996_));
 sg13g2_o21ai_1 _5506_ (.B1(_1987_),
    .Y(_1997_),
    .A1(net1125),
    .A2(_1996_));
 sg13g2_mux2_1 _5507_ (.A0(net437),
    .A1(_1997_),
    .S(net1068),
    .X(_0198_));
 sg13g2_a21oi_1 _5508_ (.A1(net1184),
    .A2(_1958_),
    .Y(_1998_),
    .B1(_1980_));
 sg13g2_nand2_1 _5509_ (.Y(_1999_),
    .A(_1025_),
    .B(_1998_));
 sg13g2_inv_1 _5510_ (.Y(_2000_),
    .A(_1999_));
 sg13g2_xor2_1 _5511_ (.B(_1998_),
    .A(_1025_),
    .X(_2001_));
 sg13g2_o21ai_1 _5512_ (.B1(_1983_),
    .Y(_2002_),
    .A1(_1979_),
    .A2(_1984_));
 sg13g2_xnor2_1 _5513_ (.Y(_2003_),
    .A(_2001_),
    .B(_2002_));
 sg13g2_a21oi_1 _5514_ (.A1(_1988_),
    .A2(_1994_),
    .Y(_2004_),
    .B1(_1993_));
 sg13g2_nand2_1 _5515_ (.Y(_2005_),
    .A(net1166),
    .B(net1080));
 sg13g2_mux4_1 _5516_ (.S0(_1823_),
    .A0(net1231),
    .A1(\dtop.detune_counter[9] ),
    .A2(_0070_),
    .A3(net1233),
    .S1(net1064),
    .X(_2006_));
 sg13g2_nand2_1 _5517_ (.Y(_2007_),
    .A(net1102),
    .B(_2006_));
 sg13g2_o21ai_1 _5518_ (.B1(_2007_),
    .Y(_2008_),
    .A1(net1101),
    .A2(_1927_));
 sg13g2_or2_1 _5519_ (.X(_2009_),
    .B(_2008_),
    .A(_2005_));
 sg13g2_xnor2_1 _5520_ (.Y(_2010_),
    .A(_2005_),
    .B(_2008_));
 sg13g2_xor2_1 _5521_ (.B(_2010_),
    .A(_2004_),
    .X(_2011_));
 sg13g2_nor2_1 _5522_ (.A(net1122),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_a21oi_2 _5523_ (.B1(_2012_),
    .Y(_2013_),
    .A2(_2003_),
    .A1(net1125));
 sg13g2_mux2_1 _5524_ (.A0(net427),
    .A1(_2013_),
    .S(net1067),
    .X(_0199_));
 sg13g2_o21ai_1 _5525_ (.B1(_2009_),
    .Y(_2014_),
    .A1(_2004_),
    .A2(_2010_));
 sg13g2_nand2_1 _5526_ (.Y(_2015_),
    .A(\dtop.vtop.logo.addr[9] ),
    .B(_1857_));
 sg13g2_nand2_1 _5527_ (.Y(_2016_),
    .A(_0087_),
    .B(net1065));
 sg13g2_o21ai_1 _5528_ (.B1(_2016_),
    .Y(_2017_),
    .A1(_2659_),
    .A2(net1065));
 sg13g2_mux4_1 _5529_ (.S0(_1824_),
    .A0(_1902_),
    .A1(_1935_),
    .A2(_1990_),
    .A3(_2017_),
    .S1(net1102),
    .X(_2018_));
 sg13g2_nor2_1 _5530_ (.A(_2015_),
    .B(_2018_),
    .Y(_2019_));
 sg13g2_xnor2_1 _5531_ (.Y(_2020_),
    .A(_2015_),
    .B(_2018_));
 sg13g2_inv_1 _5532_ (.Y(_2021_),
    .A(_2020_));
 sg13g2_xnor2_1 _5533_ (.Y(_2022_),
    .A(_2014_),
    .B(_2020_));
 sg13g2_nor2_1 _5534_ (.A(net1123),
    .B(_2022_),
    .Y(_2023_));
 sg13g2_a21o_2 _5535_ (.A2(_2002_),
    .A1(_2001_),
    .B1(_2000_),
    .X(_2024_));
 sg13g2_nand2_1 _5536_ (.Y(_2025_),
    .A(_1031_),
    .B(_1956_));
 sg13g2_nor2_1 _5537_ (.A(_1031_),
    .B(_1956_),
    .Y(_2026_));
 sg13g2_xnor2_1 _5538_ (.Y(_2027_),
    .A(_1031_),
    .B(_1955_));
 sg13g2_xnor2_1 _5539_ (.Y(_2028_),
    .A(_2024_),
    .B(_2027_));
 sg13g2_a21oi_2 _5540_ (.B1(_2023_),
    .Y(_2029_),
    .A2(_2028_),
    .A1(net1123));
 sg13g2_mux2_1 _5541_ (.A0(net409),
    .A1(_2029_),
    .S(net1068),
    .X(_0200_));
 sg13g2_nand2b_1 _5542_ (.Y(_2030_),
    .B(_1955_),
    .A_N(_1014_));
 sg13g2_xor2_1 _5543_ (.B(_1955_),
    .A(_1014_),
    .X(_2031_));
 sg13g2_a21oi_1 _5544_ (.A1(_2024_),
    .A2(_2025_),
    .Y(_2032_),
    .B1(_2026_));
 sg13g2_xnor2_1 _5545_ (.Y(_2033_),
    .A(_2031_),
    .B(_2032_));
 sg13g2_a21oi_2 _5546_ (.B1(_2019_),
    .Y(_2034_),
    .A2(_2021_),
    .A1(_2014_));
 sg13g2_mux4_1 _5547_ (.S0(_1823_),
    .A0(net1230),
    .A1(net1231),
    .A2(_0061_),
    .A3(_0070_),
    .S1(net1064),
    .X(_2035_));
 sg13g2_mux2_1 _5548_ (.A0(_1970_),
    .A1(_2035_),
    .S(net1102),
    .X(_2036_));
 sg13g2_nand4_1 _5549_ (.B(net1208),
    .C(net1112),
    .A(net1220),
    .Y(_2037_),
    .D(_1857_));
 sg13g2_and2_1 _5550_ (.A(_2036_),
    .B(_2037_),
    .X(_2038_));
 sg13g2_or2_1 _5551_ (.X(_2039_),
    .B(_2037_),
    .A(_2036_));
 sg13g2_nor2b_1 _5552_ (.A(_2038_),
    .B_N(_2039_),
    .Y(_2040_));
 sg13g2_xnor2_1 _5553_ (.Y(_2041_),
    .A(_2034_),
    .B(_2040_));
 sg13g2_nand2_1 _5554_ (.Y(_2042_),
    .A(net1111),
    .B(_2041_));
 sg13g2_o21ai_1 _5555_ (.B1(_2042_),
    .Y(_2043_),
    .A1(net1112),
    .A2(_2033_));
 sg13g2_mux2_1 _5556_ (.A0(net497),
    .A1(_2043_),
    .S(net1068),
    .X(_0201_));
 sg13g2_o21ai_1 _5557_ (.B1(_2039_),
    .Y(_2044_),
    .A1(_2034_),
    .A2(_2038_));
 sg13g2_nand2_1 _5558_ (.Y(_2045_),
    .A(_0000_),
    .B(net1065));
 sg13g2_o21ai_1 _5559_ (.B1(_2045_),
    .Y(_2046_),
    .A1(_2658_),
    .A2(net1065));
 sg13g2_nand2_1 _5560_ (.Y(_2047_),
    .A(_1824_),
    .B(_2046_));
 sg13g2_a21oi_1 _5561_ (.A1(_1823_),
    .A2(_2017_),
    .Y(_2048_),
    .B1(_1794_));
 sg13g2_nor2_1 _5562_ (.A(net1102),
    .B(_1991_),
    .Y(_2049_));
 sg13g2_a21oi_1 _5563_ (.A1(_2047_),
    .A2(_2048_),
    .Y(_2050_),
    .B1(_2049_));
 sg13g2_xnor2_1 _5564_ (.Y(_2051_),
    .A(_2044_),
    .B(_2050_));
 sg13g2_nor2_1 _5565_ (.A(net1124),
    .B(_2051_),
    .Y(_2052_));
 sg13g2_o21ai_1 _5566_ (.B1(_2030_),
    .Y(_2053_),
    .A1(_2031_),
    .A2(_2032_));
 sg13g2_xnor2_1 _5567_ (.Y(_2054_),
    .A(_0998_),
    .B(_1955_));
 sg13g2_xnor2_1 _5568_ (.Y(_2055_),
    .A(_2053_),
    .B(_2054_));
 sg13g2_a21oi_2 _5569_ (.B1(_2052_),
    .Y(_2056_),
    .A2(_2055_),
    .A1(net1123));
 sg13g2_mux2_1 _5570_ (.A0(net466),
    .A1(_2056_),
    .S(net1068),
    .X(_0202_));
 sg13g2_a22oi_1 _5571_ (.Y(_2057_),
    .B1(_0979_),
    .B2(_1479_),
    .A2(_0977_),
    .A1(net1215));
 sg13g2_mux2_1 _5572_ (.A0(_1767_),
    .A1(net494),
    .S(net983),
    .X(_0203_));
 sg13g2_mux2_1 _5573_ (.A0(_1797_),
    .A1(net480),
    .S(net983),
    .X(_0204_));
 sg13g2_mux2_1 _5574_ (.A0(_1808_),
    .A1(net509),
    .S(net983),
    .X(_0205_));
 sg13g2_mux2_1 _5575_ (.A0(_1822_),
    .A1(net502),
    .S(net984),
    .X(_0206_));
 sg13g2_mux2_1 _5576_ (.A0(_1839_),
    .A1(net477),
    .S(net983),
    .X(_0207_));
 sg13g2_mux2_1 _5577_ (.A0(_1868_),
    .A1(net489),
    .S(net983),
    .X(_0208_));
 sg13g2_mux2_1 _5578_ (.A0(_1890_),
    .A1(net513),
    .S(net983),
    .X(_0209_));
 sg13g2_mux2_1 _5579_ (.A0(_1909_),
    .A1(net496),
    .S(_2057_),
    .X(_0210_));
 sg13g2_mux2_1 _5580_ (.A0(_1932_),
    .A1(net465),
    .S(net984),
    .X(_0211_));
 sg13g2_mux2_1 _5581_ (.A0(_1952_),
    .A1(net479),
    .S(net984),
    .X(_0212_));
 sg13g2_mux2_1 _5582_ (.A0(_1978_),
    .A1(net481),
    .S(net983),
    .X(_0213_));
 sg13g2_mux2_1 _5583_ (.A0(_1997_),
    .A1(net482),
    .S(net984),
    .X(_0214_));
 sg13g2_mux2_1 _5584_ (.A0(_2013_),
    .A1(net459),
    .S(net983),
    .X(_0215_));
 sg13g2_mux2_1 _5585_ (.A0(_2029_),
    .A1(net498),
    .S(net984),
    .X(_0216_));
 sg13g2_mux2_1 _5586_ (.A0(_2043_),
    .A1(net483),
    .S(net984),
    .X(_0217_));
 sg13g2_mux2_1 _5587_ (.A0(_2056_),
    .A1(net532),
    .S(net984),
    .X(_0218_));
 sg13g2_and2_1 _5588_ (.A(net557),
    .B(net1250),
    .X(_0219_));
 sg13g2_nor2_2 _5589_ (.A(\dtop.vtop.pipeline.wave_index[0] ),
    .B(\dtop.vtop.pipeline.wave_index[1] ),
    .Y(_2058_));
 sg13g2_or2_2 _5590_ (.X(_2059_),
    .B(\dtop.vtop.pipeline.wave_index[1] ),
    .A(\dtop.vtop.pipeline.wave_index[0] ));
 sg13g2_a22oi_1 _5591_ (.Y(_2060_),
    .B1(_2058_),
    .B2(net1124),
    .A2(_0977_),
    .A1(net1162));
 sg13g2_mux2_1 _5592_ (.A0(_1767_),
    .A1(net424),
    .S(net1078),
    .X(_0220_));
 sg13g2_mux2_1 _5593_ (.A0(_1797_),
    .A1(net431),
    .S(net1078),
    .X(_0221_));
 sg13g2_mux2_1 _5594_ (.A0(_1808_),
    .A1(net432),
    .S(net1078),
    .X(_0222_));
 sg13g2_mux2_1 _5595_ (.A0(_1822_),
    .A1(net440),
    .S(net1079),
    .X(_0223_));
 sg13g2_mux2_1 _5596_ (.A0(_1839_),
    .A1(net426),
    .S(net1078),
    .X(_0224_));
 sg13g2_mux2_1 _5597_ (.A0(_1868_),
    .A1(net412),
    .S(net1078),
    .X(_0225_));
 sg13g2_mux2_1 _5598_ (.A0(_1890_),
    .A1(net423),
    .S(net1078),
    .X(_0226_));
 sg13g2_mux2_1 _5599_ (.A0(_1909_),
    .A1(net404),
    .S(_2060_),
    .X(_0227_));
 sg13g2_mux2_1 _5600_ (.A0(_1932_),
    .A1(net438),
    .S(net1079),
    .X(_0228_));
 sg13g2_mux2_1 _5601_ (.A0(_1952_),
    .A1(net415),
    .S(net1079),
    .X(_0229_));
 sg13g2_mux2_1 _5602_ (.A0(_1978_),
    .A1(net464),
    .S(net1078),
    .X(_0230_));
 sg13g2_mux2_1 _5603_ (.A0(_1997_),
    .A1(net455),
    .S(net1079),
    .X(_0231_));
 sg13g2_mux2_1 _5604_ (.A0(_2013_),
    .A1(net422),
    .S(net1078),
    .X(_0232_));
 sg13g2_mux2_1 _5605_ (.A0(_2029_),
    .A1(net434),
    .S(net1079),
    .X(_0233_));
 sg13g2_mux2_1 _5606_ (.A0(_2043_),
    .A1(net456),
    .S(net1079),
    .X(_0234_));
 sg13g2_mux2_1 _5607_ (.A0(_2056_),
    .A1(net435),
    .S(net1079),
    .X(_0235_));
 sg13g2_nor2_2 _5608_ (.A(_0994_),
    .B(_2058_),
    .Y(_2061_));
 sg13g2_nand2_1 _5609_ (.Y(_2062_),
    .A(\dtop.vtop.pipeline.zg_acc[0] ),
    .B(net1063));
 sg13g2_nor2_1 _5610_ (.A(_1272_),
    .B(_2062_),
    .Y(_2063_));
 sg13g2_xor2_1 _5611_ (.B(_2062_),
    .A(_1272_),
    .X(_2064_));
 sg13g2_mux2_1 _5612_ (.A0(net503),
    .A1(_2064_),
    .S(net1039),
    .X(_0236_));
 sg13g2_nand2_1 _5613_ (.Y(_2065_),
    .A(_2697_),
    .B(net1063));
 sg13g2_nor2_1 _5614_ (.A(_1294_),
    .B(_2065_),
    .Y(_2066_));
 sg13g2_xor2_1 _5615_ (.B(_2065_),
    .A(_1294_),
    .X(_2067_));
 sg13g2_xor2_1 _5616_ (.B(_2067_),
    .A(_2063_),
    .X(_2068_));
 sg13g2_mux2_1 _5617_ (.A0(net330),
    .A1(_2068_),
    .S(net1039),
    .X(_0237_));
 sg13g2_a21o_1 _5618_ (.A2(_2067_),
    .A1(_2063_),
    .B1(_2066_),
    .X(_2069_));
 sg13g2_nand2_1 _5619_ (.Y(_2070_),
    .A(\dtop.vtop.pipeline.zg_acc[2] ),
    .B(net1063));
 sg13g2_and3_1 _5620_ (.X(_2071_),
    .A(\dtop.vtop.pipeline.zg_acc[2] ),
    .B(_1304_),
    .C(net1063));
 sg13g2_xnor2_1 _5621_ (.Y(_2072_),
    .A(_1304_),
    .B(_2070_));
 sg13g2_xor2_1 _5622_ (.B(_2072_),
    .A(_2069_),
    .X(_2073_));
 sg13g2_mux2_1 _5623_ (.A0(net504),
    .A1(_2073_),
    .S(net1039),
    .X(_0238_));
 sg13g2_a21oi_1 _5624_ (.A1(_2069_),
    .A2(_2072_),
    .Y(_2074_),
    .B1(_2071_));
 sg13g2_nand2_1 _5625_ (.Y(_2075_),
    .A(\dtop.vtop.pipeline.zg_acc[3] ),
    .B(net1063));
 sg13g2_nand3_1 _5626_ (.B(_1311_),
    .C(net1063),
    .A(\dtop.vtop.pipeline.zg_acc[3] ),
    .Y(_2076_));
 sg13g2_xor2_1 _5627_ (.B(_2075_),
    .A(_1311_),
    .X(_2077_));
 sg13g2_xor2_1 _5628_ (.B(_2077_),
    .A(_2074_),
    .X(_2078_));
 sg13g2_mux2_1 _5629_ (.A0(net545),
    .A1(_2078_),
    .S(net1039),
    .X(_0239_));
 sg13g2_o21ai_1 _5630_ (.B1(_2076_),
    .Y(_2079_),
    .A1(_2074_),
    .A2(_2077_));
 sg13g2_nand2_1 _5631_ (.Y(_2080_),
    .A(\dtop.vtop.pipeline.zg_acc[4] ),
    .B(net1063));
 sg13g2_nor2_1 _5632_ (.A(_1318_),
    .B(_2080_),
    .Y(_2081_));
 sg13g2_xor2_1 _5633_ (.B(_2080_),
    .A(_1318_),
    .X(_2082_));
 sg13g2_xor2_1 _5634_ (.B(_2082_),
    .A(_2079_),
    .X(_2083_));
 sg13g2_mux2_1 _5635_ (.A0(net510),
    .A1(_2083_),
    .S(net1039),
    .X(_0240_));
 sg13g2_a21oi_1 _5636_ (.A1(_2079_),
    .A2(_2082_),
    .Y(_2084_),
    .B1(_2081_));
 sg13g2_and2_1 _5637_ (.A(\dtop.vtop.pipeline.zg_acc[5] ),
    .B(net1063),
    .X(_2085_));
 sg13g2_nor2_1 _5638_ (.A(_1323_),
    .B(_2085_),
    .Y(_2086_));
 sg13g2_xor2_1 _5639_ (.B(_2085_),
    .A(_1323_),
    .X(_2087_));
 sg13g2_xnor2_1 _5640_ (.Y(_2088_),
    .A(_2084_),
    .B(_2087_));
 sg13g2_mux2_1 _5641_ (.A0(net505),
    .A1(_2088_),
    .S(net1039),
    .X(_0241_));
 sg13g2_nor3_1 _5642_ (.A(_0034_),
    .B(net1094),
    .C(_2058_),
    .Y(_2089_));
 sg13g2_nor2_1 _5643_ (.A(_1326_),
    .B(_2089_),
    .Y(_2090_));
 sg13g2_nand2_1 _5644_ (.Y(_2091_),
    .A(_1326_),
    .B(_2089_));
 sg13g2_nand2b_1 _5645_ (.Y(_2092_),
    .B(_2091_),
    .A_N(_2090_));
 sg13g2_a221oi_1 _5646_ (.B2(_1323_),
    .C1(_2081_),
    .B1(_2085_),
    .A1(_2079_),
    .Y(_2093_),
    .A2(_2082_));
 sg13g2_nor2_1 _5647_ (.A(_2086_),
    .B(_2093_),
    .Y(_2094_));
 sg13g2_xnor2_1 _5648_ (.Y(_2095_),
    .A(_2092_),
    .B(_2094_));
 sg13g2_mux2_1 _5649_ (.A0(net363),
    .A1(_2095_),
    .S(net1040),
    .X(_0242_));
 sg13g2_o21ai_1 _5650_ (.B1(_2091_),
    .Y(_2096_),
    .A1(_2086_),
    .A2(_2093_));
 sg13g2_nand2b_1 _5651_ (.Y(_2097_),
    .B(_2096_),
    .A_N(_2090_));
 sg13g2_nand2b_1 _5652_ (.Y(_2098_),
    .B(_2061_),
    .A_N(_0036_));
 sg13g2_nor2_1 _5653_ (.A(_1329_),
    .B(_2098_),
    .Y(_2099_));
 sg13g2_xor2_1 _5654_ (.B(_2098_),
    .A(_1329_),
    .X(_2100_));
 sg13g2_xnor2_1 _5655_ (.Y(_2101_),
    .A(_2097_),
    .B(_2100_));
 sg13g2_mux2_1 _5656_ (.A0(net351),
    .A1(_2101_),
    .S(net1040),
    .X(_0243_));
 sg13g2_a21oi_1 _5657_ (.A1(_1329_),
    .A2(_2098_),
    .Y(_2102_),
    .B1(_2090_));
 sg13g2_a21oi_1 _5658_ (.A1(_2096_),
    .A2(_2102_),
    .Y(_2103_),
    .B1(_2099_));
 sg13g2_nand2_1 _5659_ (.Y(_2104_),
    .A(_0038_),
    .B(_2061_));
 sg13g2_o21ai_1 _5660_ (.B1(_2104_),
    .Y(_2105_),
    .A1(_0984_),
    .A2(_2061_));
 sg13g2_nand2b_1 _5661_ (.Y(_2106_),
    .B(_0997_),
    .A_N(_2105_));
 sg13g2_and2_1 _5662_ (.A(_0998_),
    .B(_2105_),
    .X(_2107_));
 sg13g2_xnor2_1 _5663_ (.Y(_2108_),
    .A(_0997_),
    .B(_2105_));
 sg13g2_xnor2_1 _5664_ (.Y(_2109_),
    .A(_2103_),
    .B(_2108_));
 sg13g2_nor2_1 _5665_ (.A(net1059),
    .B(_2109_),
    .Y(_2110_));
 sg13g2_a21oi_1 _5666_ (.A1(_2687_),
    .A2(net1059),
    .Y(_0244_),
    .B1(_2110_));
 sg13g2_o21ai_1 _5667_ (.B1(_2106_),
    .Y(_2111_),
    .A1(_2103_),
    .A2(_2107_));
 sg13g2_nor3_1 _5668_ (.A(\dtop.vtop.pipeline.zg_acc[9] ),
    .B(net1094),
    .C(_2058_),
    .Y(_2112_));
 sg13g2_xnor2_1 _5669_ (.Y(_2113_),
    .A(_0998_),
    .B(_2112_));
 sg13g2_xnor2_1 _5670_ (.Y(_2114_),
    .A(_2111_),
    .B(_2113_));
 sg13g2_mux2_1 _5671_ (.A0(net452),
    .A1(_2114_),
    .S(net1039),
    .X(_0245_));
 sg13g2_a21oi_1 _5672_ (.A1(_1479_),
    .A2(net1039),
    .Y(_0246_),
    .B1(net1113));
 sg13g2_mux2_1 _5673_ (.A0(_2064_),
    .A1(net467),
    .S(_1487_),
    .X(_0247_));
 sg13g2_mux2_1 _5674_ (.A0(_2068_),
    .A1(net523),
    .S(net993),
    .X(_0248_));
 sg13g2_mux2_1 _5675_ (.A0(_2073_),
    .A1(net540),
    .S(net991),
    .X(_0249_));
 sg13g2_nor2_1 _5676_ (.A(net991),
    .B(_2078_),
    .Y(_2115_));
 sg13g2_a21oi_1 _5677_ (.A1(_2679_),
    .A2(net991),
    .Y(_0250_),
    .B1(_2115_));
 sg13g2_nor2_1 _5678_ (.A(net991),
    .B(_2083_),
    .Y(_2116_));
 sg13g2_a21oi_1 _5679_ (.A1(_2678_),
    .A2(net991),
    .Y(_0251_),
    .B1(_2116_));
 sg13g2_nor2_1 _5680_ (.A(net991),
    .B(_2088_),
    .Y(_2117_));
 sg13g2_a21oi_1 _5681_ (.A1(_2677_),
    .A2(net993),
    .Y(_0252_),
    .B1(_2117_));
 sg13g2_mux2_1 _5682_ (.A0(_2095_),
    .A1(net625),
    .S(net992),
    .X(_0253_));
 sg13g2_mux2_1 _5683_ (.A0(_2101_),
    .A1(net624),
    .S(net992),
    .X(_0254_));
 sg13g2_nor2_1 _5684_ (.A(net992),
    .B(_2109_),
    .Y(_2118_));
 sg13g2_a21oi_1 _5685_ (.A1(_2676_),
    .A2(net991),
    .Y(_0255_),
    .B1(_2118_));
 sg13g2_mux2_1 _5686_ (.A0(_2114_),
    .A1(net645),
    .S(net991),
    .X(_0256_));
 sg13g2_nand2_1 _5687_ (.Y(_2119_),
    .A(net394),
    .B(net1140));
 sg13g2_nand2b_1 _5688_ (.Y(_2120_),
    .B(_1066_),
    .A_N(_2119_));
 sg13g2_a21oi_1 _5689_ (.A1(_1065_),
    .A2(_2119_),
    .Y(_2121_),
    .B1(net1059));
 sg13g2_a22oi_1 _5690_ (.Y(_2122_),
    .B1(_2120_),
    .B2(_2121_),
    .A2(net1059),
    .A1(net394));
 sg13g2_inv_1 _5691_ (.Y(_0257_),
    .A(_2122_));
 sg13g2_nand2_1 _5692_ (.Y(_2123_),
    .A(\dtop.vtop.pipeline.cosappr_acc[1] ),
    .B(net1140));
 sg13g2_inv_1 _5693_ (.Y(_2124_),
    .A(_2123_));
 sg13g2_xnor2_1 _5694_ (.Y(_2125_),
    .A(_1093_),
    .B(_2124_));
 sg13g2_nor2_1 _5695_ (.A(_2120_),
    .B(_2125_),
    .Y(_2126_));
 sg13g2_xnor2_1 _5696_ (.Y(_2127_),
    .A(_2120_),
    .B(_2125_));
 sg13g2_nand2_1 _5697_ (.Y(_2128_),
    .A(net333),
    .B(net1058));
 sg13g2_o21ai_1 _5698_ (.B1(_2128_),
    .Y(_0258_),
    .A1(net1058),
    .A2(_2127_));
 sg13g2_nand2_1 _5699_ (.Y(_2129_),
    .A(\dtop.vtop.pipeline.cosappr_acc[2] ),
    .B(net1140));
 sg13g2_nand2b_1 _5700_ (.Y(_2130_),
    .B(net1015),
    .A_N(_2129_));
 sg13g2_xnor2_1 _5701_ (.Y(_2131_),
    .A(net1019),
    .B(_2129_));
 sg13g2_a21oi_1 _5702_ (.A1(_1093_),
    .A2(_2124_),
    .Y(_2132_),
    .B1(_2126_));
 sg13g2_xnor2_1 _5703_ (.Y(_2133_),
    .A(_2131_),
    .B(_2132_));
 sg13g2_nand2_1 _5704_ (.Y(_2134_),
    .A(net328),
    .B(net1058));
 sg13g2_o21ai_1 _5705_ (.B1(_2134_),
    .Y(_0259_),
    .A1(net1058),
    .A2(_2133_));
 sg13g2_and3_1 _5706_ (.X(_2135_),
    .A(\dtop.vtop.pipeline.cosappr_acc[3] ),
    .B(net1029),
    .C(net1140));
 sg13g2_a21o_1 _5707_ (.A2(net1140),
    .A1(\dtop.vtop.pipeline.cosappr_acc[3] ),
    .B1(net1029),
    .X(_2136_));
 sg13g2_nand2b_1 _5708_ (.Y(_2137_),
    .B(_2136_),
    .A_N(_2135_));
 sg13g2_o21ai_1 _5709_ (.B1(_2130_),
    .Y(_2138_),
    .A1(_2131_),
    .A2(_2132_));
 sg13g2_xor2_1 _5710_ (.B(_2138_),
    .A(_2137_),
    .X(_2139_));
 sg13g2_nand2_1 _5711_ (.Y(_2140_),
    .A(net457),
    .B(net1058));
 sg13g2_o21ai_1 _5712_ (.B1(_2140_),
    .Y(_0260_),
    .A1(net1058),
    .A2(_2139_));
 sg13g2_a21oi_1 _5713_ (.A1(_2136_),
    .A2(_2138_),
    .Y(_2141_),
    .B1(_2135_));
 sg13g2_nand2_1 _5714_ (.Y(_2142_),
    .A(\dtop.vtop.pipeline.cosappr_acc[4] ),
    .B(net1140));
 sg13g2_nor2_1 _5715_ (.A(_1044_),
    .B(_2142_),
    .Y(_2143_));
 sg13g2_xnor2_1 _5716_ (.Y(_2144_),
    .A(_1044_),
    .B(_2142_));
 sg13g2_nor2_1 _5717_ (.A(_2141_),
    .B(_2144_),
    .Y(_2145_));
 sg13g2_xnor2_1 _5718_ (.Y(_2146_),
    .A(_2141_),
    .B(_2144_));
 sg13g2_nand2_1 _5719_ (.Y(_2147_),
    .A(net359),
    .B(net1058));
 sg13g2_o21ai_1 _5720_ (.B1(_2147_),
    .Y(_0261_),
    .A1(net1058),
    .A2(_2146_));
 sg13g2_nand2_1 _5721_ (.Y(_2148_),
    .A(\dtop.vtop.pipeline.cosappr_acc[5] ),
    .B(_2059_));
 sg13g2_nor2_1 _5722_ (.A(_1026_),
    .B(_2148_),
    .Y(_2149_));
 sg13g2_xnor2_1 _5723_ (.Y(_2150_),
    .A(_1026_),
    .B(_2148_));
 sg13g2_nor2_1 _5724_ (.A(_2143_),
    .B(_2145_),
    .Y(_2151_));
 sg13g2_nor2_1 _5725_ (.A(_2150_),
    .B(_2151_),
    .Y(_2152_));
 sg13g2_xor2_1 _5726_ (.B(_2151_),
    .A(_2150_),
    .X(_2153_));
 sg13g2_mux2_1 _5727_ (.A0(net400),
    .A1(_2153_),
    .S(net1040),
    .X(_0262_));
 sg13g2_nand2_1 _5728_ (.Y(_2154_),
    .A(\dtop.vtop.pipeline.cosappr_acc[6] ),
    .B(_2059_));
 sg13g2_nor2_1 _5729_ (.A(_1032_),
    .B(_2154_),
    .Y(_2155_));
 sg13g2_xnor2_1 _5730_ (.Y(_2156_),
    .A(_1032_),
    .B(_2154_));
 sg13g2_nor2_1 _5731_ (.A(_2149_),
    .B(_2152_),
    .Y(_2157_));
 sg13g2_nor2_1 _5732_ (.A(_2156_),
    .B(_2157_),
    .Y(_2158_));
 sg13g2_xor2_1 _5733_ (.B(_2157_),
    .A(_2156_),
    .X(_2159_));
 sg13g2_mux2_1 _5734_ (.A0(net408),
    .A1(_2159_),
    .S(net1040),
    .X(_0263_));
 sg13g2_nand2_1 _5735_ (.Y(_2160_),
    .A(net414),
    .B(net1140));
 sg13g2_nor2_1 _5736_ (.A(_2155_),
    .B(_2158_),
    .Y(_2161_));
 sg13g2_or2_1 _5737_ (.X(_2162_),
    .B(_2161_),
    .A(_2160_));
 sg13g2_xor2_1 _5738_ (.B(_2161_),
    .A(_2160_),
    .X(_2163_));
 sg13g2_mux2_1 _5739_ (.A0(net414),
    .A1(_2163_),
    .S(net1040),
    .X(_0264_));
 sg13g2_nand3_1 _5740_ (.B(net1140),
    .C(_2162_),
    .A(net475),
    .Y(_2164_));
 sg13g2_o21ai_1 _5741_ (.B1(_2164_),
    .Y(_2165_),
    .A1(net475),
    .A2(_2162_));
 sg13g2_mux2_1 _5742_ (.A0(net475),
    .A1(_2165_),
    .S(net1040),
    .X(_0265_));
 sg13g2_o21ai_1 _5743_ (.B1(_1483_),
    .Y(_2166_),
    .A1(\dtop.vtop.pipeline.wave_index[1] ),
    .A2(_2686_));
 sg13g2_nand2_1 _5744_ (.Y(_2167_),
    .A(net1129),
    .B(net992));
 sg13g2_nor2b_1 _5745_ (.A(_2167_),
    .B_N(net608),
    .Y(_0266_));
 sg13g2_a21oi_1 _5746_ (.A1(_1484_),
    .A2(net611),
    .Y(_0267_),
    .B1(_2167_));
 sg13g2_or3_1 _5747_ (.A(net537),
    .B(\dtop.vtop.pipeline.nstep_counter[0] ),
    .C(net992),
    .X(_2168_));
 sg13g2_or2_1 _5748_ (.X(_2169_),
    .B(_2168_),
    .A(net527));
 sg13g2_or2_2 _5749_ (.X(_2170_),
    .B(_2169_),
    .A(net484));
 sg13g2_nor2_1 _5750_ (.A(\dtop.detune_counter[12] ),
    .B(_0983_),
    .Y(_2171_));
 sg13g2_xor2_1 _5751_ (.B(_2171_),
    .A(_0008_),
    .X(_2172_));
 sg13g2_nor2_1 _5752_ (.A(net1231),
    .B(_0983_),
    .Y(_2173_));
 sg13g2_xnor2_1 _5753_ (.Y(_2174_),
    .A(net1189),
    .B(_2173_));
 sg13g2_nor2_1 _5754_ (.A(_2172_),
    .B(_2174_),
    .Y(_2175_));
 sg13g2_nor3_1 _5755_ (.A(net528),
    .B(_2170_),
    .C(_2175_),
    .Y(_2176_));
 sg13g2_nor2_1 _5756_ (.A(net1189),
    .B(_2176_),
    .Y(_2177_));
 sg13g2_nor4_2 _5757_ (.A(net528),
    .B(_2691_),
    .C(_2170_),
    .Y(_2178_),
    .D(_2175_));
 sg13g2_nor3_1 _5758_ (.A(net1111),
    .B(_2177_),
    .C(_2178_),
    .Y(_0268_));
 sg13g2_xnor2_1 _5759_ (.Y(_2179_),
    .A(net1186),
    .B(_2178_));
 sg13g2_nor2_1 _5760_ (.A(net1111),
    .B(_2179_),
    .Y(_0269_));
 sg13g2_nor2_1 _5761_ (.A(\dtop.vtop.pipeline.nstep_counter[0] ),
    .B(_2167_),
    .Y(_2180_));
 sg13g2_nor2_1 _5762_ (.A(net306),
    .B(_1488_),
    .Y(_2181_));
 sg13g2_nor2_1 _5763_ (.A(_2180_),
    .B(_2181_),
    .Y(_0270_));
 sg13g2_o21ai_1 _5764_ (.B1(net537),
    .Y(_2182_),
    .A1(\dtop.vtop.pipeline.nstep_counter[0] ),
    .A2(net992));
 sg13g2_nand3_1 _5765_ (.B(_2168_),
    .C(net538),
    .A(net1129),
    .Y(_0271_));
 sg13g2_a21oi_1 _5766_ (.A1(net527),
    .A2(_2168_),
    .Y(_2183_),
    .B1(net1114));
 sg13g2_nand2_1 _5767_ (.Y(_0272_),
    .A(_2169_),
    .B(_2183_));
 sg13g2_a21oi_1 _5768_ (.A1(net484),
    .A2(_2169_),
    .Y(_2184_),
    .B1(net1112));
 sg13g2_nand2_1 _5769_ (.Y(_0273_),
    .A(_2170_),
    .B(net485));
 sg13g2_a21o_1 _5770_ (.A2(_2170_),
    .A1(net528),
    .B1(net1111),
    .X(_0274_));
 sg13g2_mux2_1 _5771_ (.A0(_2153_),
    .A1(net541),
    .S(net993),
    .X(_0275_));
 sg13g2_mux2_1 _5772_ (.A0(_2159_),
    .A1(net443),
    .S(net993),
    .X(_0276_));
 sg13g2_mux2_1 _5773_ (.A0(_2163_),
    .A1(net565),
    .S(net993),
    .X(_0277_));
 sg13g2_mux2_1 _5774_ (.A0(_2165_),
    .A1(net595),
    .S(net993),
    .X(_0278_));
 sg13g2_nand2b_1 _5775_ (.Y(_2185_),
    .B(net429),
    .A_N(net1190));
 sg13g2_nor2_1 _5776_ (.A(_2011_),
    .B(_2022_),
    .Y(_2186_));
 sg13g2_nor2_1 _5777_ (.A(_1590_),
    .B(_2186_),
    .Y(_2187_));
 sg13g2_mux2_1 _5778_ (.A0(_1590_),
    .A1(_2187_),
    .S(_2041_),
    .X(_2188_));
 sg13g2_xnor2_1 _5779_ (.Y(_2189_),
    .A(net1141),
    .B(_2051_));
 sg13g2_nor2_1 _5780_ (.A(_2909_),
    .B(_0596_),
    .Y(_2190_));
 sg13g2_nor2_1 _5781_ (.A(_1854_),
    .B(_2190_),
    .Y(_2191_));
 sg13g2_xnor2_1 _5782_ (.Y(_2192_),
    .A(_2188_),
    .B(_2189_));
 sg13g2_a22oi_1 _5783_ (.Y(_2193_),
    .B1(_2191_),
    .B2(_2192_),
    .A2(_0598_),
    .A1(_0557_));
 sg13g2_nor2_1 _5784_ (.A(net1235),
    .B(_2884_),
    .Y(_2194_));
 sg13g2_and3_2 _5785_ (.X(_2195_),
    .A(_2662_),
    .B(_1550_),
    .C(_1581_));
 sg13g2_a21o_2 _5786_ (.A2(_2889_),
    .A1(_0086_),
    .B1(_0559_),
    .X(_2196_));
 sg13g2_nor2_1 _5787_ (.A(_2195_),
    .B(_2196_),
    .Y(_2197_));
 sg13g2_nor3_1 _5788_ (.A(_0083_),
    .B(_2195_),
    .C(_2196_),
    .Y(_2198_));
 sg13g2_o21ai_1 _5789_ (.B1(_0083_),
    .Y(_2199_),
    .A1(_2195_),
    .A2(_2196_));
 sg13g2_nand3b_1 _5790_ (.B(_2199_),
    .C(_2194_),
    .Y(_2200_),
    .A_N(_2198_));
 sg13g2_nor2b_1 _5791_ (.A(_2200_),
    .B_N(_1592_),
    .Y(_2201_));
 sg13g2_xnor2_1 _5792_ (.Y(_2202_),
    .A(_1592_),
    .B(_2200_));
 sg13g2_a21oi_1 _5793_ (.A1(net1177),
    .A2(_2202_),
    .Y(_2203_),
    .B1(_2201_));
 sg13g2_nor3_1 _5794_ (.A(_0051_),
    .B(_2195_),
    .C(_2196_),
    .Y(_2204_));
 sg13g2_o21ai_1 _5795_ (.B1(_0051_),
    .Y(_2205_),
    .A1(_2195_),
    .A2(_2196_));
 sg13g2_nand3b_1 _5796_ (.B(_2205_),
    .C(_2194_),
    .Y(_2206_),
    .A_N(_2204_));
 sg13g2_nand2b_1 _5797_ (.Y(_2207_),
    .B(_1590_),
    .A_N(_2206_));
 sg13g2_xnor2_1 _5798_ (.Y(_2208_),
    .A(_1590_),
    .B(_2206_));
 sg13g2_nand2_1 _5799_ (.Y(_2209_),
    .A(net1176),
    .B(_2208_));
 sg13g2_xnor2_1 _5800_ (.Y(_2210_),
    .A(net1176),
    .B(_2208_));
 sg13g2_nor2_1 _5801_ (.A(_2203_),
    .B(_2210_),
    .Y(_2211_));
 sg13g2_xnor2_1 _5802_ (.Y(_2212_),
    .A(net1177),
    .B(_2202_));
 sg13g2_nor4_2 _5803_ (.A(net1235),
    .B(_2884_),
    .C(_2195_),
    .Y(_2213_),
    .D(_2196_));
 sg13g2_nand2_1 _5804_ (.Y(_2214_),
    .A(_2194_),
    .B(_2197_));
 sg13g2_xnor2_1 _5805_ (.Y(_2215_),
    .A(net1220),
    .B(_2213_));
 sg13g2_a22oi_1 _5806_ (.Y(_2216_),
    .B1(_2215_),
    .B2(\dtop.oct_counter[4] ),
    .A2(_2213_),
    .A1(_0088_));
 sg13g2_or3_1 _5807_ (.A(\dtop.oct_counter[3] ),
    .B(_2668_),
    .C(_2213_),
    .X(_2217_));
 sg13g2_nor2_1 _5808_ (.A(\dtop.player_inst.program_addr[0] ),
    .B(_2214_),
    .Y(_2218_));
 sg13g2_xor2_1 _5809_ (.B(_2215_),
    .A(\dtop.oct_counter[4] ),
    .X(_2219_));
 sg13g2_a22oi_1 _5810_ (.Y(_2220_),
    .B1(_2219_),
    .B2(_2217_),
    .A2(_2218_),
    .A1(\dtop.oct_counter[3] ));
 sg13g2_o21ai_1 _5811_ (.B1(_2212_),
    .Y(_2221_),
    .A1(_2216_),
    .A2(_2220_));
 sg13g2_a22oi_1 _5812_ (.Y(_2222_),
    .B1(_2216_),
    .B2(_2220_),
    .A2(_2210_),
    .A1(_2203_));
 sg13g2_a21oi_1 _5813_ (.A1(_2221_),
    .A2(_2222_),
    .Y(_2223_),
    .B1(_2211_));
 sg13g2_nand2_1 _5814_ (.Y(_2224_),
    .A(_2207_),
    .B(_2209_));
 sg13g2_xor2_1 _5815_ (.B(_2197_),
    .A(\dtop.detune_counter[6] ),
    .X(_2225_));
 sg13g2_nand2_1 _5816_ (.Y(_2226_),
    .A(_2194_),
    .B(_2225_));
 sg13g2_xor2_1 _5817_ (.B(_2226_),
    .A(_2224_),
    .X(_2227_));
 sg13g2_xnor2_1 _5818_ (.Y(_2228_),
    .A(_2223_),
    .B(_2227_));
 sg13g2_nand2_1 _5819_ (.Y(_2229_),
    .A(net1055),
    .B(net959));
 sg13g2_nor2_2 _5820_ (.A(net1056),
    .B(_1583_),
    .Y(_2230_));
 sg13g2_nand2b_1 _5821_ (.Y(_2231_),
    .B(net1005),
    .A_N(_2230_));
 sg13g2_a21oi_1 _5822_ (.A1(net1055),
    .A2(net960),
    .Y(_2232_),
    .B1(_2231_));
 sg13g2_inv_1 _5823_ (.Y(_2233_),
    .A(_2232_));
 sg13g2_and2_1 _5824_ (.A(net1069),
    .B(net959),
    .X(_2234_));
 sg13g2_nand2_1 _5825_ (.Y(_2235_),
    .A(net1069),
    .B(net959));
 sg13g2_nand2b_1 _5826_ (.Y(_2236_),
    .B(_1583_),
    .A_N(net959));
 sg13g2_xnor2_1 _5827_ (.Y(_2237_),
    .A(_1583_),
    .B(net959));
 sg13g2_xnor2_1 _5828_ (.Y(_2238_),
    .A(net1069),
    .B(net959));
 sg13g2_o21ai_1 _5829_ (.B1(net1003),
    .Y(_2239_),
    .A1(_1579_),
    .A2(_2238_));
 sg13g2_nor2_1 _5830_ (.A(_2230_),
    .B(_2239_),
    .Y(_2240_));
 sg13g2_o21ai_1 _5831_ (.B1(_2233_),
    .Y(_2241_),
    .A1(_2230_),
    .A2(_2239_));
 sg13g2_nor2_1 _5832_ (.A(net1056),
    .B(_2235_),
    .Y(_2242_));
 sg13g2_nor2_1 _5833_ (.A(net990),
    .B(net1002),
    .Y(_2243_));
 sg13g2_nand3_1 _5834_ (.B(net1055),
    .C(_2234_),
    .A(net1005),
    .Y(_2244_));
 sg13g2_mux2_1 _5835_ (.A0(_2241_),
    .A1(_2244_),
    .S(net985),
    .X(_2245_));
 sg13g2_nor2_2 _5836_ (.A(net1004),
    .B(_2230_),
    .Y(_2246_));
 sg13g2_o21ai_1 _5837_ (.B1(_2246_),
    .Y(_2247_),
    .A1(net1055),
    .A2(_2237_));
 sg13g2_nand2_2 _5838_ (.Y(_2248_),
    .A(net1004),
    .B(net1057));
 sg13g2_and2_1 _5839_ (.A(_2247_),
    .B(_2248_),
    .X(_2249_));
 sg13g2_nor2_1 _5840_ (.A(_1578_),
    .B(net1069),
    .Y(_2250_));
 sg13g2_nand2_1 _5841_ (.Y(_2251_),
    .A(net1055),
    .B(_1583_));
 sg13g2_a21oi_1 _5842_ (.A1(net1056),
    .A2(_2235_),
    .Y(_2252_),
    .B1(_2230_));
 sg13g2_nand2_1 _5843_ (.Y(_2253_),
    .A(net1003),
    .B(_2252_));
 sg13g2_a21o_2 _5844_ (.A2(_2234_),
    .A1(net1005),
    .B1(_2232_),
    .X(_2254_));
 sg13g2_nor2_1 _5845_ (.A(net989),
    .B(_2254_),
    .Y(_2255_));
 sg13g2_a221oi_1 _5846_ (.B2(_2255_),
    .C1(net1172),
    .B1(_2253_),
    .A1(net990),
    .Y(_2256_),
    .A2(_2249_));
 sg13g2_nor2_1 _5847_ (.A(net1163),
    .B(net987),
    .Y(_2257_));
 sg13g2_a21oi_1 _5848_ (.A1(net1172),
    .A2(_2245_),
    .Y(_2258_),
    .B1(_2256_));
 sg13g2_nand2_1 _5849_ (.Y(_2259_),
    .A(net1168),
    .B(_2258_));
 sg13g2_nand2_2 _5850_ (.Y(_2260_),
    .A(net1055),
    .B(_2238_));
 sg13g2_o21ai_1 _5851_ (.B1(net1004),
    .Y(_2261_),
    .A1(net960),
    .A2(_2251_));
 sg13g2_nand2_1 _5852_ (.Y(_2262_),
    .A(net1005),
    .B(_2260_));
 sg13g2_nor2_2 _5853_ (.A(net1056),
    .B(net959),
    .Y(_2263_));
 sg13g2_o21ai_1 _5854_ (.B1(net1003),
    .Y(_2264_),
    .A1(_2237_),
    .A2(_2263_));
 sg13g2_inv_1 _5855_ (.Y(_2265_),
    .A(_2264_));
 sg13g2_nor2_1 _5856_ (.A(net989),
    .B(_2265_),
    .Y(_2266_));
 sg13g2_nor2_1 _5857_ (.A(net985),
    .B(_2254_),
    .Y(_2267_));
 sg13g2_a22oi_1 _5858_ (.Y(_2268_),
    .B1(_2267_),
    .B2(_2239_),
    .A2(_2266_),
    .A1(_2262_));
 sg13g2_a21oi_2 _5859_ (.B1(net987),
    .Y(_2269_),
    .A2(_2260_),
    .A1(net1005));
 sg13g2_nand2_2 _5860_ (.Y(_2270_),
    .A(net1056),
    .B(net960));
 sg13g2_nand2_1 _5861_ (.Y(_2271_),
    .A(net1056),
    .B(_1583_));
 sg13g2_nand3_1 _5862_ (.B(_2270_),
    .C(_2271_),
    .A(_2246_),
    .Y(_2272_));
 sg13g2_and2_1 _5863_ (.A(_2229_),
    .B(_2236_),
    .X(_2273_));
 sg13g2_nor2_1 _5864_ (.A(net1006),
    .B(_2273_),
    .Y(_2274_));
 sg13g2_nand2_1 _5865_ (.Y(_2275_),
    .A(_1583_),
    .B(net959));
 sg13g2_nand2_1 _5866_ (.Y(_2276_),
    .A(net1069),
    .B(_2263_));
 sg13g2_nand3_1 _5867_ (.B(_2275_),
    .C(_2276_),
    .A(net1004),
    .Y(_2277_));
 sg13g2_nor2_1 _5868_ (.A(net990),
    .B(_2274_),
    .Y(_2278_));
 sg13g2_a221oi_1 _5869_ (.B2(_2278_),
    .C1(net1170),
    .B1(_2277_),
    .A1(_2269_),
    .Y(_2279_),
    .A2(_2272_));
 sg13g2_a21oi_1 _5870_ (.A1(net1172),
    .A2(_2268_),
    .Y(_2280_),
    .B1(_2279_));
 sg13g2_a21oi_1 _5871_ (.A1(net1163),
    .A2(_2280_),
    .Y(_2281_),
    .B1(net1167));
 sg13g2_nor2_1 _5872_ (.A(net990),
    .B(_2241_),
    .Y(_2282_));
 sg13g2_nand3_1 _5873_ (.B(net1057),
    .C(_2238_),
    .A(net1002),
    .Y(_2283_));
 sg13g2_nand3_1 _5874_ (.B(net1055),
    .C(_2235_),
    .A(net1002),
    .Y(_2284_));
 sg13g2_nand2_1 _5875_ (.Y(_2285_),
    .A(net989),
    .B(_2284_));
 sg13g2_nand3b_1 _5876_ (.B(_2283_),
    .C(_2284_),
    .Y(_2286_),
    .A_N(_2254_));
 sg13g2_o21ai_1 _5877_ (.B1(net1168),
    .Y(_2287_),
    .A1(net985),
    .A2(_2286_));
 sg13g2_nand3_1 _5878_ (.B(_2231_),
    .C(_2239_),
    .A(net985),
    .Y(_2288_));
 sg13g2_o21ai_1 _5879_ (.B1(net1002),
    .Y(_2289_),
    .A1(_2238_),
    .A2(_2250_));
 sg13g2_a21oi_1 _5880_ (.A1(_2267_),
    .A2(_2289_),
    .Y(_2290_),
    .B1(net1168));
 sg13g2_nor2_1 _5881_ (.A(net1163),
    .B(net989),
    .Y(_2291_));
 sg13g2_o21ai_1 _5882_ (.B1(net1173),
    .Y(_2292_),
    .A1(_2282_),
    .A2(_2287_));
 sg13g2_a21oi_1 _5883_ (.A1(_2288_),
    .A2(_2290_),
    .Y(_2293_),
    .B1(_2292_));
 sg13g2_and2_1 _5884_ (.A(net985),
    .B(_2248_),
    .X(_2294_));
 sg13g2_a221oi_1 _5885_ (.B2(_2247_),
    .C1(net1163),
    .B1(_2269_),
    .A1(net985),
    .Y(_2295_),
    .A2(_2249_));
 sg13g2_nor2_2 _5886_ (.A(net1168),
    .B(net986),
    .Y(_2296_));
 sg13g2_nand2_1 _5887_ (.Y(_2297_),
    .A(_2261_),
    .B(_2264_));
 sg13g2_nand2_1 _5888_ (.Y(_2298_),
    .A(net1163),
    .B(net987));
 sg13g2_inv_1 _5889_ (.Y(_2299_),
    .A(_2298_));
 sg13g2_o21ai_1 _5890_ (.B1(net1004),
    .Y(_2300_),
    .A1(net1057),
    .A2(_2234_));
 sg13g2_nand2_1 _5891_ (.Y(_2301_),
    .A(_2284_),
    .B(_2300_));
 sg13g2_a22oi_1 _5892_ (.Y(_2302_),
    .B1(_2299_),
    .B2(_2301_),
    .A2(_2297_),
    .A1(_2296_));
 sg13g2_nand2_1 _5893_ (.Y(_2303_),
    .A(_2667_),
    .B(_2302_));
 sg13g2_o21ai_1 _5894_ (.B1(net1167),
    .Y(_2304_),
    .A1(_2295_),
    .A2(_2303_));
 sg13g2_nor2_1 _5895_ (.A(_2293_),
    .B(_2304_),
    .Y(_2305_));
 sg13g2_a21oi_1 _5896_ (.A1(_2259_),
    .A2(_2281_),
    .Y(_2306_),
    .B1(_2305_));
 sg13g2_and2_1 _5897_ (.A(net989),
    .B(_2231_),
    .X(_2307_));
 sg13g2_o21ai_1 _5898_ (.B1(_2307_),
    .Y(_2308_),
    .A1(_2230_),
    .A2(_2239_));
 sg13g2_nand2_1 _5899_ (.Y(_2309_),
    .A(net1004),
    .B(_2271_));
 sg13g2_nand2b_1 _5900_ (.Y(_2310_),
    .B(_2260_),
    .A_N(_2309_));
 sg13g2_nand2b_1 _5901_ (.Y(_2311_),
    .B(_2275_),
    .A_N(_2263_));
 sg13g2_a21oi_1 _5902_ (.A1(net1003),
    .A2(_2311_),
    .Y(_2312_),
    .B1(net990));
 sg13g2_a21oi_1 _5903_ (.A1(_2310_),
    .A2(_2312_),
    .Y(_2313_),
    .B1(_2667_));
 sg13g2_and2_1 _5904_ (.A(net987),
    .B(_2309_),
    .X(_2314_));
 sg13g2_nand3_1 _5905_ (.B(_2247_),
    .C(_2277_),
    .A(net990),
    .Y(_2315_));
 sg13g2_a21oi_1 _5906_ (.A1(_2289_),
    .A2(_2314_),
    .Y(_2316_),
    .B1(net1171));
 sg13g2_a22oi_1 _5907_ (.Y(_2317_),
    .B1(_2315_),
    .B2(_2316_),
    .A2(_2313_),
    .A1(_2308_));
 sg13g2_nand2_1 _5908_ (.Y(_2318_),
    .A(_2289_),
    .B(_2300_));
 sg13g2_nand3_1 _5909_ (.B(_2289_),
    .C(_2300_),
    .A(net987),
    .Y(_2319_));
 sg13g2_nand4_1 _5910_ (.B(_2283_),
    .C(_2284_),
    .A(net989),
    .Y(_2320_),
    .D(_2309_));
 sg13g2_and2_1 _5911_ (.A(_0930_),
    .B(_2320_),
    .X(_2321_));
 sg13g2_nand2_1 _5912_ (.Y(_2322_),
    .A(net1004),
    .B(_2273_));
 sg13g2_a21oi_2 _5913_ (.B1(net1004),
    .Y(_2323_),
    .A2(net1069),
    .A1(net1056));
 sg13g2_nor2_1 _5914_ (.A(net987),
    .B(_2323_),
    .Y(_2324_));
 sg13g2_a221oi_1 _5915_ (.B2(_2310_),
    .C1(_1428_),
    .B1(_2324_),
    .A1(_2266_),
    .Y(_2325_),
    .A2(_2322_));
 sg13g2_a21oi_1 _5916_ (.A1(_2319_),
    .A2(_2321_),
    .Y(_2326_),
    .B1(_2325_));
 sg13g2_o21ai_1 _5917_ (.B1(_2326_),
    .Y(_2327_),
    .A1(net1163),
    .A2(_2317_));
 sg13g2_nand3_1 _5918_ (.B(_2247_),
    .C(_2322_),
    .A(net1171),
    .Y(_2328_));
 sg13g2_o21ai_1 _5919_ (.B1(_2328_),
    .Y(_2329_),
    .A1(net1170),
    .A2(_2318_));
 sg13g2_nand3b_1 _5920_ (.B(net1002),
    .C(_2667_),
    .Y(_2330_),
    .A_N(_2252_));
 sg13g2_o21ai_1 _5921_ (.B1(_2236_),
    .Y(_2331_),
    .A1(net1006),
    .A2(net1056));
 sg13g2_nand4_1 _5922_ (.B(_2248_),
    .C(_2284_),
    .A(net1170),
    .Y(_2332_),
    .D(_2331_));
 sg13g2_a21oi_1 _5923_ (.A1(_2330_),
    .A2(_2332_),
    .Y(_2333_),
    .B1(_2257_));
 sg13g2_nand4_1 _5924_ (.B(net1002),
    .C(net1069),
    .A(_2667_),
    .Y(_2334_),
    .D(_2263_));
 sg13g2_nand2_1 _5925_ (.Y(_2335_),
    .A(_2270_),
    .B(_2323_));
 sg13g2_nand4_1 _5926_ (.B(_2251_),
    .C(_2270_),
    .A(net1170),
    .Y(_2336_),
    .D(_2323_));
 sg13g2_a21oi_1 _5927_ (.A1(_2334_),
    .A2(_2336_),
    .Y(_2337_),
    .B1(_2298_));
 sg13g2_a221oi_1 _5928_ (.B2(_2298_),
    .C1(_2337_),
    .B1(_2333_),
    .A1(_2257_),
    .Y(_2338_),
    .A2(_2329_));
 sg13g2_nand2_1 _5929_ (.Y(_2339_),
    .A(_2665_),
    .B(_2338_));
 sg13g2_a21oi_1 _5930_ (.A1(net1167),
    .A2(_2327_),
    .Y(_2340_),
    .B1(net1166));
 sg13g2_a221oi_1 _5931_ (.B2(_2340_),
    .C1(\dtop.vtop.logo.addr[9] ),
    .B1(_2339_),
    .A1(net1166),
    .Y(_2341_),
    .A2(_2306_));
 sg13g2_o21ai_1 _5932_ (.B1(_2299_),
    .Y(_2342_),
    .A1(_2240_),
    .A2(_2254_));
 sg13g2_nor3_1 _5933_ (.A(net1005),
    .B(_2237_),
    .C(_2263_),
    .Y(_2343_));
 sg13g2_o21ai_1 _5934_ (.B1(_2291_),
    .Y(_2344_),
    .A1(_2254_),
    .A2(_2343_));
 sg13g2_nor2_1 _5935_ (.A(_2231_),
    .B(_2263_),
    .Y(_2345_));
 sg13g2_o21ai_1 _5936_ (.B1(net989),
    .Y(_2346_),
    .A1(_2265_),
    .A2(_2345_));
 sg13g2_nand3b_1 _5937_ (.B(_2296_),
    .C(net1005),
    .Y(_2347_),
    .A_N(_2263_));
 sg13g2_and4_1 _5938_ (.A(net1172),
    .B(_2344_),
    .C(_2346_),
    .D(_2347_),
    .X(_2348_));
 sg13g2_nand2_1 _5939_ (.Y(_2349_),
    .A(_2247_),
    .B(_2261_));
 sg13g2_o21ai_1 _5940_ (.B1(_2289_),
    .Y(_2350_),
    .A1(net1003),
    .A2(_2242_));
 sg13g2_a22oi_1 _5941_ (.Y(_2351_),
    .B1(_2350_),
    .B2(_2296_),
    .A2(_2349_),
    .A1(_2299_));
 sg13g2_a22oi_1 _5942_ (.Y(_2352_),
    .B1(_2307_),
    .B2(_2289_),
    .A2(_2294_),
    .A1(_2238_));
 sg13g2_a21oi_1 _5943_ (.A1(net1168),
    .A2(_2352_),
    .Y(_2353_),
    .B1(net1172));
 sg13g2_a221oi_1 _5944_ (.B2(_2353_),
    .C1(_2665_),
    .B1(_2351_),
    .A1(_2342_),
    .Y(_2354_),
    .A2(_2348_));
 sg13g2_o21ai_1 _5945_ (.B1(net1172),
    .Y(_2355_),
    .A1(_2285_),
    .A2(_2345_));
 sg13g2_or2_1 _5946_ (.X(_2356_),
    .B(_2355_),
    .A(_2282_));
 sg13g2_a221oi_1 _5947_ (.B2(_2239_),
    .C1(net1172),
    .B1(_2307_),
    .A1(_2247_),
    .Y(_2357_),
    .A2(_2294_));
 sg13g2_nor2_1 _5948_ (.A(net1163),
    .B(_2357_),
    .Y(_2358_));
 sg13g2_nand2_1 _5949_ (.Y(_2359_),
    .A(_2276_),
    .B(_2323_));
 sg13g2_nand2_1 _5950_ (.Y(_2360_),
    .A(_2269_),
    .B(_2359_));
 sg13g2_o21ai_1 _5951_ (.B1(_2360_),
    .Y(_2361_),
    .A1(net989),
    .A2(_2297_));
 sg13g2_a22oi_1 _5952_ (.Y(_2362_),
    .B1(_2264_),
    .B2(_2267_),
    .A2(_2255_),
    .A1(_2239_));
 sg13g2_o21ai_1 _5953_ (.B1(_2665_),
    .Y(_2363_),
    .A1(_1428_),
    .A2(_2362_));
 sg13g2_a221oi_1 _5954_ (.B2(_0930_),
    .C1(_2363_),
    .B1(_2361_),
    .A1(_2356_),
    .Y(_2364_),
    .A2(_2358_));
 sg13g2_nor3_1 _5955_ (.A(net1166),
    .B(_2354_),
    .C(_2364_),
    .Y(_2365_));
 sg13g2_nand3_1 _5956_ (.B(_2239_),
    .C(_2260_),
    .A(net986),
    .Y(_2366_));
 sg13g2_a21oi_1 _5957_ (.A1(_2233_),
    .A2(_2289_),
    .Y(_2367_),
    .B1(net986));
 sg13g2_nor2b_1 _5958_ (.A(_2367_),
    .B_N(_0930_),
    .Y(_2368_));
 sg13g2_a221oi_1 _5959_ (.B2(_2262_),
    .C1(net1170),
    .B1(_2312_),
    .A1(_2253_),
    .Y(_2369_),
    .A2(_2307_));
 sg13g2_o21ai_1 _5960_ (.B1(net1172),
    .Y(_2370_),
    .A1(net985),
    .A2(_2244_));
 sg13g2_a21oi_1 _5961_ (.A1(_2255_),
    .A2(_2335_),
    .Y(_2371_),
    .B1(_2370_));
 sg13g2_or3_1 _5962_ (.A(net1163),
    .B(_2369_),
    .C(_2371_),
    .X(_2372_));
 sg13g2_nand3_1 _5963_ (.B(_2248_),
    .C(_2270_),
    .A(_2237_),
    .Y(_2373_));
 sg13g2_a21oi_1 _5964_ (.A1(net985),
    .A2(_2373_),
    .Y(_2374_),
    .B1(_1428_));
 sg13g2_a221oi_1 _5965_ (.B2(_2346_),
    .C1(net1167),
    .B1(_2374_),
    .A1(_2366_),
    .Y(_2375_),
    .A2(_2368_));
 sg13g2_a21oi_1 _5966_ (.A1(net1002),
    .A2(_2250_),
    .Y(_2376_),
    .B1(net988));
 sg13g2_a221oi_1 _5967_ (.B2(_2376_),
    .C1(net1170),
    .B1(_2300_),
    .A1(_2230_),
    .Y(_2377_),
    .A2(_2243_));
 sg13g2_nor2_1 _5968_ (.A(net988),
    .B(_2246_),
    .Y(_2378_));
 sg13g2_o21ai_1 _5969_ (.B1(_2378_),
    .Y(_2379_),
    .A1(net1002),
    .A2(_2242_));
 sg13g2_nand3_1 _5970_ (.B(_2236_),
    .C(_2243_),
    .A(net1055),
    .Y(_2380_));
 sg13g2_nand3_1 _5971_ (.B(_2379_),
    .C(_2380_),
    .A(net1170),
    .Y(_2381_));
 sg13g2_nand2b_1 _5972_ (.Y(_2382_),
    .B(_2381_),
    .A_N(_2377_));
 sg13g2_a221oi_1 _5973_ (.B2(net1167),
    .C1(_2664_),
    .B1(_2382_),
    .A1(_2372_),
    .Y(_2383_),
    .A2(_2375_));
 sg13g2_nor3_2 _5974_ (.A(_2663_),
    .B(_2365_),
    .C(_2383_),
    .Y(_2384_));
 sg13g2_or4_2 _5975_ (.A(_1587_),
    .B(_2193_),
    .C(_2341_),
    .D(_2384_),
    .X(_2385_));
 sg13g2_nand2_1 _5976_ (.Y(_2386_),
    .A(net1225),
    .B(\dtop.vtop.color[4] ));
 sg13g2_nor2_1 _5977_ (.A(_0005_),
    .B(_2386_),
    .Y(_2387_));
 sg13g2_xor2_1 _5978_ (.B(net1219),
    .A(\dtop.oct_counter[3] ),
    .X(_2388_));
 sg13g2_nor2_1 _5979_ (.A(_2387_),
    .B(_2388_),
    .Y(_2389_));
 sg13g2_a21oi_2 _5980_ (.B1(_2389_),
    .Y(_2390_),
    .A2(_2386_),
    .A1(_0005_));
 sg13g2_nand3_1 _5981_ (.B(\dtop.vtop.color[6] ),
    .C(_2390_),
    .A(\dtop.vtop.color[7] ),
    .Y(_2391_));
 sg13g2_o21ai_1 _5982_ (.B1(_2385_),
    .Y(_2392_),
    .A1(_2881_),
    .A2(_2391_));
 sg13g2_nand2b_1 _5983_ (.Y(_2393_),
    .B(\dtop.player_inst.program_addr[6] ),
    .A_N(\dtop.out_sample[6] ));
 sg13g2_nand2b_1 _5984_ (.Y(_2394_),
    .B(net1215),
    .A_N(\dtop.out_sample[2] ));
 sg13g2_a22oi_1 _5985_ (.Y(_2395_),
    .B1(_2669_),
    .B2(\dtop.out_sample[1] ),
    .A2(_2668_),
    .A1(\dtop.out_sample[0] ));
 sg13g2_o21ai_1 _5986_ (.B1(_2394_),
    .Y(_2396_),
    .A1(\dtop.out_sample[1] ),
    .A2(_2669_));
 sg13g2_nor2_1 _5987_ (.A(_2395_),
    .B(_2396_),
    .Y(_2397_));
 sg13g2_a221oi_1 _5988_ (.B2(\dtop.out_sample[2] ),
    .C1(_2397_),
    .B1(net1162),
    .A1(\dtop.out_sample[3] ),
    .Y(_2398_),
    .A2(_2670_));
 sg13g2_nand2b_1 _5989_ (.Y(_2399_),
    .B(net1207),
    .A_N(\dtop.out_sample[4] ));
 sg13g2_o21ai_1 _5990_ (.B1(_2399_),
    .Y(_2400_),
    .A1(\dtop.out_sample[3] ),
    .A2(_2670_));
 sg13g2_nor2_1 _5991_ (.A(_2398_),
    .B(_2400_),
    .Y(_2401_));
 sg13g2_a221oi_1 _5992_ (.B2(\dtop.out_sample[4] ),
    .C1(_2401_),
    .B1(_2656_),
    .A1(\dtop.out_sample[5] ),
    .Y(_2402_),
    .A2(_2655_));
 sg13g2_o21ai_1 _5993_ (.B1(_2393_),
    .Y(_2403_),
    .A1(\dtop.out_sample[5] ),
    .A2(_2655_));
 sg13g2_nor2_1 _5994_ (.A(_2402_),
    .B(_2403_),
    .Y(_2404_));
 sg13g2_a21oi_1 _5995_ (.A1(\dtop.out_sample[6] ),
    .A2(_2654_),
    .Y(_2405_),
    .B1(_2404_));
 sg13g2_xor2_1 _5996_ (.B(_2405_),
    .A(net1182),
    .X(_2406_));
 sg13g2_and2_1 _5997_ (.A(net1120),
    .B(_2406_),
    .X(_2407_));
 sg13g2_a21o_1 _5998_ (.A2(_2390_),
    .A1(\dtop.vtop.color[6] ),
    .B1(\dtop.vtop.color[7] ),
    .X(_2408_));
 sg13g2_and2_1 _5999_ (.A(_2391_),
    .B(_2408_),
    .X(_2409_));
 sg13g2_a221oi_1 _6000_ (.B2(_2882_),
    .C1(_2392_),
    .B1(_2409_),
    .A1(_0049_),
    .Y(_2410_),
    .A2(_2407_));
 sg13g2_nor2b_1 _6001_ (.A(_2190_),
    .B_N(_0556_),
    .Y(_2411_));
 sg13g2_nand2_1 _6002_ (.Y(_2412_),
    .A(_0070_),
    .B(net1076));
 sg13g2_a21oi_1 _6003_ (.A1(_0072_),
    .A2(net1077),
    .Y(_2413_),
    .B1(\dtop.vtop.pipeline.neg_t[7] ));
 sg13g2_o21ai_1 _6004_ (.B1(\dtop.vtop.pipeline.neg_t[9] ),
    .Y(_2414_),
    .A1(_0071_),
    .A2(_2412_));
 sg13g2_a21oi_1 _6005_ (.A1(_0071_),
    .A2(_2412_),
    .Y(_2415_),
    .B1(_2413_));
 sg13g2_nand2b_1 _6006_ (.Y(_2416_),
    .B(_2415_),
    .A_N(_2414_));
 sg13g2_nand3_1 _6007_ (.B(_0079_),
    .C(net1077),
    .A(\dtop.vtop.pipeline.neg_t[3] ),
    .Y(_2417_));
 sg13g2_nand2_1 _6008_ (.Y(_2418_),
    .A(_0078_),
    .B(net1076));
 sg13g2_o21ai_1 _6009_ (.B1(_2417_),
    .Y(_2419_),
    .A1(_0077_),
    .A2(_2418_));
 sg13g2_a21oi_1 _6010_ (.A1(_0079_),
    .A2(net1077),
    .Y(_2420_),
    .B1(\dtop.vtop.pipeline.neg_t[3] ));
 sg13g2_nand2_1 _6011_ (.Y(_2421_),
    .A(_0051_),
    .B(net1077));
 sg13g2_nand3_1 _6012_ (.B(_0051_),
    .C(net1077),
    .A(\dtop.vtop.pipeline.neg_t[1] ),
    .Y(_2422_));
 sg13g2_nand2_1 _6013_ (.Y(_2423_),
    .A(_0083_),
    .B(net1077));
 sg13g2_a21oi_1 _6014_ (.A1(_0083_),
    .A2(net1077),
    .Y(_2424_),
    .B1(\dtop.vtop.pipeline.neg_t[0] ));
 sg13g2_xnor2_1 _6015_ (.Y(_2425_),
    .A(_0082_),
    .B(_2421_));
 sg13g2_o21ai_1 _6016_ (.B1(_2422_),
    .Y(_2426_),
    .A1(_2424_),
    .A2(_2425_));
 sg13g2_and2_1 _6017_ (.A(_0080_),
    .B(net1076),
    .X(_2427_));
 sg13g2_xnor2_1 _6018_ (.Y(_2428_),
    .A(_0081_),
    .B(_2427_));
 sg13g2_a22oi_1 _6019_ (.Y(_2429_),
    .B1(_2428_),
    .B2(_2426_),
    .A2(_2427_),
    .A1(\dtop.vtop.pipeline.neg_t[2] ));
 sg13g2_nor2_1 _6020_ (.A(_2420_),
    .B(_2429_),
    .Y(_2430_));
 sg13g2_nor2_1 _6021_ (.A(_2419_),
    .B(_2430_),
    .Y(_2431_));
 sg13g2_nand2_1 _6022_ (.Y(_2432_),
    .A(_0073_),
    .B(net1076));
 sg13g2_xor2_1 _6023_ (.B(_2432_),
    .A(_0074_),
    .X(_2433_));
 sg13g2_nand2_1 _6024_ (.Y(_2434_),
    .A(_0075_),
    .B(net1076));
 sg13g2_xnor2_1 _6025_ (.Y(_2435_),
    .A(_0076_),
    .B(_2434_));
 sg13g2_a21o_1 _6026_ (.A2(_2418_),
    .A1(_0077_),
    .B1(_2435_),
    .X(_2436_));
 sg13g2_nand3_1 _6027_ (.B(_0072_),
    .C(net1076),
    .A(\dtop.vtop.pipeline.neg_t[7] ),
    .Y(_2437_));
 sg13g2_o21ai_1 _6028_ (.B1(_2437_),
    .Y(_2438_),
    .A1(_2652_),
    .A2(_2432_));
 sg13g2_nand3_1 _6029_ (.B(_0075_),
    .C(net1076),
    .A(\dtop.vtop.pipeline.neg_t[5] ),
    .Y(_2439_));
 sg13g2_o21ai_1 _6030_ (.B1(_2439_),
    .Y(_2440_),
    .A1(_2431_),
    .A2(_2436_));
 sg13g2_a21oi_1 _6031_ (.A1(_2433_),
    .A2(_2440_),
    .Y(_2441_),
    .B1(_2438_));
 sg13g2_nand4_1 _6032_ (.B(\dtop.vtop.pipeline.neg_t[8] ),
    .C(_0070_),
    .A(\dtop.vtop.pipeline.neg_t[9] ),
    .Y(_2442_),
    .D(net1076));
 sg13g2_o21ai_1 _6033_ (.B1(_2442_),
    .Y(_2443_),
    .A1(_2416_),
    .A2(_2441_));
 sg13g2_nand2b_1 _6034_ (.Y(_2444_),
    .B(_2437_),
    .A_N(_2420_));
 sg13g2_xnor2_1 _6035_ (.Y(_2445_),
    .A(_0059_),
    .B(_2423_));
 sg13g2_nor2_1 _6036_ (.A(_2419_),
    .B(_2425_),
    .Y(_2446_));
 sg13g2_nor4_1 _6037_ (.A(_2416_),
    .B(_2436_),
    .C(_2444_),
    .D(_2445_),
    .Y(_2447_));
 sg13g2_nand4_1 _6038_ (.B(_2433_),
    .C(_2446_),
    .A(_2428_),
    .Y(_2448_),
    .D(_2447_));
 sg13g2_nand2_1 _6039_ (.Y(_2449_),
    .A(_2443_),
    .B(_2448_));
 sg13g2_xnor2_1 _6040_ (.Y(_2450_),
    .A(_2909_),
    .B(_2449_));
 sg13g2_nor2_1 _6041_ (.A(_0062_),
    .B(_2450_),
    .Y(_2451_));
 sg13g2_o21ai_1 _6042_ (.B1(_2451_),
    .Y(_2452_),
    .A1(_1601_),
    .A2(_1612_));
 sg13g2_nand3_1 _6043_ (.B(_1568_),
    .C(_2452_),
    .A(_0983_),
    .Y(_2453_));
 sg13g2_and2_1 _6044_ (.A(_0557_),
    .B(_2453_),
    .X(_2454_));
 sg13g2_nand2_1 _6045_ (.Y(_2455_),
    .A(_0983_),
    .B(_1569_));
 sg13g2_a21oi_1 _6046_ (.A1(_2454_),
    .A2(_2455_),
    .Y(_2456_),
    .B1(_2881_));
 sg13g2_nor3_1 _6047_ (.A(\dtop.vtop.rs.x_scan.phase[1] ),
    .B(\dtop.vtop.rs.x_scan.phase[0] ),
    .C(_1425_),
    .Y(_2457_));
 sg13g2_nand2_1 _6048_ (.Y(_2458_),
    .A(net1191),
    .B(_2457_));
 sg13g2_a21oi_2 _6049_ (.B1(_2458_),
    .Y(_2459_),
    .A2(_2456_),
    .A1(_2385_));
 sg13g2_inv_1 _6050_ (.Y(_2460_),
    .A(_2459_));
 sg13g2_o21ai_1 _6051_ (.B1(_2185_),
    .Y(_0279_),
    .A1(_2410_),
    .A2(_2460_));
 sg13g2_nand2b_1 _6052_ (.Y(_2461_),
    .B(net461),
    .A_N(net1191));
 sg13g2_nand2b_1 _6053_ (.Y(_2462_),
    .B(net1225),
    .A_N(\dtop.vtop.pipeline.zg[6] ));
 sg13g2_nand2_1 _6054_ (.Y(_2463_),
    .A(\dtop.vtop.pipeline.zg[7] ),
    .B(_2462_));
 sg13g2_nor2_1 _6055_ (.A(\dtop.vtop.pipeline.zg[7] ),
    .B(_2462_),
    .Y(_2464_));
 sg13g2_a21oi_1 _6056_ (.A1(_2388_),
    .A2(_2463_),
    .Y(_2465_),
    .B1(_2464_));
 sg13g2_nand2b_1 _6057_ (.Y(_2466_),
    .B(_2676_),
    .A_N(_2465_));
 sg13g2_nand2b_1 _6058_ (.Y(_2467_),
    .B(_2675_),
    .A_N(_2466_));
 sg13g2_o21ai_1 _6059_ (.B1(_2385_),
    .Y(_2468_),
    .A1(net1120),
    .A2(_2467_));
 sg13g2_xnor2_1 _6060_ (.Y(_2469_),
    .A(_2675_),
    .B(_2466_));
 sg13g2_a221oi_1 _6061_ (.B2(_2882_),
    .C1(_2468_),
    .B1(_2469_),
    .A1(net1178),
    .Y(_2470_),
    .A2(_2407_));
 sg13g2_o21ai_1 _6062_ (.B1(_2461_),
    .Y(_0280_),
    .A1(_2460_),
    .A2(_2470_));
 sg13g2_nand2_1 _6063_ (.Y(_2471_),
    .A(_0055_),
    .B(_2407_));
 sg13g2_xor2_1 _6064_ (.B(_2390_),
    .A(_0006_),
    .X(_2472_));
 sg13g2_o21ai_1 _6065_ (.B1(_2471_),
    .Y(_2473_),
    .A1(net1120),
    .A2(_2472_));
 sg13g2_o21ai_1 _6066_ (.B1(_2459_),
    .Y(_2474_),
    .A1(_2392_),
    .A2(_2473_));
 sg13g2_o21ai_1 _6067_ (.B1(_2474_),
    .Y(_0281_),
    .A1(net1190),
    .A2(_2700_));
 sg13g2_xnor2_1 _6068_ (.Y(_2475_),
    .A(\dtop.vtop.pipeline.zg[8] ),
    .B(_2465_));
 sg13g2_o21ai_1 _6069_ (.B1(_2471_),
    .Y(_2476_),
    .A1(net1120),
    .A2(_2475_));
 sg13g2_o21ai_1 _6070_ (.B1(_2459_),
    .Y(_2477_),
    .A1(_2468_),
    .A2(_2476_));
 sg13g2_o21ai_1 _6071_ (.B1(_2477_),
    .Y(_0282_),
    .A1(net1190),
    .A2(_2701_));
 sg13g2_o21ai_1 _6072_ (.B1(net1250),
    .Y(_2478_),
    .A1(net1182),
    .A2(_0922_));
 sg13g2_a21oi_1 _6073_ (.A1(net1183),
    .A2(_0922_),
    .Y(_0283_),
    .B1(_2478_));
 sg13g2_o21ai_1 _6074_ (.B1(net1251),
    .Y(_2479_),
    .A1(net1180),
    .A2(_0923_));
 sg13g2_a21oi_1 _6075_ (.A1(net1180),
    .A2(_0923_),
    .Y(_0284_),
    .B1(net618));
 sg13g2_o21ai_1 _6076_ (.B1(net1250),
    .Y(_2480_),
    .A1(net1179),
    .A2(net605));
 sg13g2_a21oi_1 _6077_ (.A1(net1179),
    .A2(net605),
    .Y(_0285_),
    .B1(_2480_));
 sg13g2_nor2b_1 _6078_ (.A(net1190),
    .B_N(net609),
    .Y(_2481_));
 sg13g2_nand4_1 _6079_ (.B(_2676_),
    .C(\dtop.vtop.color[7] ),
    .A(_2675_),
    .Y(_2482_),
    .D(_2882_));
 sg13g2_o21ai_1 _6080_ (.B1(\dtop.vtop.color[7] ),
    .Y(_2483_),
    .A1(\dtop.vtop.pipeline.zg[9] ),
    .A2(\dtop.vtop.pipeline.zg[8] ));
 sg13g2_nor3_1 _6081_ (.A(\dtop.vtop.pipeline.zg[9] ),
    .B(\dtop.vtop.pipeline.zg[8] ),
    .C(\dtop.vtop.color[7] ),
    .Y(_2484_));
 sg13g2_or2_1 _6082_ (.X(_2485_),
    .B(\dtop.vtop.pipeline.zg[7] ),
    .A(\dtop.vtop.pipeline.zg[9] ));
 sg13g2_nor2_1 _6083_ (.A(\dtop.vtop.color[6] ),
    .B(_2485_),
    .Y(_2486_));
 sg13g2_nor2_1 _6084_ (.A(\dtop.vtop.pipeline.zg[9] ),
    .B(\dtop.vtop.pipeline.zg[6] ),
    .Y(_2487_));
 sg13g2_o21ai_1 _6085_ (.B1(\dtop.vtop.color[4] ),
    .Y(_2488_),
    .A1(\dtop.vtop.pipeline.zg[9] ),
    .A2(\dtop.vtop.pipeline.zg[5] ));
 sg13g2_o21ai_1 _6086_ (.B1(_2488_),
    .Y(_2489_),
    .A1(_0005_),
    .A2(_2487_));
 sg13g2_a21oi_1 _6087_ (.A1(_0005_),
    .A2(_2487_),
    .Y(_2490_),
    .B1(_2486_));
 sg13g2_a22oi_1 _6088_ (.Y(_2491_),
    .B1(_2489_),
    .B2(_2490_),
    .A2(_2485_),
    .A1(\dtop.vtop.color[6] ));
 sg13g2_o21ai_1 _6089_ (.B1(_2483_),
    .Y(_2492_),
    .A1(_2484_),
    .A2(_2491_));
 sg13g2_nand3_1 _6090_ (.B(_2675_),
    .C(_2677_),
    .A(net1225),
    .Y(_2493_));
 sg13g2_nand2b_1 _6091_ (.Y(_2494_),
    .B(_2493_),
    .A_N(_2487_));
 sg13g2_nor2_1 _6092_ (.A(\dtop.vtop.pipeline.zg[6] ),
    .B(_2493_),
    .Y(_2495_));
 sg13g2_a21oi_1 _6093_ (.A1(_2388_),
    .A2(_2494_),
    .Y(_2496_),
    .B1(_2495_));
 sg13g2_nand2_1 _6094_ (.Y(_2497_),
    .A(_2492_),
    .B(_2496_));
 sg13g2_o21ai_1 _6095_ (.B1(_2497_),
    .Y(_2498_),
    .A1(_2390_),
    .A2(_2492_));
 sg13g2_mux2_1 _6096_ (.A0(_0006_),
    .A1(_2485_),
    .S(_2492_),
    .X(_2499_));
 sg13g2_or2_1 _6097_ (.X(_2500_),
    .B(_2499_),
    .A(_2498_));
 sg13g2_o21ai_1 _6098_ (.B1(_2385_),
    .Y(_2501_),
    .A1(_2482_),
    .A2(_2500_));
 sg13g2_o21ai_1 _6099_ (.B1(_2482_),
    .Y(_2502_),
    .A1(net1120),
    .A2(_2500_));
 sg13g2_or3_1 _6100_ (.A(_2407_),
    .B(_2501_),
    .C(_2502_),
    .X(_2503_));
 sg13g2_nor2_1 _6101_ (.A(_1001_),
    .B(_2458_),
    .Y(_2504_));
 sg13g2_a21o_1 _6102_ (.A2(_2504_),
    .A1(_2454_),
    .B1(_2459_),
    .X(_2505_));
 sg13g2_a21o_1 _6103_ (.A2(_2505_),
    .A1(_2503_),
    .B1(_2481_),
    .X(_0286_));
 sg13g2_nor2b_1 _6104_ (.A(net1190),
    .B_N(net594),
    .Y(_2506_));
 sg13g2_nand2_1 _6105_ (.Y(_2507_),
    .A(_2882_),
    .B(_2500_));
 sg13g2_a21oi_1 _6106_ (.A1(_2498_),
    .A2(_2499_),
    .Y(_2508_),
    .B1(_2507_));
 sg13g2_or3_1 _6107_ (.A(_2407_),
    .B(_2501_),
    .C(_2508_),
    .X(_2509_));
 sg13g2_a21o_1 _6108_ (.A2(_2509_),
    .A1(_2505_),
    .B1(_2506_),
    .X(_0287_));
 sg13g2_mux2_1 _6109_ (.A0(net471),
    .A1(net390),
    .S(net1192),
    .X(_0288_));
 sg13g2_mux2_1 _6110_ (.A0(net506),
    .A1(_1411_),
    .S(net1190),
    .X(_0289_));
 sg13g2_xnor2_1 _6111_ (.Y(_2510_),
    .A(\dtop.oct_counter[3] ),
    .B(_0925_));
 sg13g2_nor2_1 _6112_ (.A(_0935_),
    .B(_2510_),
    .Y(_0290_));
 sg13g2_xnor2_1 _6113_ (.Y(_2511_),
    .A(net601),
    .B(_0926_));
 sg13g2_nor2_1 _6114_ (.A(net1050),
    .B(net602),
    .Y(_0291_));
 sg13g2_a21oi_1 _6115_ (.A1(_2672_),
    .A2(_0926_),
    .Y(_2512_),
    .B1(net1177));
 sg13g2_nor3_1 _6116_ (.A(_0927_),
    .B(_0935_),
    .C(net576),
    .Y(_0292_));
 sg13g2_nor2_1 _6117_ (.A(net1176),
    .B(_0927_),
    .Y(_2513_));
 sg13g2_nor3_1 _6118_ (.A(_0928_),
    .B(net1050),
    .C(_2513_),
    .Y(_0293_));
 sg13g2_xnor2_1 _6119_ (.Y(_2514_),
    .A(net1175),
    .B(_0928_));
 sg13g2_nor2_1 _6120_ (.A(net1050),
    .B(_2514_),
    .Y(_0294_));
 sg13g2_nor2b_1 _6121_ (.A(net613),
    .B_N(_0928_),
    .Y(_2515_));
 sg13g2_xnor2_1 _6122_ (.Y(_2516_),
    .A(net1169),
    .B(_2515_));
 sg13g2_nor2_1 _6123_ (.A(net1050),
    .B(net614),
    .Y(_0295_));
 sg13g2_xnor2_1 _6124_ (.Y(_2517_),
    .A(net580),
    .B(_0929_));
 sg13g2_nor2_1 _6125_ (.A(net1050),
    .B(_2517_),
    .Y(_0296_));
 sg13g2_nor2b_1 _6126_ (.A(net550),
    .B_N(_0929_),
    .Y(_2518_));
 sg13g2_xnor2_1 _6127_ (.Y(_2519_),
    .A(net1166),
    .B(_2518_));
 sg13g2_nor2_1 _6128_ (.A(net1050),
    .B(net551),
    .Y(_0297_));
 sg13g2_xnor2_1 _6129_ (.Y(_2520_),
    .A(_2663_),
    .B(_0936_));
 sg13g2_nor2_1 _6130_ (.A(net1050),
    .B(_2520_),
    .Y(_0298_));
 sg13g2_nor2b_1 _6131_ (.A(_2843_),
    .B_N(net1001),
    .Y(_2521_));
 sg13g2_o21ai_1 _6132_ (.B1(net1249),
    .Y(_2522_),
    .A1(net630),
    .A2(net981));
 sg13g2_xnor2_1 _6133_ (.Y(_2523_),
    .A(_0896_),
    .B(_0899_));
 sg13g2_a21oi_1 _6134_ (.A1(net981),
    .A2(_2523_),
    .Y(_0299_),
    .B1(_2522_));
 sg13g2_xnor2_1 _6135_ (.Y(_2524_),
    .A(_0900_),
    .B(_0901_));
 sg13g2_o21ai_1 _6136_ (.B1(net1248),
    .Y(_2525_),
    .A1(net638),
    .A2(net980));
 sg13g2_a21oi_1 _6137_ (.A1(net980),
    .A2(_2524_),
    .Y(_0300_),
    .B1(_2525_));
 sg13g2_xnor2_1 _6138_ (.Y(_2526_),
    .A(_0902_),
    .B(_0903_));
 sg13g2_o21ai_1 _6139_ (.B1(net1248),
    .Y(_2527_),
    .A1(net646),
    .A2(net980));
 sg13g2_a21oi_1 _6140_ (.A1(net980),
    .A2(_2526_),
    .Y(_0301_),
    .B1(_2527_));
 sg13g2_xnor2_1 _6141_ (.Y(_2528_),
    .A(_0905_),
    .B(_0908_));
 sg13g2_o21ai_1 _6142_ (.B1(net1249),
    .Y(_2529_),
    .A1(net642),
    .A2(net980));
 sg13g2_a21oi_1 _6143_ (.A1(net980),
    .A2(_2528_),
    .Y(_0302_),
    .B1(_2529_));
 sg13g2_xnor2_1 _6144_ (.Y(_2530_),
    .A(_0909_),
    .B(_0910_));
 sg13g2_o21ai_1 _6145_ (.B1(net1252),
    .Y(_2531_),
    .A1(net635),
    .A2(net980));
 sg13g2_a21oi_1 _6146_ (.A1(net980),
    .A2(_2530_),
    .Y(_0303_),
    .B1(_2531_));
 sg13g2_a21oi_1 _6147_ (.A1(net599),
    .A2(net1248),
    .Y(_2532_),
    .B1(net981));
 sg13g2_and2_1 _6148_ (.A(_0798_),
    .B(_0799_),
    .X(_2533_));
 sg13g2_xnor2_1 _6149_ (.Y(_2534_),
    .A(_0911_),
    .B(_2533_));
 sg13g2_a21oi_1 _6150_ (.A1(net981),
    .A2(_2534_),
    .Y(_0304_),
    .B1(_2532_));
 sg13g2_nand3b_1 _6151_ (.B(_0798_),
    .C(_0912_),
    .Y(_2535_),
    .A_N(_0775_));
 sg13g2_nand3_1 _6152_ (.B(net982),
    .C(_2535_),
    .A(_0914_),
    .Y(_2536_));
 sg13g2_nand2_1 _6153_ (.Y(_2537_),
    .A(net620),
    .B(net1251));
 sg13g2_o21ai_1 _6154_ (.B1(_2536_),
    .Y(_0305_),
    .A1(net982),
    .A2(_2537_));
 sg13g2_a21oi_1 _6155_ (.A1(net636),
    .A2(net1251),
    .Y(_2538_),
    .B1(net982));
 sg13g2_nor2_1 _6156_ (.A(_0744_),
    .B(_0745_),
    .Y(_2539_));
 sg13g2_xnor2_1 _6157_ (.Y(_2540_),
    .A(_0915_),
    .B(_2539_));
 sg13g2_a21oi_1 _6158_ (.A1(net982),
    .A2(_2540_),
    .Y(_0306_),
    .B1(_2538_));
 sg13g2_nor3_1 _6159_ (.A(_0720_),
    .B(_0745_),
    .C(_0916_),
    .Y(_2541_));
 sg13g2_nand2_1 _6160_ (.Y(_2542_),
    .A(_0917_),
    .B(_2521_));
 sg13g2_nand3b_1 _6161_ (.B(net1251),
    .C(net586),
    .Y(_2543_),
    .A_N(net982));
 sg13g2_o21ai_1 _6162_ (.B1(_2543_),
    .Y(_0307_),
    .A1(_2541_),
    .A2(_2542_));
 sg13g2_and2_1 _6163_ (.A(\dtop.player_inst.synth.alu.acc[9] ),
    .B(net1252),
    .X(_2544_));
 sg13g2_nor2b_1 _6164_ (.A(_0697_),
    .B_N(_0698_),
    .Y(_2545_));
 sg13g2_xnor2_1 _6165_ (.Y(_2546_),
    .A(_0918_),
    .B(_2545_));
 sg13g2_mux2_1 _6166_ (.A0(_2544_),
    .A1(_2546_),
    .S(net982),
    .X(_0308_));
 sg13g2_xnor2_1 _6167_ (.Y(_2547_),
    .A(_0549_),
    .B(_0919_));
 sg13g2_o21ai_1 _6168_ (.B1(net1251),
    .Y(_2548_),
    .A1(net1165),
    .A2(net982));
 sg13g2_a21oi_1 _6169_ (.A1(net982),
    .A2(_2547_),
    .Y(_0309_),
    .B1(_2548_));
 sg13g2_nand2_1 _6170_ (.Y(_2549_),
    .A(_2853_),
    .B(net1001));
 sg13g2_nand3_1 _6171_ (.B(net1248),
    .C(net979),
    .A(net373),
    .Y(_2550_));
 sg13g2_o21ai_1 _6172_ (.B1(_2550_),
    .Y(_0310_),
    .A1(_2636_),
    .A2(net979));
 sg13g2_nand3_1 _6173_ (.B(net1248),
    .C(net979),
    .A(net500),
    .Y(_2551_));
 sg13g2_o21ai_1 _6174_ (.B1(_2551_),
    .Y(_0311_),
    .A1(_2635_),
    .A2(net979));
 sg13g2_nand3_1 _6175_ (.B(net1249),
    .C(net979),
    .A(net442),
    .Y(_2552_));
 sg13g2_o21ai_1 _6176_ (.B1(_2552_),
    .Y(_0312_),
    .A1(_2634_),
    .A2(net979));
 sg13g2_nand3_1 _6177_ (.B(net1249),
    .C(net978),
    .A(net449),
    .Y(_2553_));
 sg13g2_o21ai_1 _6178_ (.B1(_2553_),
    .Y(_0313_),
    .A1(_2633_),
    .A2(net978));
 sg13g2_nand3_1 _6179_ (.B(net1249),
    .C(net978),
    .A(net395),
    .Y(_2554_));
 sg13g2_o21ai_1 _6180_ (.B1(_2554_),
    .Y(_0314_),
    .A1(_2632_),
    .A2(net978));
 sg13g2_nand3_1 _6181_ (.B(net1249),
    .C(net978),
    .A(net445),
    .Y(_2555_));
 sg13g2_o21ai_1 _6182_ (.B1(_2555_),
    .Y(_0315_),
    .A1(_2631_),
    .A2(net978));
 sg13g2_nand3_1 _6183_ (.B(net1249),
    .C(net978),
    .A(net417),
    .Y(_2556_));
 sg13g2_o21ai_1 _6184_ (.B1(_2556_),
    .Y(_0316_),
    .A1(_2630_),
    .A2(net978));
 sg13g2_nor3_1 _6185_ (.A(_2857_),
    .B(_2943_),
    .C(_0472_),
    .Y(_2557_));
 sg13g2_nand2_1 _6186_ (.Y(_2558_),
    .A(_0428_),
    .B(_0463_));
 sg13g2_nor2_1 _6187_ (.A(_2856_),
    .B(_2868_),
    .Y(_2559_));
 sg13g2_nand3_1 _6188_ (.B(_2831_),
    .C(_0416_),
    .A(net1250),
    .Y(_2560_));
 sg13g2_nor4_1 _6189_ (.A(_2810_),
    .B(_2852_),
    .C(_2866_),
    .D(_2560_),
    .Y(_2561_));
 sg13g2_nor4_1 _6190_ (.A(_2942_),
    .B(_2944_),
    .C(_2946_),
    .D(_0432_),
    .Y(_2562_));
 sg13g2_a21oi_1 _6191_ (.A1(net1136),
    .A2(net1130),
    .Y(_2563_),
    .B1(_2863_));
 sg13g2_nand2_1 _6192_ (.Y(_2564_),
    .A(_2562_),
    .B(_2563_));
 sg13g2_nand4_1 _6193_ (.B(_2557_),
    .C(_2559_),
    .A(_2834_),
    .Y(_2565_),
    .D(_2561_));
 sg13g2_or4_1 _6194_ (.A(_0474_),
    .B(_2558_),
    .C(_2564_),
    .D(_2565_),
    .X(_2566_));
 sg13g2_nor4_2 _6195_ (.A(_2799_),
    .B(_2905_),
    .C(_2930_),
    .Y(_2567_),
    .D(_2566_));
 sg13g2_o21ai_1 _6196_ (.B1(net1241),
    .Y(_2568_),
    .A1(net507),
    .A2(net975));
 sg13g2_a21oi_1 _6197_ (.A1(_2636_),
    .A2(net975),
    .Y(_0317_),
    .B1(_2568_));
 sg13g2_o21ai_1 _6198_ (.B1(net1244),
    .Y(_2569_),
    .A1(net529),
    .A2(net977));
 sg13g2_a21oi_1 _6199_ (.A1(_2635_),
    .A2(net977),
    .Y(_0318_),
    .B1(_2569_));
 sg13g2_o21ai_1 _6200_ (.B1(net1241),
    .Y(_2570_),
    .A1(net524),
    .A2(net976));
 sg13g2_a21oi_1 _6201_ (.A1(_2634_),
    .A2(net976),
    .Y(_0319_),
    .B1(_2570_));
 sg13g2_o21ai_1 _6202_ (.B1(net1241),
    .Y(_2571_),
    .A1(net511),
    .A2(net975));
 sg13g2_a21oi_1 _6203_ (.A1(_2633_),
    .A2(net975),
    .Y(_0320_),
    .B1(_2571_));
 sg13g2_o21ai_1 _6204_ (.B1(net1242),
    .Y(_2572_),
    .A1(net552),
    .A2(net976));
 sg13g2_a21oi_1 _6205_ (.A1(_2632_),
    .A2(net976),
    .Y(_0321_),
    .B1(_2572_));
 sg13g2_o21ai_1 _6206_ (.B1(net1241),
    .Y(_2573_),
    .A1(net559),
    .A2(net975));
 sg13g2_a21oi_1 _6207_ (.A1(_2631_),
    .A2(net975),
    .Y(_0322_),
    .B1(_2573_));
 sg13g2_o21ai_1 _6208_ (.B1(net1241),
    .Y(_2574_),
    .A1(net521),
    .A2(net975));
 sg13g2_a21oi_1 _6209_ (.A1(_2630_),
    .A2(net975),
    .Y(_0323_),
    .B1(_2574_));
 sg13g2_o21ai_1 _6210_ (.B1(net1244),
    .Y(_2575_),
    .A1(net534),
    .A2(_2567_));
 sg13g2_a21oi_1 _6211_ (.A1(_2637_),
    .A2(_2567_),
    .Y(_0324_),
    .B1(_2575_));
 sg13g2_o21ai_1 _6212_ (.B1(net1246),
    .Y(_2576_),
    .A1(net514),
    .A2(net977));
 sg13g2_a21oi_1 _6213_ (.A1(_2640_),
    .A2(_2567_),
    .Y(_0325_),
    .B1(_2576_));
 sg13g2_o21ai_1 _6214_ (.B1(net1246),
    .Y(_2577_),
    .A1(net553),
    .A2(net977));
 sg13g2_a21oi_1 _6215_ (.A1(_2639_),
    .A2(net977),
    .Y(_0326_),
    .B1(_2577_));
 sg13g2_o21ai_1 _6216_ (.B1(net1248),
    .Y(_2578_),
    .A1(net525),
    .A2(net977));
 sg13g2_a21oi_1 _6217_ (.A1(_2638_),
    .A2(net977),
    .Y(_0327_),
    .B1(_2578_));
 sg13g2_nand3_1 _6218_ (.B(_2852_),
    .C(net1001),
    .A(net1224),
    .Y(_2579_));
 sg13g2_nand3_1 _6219_ (.B(net1239),
    .C(net971),
    .A(net382),
    .Y(_2580_));
 sg13g2_o21ai_1 _6220_ (.B1(_2580_),
    .Y(_0328_),
    .A1(_2636_),
    .A2(net971));
 sg13g2_nand3_1 _6221_ (.B(net1244),
    .C(net973),
    .A(net344),
    .Y(_2581_));
 sg13g2_o21ai_1 _6222_ (.B1(_2581_),
    .Y(_0329_),
    .A1(_2635_),
    .A2(net973));
 sg13g2_nand3_1 _6223_ (.B(net1240),
    .C(net971),
    .A(net381),
    .Y(_2582_));
 sg13g2_o21ai_1 _6224_ (.B1(_2582_),
    .Y(_0330_),
    .A1(_2634_),
    .A2(net971));
 sg13g2_nand3_1 _6225_ (.B(net1240),
    .C(net971),
    .A(net348),
    .Y(_2583_));
 sg13g2_o21ai_1 _6226_ (.B1(_2583_),
    .Y(_0331_),
    .A1(_2633_),
    .A2(net971));
 sg13g2_nand3_1 _6227_ (.B(net1242),
    .C(net972),
    .A(net380),
    .Y(_2584_));
 sg13g2_o21ai_1 _6228_ (.B1(_2584_),
    .Y(_0332_),
    .A1(_2632_),
    .A2(net972));
 sg13g2_nand3_1 _6229_ (.B(net1240),
    .C(net971),
    .A(net386),
    .Y(_2585_));
 sg13g2_o21ai_1 _6230_ (.B1(_2585_),
    .Y(_0333_),
    .A1(_2631_),
    .A2(net971));
 sg13g2_nand3_1 _6231_ (.B(net1239),
    .C(net972),
    .A(net346),
    .Y(_2586_));
 sg13g2_o21ai_1 _6232_ (.B1(_2586_),
    .Y(_0334_),
    .A1(_2630_),
    .A2(net972));
 sg13g2_nand3_1 _6233_ (.B(net1244),
    .C(net973),
    .A(net377),
    .Y(_2587_));
 sg13g2_o21ai_1 _6234_ (.B1(_2587_),
    .Y(_0335_),
    .A1(_2637_),
    .A2(net973));
 sg13g2_nand3_1 _6235_ (.B(net1244),
    .C(net973),
    .A(net392),
    .Y(_2588_));
 sg13g2_o21ai_1 _6236_ (.B1(_2588_),
    .Y(_0336_),
    .A1(_2640_),
    .A2(net973));
 sg13g2_nand3_1 _6237_ (.B(net1246),
    .C(net974),
    .A(net353),
    .Y(_2589_));
 sg13g2_o21ai_1 _6238_ (.B1(_2589_),
    .Y(_0337_),
    .A1(_2639_),
    .A2(net974));
 sg13g2_nand3_1 _6239_ (.B(net1248),
    .C(net973),
    .A(net418),
    .Y(_2590_));
 sg13g2_o21ai_1 _6240_ (.B1(_2590_),
    .Y(_0338_),
    .A1(_2638_),
    .A2(net973));
 sg13g2_nand3b_1 _6241_ (.B(_2406_),
    .C(net1190),
    .Y(_2591_),
    .A_N(net4));
 sg13g2_o21ai_1 _6242_ (.B1(_2591_),
    .Y(_0339_),
    .A1(net1190),
    .A2(_2702_));
 sg13g2_nand2_2 _6243_ (.Y(_2592_),
    .A(_2856_),
    .B(net1001));
 sg13g2_nand3_1 _6244_ (.B(net1239),
    .C(net969),
    .A(net368),
    .Y(_2593_));
 sg13g2_o21ai_1 _6245_ (.B1(_2593_),
    .Y(_0340_),
    .A1(_2636_),
    .A2(net969));
 sg13g2_nand3_1 _6246_ (.B(net1244),
    .C(net970),
    .A(net331),
    .Y(_2594_));
 sg13g2_o21ai_1 _6247_ (.B1(_2594_),
    .Y(_0341_),
    .A1(_2635_),
    .A2(net970));
 sg13g2_nand3_1 _6248_ (.B(net1238),
    .C(net969),
    .A(net327),
    .Y(_2595_));
 sg13g2_o21ai_1 _6249_ (.B1(_2595_),
    .Y(_0342_),
    .A1(_2634_),
    .A2(net969));
 sg13g2_nand3_1 _6250_ (.B(net1238),
    .C(net969),
    .A(net372),
    .Y(_2596_));
 sg13g2_o21ai_1 _6251_ (.B1(_2596_),
    .Y(_0343_),
    .A1(_2633_),
    .A2(net969));
 sg13g2_nand3_1 _6252_ (.B(net1242),
    .C(net970),
    .A(net352),
    .Y(_2597_));
 sg13g2_o21ai_1 _6253_ (.B1(_2597_),
    .Y(_0344_),
    .A1(_2632_),
    .A2(_2592_));
 sg13g2_nand3_1 _6254_ (.B(net1239),
    .C(net969),
    .A(net342),
    .Y(_2598_));
 sg13g2_o21ai_1 _6255_ (.B1(_2598_),
    .Y(_0345_),
    .A1(_2631_),
    .A2(net969));
 sg13g2_nand3_1 _6256_ (.B(net1239),
    .C(net970),
    .A(net371),
    .Y(_2599_));
 sg13g2_o21ai_1 _6257_ (.B1(_2599_),
    .Y(_0346_),
    .A1(_2630_),
    .A2(net970));
 sg13g2_nand3_1 _6258_ (.B(net1244),
    .C(net970),
    .A(net383),
    .Y(_2600_));
 sg13g2_o21ai_1 _6259_ (.B1(_2600_),
    .Y(_0347_),
    .A1(_2637_),
    .A2(net970));
 sg13g2_nand2b_2 _6260_ (.Y(_2601_),
    .B(net1001),
    .A_N(_2557_));
 sg13g2_nand3_1 _6261_ (.B(net1245),
    .C(net965),
    .A(net447),
    .Y(_2602_));
 sg13g2_o21ai_1 _6262_ (.B1(_2602_),
    .Y(_0348_),
    .A1(_2636_),
    .A2(net965));
 sg13g2_nand3_1 _6263_ (.B(net1245),
    .C(net966),
    .A(net349),
    .Y(_2603_));
 sg13g2_o21ai_1 _6264_ (.B1(_2603_),
    .Y(_0349_),
    .A1(_2635_),
    .A2(net966));
 sg13g2_nand3_1 _6265_ (.B(net1247),
    .C(net965),
    .A(net411),
    .Y(_2604_));
 sg13g2_o21ai_1 _6266_ (.B1(_2604_),
    .Y(_0350_),
    .A1(_2634_),
    .A2(net965));
 sg13g2_nand3_1 _6267_ (.B(net1247),
    .C(net965),
    .A(net338),
    .Y(_2605_));
 sg13g2_o21ai_1 _6268_ (.B1(_2605_),
    .Y(_0351_),
    .A1(_2633_),
    .A2(net966));
 sg13g2_nand3_1 _6269_ (.B(net1246),
    .C(net967),
    .A(net450),
    .Y(_2606_));
 sg13g2_o21ai_1 _6270_ (.B1(_2606_),
    .Y(_0352_),
    .A1(_2632_),
    .A2(net967));
 sg13g2_nand3_1 _6271_ (.B(net1247),
    .C(net965),
    .A(net354),
    .Y(_2607_));
 sg13g2_o21ai_1 _6272_ (.B1(_2607_),
    .Y(_0353_),
    .A1(_2631_),
    .A2(net965));
 sg13g2_nand3_1 _6273_ (.B(net1247),
    .C(net965),
    .A(net317),
    .Y(_2608_));
 sg13g2_o21ai_1 _6274_ (.B1(_2608_),
    .Y(_0354_),
    .A1(_2630_),
    .A2(net966));
 sg13g2_nand3_1 _6275_ (.B(net1246),
    .C(net968),
    .A(net324),
    .Y(_2609_));
 sg13g2_o21ai_1 _6276_ (.B1(_2609_),
    .Y(_0355_),
    .A1(_2637_),
    .A2(net968));
 sg13g2_nand3_1 _6277_ (.B(net1245),
    .C(net967),
    .A(net313),
    .Y(_2610_));
 sg13g2_o21ai_1 _6278_ (.B1(_2610_),
    .Y(_0356_),
    .A1(_2640_),
    .A2(net967));
 sg13g2_nand3_1 _6279_ (.B(net1246),
    .C(net967),
    .A(net319),
    .Y(_2611_));
 sg13g2_o21ai_1 _6280_ (.B1(_2611_),
    .Y(_0357_),
    .A1(_2639_),
    .A2(net967));
 sg13g2_nand3_1 _6281_ (.B(net1246),
    .C(net967),
    .A(net339),
    .Y(_2612_));
 sg13g2_o21ai_1 _6282_ (.B1(_2612_),
    .Y(_0358_),
    .A1(_2638_),
    .A2(net967));
 sg13g2_nand2_2 _6283_ (.Y(_2613_),
    .A(_2868_),
    .B(net1001));
 sg13g2_nand3_1 _6284_ (.B(net1238),
    .C(net963),
    .A(net379),
    .Y(_2614_));
 sg13g2_o21ai_1 _6285_ (.B1(_2614_),
    .Y(_0359_),
    .A1(_2636_),
    .A2(net963));
 sg13g2_nand3_1 _6286_ (.B(net1241),
    .C(_2613_),
    .A(net364),
    .Y(_2615_));
 sg13g2_o21ai_1 _6287_ (.B1(_2615_),
    .Y(_0360_),
    .A1(_2635_),
    .A2(net964));
 sg13g2_nand3_1 _6288_ (.B(net1240),
    .C(net963),
    .A(net441),
    .Y(_2616_));
 sg13g2_o21ai_1 _6289_ (.B1(_2616_),
    .Y(_0361_),
    .A1(_2634_),
    .A2(net963));
 sg13g2_nand3_1 _6290_ (.B(net1238),
    .C(net963),
    .A(net439),
    .Y(_2617_));
 sg13g2_o21ai_1 _6291_ (.B1(_2617_),
    .Y(_0362_),
    .A1(_2633_),
    .A2(net963));
 sg13g2_nand3_1 _6292_ (.B(net1241),
    .C(net964),
    .A(net375),
    .Y(_2618_));
 sg13g2_o21ai_1 _6293_ (.B1(_2618_),
    .Y(_0363_),
    .A1(_2632_),
    .A2(net964));
 sg13g2_nand3_1 _6294_ (.B(net1239),
    .C(net963),
    .A(net360),
    .Y(_2619_));
 sg13g2_o21ai_1 _6295_ (.B1(_2619_),
    .Y(_0364_),
    .A1(_2631_),
    .A2(net963));
 sg13g2_nand3_1 _6296_ (.B(net1241),
    .C(net964),
    .A(net410),
    .Y(_2620_));
 sg13g2_o21ai_1 _6297_ (.B1(_2620_),
    .Y(_0365_),
    .A1(_2630_),
    .A2(net964));
 sg13g2_nand3_1 _6298_ (.B(net1244),
    .C(net964),
    .A(net361),
    .Y(_2621_));
 sg13g2_o21ai_1 _6299_ (.B1(_2621_),
    .Y(_0366_),
    .A1(_2637_),
    .A2(net964));
 sg13g2_nand2_2 _6300_ (.Y(_2622_),
    .A(net1001),
    .B(_2564_));
 sg13g2_nand3_1 _6301_ (.B(net1238),
    .C(net961),
    .A(net420),
    .Y(_2623_));
 sg13g2_o21ai_1 _6302_ (.B1(_2623_),
    .Y(_0367_),
    .A1(_2636_),
    .A2(net961));
 sg13g2_nand3_1 _6303_ (.B(net1245),
    .C(net962),
    .A(net336),
    .Y(_2624_));
 sg13g2_o21ai_1 _6304_ (.B1(_2624_),
    .Y(_0368_),
    .A1(_2635_),
    .A2(net962));
 sg13g2_nand3_1 _6305_ (.B(net1238),
    .C(net961),
    .A(net398),
    .Y(_2625_));
 sg13g2_o21ai_1 _6306_ (.B1(_2625_),
    .Y(_0369_),
    .A1(_2634_),
    .A2(net961));
 sg13g2_nand3_1 _6307_ (.B(net1238),
    .C(net961),
    .A(net397),
    .Y(_2626_));
 sg13g2_o21ai_1 _6308_ (.B1(_2626_),
    .Y(_0370_),
    .A1(_2633_),
    .A2(net961));
 sg13g2_nand3_1 _6309_ (.B(net1243),
    .C(net962),
    .A(net356),
    .Y(_2627_));
 sg13g2_o21ai_1 _6310_ (.B1(_2627_),
    .Y(_0371_),
    .A1(_2632_),
    .A2(net962));
 sg13g2_nand3_1 _6311_ (.B(net1238),
    .C(net961),
    .A(net326),
    .Y(_2628_));
 sg13g2_o21ai_1 _6312_ (.B1(_2628_),
    .Y(_0372_),
    .A1(_2631_),
    .A2(net961));
 sg13g2_nand3_1 _6313_ (.B(net1239),
    .C(net962),
    .A(net347),
    .Y(_2629_));
 sg13g2_o21ai_1 _6314_ (.B1(_2629_),
    .Y(_0373_),
    .A1(_2630_),
    .A2(net962));
 sg13g2_dfrbp_1 _6315_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net213),
    .D(_0089_),
    .Q_N(_3156_),
    .Q(\dtop.player_inst.synth.alu.carry ));
 sg13g2_dfrbp_1 _6316_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net204),
    .D(_0090_),
    .Q_N(_0083_),
    .Q(\dtop.detune_counter[4] ));
 sg13g2_dfrbp_1 _6317_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net203),
    .D(_0091_),
    .Q_N(_0051_),
    .Q(\dtop.detune_counter[5] ));
 sg13g2_dfrbp_1 _6318_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net202),
    .D(_0092_),
    .Q_N(_0080_),
    .Q(\dtop.detune_counter[6] ));
 sg13g2_dfrbp_1 _6319_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net201),
    .D(_0093_),
    .Q_N(_0079_),
    .Q(\dtop.detune_counter[7] ));
 sg13g2_dfrbp_1 _6320_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net200),
    .D(_0094_),
    .Q_N(_0078_),
    .Q(\dtop.detune_counter[8] ));
 sg13g2_dfrbp_1 _6321_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net199),
    .D(_0095_),
    .Q_N(_0075_),
    .Q(\dtop.detune_counter[9] ));
 sg13g2_dfrbp_1 _6322_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net198),
    .D(_0096_),
    .Q_N(_0073_),
    .Q(\dtop.detune_counter[10] ));
 sg13g2_dfrbp_1 _6323_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net197),
    .D(_0097_),
    .Q_N(_0072_),
    .Q(\dtop.detune_counter[11] ));
 sg13g2_dfrbp_1 _6324_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net196),
    .D(_0098_),
    .Q_N(_0070_),
    .Q(\dtop.detune_counter[12] ));
 sg13g2_dfrbp_1 _6325_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net195),
    .D(_0099_),
    .Q_N(_0087_),
    .Q(\dtop.detune_counter[13] ));
 sg13g2_dfrbp_1 _6326_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net194),
    .D(_0100_),
    .Q_N(_0061_),
    .Q(\dtop.detune_counter[14] ));
 sg13g2_dfrbp_1 _6327_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net193),
    .D(_0101_),
    .Q_N(_0000_),
    .Q(\dtop.detune_counter[15] ));
 sg13g2_dfrbp_1 _6328_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net192),
    .D(_0102_),
    .Q_N(_0058_),
    .Q(\dtop.detune_counter[16] ));
 sg13g2_dfrbp_1 _6329_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net191),
    .D(_0103_),
    .Q_N(_0057_),
    .Q(\dtop.detune_counter[17] ));
 sg13g2_dfrbp_1 _6330_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net190),
    .D(_0104_),
    .Q_N(_0009_),
    .Q(\dtop.vtop.dphases[0][0] ));
 sg13g2_dfrbp_1 _6331_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net189),
    .D(_0105_),
    .Q_N(_0011_),
    .Q(\dtop.vtop.dphases[0][1] ));
 sg13g2_dfrbp_1 _6332_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net188),
    .D(_0106_),
    .Q_N(_0013_),
    .Q(\dtop.vtop.dphases[0][2] ));
 sg13g2_dfrbp_1 _6333_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net187),
    .D(_0107_),
    .Q_N(_0015_),
    .Q(\dtop.vtop.dphases[0][3] ));
 sg13g2_dfrbp_1 _6334_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net186),
    .D(_0108_),
    .Q_N(_0017_),
    .Q(\dtop.vtop.dphases[0][4] ));
 sg13g2_dfrbp_1 _6335_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net185),
    .D(_0109_),
    .Q_N(_0019_),
    .Q(\dtop.vtop.dphases[0][5] ));
 sg13g2_dfrbp_1 _6336_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net184),
    .D(_0110_),
    .Q_N(_0021_),
    .Q(\dtop.vtop.dphases[0][6] ));
 sg13g2_dfrbp_1 _6337_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net183),
    .D(_0111_),
    .Q_N(_0023_),
    .Q(\dtop.vtop.dphases[0][7] ));
 sg13g2_dfrbp_1 _6338_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net182),
    .D(_0112_),
    .Q_N(_0026_),
    .Q(\dtop.vtop.dphases[0][8] ));
 sg13g2_dfrbp_1 _6339_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net181),
    .D(_0113_),
    .Q_N(_0028_),
    .Q(\dtop.vtop.dphases[0][9] ));
 sg13g2_dfrbp_1 _6340_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net180),
    .D(_0114_),
    .Q_N(_0030_),
    .Q(\dtop.vtop.dphases[0][10] ));
 sg13g2_dfrbp_1 _6341_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net179),
    .D(_0115_),
    .Q_N(_3155_),
    .Q(\dtop.vtop.dphases[1][0] ));
 sg13g2_dfrbp_1 _6342_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net178),
    .D(_0116_),
    .Q_N(_3154_),
    .Q(\dtop.vtop.dphases[1][1] ));
 sg13g2_dfrbp_1 _6343_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net177),
    .D(_0117_),
    .Q_N(_3153_),
    .Q(\dtop.vtop.dphases[1][2] ));
 sg13g2_dfrbp_1 _6344_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net176),
    .D(_0118_),
    .Q_N(_3152_),
    .Q(\dtop.vtop.dphases[1][3] ));
 sg13g2_dfrbp_1 _6345_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net175),
    .D(_0119_),
    .Q_N(_3151_),
    .Q(\dtop.vtop.dphases[1][4] ));
 sg13g2_dfrbp_1 _6346_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net174),
    .D(_0120_),
    .Q_N(_3150_),
    .Q(\dtop.vtop.dphases[1][5] ));
 sg13g2_dfrbp_1 _6347_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net173),
    .D(_0121_),
    .Q_N(_3149_),
    .Q(\dtop.vtop.dphases[1][6] ));
 sg13g2_dfrbp_1 _6348_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net172),
    .D(_0122_),
    .Q_N(_3148_),
    .Q(\dtop.vtop.dphases[1][7] ));
 sg13g2_dfrbp_1 _6349_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net171),
    .D(_0123_),
    .Q_N(_3147_),
    .Q(\dtop.vtop.dphases[1][8] ));
 sg13g2_dfrbp_1 _6350_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net170),
    .D(_0124_),
    .Q_N(_3146_),
    .Q(\dtop.vtop.dphases[1][9] ));
 sg13g2_dfrbp_1 _6351_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net169),
    .D(_0125_),
    .Q_N(_3145_),
    .Q(\dtop.vtop.dphases[1][10] ));
 sg13g2_dfrbp_1 _6352_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net168),
    .D(_0126_),
    .Q_N(_3144_),
    .Q(\dtop.vtop.dphases[2][0] ));
 sg13g2_dfrbp_1 _6353_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net167),
    .D(_0127_),
    .Q_N(_3143_),
    .Q(\dtop.vtop.dphases[2][1] ));
 sg13g2_dfrbp_1 _6354_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net166),
    .D(_0128_),
    .Q_N(_3142_),
    .Q(\dtop.vtop.dphases[2][2] ));
 sg13g2_dfrbp_1 _6355_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net165),
    .D(_0129_),
    .Q_N(_3141_),
    .Q(\dtop.vtop.dphases[2][3] ));
 sg13g2_dfrbp_1 _6356_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net164),
    .D(_0130_),
    .Q_N(_3140_),
    .Q(\dtop.vtop.dphases[2][4] ));
 sg13g2_dfrbp_1 _6357_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net163),
    .D(_0131_),
    .Q_N(_3139_),
    .Q(\dtop.vtop.dphases[2][5] ));
 sg13g2_dfrbp_1 _6358_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net162),
    .D(_0132_),
    .Q_N(_3138_),
    .Q(\dtop.vtop.dphases[2][6] ));
 sg13g2_dfrbp_1 _6359_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net161),
    .D(_0133_),
    .Q_N(_3137_),
    .Q(\dtop.vtop.dphases[2][7] ));
 sg13g2_dfrbp_1 _6360_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net160),
    .D(_0134_),
    .Q_N(_3136_),
    .Q(\dtop.vtop.dphases[2][8] ));
 sg13g2_dfrbp_1 _6361_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net159),
    .D(_0135_),
    .Q_N(_3135_),
    .Q(\dtop.vtop.dphases[2][9] ));
 sg13g2_dfrbp_1 _6362_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net158),
    .D(_0136_),
    .Q_N(_3134_),
    .Q(\dtop.vtop.dphases[2][10] ));
 sg13g2_dfrbp_1 _6363_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net157),
    .D(_0137_),
    .Q_N(_3133_),
    .Q(\dtop.player_inst.synth.alu.oct_en ));
 sg13g2_dfrbp_1 _6364_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net156),
    .D(_0138_),
    .Q_N(_3132_),
    .Q(\dtop.vtop.rs.saturated ));
 sg13g2_dfrbp_1 _6365_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net155),
    .D(net391),
    .Q_N(_3131_),
    .Q(\dtop.vsync ));
 sg13g2_dfrbp_1 _6366_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net154),
    .D(_0140_),
    .Q_N(_3130_),
    .Q(\dtop.vtop.rs.scan_y.phase[0] ));
 sg13g2_dfrbp_1 _6367_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net153),
    .D(_0141_),
    .Q_N(_3129_),
    .Q(\dtop.vtop.rs.scan_y.phase[1] ));
 sg13g2_dfrbp_1 _6368_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net152),
    .D(_0142_),
    .Q_N(_3128_),
    .Q(\dtop.vtop.rs.x_scan.phase[0] ));
 sg13g2_dfrbp_1 _6369_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net151),
    .D(_0143_),
    .Q_N(_3127_),
    .Q(\dtop.vtop.rs.x_scan.phase[1] ));
 sg13g2_dfrbp_1 _6370_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net150),
    .D(_0144_),
    .Q_N(_3126_),
    .Q(\dtop.player_inst.program_addr[0] ));
 sg13g2_dfrbp_1 _6371_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net149),
    .D(_0145_),
    .Q_N(_0088_),
    .Q(\dtop.player_inst.program_addr[1] ));
 sg13g2_dfrbp_1 _6372_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net148),
    .D(_0146_),
    .Q_N(_0001_),
    .Q(\dtop.player_inst.program_addr[2] ));
 sg13g2_dfrbp_1 _6373_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net147),
    .D(_0147_),
    .Q_N(_0063_),
    .Q(\dtop.player_inst.program_addr[3] ));
 sg13g2_dfrbp_1 _6374_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0148_),
    .Q_N(_3125_),
    .Q(\dtop.player_inst.program_addr[4] ));
 sg13g2_dfrbp_1 _6375_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net145),
    .D(_0149_),
    .Q_N(_3124_),
    .Q(\dtop.player_inst.program_addr[5] ));
 sg13g2_dfrbp_1 _6376_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net144),
    .D(_0150_),
    .Q_N(_0050_),
    .Q(\dtop.player_inst.program_addr[6] ));
 sg13g2_dfrbp_1 _6377_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net143),
    .D(_0151_),
    .Q_N(_3123_),
    .Q(\dtop.vtop.pipeline.nstep_zg[0] ));
 sg13g2_dfrbp_1 _6378_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net142),
    .D(_0152_),
    .Q_N(_3122_),
    .Q(\dtop.vtop.pipeline.nstep_zg[1] ));
 sg13g2_dfrbp_1 _6379_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net141),
    .D(_0153_),
    .Q_N(_0059_),
    .Q(\dtop.vtop.pipeline.neg_t[0] ));
 sg13g2_dfrbp_1 _6380_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net139),
    .D(_0154_),
    .Q_N(_0082_),
    .Q(\dtop.vtop.pipeline.neg_t[1] ));
 sg13g2_dfrbp_1 _6381_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net137),
    .D(_0155_),
    .Q_N(_0081_),
    .Q(\dtop.vtop.pipeline.neg_t[2] ));
 sg13g2_dfrbp_1 _6382_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net135),
    .D(_0156_),
    .Q_N(_0040_),
    .Q(\dtop.vtop.pipeline.neg_t[3] ));
 sg13g2_dfrbp_1 _6383_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net133),
    .D(net520),
    .Q_N(_0077_),
    .Q(\dtop.vtop.pipeline.neg_t[4] ));
 sg13g2_dfrbp_1 _6384_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net131),
    .D(_0158_),
    .Q_N(_0076_),
    .Q(\dtop.vtop.pipeline.neg_t[5] ));
 sg13g2_dfrbp_1 _6385_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net129),
    .D(_0159_),
    .Q_N(_0074_),
    .Q(\dtop.vtop.pipeline.neg_t[6] ));
 sg13g2_dfrbp_1 _6386_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net127),
    .D(net589),
    .Q_N(_0043_),
    .Q(\dtop.vtop.pipeline.neg_t[7] ));
 sg13g2_dfrbp_1 _6387_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net125),
    .D(_0161_),
    .Q_N(_0071_),
    .Q(\dtop.vtop.pipeline.neg_t[8] ));
 sg13g2_dfrbp_1 _6388_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net123),
    .D(_0162_),
    .Q_N(_0041_),
    .Q(\dtop.vtop.pipeline.neg_t[9] ));
 sg13g2_dfrbp_1 _6389_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net121),
    .D(net555),
    .Q_N(_0060_),
    .Q(\dtop.vtop.pipeline.dz[0] ));
 sg13g2_dfrbp_1 _6390_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net119),
    .D(_0164_),
    .Q_N(_0039_),
    .Q(\dtop.vtop.pipeline.dz[1] ));
 sg13g2_dfrbp_1 _6391_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net117),
    .D(_0165_),
    .Q_N(_0069_),
    .Q(\dtop.vtop.pipeline.dz[2] ));
 sg13g2_dfrbp_1 _6392_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net115),
    .D(_0166_),
    .Q_N(_0068_),
    .Q(\dtop.vtop.pipeline.dz[3] ));
 sg13g2_dfrbp_1 _6393_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net113),
    .D(_0167_),
    .Q_N(_0042_),
    .Q(\dtop.vtop.pipeline.dz[4] ));
 sg13g2_dfrbp_1 _6394_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net111),
    .D(_0168_),
    .Q_N(_0067_),
    .Q(\dtop.vtop.pipeline.dz[5] ));
 sg13g2_dfrbp_1 _6395_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net109),
    .D(_0169_),
    .Q_N(_0066_),
    .Q(\dtop.vtop.pipeline.dz[6] ));
 sg13g2_dfrbp_1 _6396_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net107),
    .D(_0170_),
    .Q_N(_0065_),
    .Q(\dtop.vtop.pipeline.dz[7] ));
 sg13g2_dfrbp_1 _6397_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net105),
    .D(_0171_),
    .Q_N(_0064_),
    .Q(\dtop.vtop.pipeline.dz[8] ));
 sg13g2_dfrbp_1 _6398_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net103),
    .D(_0172_),
    .Q_N(_3121_),
    .Q(\dtop.vtop.pipeline.z[0] ));
 sg13g2_dfrbp_1 _6399_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net101),
    .D(_0173_),
    .Q_N(_3120_),
    .Q(\dtop.vtop.pipeline.z[1] ));
 sg13g2_dfrbp_1 _6400_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net99),
    .D(_0174_),
    .Q_N(_3119_),
    .Q(\dtop.vtop.pipeline.z[2] ));
 sg13g2_dfrbp_1 _6401_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net97),
    .D(_0175_),
    .Q_N(_3118_),
    .Q(\dtop.vtop.pipeline.z[3] ));
 sg13g2_dfrbp_1 _6402_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net95),
    .D(net492),
    .Q_N(_3117_),
    .Q(\dtop.vtop.pipeline.z[4] ));
 sg13g2_dfrbp_1 _6403_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net93),
    .D(net593),
    .Q_N(_3116_),
    .Q(\dtop.vtop.pipeline.z[5] ));
 sg13g2_dfrbp_1 _6404_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net91),
    .D(net563),
    .Q_N(_3115_),
    .Q(\dtop.vtop.pipeline.z[6] ));
 sg13g2_dfrbp_1 _6405_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net89),
    .D(_0179_),
    .Q_N(_3114_),
    .Q(\dtop.vtop.pipeline.z[7] ));
 sg13g2_dfrbp_1 _6406_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net87),
    .D(net548),
    .Q_N(_3113_),
    .Q(\dtop.vtop.pipeline.z[8] ));
 sg13g2_dfrbp_1 _6407_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net85),
    .D(_0181_),
    .Q_N(_3112_),
    .Q(\dtop.vtop.pipeline.z[9] ));
 sg13g2_dfrbp_1 _6408_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net83),
    .D(_0182_),
    .Q_N(_3111_),
    .Q(\dtop.vtop.pipeline.z[10] ));
 sg13g2_dfrbp_1 _6409_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net81),
    .D(_0183_),
    .Q_N(_3110_),
    .Q(\dtop.vtop.pipeline.z[11] ));
 sg13g2_dfrbp_1 _6410_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net79),
    .D(_0184_),
    .Q_N(_3109_),
    .Q(\dtop.vtop.pipeline.z[12] ));
 sg13g2_dfrbp_1 _6411_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net77),
    .D(_0185_),
    .Q_N(_3108_),
    .Q(\dtop.vtop.pipeline.z[13] ));
 sg13g2_dfrbp_1 _6412_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net75),
    .D(_0186_),
    .Q_N(_3107_),
    .Q(\dtop.vtop.pipeline.z[14] ));
 sg13g2_dfrbp_1 _6413_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net73),
    .D(net406),
    .Q_N(_3106_),
    .Q(\dtop.vtop.pipeline.phases[1][0] ));
 sg13g2_dfrbp_1 _6414_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net72),
    .D(_0188_),
    .Q_N(_3105_),
    .Q(\dtop.vtop.pipeline.phases[1][1] ));
 sg13g2_dfrbp_1 _6415_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net71),
    .D(_0189_),
    .Q_N(_3104_),
    .Q(\dtop.vtop.pipeline.phases[1][2] ));
 sg13g2_dfrbp_1 _6416_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net70),
    .D(_0190_),
    .Q_N(_3103_),
    .Q(\dtop.vtop.pipeline.phases[1][3] ));
 sg13g2_dfrbp_1 _6417_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net69),
    .D(_0191_),
    .Q_N(_3102_),
    .Q(\dtop.vtop.pipeline.phases[1][4] ));
 sg13g2_dfrbp_1 _6418_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net68),
    .D(_0192_),
    .Q_N(_3101_),
    .Q(\dtop.vtop.pipeline.phases[1][5] ));
 sg13g2_dfrbp_1 _6419_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net67),
    .D(_0193_),
    .Q_N(_3100_),
    .Q(\dtop.vtop.pipeline.phases[1][6] ));
 sg13g2_dfrbp_1 _6420_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net66),
    .D(_0194_),
    .Q_N(_3099_),
    .Q(\dtop.vtop.pipeline.phases[1][7] ));
 sg13g2_dfrbp_1 _6421_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net65),
    .D(_0195_),
    .Q_N(_3098_),
    .Q(\dtop.vtop.pipeline.phases[1][8] ));
 sg13g2_dfrbp_1 _6422_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net64),
    .D(_0196_),
    .Q_N(_3097_),
    .Q(\dtop.vtop.pipeline.phases[1][9] ));
 sg13g2_dfrbp_1 _6423_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net63),
    .D(_0197_),
    .Q_N(_3096_),
    .Q(\dtop.vtop.pipeline.phases[1][10] ));
 sg13g2_dfrbp_1 _6424_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net62),
    .D(_0198_),
    .Q_N(_3095_),
    .Q(\dtop.vtop.pipeline.phases[1][11] ));
 sg13g2_dfrbp_1 _6425_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net61),
    .D(_0199_),
    .Q_N(_3094_),
    .Q(\dtop.vtop.pipeline.phases[1][12] ));
 sg13g2_dfrbp_1 _6426_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net60),
    .D(_0200_),
    .Q_N(_3093_),
    .Q(\dtop.vtop.pipeline.phases[1][13] ));
 sg13g2_dfrbp_1 _6427_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net59),
    .D(_0201_),
    .Q_N(_3092_),
    .Q(\dtop.vtop.pipeline.phases[1][14] ));
 sg13g2_dfrbp_1 _6428_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net58),
    .D(_0202_),
    .Q_N(_3091_),
    .Q(\dtop.vtop.pipeline.phases[1][15] ));
 sg13g2_dfrbp_1 _6429_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net57),
    .D(net495),
    .Q_N(_3090_),
    .Q(\dtop.vtop.pipeline.phases[2][0] ));
 sg13g2_dfrbp_1 _6430_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net56),
    .D(_0204_),
    .Q_N(_3089_),
    .Q(\dtop.vtop.pipeline.phases[2][1] ));
 sg13g2_dfrbp_1 _6431_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net55),
    .D(_0205_),
    .Q_N(_3088_),
    .Q(\dtop.vtop.pipeline.phases[2][2] ));
 sg13g2_dfrbp_1 _6432_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net54),
    .D(_0206_),
    .Q_N(_3087_),
    .Q(\dtop.vtop.pipeline.phases[2][3] ));
 sg13g2_dfrbp_1 _6433_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net53),
    .D(_0207_),
    .Q_N(_3086_),
    .Q(\dtop.vtop.pipeline.phases[2][4] ));
 sg13g2_dfrbp_1 _6434_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net52),
    .D(_0208_),
    .Q_N(_3085_),
    .Q(\dtop.vtop.pipeline.phases[2][5] ));
 sg13g2_dfrbp_1 _6435_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net51),
    .D(_0209_),
    .Q_N(_3084_),
    .Q(\dtop.vtop.pipeline.phases[2][6] ));
 sg13g2_dfrbp_1 _6436_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net50),
    .D(_0210_),
    .Q_N(_3083_),
    .Q(\dtop.vtop.pipeline.phases[2][7] ));
 sg13g2_dfrbp_1 _6437_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net49),
    .D(_0211_),
    .Q_N(_3082_),
    .Q(\dtop.vtop.pipeline.phases[2][8] ));
 sg13g2_dfrbp_1 _6438_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net48),
    .D(_0212_),
    .Q_N(_3081_),
    .Q(\dtop.vtop.pipeline.phases[2][9] ));
 sg13g2_dfrbp_1 _6439_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net47),
    .D(_0213_),
    .Q_N(_3080_),
    .Q(\dtop.vtop.pipeline.phases[2][10] ));
 sg13g2_dfrbp_1 _6440_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net46),
    .D(_0214_),
    .Q_N(_3079_),
    .Q(\dtop.vtop.pipeline.phases[2][11] ));
 sg13g2_dfrbp_1 _6441_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net45),
    .D(_0215_),
    .Q_N(_3078_),
    .Q(\dtop.vtop.pipeline.phases[2][12] ));
 sg13g2_dfrbp_1 _6442_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net44),
    .D(_0216_),
    .Q_N(_3077_),
    .Q(\dtop.vtop.pipeline.phases[2][13] ));
 sg13g2_dfrbp_1 _6443_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net43),
    .D(_0217_),
    .Q_N(_3076_),
    .Q(\dtop.vtop.pipeline.phases[2][14] ));
 sg13g2_dfrbp_1 _6444_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net42),
    .D(_0218_),
    .Q_N(_3075_),
    .Q(\dtop.vtop.pipeline.phases[2][15] ));
 sg13g2_dfrbp_1 _6445_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net41),
    .D(_0219_),
    .Q_N(_2962_),
    .Q(\dtop.enable ));
 sg13g2_dfrbp_1 _6446_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net40),
    .D(net425),
    .Q_N(_0007_),
    .Q(\dtop.vtop.pipeline.phases[0][0] ));
 sg13g2_dfrbp_1 _6447_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net39),
    .D(_0221_),
    .Q_N(_0010_),
    .Q(\dtop.vtop.pipeline.phases[0][1] ));
 sg13g2_dfrbp_1 _6448_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net38),
    .D(_0222_),
    .Q_N(_0012_),
    .Q(\dtop.vtop.pipeline.phases[0][2] ));
 sg13g2_dfrbp_1 _6449_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net37),
    .D(_0223_),
    .Q_N(_0014_),
    .Q(\dtop.vtop.pipeline.phases[0][3] ));
 sg13g2_dfrbp_1 _6450_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net36),
    .D(_0224_),
    .Q_N(_0016_),
    .Q(\dtop.vtop.pipeline.phases[0][4] ));
 sg13g2_dfrbp_1 _6451_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net35),
    .D(_0225_),
    .Q_N(_0018_),
    .Q(\dtop.vtop.pipeline.phases[0][5] ));
 sg13g2_dfrbp_1 _6452_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net34),
    .D(_0226_),
    .Q_N(_0020_),
    .Q(\dtop.vtop.pipeline.phases[0][6] ));
 sg13g2_dfrbp_1 _6453_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net33),
    .D(_0227_),
    .Q_N(_0022_),
    .Q(\dtop.vtop.pipeline.phases[0][7] ));
 sg13g2_dfrbp_1 _6454_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net32),
    .D(_0228_),
    .Q_N(_0024_),
    .Q(\dtop.vtop.pipeline.phases[0][8] ));
 sg13g2_dfrbp_1 _6455_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net31),
    .D(_0229_),
    .Q_N(_0027_),
    .Q(\dtop.vtop.pipeline.phases[0][9] ));
 sg13g2_dfrbp_1 _6456_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net30),
    .D(_0230_),
    .Q_N(_0029_),
    .Q(\dtop.vtop.pipeline.phases[0][10] ));
 sg13g2_dfrbp_1 _6457_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net29),
    .D(_0231_),
    .Q_N(_0031_),
    .Q(\dtop.vtop.pipeline.phases[0][11] ));
 sg13g2_dfrbp_1 _6458_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net28),
    .D(_0232_),
    .Q_N(_0032_),
    .Q(\dtop.vtop.pipeline.phases[0][12] ));
 sg13g2_dfrbp_1 _6459_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net27),
    .D(_0233_),
    .Q_N(_0033_),
    .Q(\dtop.vtop.pipeline.phases[0][13] ));
 sg13g2_dfrbp_1 _6460_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net26),
    .D(_0234_),
    .Q_N(_0035_),
    .Q(\dtop.vtop.pipeline.phases[0][14] ));
 sg13g2_dfrbp_1 _6461_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net25),
    .D(_0235_),
    .Q_N(_0002_),
    .Q(\dtop.vtop.pipeline.phases[0][15] ));
 sg13g2_dfrbp_1 _6462_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net24),
    .D(_0236_),
    .Q_N(_3074_),
    .Q(\dtop.vtop.pipeline.zg_acc[0] ));
 sg13g2_dfrbp_1 _6463_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net23),
    .D(_0237_),
    .Q_N(_0025_),
    .Q(\dtop.vtop.pipeline.zg_acc[1] ));
 sg13g2_dfrbp_1 _6464_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net22),
    .D(_0238_),
    .Q_N(_3073_),
    .Q(\dtop.vtop.pipeline.zg_acc[2] ));
 sg13g2_dfrbp_1 _6465_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net21),
    .D(_0239_),
    .Q_N(_3072_),
    .Q(\dtop.vtop.pipeline.zg_acc[3] ));
 sg13g2_dfrbp_1 _6466_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net20),
    .D(_0240_),
    .Q_N(_3071_),
    .Q(\dtop.vtop.pipeline.zg_acc[4] ));
 sg13g2_dfrbp_1 _6467_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net304),
    .D(_0241_),
    .Q_N(_3070_),
    .Q(\dtop.vtop.pipeline.zg_acc[5] ));
 sg13g2_dfrbp_1 _6468_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net303),
    .D(_0242_),
    .Q_N(_0034_),
    .Q(\dtop.vtop.pipeline.zg_acc[6] ));
 sg13g2_dfrbp_1 _6469_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net302),
    .D(_0243_),
    .Q_N(_0036_),
    .Q(\dtop.vtop.pipeline.zg_acc[7] ));
 sg13g2_dfrbp_1 _6470_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net301),
    .D(_0244_),
    .Q_N(_0038_),
    .Q(\dtop.vtop.pipeline.zg_acc[8] ));
 sg13g2_dfrbp_1 _6471_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net300),
    .D(_0245_),
    .Q_N(_3069_),
    .Q(\dtop.vtop.pipeline.zg_acc[9] ));
 sg13g2_dfrbp_1 _6472_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net299),
    .D(_0246_),
    .Q_N(_0062_),
    .Q(\dtop.vtop.pipeline.zg_valid ));
 sg13g2_dfrbp_1 _6473_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net297),
    .D(_0247_),
    .Q_N(_3068_),
    .Q(\dtop.vtop.pipeline.zg[0] ));
 sg13g2_dfrbp_1 _6474_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net296),
    .D(_0248_),
    .Q_N(_3067_),
    .Q(\dtop.vtop.pipeline.zg[1] ));
 sg13g2_dfrbp_1 _6475_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net295),
    .D(_0249_),
    .Q_N(_3066_),
    .Q(\dtop.vtop.pipeline.zg[2] ));
 sg13g2_dfrbp_1 _6476_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net294),
    .D(_0250_),
    .Q_N(_3065_),
    .Q(\dtop.vtop.pipeline.zg[3] ));
 sg13g2_dfrbp_1 _6477_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net293),
    .D(_0251_),
    .Q_N(_3064_),
    .Q(\dtop.vtop.pipeline.zg[4] ));
 sg13g2_dfrbp_1 _6478_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net292),
    .D(_0252_),
    .Q_N(_3063_),
    .Q(\dtop.vtop.pipeline.zg[5] ));
 sg13g2_dfrbp_1 _6479_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net291),
    .D(_0253_),
    .Q_N(_3062_),
    .Q(\dtop.vtop.pipeline.zg[6] ));
 sg13g2_dfrbp_1 _6480_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net290),
    .D(_0254_),
    .Q_N(_3061_),
    .Q(\dtop.vtop.pipeline.zg[7] ));
 sg13g2_dfrbp_1 _6481_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net289),
    .D(_0255_),
    .Q_N(_3060_),
    .Q(\dtop.vtop.pipeline.zg[8] ));
 sg13g2_dfrbp_1 _6482_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net288),
    .D(_0256_),
    .Q_N(_3059_),
    .Q(\dtop.vtop.pipeline.zg[9] ));
 sg13g2_dfrbp_1 _6483_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net287),
    .D(_0257_),
    .Q_N(_3058_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[0] ));
 sg13g2_dfrbp_1 _6484_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net286),
    .D(_0258_),
    .Q_N(_3057_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[1] ));
 sg13g2_dfrbp_1 _6485_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net285),
    .D(_0259_),
    .Q_N(_3056_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[2] ));
 sg13g2_dfrbp_1 _6486_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net284),
    .D(_0260_),
    .Q_N(_3055_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[3] ));
 sg13g2_dfrbp_1 _6487_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net283),
    .D(_0261_),
    .Q_N(_3054_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[4] ));
 sg13g2_dfrbp_1 _6488_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net282),
    .D(_0262_),
    .Q_N(_3053_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[5] ));
 sg13g2_dfrbp_1 _6489_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net281),
    .D(_0263_),
    .Q_N(_3052_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[6] ));
 sg13g2_dfrbp_1 _6490_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net280),
    .D(_0264_),
    .Q_N(_3051_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[7] ));
 sg13g2_dfrbp_1 _6491_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net279),
    .D(_0265_),
    .Q_N(_3050_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[8] ));
 sg13g2_dfrbp_1 _6492_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net278),
    .D(_0266_),
    .Q_N(_0003_),
    .Q(\dtop.vtop.pipeline.wave_index[0] ));
 sg13g2_dfrbp_1 _6493_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net277),
    .D(_0267_),
    .Q_N(_0004_),
    .Q(\dtop.vtop.pipeline.wave_index[1] ));
 sg13g2_dfrbp_1 _6494_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net276),
    .D(_0268_),
    .Q_N(_3049_),
    .Q(\dtop.vtop.pipeline.nstep[0] ));
 sg13g2_dfrbp_1 _6495_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net275),
    .D(_0269_),
    .Q_N(_0008_),
    .Q(\dtop.vtop.pipeline.nstep[1] ));
 sg13g2_dfrbp_1 _6496_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net274),
    .D(net307),
    .Q_N(\dtop.vtop.pipeline.next_nstep_counter[0] ),
    .Q(\dtop.vtop.pipeline.nstep_counter[0] ));
 sg13g2_dfrbp_1 _6497_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net272),
    .D(net539),
    .Q_N(_3048_),
    .Q(\dtop.vtop.pipeline.nstep_counter[1] ));
 sg13g2_dfrbp_1 _6498_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net270),
    .D(_0272_),
    .Q_N(_3047_),
    .Q(\dtop.vtop.pipeline.nstep_counter[2] ));
 sg13g2_dfrbp_1 _6499_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net268),
    .D(net486),
    .Q_N(_3046_),
    .Q(\dtop.vtop.pipeline.nstep_counter[3] ));
 sg13g2_dfrbp_1 _6500_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net266),
    .D(_0274_),
    .Q_N(_3045_),
    .Q(\dtop.vtop.pipeline.nstep_counter[4] ));
 sg13g2_dfrbp_1 _6501_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net264),
    .D(_0275_),
    .Q_N(_3044_),
    .Q(\dtop.vtop.color[4] ));
 sg13g2_dfrbp_1 _6502_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net263),
    .D(_0276_),
    .Q_N(_0005_),
    .Q(\dtop.vtop.color[5] ));
 sg13g2_dfrbp_1 _6503_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net262),
    .D(_0277_),
    .Q_N(_0006_),
    .Q(\dtop.vtop.color[6] ));
 sg13g2_dfrbp_1 _6504_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net261),
    .D(_0278_),
    .Q_N(_3043_),
    .Q(\dtop.vtop.color[7] ));
 sg13g2_dfrbp_1 _6505_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net260),
    .D(net430),
    .Q_N(_3042_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _6506_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net258),
    .D(net462),
    .Q_N(_3041_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _6507_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net256),
    .D(net474),
    .Q_N(_3040_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _6508_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net254),
    .D(net470),
    .Q_N(_3039_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _6509_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net252),
    .D(_0283_),
    .Q_N(_0056_),
    .Q(\dtop.oct_counter[0] ));
 sg13g2_dfrbp_1 _6510_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net251),
    .D(net619),
    .Q_N(_0055_),
    .Q(\dtop.oct_counter[1] ));
 sg13g2_dfrbp_1 _6511_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net250),
    .D(net606),
    .Q_N(_0049_),
    .Q(\dtop.oct_counter[2] ));
 sg13g2_dfrbp_1 _6512_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net249),
    .D(_0286_),
    .Q_N(_3038_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _6513_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net247),
    .D(_0287_),
    .Q_N(_3037_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _6514_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net245),
    .D(net472),
    .Q_N(_3036_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _6515_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net244),
    .D(_0289_),
    .Q_N(_3035_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _6516_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net243),
    .D(_0290_),
    .Q_N(_0054_),
    .Q(\dtop.oct_counter[3] ));
 sg13g2_dfrbp_1 _6517_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net242),
    .D(_0291_),
    .Q_N(_0053_),
    .Q(\dtop.oct_counter[4] ));
 sg13g2_dfrbp_1 _6518_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net241),
    .D(_0292_),
    .Q_N(_3034_),
    .Q(\dtop.oct_counter[5] ));
 sg13g2_dfrbp_1 _6519_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net240),
    .D(_0293_),
    .Q_N(_3033_),
    .Q(\dtop.oct_counter[6] ));
 sg13g2_dfrbp_1 _6520_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net239),
    .D(_0294_),
    .Q_N(_0086_),
    .Q(\dtop.vtop.logo.addr[5] ));
 sg13g2_dfrbp_1 _6521_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net238),
    .D(_0295_),
    .Q_N(_3032_),
    .Q(\dtop.vtop.logo.addr[6] ));
 sg13g2_dfrbp_1 _6522_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net237),
    .D(_0296_),
    .Q_N(_0085_),
    .Q(\dtop.vtop.logo.addr[7] ));
 sg13g2_dfrbp_1 _6523_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net236),
    .D(_0297_),
    .Q_N(_0084_),
    .Q(\dtop.vtop.logo.addr[8] ));
 sg13g2_dfrbp_1 _6524_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net235),
    .D(_0298_),
    .Q_N(_0052_),
    .Q(\dtop.vtop.logo.addr[9] ));
 sg13g2_dfrbp_1 _6525_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net234),
    .D(_0299_),
    .Q_N(_3031_),
    .Q(\dtop.player_inst.synth.alu.acc[0] ));
 sg13g2_dfrbp_1 _6526_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net232),
    .D(_0300_),
    .Q_N(_3030_),
    .Q(\dtop.player_inst.synth.alu.acc[1] ));
 sg13g2_dfrbp_1 _6527_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net230),
    .D(_0301_),
    .Q_N(_3029_),
    .Q(\dtop.player_inst.synth.alu.acc[2] ));
 sg13g2_dfrbp_1 _6528_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net228),
    .D(_0302_),
    .Q_N(_3028_),
    .Q(\dtop.player_inst.synth.alu.acc[3] ));
 sg13g2_dfrbp_1 _6529_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net226),
    .D(_0303_),
    .Q_N(_3027_),
    .Q(\dtop.player_inst.synth.alu.acc[4] ));
 sg13g2_dfrbp_1 _6530_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net224),
    .D(_0304_),
    .Q_N(_3026_),
    .Q(\dtop.player_inst.synth.alu.acc[5] ));
 sg13g2_dfrbp_1 _6531_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net222),
    .D(_0305_),
    .Q_N(_3025_),
    .Q(\dtop.player_inst.synth.alu.acc[6] ));
 sg13g2_dfrbp_1 _6532_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net220),
    .D(_0306_),
    .Q_N(_3024_),
    .Q(\dtop.player_inst.synth.alu.acc[7] ));
 sg13g2_dfrbp_1 _6533_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net218),
    .D(_0307_),
    .Q_N(_3023_),
    .Q(\dtop.player_inst.synth.alu.acc[8] ));
 sg13g2_dfrbp_1 _6534_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net216),
    .D(_0308_),
    .Q_N(_3022_),
    .Q(\dtop.player_inst.synth.alu.acc[9] ));
 sg13g2_dfrbp_1 _6535_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net214),
    .D(_0309_),
    .Q_N(_0037_),
    .Q(\dtop.player_inst.synth.alu.acc[10] ));
 sg13g2_dfrbp_1 _6536_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net212),
    .D(net374),
    .Q_N(_3021_),
    .Q(\dtop.out_sample[0] ));
 sg13g2_dfrbp_1 _6537_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net210),
    .D(net501),
    .Q_N(_3020_),
    .Q(\dtop.out_sample[1] ));
 sg13g2_dfrbp_1 _6538_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net208),
    .D(_0312_),
    .Q_N(_3019_),
    .Q(\dtop.out_sample[2] ));
 sg13g2_dfrbp_1 _6539_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net206),
    .D(_0313_),
    .Q_N(_3018_),
    .Q(\dtop.out_sample[3] ));
 sg13g2_dfrbp_1 _6540_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net140),
    .D(net396),
    .Q_N(_3017_),
    .Q(\dtop.out_sample[4] ));
 sg13g2_dfrbp_1 _6541_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net136),
    .D(net446),
    .Q_N(_3016_),
    .Q(\dtop.out_sample[5] ));
 sg13g2_dfrbp_1 _6542_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net132),
    .D(_0316_),
    .Q_N(_3015_),
    .Q(\dtop.out_sample[6] ));
 sg13g2_dfrbp_1 _6543_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net128),
    .D(net508),
    .Q_N(_3014_),
    .Q(\dtop.player_inst.synth.alu.registers[0][0] ));
 sg13g2_dfrbp_1 _6544_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net124),
    .D(net530),
    .Q_N(_3013_),
    .Q(\dtop.player_inst.synth.alu.registers[0][1] ));
 sg13g2_dfrbp_1 _6545_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net120),
    .D(_0319_),
    .Q_N(_3012_),
    .Q(\dtop.player_inst.synth.alu.registers[0][2] ));
 sg13g2_dfrbp_1 _6546_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net116),
    .D(_0320_),
    .Q_N(_3011_),
    .Q(\dtop.player_inst.synth.alu.registers[0][3] ));
 sg13g2_dfrbp_1 _6547_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net112),
    .D(_0321_),
    .Q_N(_3010_),
    .Q(\dtop.player_inst.synth.alu.registers[0][4] ));
 sg13g2_dfrbp_1 _6548_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net108),
    .D(_0322_),
    .Q_N(_3009_),
    .Q(\dtop.player_inst.synth.alu.registers[0][5] ));
 sg13g2_dfrbp_1 _6549_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net104),
    .D(_0323_),
    .Q_N(_3008_),
    .Q(\dtop.player_inst.synth.alu.registers[0][6] ));
 sg13g2_dfrbp_1 _6550_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net100),
    .D(net535),
    .Q_N(_3007_),
    .Q(\dtop.player_inst.synth.alu.registers[0][7] ));
 sg13g2_dfrbp_1 _6551_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net96),
    .D(net515),
    .Q_N(_3006_),
    .Q(\dtop.player_inst.synth.alu.registers[0][8] ));
 sg13g2_dfrbp_1 _6552_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net92),
    .D(_0326_),
    .Q_N(_3005_),
    .Q(\dtop.player_inst.synth.alu.registers[0][9] ));
 sg13g2_dfrbp_1 _6553_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net88),
    .D(net526),
    .Q_N(_3004_),
    .Q(\dtop.player_inst.synth.alu.registers[0][10] ));
 sg13g2_dfrbp_1 _6554_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net84),
    .D(_0328_),
    .Q_N(_3003_),
    .Q(\dtop.player_inst.synth.alu.registers[1][0] ));
 sg13g2_dfrbp_1 _6555_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net80),
    .D(net345),
    .Q_N(_3002_),
    .Q(\dtop.player_inst.synth.alu.registers[1][1] ));
 sg13g2_dfrbp_1 _6556_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net76),
    .D(_0330_),
    .Q_N(_3001_),
    .Q(\dtop.player_inst.synth.alu.registers[1][2] ));
 sg13g2_dfrbp_1 _6557_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net298),
    .D(_0331_),
    .Q_N(_3000_),
    .Q(\dtop.player_inst.synth.alu.registers[1][3] ));
 sg13g2_dfrbp_1 _6558_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net271),
    .D(_0332_),
    .Q_N(_2999_),
    .Q(\dtop.player_inst.synth.alu.registers[1][4] ));
 sg13g2_dfrbp_1 _6559_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net267),
    .D(_0333_),
    .Q_N(_2998_),
    .Q(\dtop.player_inst.synth.alu.registers[1][5] ));
 sg13g2_dfrbp_1 _6560_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net259),
    .D(_0334_),
    .Q_N(_2997_),
    .Q(\dtop.player_inst.synth.alu.registers[1][6] ));
 sg13g2_dfrbp_1 _6561_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net255),
    .D(net378),
    .Q_N(_2996_),
    .Q(\dtop.player_inst.synth.alu.registers[1][7] ));
 sg13g2_dfrbp_1 _6562_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net248),
    .D(net393),
    .Q_N(_2995_),
    .Q(\dtop.player_inst.synth.alu.registers[1][8] ));
 sg13g2_dfrbp_1 _6563_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net233),
    .D(_0337_),
    .Q_N(_2994_),
    .Q(\dtop.player_inst.synth.alu.registers[1][9] ));
 sg13g2_dfrbp_1 _6564_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net229),
    .D(net419),
    .Q_N(_2993_),
    .Q(\dtop.player_inst.synth.alu.registers[1][10] ));
 sg13g2_dfrbp_1 _6565_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net225),
    .D(_0339_),
    .Q_N(_2992_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _6566_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net223),
    .D(net369),
    .Q_N(_2991_),
    .Q(\dtop.player_inst.synth.alu.registers[2][0] ));
 sg13g2_dfrbp_1 _6567_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net219),
    .D(net332),
    .Q_N(_2990_),
    .Q(\dtop.player_inst.synth.alu.registers[2][1] ));
 sg13g2_dfrbp_1 _6568_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net215),
    .D(_0342_),
    .Q_N(_2989_),
    .Q(\dtop.player_inst.synth.alu.registers[2][2] ));
 sg13g2_dfrbp_1 _6569_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net211),
    .D(_0343_),
    .Q_N(_2988_),
    .Q(\dtop.player_inst.synth.alu.registers[2][3] ));
 sg13g2_dfrbp_1 _6570_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net207),
    .D(_0344_),
    .Q_N(_2987_),
    .Q(\dtop.player_inst.synth.alu.registers[2][4] ));
 sg13g2_dfrbp_1 _6571_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net138),
    .D(_0345_),
    .Q_N(_2986_),
    .Q(\dtop.player_inst.synth.alu.registers[2][5] ));
 sg13g2_dfrbp_1 _6572_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net130),
    .D(_0346_),
    .Q_N(_2985_),
    .Q(\dtop.player_inst.synth.alu.registers[2][6] ));
 sg13g2_dfrbp_1 _6573_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net122),
    .D(net384),
    .Q_N(_2984_),
    .Q(\dtop.player_inst.synth.alu.registers[2][7] ));
 sg13g2_dfrbp_1 _6574_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net114),
    .D(net448),
    .Q_N(_2983_),
    .Q(\dtop.player_inst.synth.alu.registers[4][0] ));
 sg13g2_dfrbp_1 _6575_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net106),
    .D(net350),
    .Q_N(_2982_),
    .Q(\dtop.player_inst.synth.alu.registers[4][1] ));
 sg13g2_dfrbp_1 _6576_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net98),
    .D(_0350_),
    .Q_N(_2981_),
    .Q(\dtop.player_inst.synth.alu.registers[4][2] ));
 sg13g2_dfrbp_1 _6577_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net90),
    .D(_0351_),
    .Q_N(_2980_),
    .Q(\dtop.player_inst.synth.alu.registers[4][3] ));
 sg13g2_dfrbp_1 _6578_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net82),
    .D(net451),
    .Q_N(_2979_),
    .Q(\dtop.player_inst.synth.alu.registers[4][4] ));
 sg13g2_dfrbp_1 _6579_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net74),
    .D(net355),
    .Q_N(_2978_),
    .Q(\dtop.player_inst.synth.alu.registers[4][5] ));
 sg13g2_dfrbp_1 _6580_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net269),
    .D(net318),
    .Q_N(_0044_),
    .Q(\dtop.player_inst.synth.alu.registers[4][6] ));
 sg13g2_dfrbp_1 _6581_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net257),
    .D(net325),
    .Q_N(_0045_),
    .Q(\dtop.player_inst.synth.alu.registers[4][7] ));
 sg13g2_dfrbp_1 _6582_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net246),
    .D(net314),
    .Q_N(_0046_),
    .Q(\dtop.player_inst.synth.alu.registers[4][8] ));
 sg13g2_dfrbp_1 _6583_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net227),
    .D(_0357_),
    .Q_N(_0047_),
    .Q(\dtop.player_inst.synth.alu.registers[4][9] ));
 sg13g2_dfrbp_1 _6584_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net217),
    .D(net340),
    .Q_N(_0048_),
    .Q(\dtop.player_inst.synth.alu.registers[4][10] ));
 sg13g2_dfrbp_1 _6585_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net209),
    .D(_0359_),
    .Q_N(_2977_),
    .Q(\dtop.player_inst.synth.alu.registers[3][0] ));
 sg13g2_dfrbp_1 _6586_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net134),
    .D(net365),
    .Q_N(_2976_),
    .Q(\dtop.player_inst.synth.alu.registers[3][1] ));
 sg13g2_dfrbp_1 _6587_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net118),
    .D(_0361_),
    .Q_N(_2975_),
    .Q(\dtop.player_inst.synth.alu.registers[3][2] ));
 sg13g2_dfrbp_1 _6588_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net102),
    .D(_0362_),
    .Q_N(_2974_),
    .Q(\dtop.player_inst.synth.alu.registers[3][3] ));
 sg13g2_dfrbp_1 _6589_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net86),
    .D(net376),
    .Q_N(_2973_),
    .Q(\dtop.player_inst.synth.alu.registers[3][4] ));
 sg13g2_dfrbp_1 _6590_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net273),
    .D(_0364_),
    .Q_N(_2972_),
    .Q(\dtop.player_inst.synth.alu.registers[3][5] ));
 sg13g2_dfrbp_1 _6591_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net253),
    .D(_0365_),
    .Q_N(_2971_),
    .Q(\dtop.player_inst.synth.alu.registers[3][6] ));
 sg13g2_dfrbp_1 _6592_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net221),
    .D(net362),
    .Q_N(_2970_),
    .Q(\dtop.player_inst.synth.alu.registers[3][7] ));
 sg13g2_dfrbp_1 _6593_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net205),
    .D(_0367_),
    .Q_N(_2969_),
    .Q(\dtop.player_inst.synth.alu.registers[5][0] ));
 sg13g2_dfrbp_1 _6594_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net110),
    .D(net337),
    .Q_N(_2968_),
    .Q(\dtop.player_inst.synth.alu.registers[5][1] ));
 sg13g2_dfrbp_1 _6595_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net78),
    .D(_0369_),
    .Q_N(_2967_),
    .Q(\dtop.player_inst.synth.alu.registers[5][2] ));
 sg13g2_dfrbp_1 _6596_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net231),
    .D(_0370_),
    .Q_N(_2966_),
    .Q(\dtop.player_inst.synth.alu.registers[5][3] ));
 sg13g2_dfrbp_1 _6597_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net126),
    .D(net357),
    .Q_N(_2965_),
    .Q(\dtop.player_inst.synth.alu.registers[5][4] ));
 sg13g2_dfrbp_1 _6598_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net265),
    .D(_0372_),
    .Q_N(_2964_),
    .Q(\dtop.player_inst.synth.alu.registers[5][5] ));
 sg13g2_dfrbp_1 _6599_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net94),
    .D(_0373_),
    .Q_N(_2963_),
    .Q(\dtop.player_inst.synth.alu.registers[5][6] ));
 sg13g2_tiehi _6465__21 (.L_HI(net21));
 sg13g2_tiehi _6464__22 (.L_HI(net22));
 sg13g2_tiehi _6463__23 (.L_HI(net23));
 sg13g2_tiehi _6462__24 (.L_HI(net24));
 sg13g2_tiehi _6461__25 (.L_HI(net25));
 sg13g2_tiehi _6460__26 (.L_HI(net26));
 sg13g2_tiehi _6459__27 (.L_HI(net27));
 sg13g2_tiehi _6458__28 (.L_HI(net28));
 sg13g2_tiehi _6457__29 (.L_HI(net29));
 sg13g2_tiehi _6456__30 (.L_HI(net30));
 sg13g2_tiehi _6455__31 (.L_HI(net31));
 sg13g2_tiehi _6454__32 (.L_HI(net32));
 sg13g2_tiehi _6453__33 (.L_HI(net33));
 sg13g2_tiehi _6452__34 (.L_HI(net34));
 sg13g2_tiehi _6451__35 (.L_HI(net35));
 sg13g2_tiehi _6450__36 (.L_HI(net36));
 sg13g2_tiehi _6449__37 (.L_HI(net37));
 sg13g2_tiehi _6448__38 (.L_HI(net38));
 sg13g2_tiehi _6447__39 (.L_HI(net39));
 sg13g2_tiehi _6446__40 (.L_HI(net40));
 sg13g2_tiehi _6445__41 (.L_HI(net41));
 sg13g2_tiehi _6444__42 (.L_HI(net42));
 sg13g2_tiehi _6443__43 (.L_HI(net43));
 sg13g2_tiehi _6442__44 (.L_HI(net44));
 sg13g2_tiehi _6441__45 (.L_HI(net45));
 sg13g2_tiehi _6440__46 (.L_HI(net46));
 sg13g2_tiehi _6439__47 (.L_HI(net47));
 sg13g2_tiehi _6438__48 (.L_HI(net48));
 sg13g2_tiehi _6437__49 (.L_HI(net49));
 sg13g2_tiehi _6436__50 (.L_HI(net50));
 sg13g2_tiehi _6435__51 (.L_HI(net51));
 sg13g2_tiehi _6434__52 (.L_HI(net52));
 sg13g2_tiehi _6433__53 (.L_HI(net53));
 sg13g2_tiehi _6432__54 (.L_HI(net54));
 sg13g2_tiehi _6431__55 (.L_HI(net55));
 sg13g2_tiehi _6430__56 (.L_HI(net56));
 sg13g2_tiehi _6429__57 (.L_HI(net57));
 sg13g2_tiehi _6428__58 (.L_HI(net58));
 sg13g2_tiehi _6427__59 (.L_HI(net59));
 sg13g2_tiehi _6426__60 (.L_HI(net60));
 sg13g2_tiehi _6425__61 (.L_HI(net61));
 sg13g2_tiehi _6424__62 (.L_HI(net62));
 sg13g2_tiehi _6423__63 (.L_HI(net63));
 sg13g2_tiehi _6422__64 (.L_HI(net64));
 sg13g2_tiehi _6421__65 (.L_HI(net65));
 sg13g2_tiehi _6420__66 (.L_HI(net66));
 sg13g2_tiehi _6419__67 (.L_HI(net67));
 sg13g2_tiehi _6418__68 (.L_HI(net68));
 sg13g2_tiehi _6417__69 (.L_HI(net69));
 sg13g2_tiehi _6416__70 (.L_HI(net70));
 sg13g2_tiehi _6415__71 (.L_HI(net71));
 sg13g2_tiehi _6414__72 (.L_HI(net72));
 sg13g2_tiehi _6413__73 (.L_HI(net73));
 sg13g2_tiehi _6579__74 (.L_HI(net74));
 sg13g2_tiehi _6412__75 (.L_HI(net75));
 sg13g2_tiehi _6556__76 (.L_HI(net76));
 sg13g2_tiehi _6411__77 (.L_HI(net77));
 sg13g2_tiehi _6595__78 (.L_HI(net78));
 sg13g2_tiehi _6410__79 (.L_HI(net79));
 sg13g2_tiehi _6555__80 (.L_HI(net80));
 sg13g2_tiehi _6409__81 (.L_HI(net81));
 sg13g2_tiehi _6578__82 (.L_HI(net82));
 sg13g2_tiehi _6408__83 (.L_HI(net83));
 sg13g2_tiehi _6554__84 (.L_HI(net84));
 sg13g2_tiehi _6407__85 (.L_HI(net85));
 sg13g2_tiehi _6589__86 (.L_HI(net86));
 sg13g2_tiehi _6406__87 (.L_HI(net87));
 sg13g2_tiehi _6553__88 (.L_HI(net88));
 sg13g2_tiehi _6405__89 (.L_HI(net89));
 sg13g2_tiehi _6577__90 (.L_HI(net90));
 sg13g2_tiehi _6404__91 (.L_HI(net91));
 sg13g2_tiehi _6552__92 (.L_HI(net92));
 sg13g2_tiehi _6403__93 (.L_HI(net93));
 sg13g2_tiehi _6599__94 (.L_HI(net94));
 sg13g2_tiehi _6402__95 (.L_HI(net95));
 sg13g2_tiehi _6551__96 (.L_HI(net96));
 sg13g2_tiehi _6401__97 (.L_HI(net97));
 sg13g2_tiehi _6576__98 (.L_HI(net98));
 sg13g2_tiehi _6400__99 (.L_HI(net99));
 sg13g2_tiehi _6550__100 (.L_HI(net100));
 sg13g2_tiehi _6399__101 (.L_HI(net101));
 sg13g2_tiehi _6588__102 (.L_HI(net102));
 sg13g2_tiehi _6398__103 (.L_HI(net103));
 sg13g2_tiehi _6549__104 (.L_HI(net104));
 sg13g2_tiehi _6397__105 (.L_HI(net105));
 sg13g2_tiehi _6575__106 (.L_HI(net106));
 sg13g2_tiehi _6396__107 (.L_HI(net107));
 sg13g2_tiehi _6548__108 (.L_HI(net108));
 sg13g2_tiehi _6395__109 (.L_HI(net109));
 sg13g2_tiehi _6594__110 (.L_HI(net110));
 sg13g2_tiehi _6394__111 (.L_HI(net111));
 sg13g2_tiehi _6547__112 (.L_HI(net112));
 sg13g2_tiehi _6393__113 (.L_HI(net113));
 sg13g2_tiehi _6574__114 (.L_HI(net114));
 sg13g2_tiehi _6392__115 (.L_HI(net115));
 sg13g2_tiehi _6546__116 (.L_HI(net116));
 sg13g2_tiehi _6391__117 (.L_HI(net117));
 sg13g2_tiehi _6587__118 (.L_HI(net118));
 sg13g2_tiehi _6390__119 (.L_HI(net119));
 sg13g2_tiehi _6545__120 (.L_HI(net120));
 sg13g2_tiehi _6389__121 (.L_HI(net121));
 sg13g2_tiehi _6573__122 (.L_HI(net122));
 sg13g2_tiehi _6388__123 (.L_HI(net123));
 sg13g2_tiehi _6544__124 (.L_HI(net124));
 sg13g2_tiehi _6387__125 (.L_HI(net125));
 sg13g2_tiehi _6597__126 (.L_HI(net126));
 sg13g2_tiehi _6386__127 (.L_HI(net127));
 sg13g2_tiehi _6543__128 (.L_HI(net128));
 sg13g2_tiehi _6385__129 (.L_HI(net129));
 sg13g2_tiehi _6572__130 (.L_HI(net130));
 sg13g2_tiehi _6384__131 (.L_HI(net131));
 sg13g2_tiehi _6542__132 (.L_HI(net132));
 sg13g2_tiehi _6383__133 (.L_HI(net133));
 sg13g2_tiehi _6586__134 (.L_HI(net134));
 sg13g2_tiehi _6382__135 (.L_HI(net135));
 sg13g2_tiehi _6541__136 (.L_HI(net136));
 sg13g2_tiehi _6381__137 (.L_HI(net137));
 sg13g2_tiehi _6571__138 (.L_HI(net138));
 sg13g2_tiehi _6380__139 (.L_HI(net139));
 sg13g2_tiehi _6540__140 (.L_HI(net140));
 sg13g2_tiehi _6379__141 (.L_HI(net141));
 sg13g2_tiehi _6378__142 (.L_HI(net142));
 sg13g2_tiehi _6377__143 (.L_HI(net143));
 sg13g2_tiehi _6376__144 (.L_HI(net144));
 sg13g2_tiehi _6375__145 (.L_HI(net145));
 sg13g2_tiehi _6374__146 (.L_HI(net146));
 sg13g2_tiehi _6373__147 (.L_HI(net147));
 sg13g2_tiehi _6372__148 (.L_HI(net148));
 sg13g2_tiehi _6371__149 (.L_HI(net149));
 sg13g2_tiehi _6370__150 (.L_HI(net150));
 sg13g2_tiehi _6369__151 (.L_HI(net151));
 sg13g2_tiehi _6368__152 (.L_HI(net152));
 sg13g2_tiehi _6367__153 (.L_HI(net153));
 sg13g2_tiehi _6366__154 (.L_HI(net154));
 sg13g2_tiehi _6365__155 (.L_HI(net155));
 sg13g2_tiehi _6364__156 (.L_HI(net156));
 sg13g2_tiehi _6363__157 (.L_HI(net157));
 sg13g2_tiehi _6362__158 (.L_HI(net158));
 sg13g2_tiehi _6361__159 (.L_HI(net159));
 sg13g2_tiehi _6360__160 (.L_HI(net160));
 sg13g2_tiehi _6359__161 (.L_HI(net161));
 sg13g2_tiehi _6358__162 (.L_HI(net162));
 sg13g2_tiehi _6357__163 (.L_HI(net163));
 sg13g2_tiehi _6356__164 (.L_HI(net164));
 sg13g2_tiehi _6355__165 (.L_HI(net165));
 sg13g2_tiehi _6354__166 (.L_HI(net166));
 sg13g2_tiehi _6353__167 (.L_HI(net167));
 sg13g2_tiehi _6352__168 (.L_HI(net168));
 sg13g2_tiehi _6351__169 (.L_HI(net169));
 sg13g2_tiehi _6350__170 (.L_HI(net170));
 sg13g2_tiehi _6349__171 (.L_HI(net171));
 sg13g2_tiehi _6348__172 (.L_HI(net172));
 sg13g2_tiehi _6347__173 (.L_HI(net173));
 sg13g2_tiehi _6346__174 (.L_HI(net174));
 sg13g2_tiehi _6345__175 (.L_HI(net175));
 sg13g2_tiehi _6344__176 (.L_HI(net176));
 sg13g2_tiehi _6343__177 (.L_HI(net177));
 sg13g2_tiehi _6342__178 (.L_HI(net178));
 sg13g2_tiehi _6341__179 (.L_HI(net179));
 sg13g2_tiehi _6340__180 (.L_HI(net180));
 sg13g2_tiehi _6339__181 (.L_HI(net181));
 sg13g2_tiehi _6338__182 (.L_HI(net182));
 sg13g2_tiehi _6337__183 (.L_HI(net183));
 sg13g2_tiehi _6336__184 (.L_HI(net184));
 sg13g2_tiehi _6335__185 (.L_HI(net185));
 sg13g2_tiehi _6334__186 (.L_HI(net186));
 sg13g2_tiehi _6333__187 (.L_HI(net187));
 sg13g2_tiehi _6332__188 (.L_HI(net188));
 sg13g2_tiehi _6331__189 (.L_HI(net189));
 sg13g2_tiehi _6330__190 (.L_HI(net190));
 sg13g2_tiehi _6329__191 (.L_HI(net191));
 sg13g2_tiehi _6328__192 (.L_HI(net192));
 sg13g2_tiehi _6327__193 (.L_HI(net193));
 sg13g2_tiehi _6326__194 (.L_HI(net194));
 sg13g2_tiehi _6325__195 (.L_HI(net195));
 sg13g2_tiehi _6324__196 (.L_HI(net196));
 sg13g2_tiehi _6323__197 (.L_HI(net197));
 sg13g2_tiehi _6322__198 (.L_HI(net198));
 sg13g2_tiehi _6321__199 (.L_HI(net199));
 sg13g2_tiehi _6320__200 (.L_HI(net200));
 sg13g2_tiehi _6319__201 (.L_HI(net201));
 sg13g2_tiehi _6318__202 (.L_HI(net202));
 sg13g2_tiehi _6317__203 (.L_HI(net203));
 sg13g2_tiehi _6316__204 (.L_HI(net204));
 sg13g2_tiehi _6593__205 (.L_HI(net205));
 sg13g2_tiehi _6539__206 (.L_HI(net206));
 sg13g2_tiehi _6570__207 (.L_HI(net207));
 sg13g2_tiehi _6538__208 (.L_HI(net208));
 sg13g2_tiehi _6585__209 (.L_HI(net209));
 sg13g2_tiehi _6537__210 (.L_HI(net210));
 sg13g2_tiehi _6569__211 (.L_HI(net211));
 sg13g2_tiehi _6536__212 (.L_HI(net212));
 sg13g2_tiehi _6315__213 (.L_HI(net213));
 sg13g2_tiehi _6535__214 (.L_HI(net214));
 sg13g2_tiehi _6568__215 (.L_HI(net215));
 sg13g2_tiehi _6534__216 (.L_HI(net216));
 sg13g2_tiehi _6584__217 (.L_HI(net217));
 sg13g2_tiehi _6533__218 (.L_HI(net218));
 sg13g2_tiehi _6567__219 (.L_HI(net219));
 sg13g2_tiehi _6532__220 (.L_HI(net220));
 sg13g2_tiehi _6592__221 (.L_HI(net221));
 sg13g2_tiehi _6531__222 (.L_HI(net222));
 sg13g2_tiehi _6566__223 (.L_HI(net223));
 sg13g2_tiehi _6530__224 (.L_HI(net224));
 sg13g2_tiehi _6565__225 (.L_HI(net225));
 sg13g2_tiehi _6529__226 (.L_HI(net226));
 sg13g2_tiehi _6583__227 (.L_HI(net227));
 sg13g2_tiehi _6528__228 (.L_HI(net228));
 sg13g2_tiehi _6564__229 (.L_HI(net229));
 sg13g2_tiehi _6527__230 (.L_HI(net230));
 sg13g2_tiehi _6596__231 (.L_HI(net231));
 sg13g2_tiehi _6526__232 (.L_HI(net232));
 sg13g2_tiehi _6563__233 (.L_HI(net233));
 sg13g2_tiehi _6525__234 (.L_HI(net234));
 sg13g2_tiehi _6524__235 (.L_HI(net235));
 sg13g2_tiehi _6523__236 (.L_HI(net236));
 sg13g2_tiehi _6522__237 (.L_HI(net237));
 sg13g2_tiehi _6521__238 (.L_HI(net238));
 sg13g2_tiehi _6520__239 (.L_HI(net239));
 sg13g2_tiehi _6519__240 (.L_HI(net240));
 sg13g2_tiehi _6518__241 (.L_HI(net241));
 sg13g2_tiehi _6517__242 (.L_HI(net242));
 sg13g2_tiehi _6516__243 (.L_HI(net243));
 sg13g2_tiehi _6515__244 (.L_HI(net244));
 sg13g2_tiehi _6514__245 (.L_HI(net245));
 sg13g2_tiehi _6582__246 (.L_HI(net246));
 sg13g2_tiehi _6513__247 (.L_HI(net247));
 sg13g2_tiehi _6562__248 (.L_HI(net248));
 sg13g2_tiehi _6512__249 (.L_HI(net249));
 sg13g2_tiehi _6511__250 (.L_HI(net250));
 sg13g2_tiehi _6510__251 (.L_HI(net251));
 sg13g2_tiehi _6509__252 (.L_HI(net252));
 sg13g2_tiehi _6591__253 (.L_HI(net253));
 sg13g2_tiehi _6508__254 (.L_HI(net254));
 sg13g2_tiehi _6561__255 (.L_HI(net255));
 sg13g2_tiehi _6507__256 (.L_HI(net256));
 sg13g2_tiehi _6581__257 (.L_HI(net257));
 sg13g2_tiehi _6506__258 (.L_HI(net258));
 sg13g2_tiehi _6560__259 (.L_HI(net259));
 sg13g2_tiehi _6505__260 (.L_HI(net260));
 sg13g2_tiehi _6504__261 (.L_HI(net261));
 sg13g2_tiehi _6503__262 (.L_HI(net262));
 sg13g2_tiehi _6502__263 (.L_HI(net263));
 sg13g2_tiehi _6501__264 (.L_HI(net264));
 sg13g2_tiehi _6598__265 (.L_HI(net265));
 sg13g2_tiehi _6500__266 (.L_HI(net266));
 sg13g2_tiehi _6559__267 (.L_HI(net267));
 sg13g2_tiehi _6499__268 (.L_HI(net268));
 sg13g2_tiehi _6580__269 (.L_HI(net269));
 sg13g2_tiehi _6498__270 (.L_HI(net270));
 sg13g2_tiehi _6558__271 (.L_HI(net271));
 sg13g2_tiehi _6497__272 (.L_HI(net272));
 sg13g2_tiehi _6590__273 (.L_HI(net273));
 sg13g2_tiehi _6496__274 (.L_HI(net274));
 sg13g2_tiehi _6495__275 (.L_HI(net275));
 sg13g2_tiehi _6494__276 (.L_HI(net276));
 sg13g2_tiehi _6493__277 (.L_HI(net277));
 sg13g2_tiehi _6492__278 (.L_HI(net278));
 sg13g2_tiehi _6491__279 (.L_HI(net279));
 sg13g2_tiehi _6490__280 (.L_HI(net280));
 sg13g2_tiehi _6489__281 (.L_HI(net281));
 sg13g2_tiehi _6488__282 (.L_HI(net282));
 sg13g2_tiehi _6487__283 (.L_HI(net283));
 sg13g2_tiehi _6486__284 (.L_HI(net284));
 sg13g2_tiehi _6485__285 (.L_HI(net285));
 sg13g2_tiehi _6484__286 (.L_HI(net286));
 sg13g2_tiehi _6483__287 (.L_HI(net287));
 sg13g2_tiehi _6482__288 (.L_HI(net288));
 sg13g2_tiehi _6481__289 (.L_HI(net289));
 sg13g2_tiehi _6480__290 (.L_HI(net290));
 sg13g2_tiehi _6479__291 (.L_HI(net291));
 sg13g2_tiehi _6478__292 (.L_HI(net292));
 sg13g2_tiehi _6477__293 (.L_HI(net293));
 sg13g2_tiehi _6476__294 (.L_HI(net294));
 sg13g2_tiehi _6475__295 (.L_HI(net295));
 sg13g2_tiehi _6474__296 (.L_HI(net296));
 sg13g2_tiehi _6473__297 (.L_HI(net297));
 sg13g2_tiehi _6557__298 (.L_HI(net298));
 sg13g2_tiehi _6472__299 (.L_HI(net299));
 sg13g2_tiehi _6471__300 (.L_HI(net300));
 sg13g2_tiehi _6470__301 (.L_HI(net301));
 sg13g2_tiehi _6469__302 (.L_HI(net302));
 sg13g2_tiehi _6468__303 (.L_HI(net303));
 sg13g2_tiehi _6467__304 (.L_HI(net304));
 sg13g2_tiehi tt_um_toivoh_demo_tt08_305 (.L_HI(net305));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_toivoh_demo_tt08_7 (.L_LO(net7));
 sg13g2_tielo tt_um_toivoh_demo_tt08_8 (.L_LO(net8));
 sg13g2_tielo tt_um_toivoh_demo_tt08_9 (.L_LO(net9));
 sg13g2_tielo tt_um_toivoh_demo_tt08_10 (.L_LO(net10));
 sg13g2_tielo tt_um_toivoh_demo_tt08_11 (.L_LO(net11));
 sg13g2_tielo tt_um_toivoh_demo_tt08_12 (.L_LO(net12));
 sg13g2_tielo tt_um_toivoh_demo_tt08_13 (.L_LO(net13));
 sg13g2_tielo tt_um_toivoh_demo_tt08_14 (.L_LO(net14));
 sg13g2_tielo tt_um_toivoh_demo_tt08_15 (.L_LO(net15));
 sg13g2_tielo tt_um_toivoh_demo_tt08_16 (.L_LO(net16));
 sg13g2_tielo tt_um_toivoh_demo_tt08_17 (.L_LO(net17));
 sg13g2_tielo tt_um_toivoh_demo_tt08_18 (.L_LO(net18));
 sg13g2_tielo tt_um_toivoh_demo_tt08_19 (.L_LO(net19));
 sg13g2_tiehi _6466__20 (.L_HI(net20));
 sg13g2_buf_2 fanout952 (.A(net953),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_0956_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(net956),
    .X(net954));
 sg13g2_buf_1 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_1623_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_1613_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_1613_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_2228_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(net962),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_2622_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(net964),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_2613_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net968),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(net968),
    .X(net967));
 sg13g2_buf_1 fanout968 (.A(_2601_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(net970),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_2592_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(net972),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(net974),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(net974),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_2579_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(net976),
    .X(net975));
 sg13g2_buf_1 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_2567_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(net979),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_2549_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(net981),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_2521_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_2521_),
    .X(net982));
 sg13g2_buf_4 fanout983 (.X(net983),
    .A(net984));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(_2057_));
 sg13g2_buf_2 fanout985 (.A(net986),
    .X(net985));
 sg13g2_buf_1 fanout986 (.A(net987),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(net988),
    .X(net987));
 sg13g2_buf_4 fanout988 (.X(net988),
    .A(_1571_));
 sg13g2_buf_2 fanout989 (.A(net990),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_1570_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(net993),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(net993),
    .X(net992));
 sg13g2_buf_4 fanout993 (.X(net993),
    .A(_1487_));
 sg13g2_buf_2 fanout994 (.A(_0488_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(net997),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(net997),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_1489_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(net999),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_0495_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_0398_),
    .X(net1000));
 sg13g2_buf_4 fanout1001 (.X(net1001),
    .A(_2931_));
 sg13g2_buf_2 fanout1002 (.A(_1574_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_1574_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(net1006),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(net1006),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_1573_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(net1008),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_1107_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(net1010),
    .X(net1009));
 sg13g2_buf_1 fanout1010 (.A(_1093_),
    .X(net1010));
 sg13g2_buf_4 fanout1011 (.X(net1011),
    .A(_1092_));
 sg13g2_buf_2 fanout1012 (.A(_1092_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_4 fanout1014 (.X(net1014),
    .A(net1015));
 sg13g2_buf_2 fanout1015 (.A(_1055_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(net1017),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(net1018),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_1054_),
    .X(net1019));
 sg13g2_buf_4 fanout1020 (.X(net1020),
    .A(_1045_));
 sg13g2_buf_2 fanout1021 (.A(_1045_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(net1023),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_1044_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(net1029),
    .X(net1025));
 sg13g2_buf_1 fanout1026 (.A(net1029),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(net1028),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_1040_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_1039_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_1039_),
    .X(net1031));
 sg13g2_buf_4 fanout1032 (.X(net1032),
    .A(_1026_));
 sg13g2_buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(net1036),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(net1036),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_0509_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(net1038),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_0502_),
    .X(net1038));
 sg13g2_buf_4 fanout1039 (.X(net1039),
    .A(_1486_));
 sg13g2_buf_4 fanout1040 (.X(net1040),
    .A(_1486_));
 sg13g2_buf_2 fanout1041 (.A(net1045),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(net1044),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(net1044),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(net1045),
    .X(net1044));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(_1477_));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(_1021_));
 sg13g2_buf_4 fanout1047 (.X(net1047),
    .A(net1048));
 sg13g2_buf_2 fanout1048 (.A(_1004_),
    .X(net1048));
 sg13g2_buf_4 fanout1049 (.X(net1049),
    .A(_0988_));
 sg13g2_buf_2 fanout1050 (.A(_0935_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(net1052),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(net1053),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_0522_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_0375_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_1579_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(net1057),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_1578_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(net1059),
    .X(net1058));
 sg13g2_buf_4 fanout1059 (.X(net1059),
    .A(_1485_));
 sg13g2_buf_2 fanout1060 (.A(_1020_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_1018_),
    .X(net1061));
 sg13g2_buf_4 fanout1062 (.X(net1062),
    .A(_0455_));
 sg13g2_buf_2 fanout1063 (.A(_2061_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(net1066),
    .X(net1064));
 sg13g2_buf_1 fanout1065 (.A(net1066),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_1787_),
    .X(net1066));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(net1068));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(_1757_));
 sg13g2_buf_4 fanout1069 (.X(net1069),
    .A(_1582_));
 sg13g2_buf_2 fanout1070 (.A(net1071),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_0980_),
    .X(net1071));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(net1074));
 sg13g2_buf_1 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_0454_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_0380_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_2411_),
    .X(net1077));
 sg13g2_buf_4 fanout1078 (.X(net1078),
    .A(net1079));
 sg13g2_buf_4 fanout1079 (.X(net1079),
    .A(_2060_));
 sg13g2_buf_2 fanout1080 (.A(_1857_),
    .X(net1080));
 sg13g2_buf_4 fanout1081 (.X(net1081),
    .A(_1760_));
 sg13g2_buf_2 fanout1082 (.A(net1083),
    .X(net1082));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(_1341_));
 sg13g2_buf_1 fanout1084 (.A(_1341_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_1332_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(net1090),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(net1090),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_1210_),
    .X(net1090));
 sg13g2_buf_4 fanout1091 (.X(net1091),
    .A(net1092));
 sg13g2_buf_4 fanout1092 (.X(net1092),
    .A(_1022_));
 sg13g2_buf_4 fanout1093 (.X(net1093),
    .A(_1010_));
 sg13g2_buf_4 fanout1094 (.X(net1094),
    .A(_0994_));
 sg13g2_buf_2 fanout1095 (.A(net1096),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_0992_),
    .X(net1096));
 sg13g2_buf_4 fanout1097 (.X(net1097),
    .A(_0992_));
 sg13g2_buf_4 fanout1098 (.X(net1098),
    .A(_0453_));
 sg13g2_buf_2 fanout1099 (.A(_2736_),
    .X(net1099));
 sg13g2_buf_1 fanout1100 (.A(_2736_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(net1102),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_1795_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_buf_4 fanout1104 (.X(net1104),
    .A(_0991_));
 sg13g2_buf_4 fanout1105 (.X(net1105),
    .A(net1106));
 sg13g2_buf_4 fanout1106 (.X(net1106),
    .A(_0989_));
 sg13g2_buf_2 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_0989_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(net1110),
    .X(net1109));
 sg13g2_buf_4 fanout1110 (.X(net1110),
    .A(net1115));
 sg13g2_buf_2 fanout1111 (.A(net1112),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(net1115),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(net1114),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(net1115),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_0975_),
    .X(net1115));
 sg13g2_buf_4 fanout1116 (.X(net1116),
    .A(_0482_));
 sg13g2_buf_4 fanout1117 (.X(net1117),
    .A(_0464_));
 sg13g2_buf_2 fanout1118 (.A(_0406_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_2913_),
    .X(net1119));
 sg13g2_buf_4 fanout1120 (.X(net1120),
    .A(_2881_));
 sg13g2_buf_4 fanout1121 (.X(net1121),
    .A(_2836_));
 sg13g2_buf_4 fanout1122 (.X(net1122),
    .A(net1125));
 sg13g2_buf_4 fanout1123 (.X(net1123),
    .A(net1125));
 sg13g2_buf_2 fanout1124 (.A(net1125),
    .X(net1124));
 sg13g2_buf_4 fanout1125 (.X(net1125),
    .A(_0976_));
 sg13g2_buf_2 fanout1126 (.A(net1127),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(net1129),
    .X(net1128));
 sg13g2_buf_4 fanout1129 (.X(net1129),
    .A(_0976_));
 sg13g2_buf_2 fanout1130 (.A(_2759_),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_2757_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(_2738_),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_2738_),
    .X(net1133));
 sg13g2_buf_4 fanout1134 (.X(net1134),
    .A(_2730_));
 sg13g2_buf_1 fanout1135 (.A(_2730_),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(_2712_),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(net1138),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(_2705_),
    .X(net1138));
 sg13g2_buf_4 fanout1139 (.X(net1139),
    .A(_2705_));
 sg13g2_buf_2 fanout1140 (.A(_2059_),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(_2910_),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(_2910_),
    .X(net1142));
 sg13g2_buf_4 fanout1143 (.X(net1143),
    .A(_2760_));
 sg13g2_buf_2 fanout1144 (.A(_2760_),
    .X(net1144));
 sg13g2_buf_4 fanout1145 (.X(net1145),
    .A(_2748_));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(net1147));
 sg13g2_buf_2 fanout1147 (.A(_2744_),
    .X(net1147));
 sg13g2_buf_4 fanout1148 (.X(net1148),
    .A(_2725_));
 sg13g2_buf_4 fanout1149 (.X(net1149),
    .A(_2724_));
 sg13g2_buf_2 fanout1150 (.A(_2724_),
    .X(net1150));
 sg13g2_buf_2 fanout1151 (.A(net1152),
    .X(net1151));
 sg13g2_buf_4 fanout1152 (.X(net1152),
    .A(_2718_));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(_2716_));
 sg13g2_buf_2 fanout1154 (.A(_2715_),
    .X(net1154));
 sg13g2_buf_2 fanout1155 (.A(_2715_),
    .X(net1155));
 sg13g2_buf_4 fanout1156 (.X(net1156),
    .A(net1157));
 sg13g2_buf_4 fanout1157 (.X(net1157),
    .A(_2711_));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(net1159));
 sg13g2_buf_2 fanout1159 (.A(net1160),
    .X(net1159));
 sg13g2_buf_2 fanout1160 (.A(_2708_),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(_2691_),
    .X(net1161));
 sg13g2_buf_4 fanout1162 (.X(net1162),
    .A(_2671_));
 sg13g2_buf_2 fanout1163 (.A(_2666_),
    .X(net1163));
 sg13g2_buf_4 fanout1164 (.X(net1164),
    .A(\dtop.player_inst.synth.alu.acc[10] ));
 sg13g2_buf_4 fanout1165 (.X(net1165),
    .A(net640));
 sg13g2_buf_4 fanout1166 (.X(net1166),
    .A(\dtop.vtop.logo.addr[8] ));
 sg13g2_buf_2 fanout1167 (.A(\dtop.vtop.logo.addr[7] ),
    .X(net1167));
 sg13g2_buf_2 fanout1168 (.A(net1169),
    .X(net1168));
 sg13g2_buf_2 fanout1169 (.A(\dtop.vtop.logo.addr[6] ),
    .X(net1169));
 sg13g2_buf_2 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_buf_1 fanout1171 (.A(net1173),
    .X(net1171));
 sg13g2_buf_2 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_1 fanout1173 (.A(net1174),
    .X(net1173));
 sg13g2_buf_1 fanout1174 (.A(net1175),
    .X(net1174));
 sg13g2_buf_2 fanout1175 (.A(net612),
    .X(net1175));
 sg13g2_buf_4 fanout1176 (.X(net1176),
    .A(net623));
 sg13g2_buf_2 fanout1177 (.A(\dtop.oct_counter[5] ),
    .X(net1177));
 sg13g2_buf_4 fanout1178 (.X(net1178),
    .A(_0049_));
 sg13g2_buf_4 fanout1179 (.X(net1179),
    .A(\dtop.oct_counter[2] ));
 sg13g2_buf_4 fanout1180 (.X(net1180),
    .A(\dtop.oct_counter[1] ));
 sg13g2_buf_1 fanout1181 (.A(\dtop.oct_counter[1] ),
    .X(net1181));
 sg13g2_buf_2 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_2 fanout1183 (.A(net579),
    .X(net1183));
 sg13g2_buf_4 fanout1184 (.X(net1184),
    .A(net1186));
 sg13g2_buf_2 fanout1185 (.A(net1186),
    .X(net1185));
 sg13g2_buf_4 fanout1186 (.X(net1186),
    .A(net598));
 sg13g2_buf_2 fanout1187 (.A(net1188),
    .X(net1187));
 sg13g2_buf_2 fanout1188 (.A(net1189),
    .X(net1188));
 sg13g2_buf_2 fanout1189 (.A(net587),
    .X(net1189));
 sg13g2_buf_2 fanout1190 (.A(net1191),
    .X(net1190));
 sg13g2_buf_2 fanout1191 (.A(net1192),
    .X(net1191));
 sg13g2_buf_2 fanout1192 (.A(\dtop.enable ),
    .X(net1192));
 sg13g2_buf_2 fanout1193 (.A(net1195),
    .X(net1193));
 sg13g2_buf_1 fanout1194 (.A(net1195),
    .X(net1194));
 sg13g2_buf_2 fanout1195 (.A(net603),
    .X(net1195));
 sg13g2_buf_2 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_buf_2 fanout1197 (.A(\dtop.vtop.pipeline.nstep_zg[0] ),
    .X(net1197));
 sg13g2_buf_2 fanout1198 (.A(net1200),
    .X(net1198));
 sg13g2_buf_1 fanout1199 (.A(net1200),
    .X(net1199));
 sg13g2_buf_2 fanout1200 (.A(_0050_),
    .X(net1200));
 sg13g2_buf_2 fanout1201 (.A(net1203),
    .X(net1201));
 sg13g2_buf_2 fanout1202 (.A(net1203),
    .X(net1202));
 sg13g2_buf_1 fanout1203 (.A(net1204),
    .X(net1203));
 sg13g2_buf_2 fanout1204 (.A(net643),
    .X(net1204));
 sg13g2_buf_2 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_buf_2 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_2 fanout1207 (.A(\dtop.player_inst.program_addr[4] ),
    .X(net1207));
 sg13g2_buf_2 fanout1208 (.A(_0063_),
    .X(net1208));
 sg13g2_buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_2 fanout1210 (.A(net1211),
    .X(net1210));
 sg13g2_buf_4 fanout1211 (.X(net1211),
    .A(net626));
 sg13g2_buf_2 fanout1212 (.A(net1213),
    .X(net1212));
 sg13g2_buf_2 fanout1213 (.A(net1214),
    .X(net1213));
 sg13g2_buf_2 fanout1214 (.A(net1215),
    .X(net1214));
 sg13g2_buf_4 fanout1215 (.X(net1215),
    .A(\dtop.player_inst.program_addr[2] ));
 sg13g2_buf_2 fanout1216 (.A(net1218),
    .X(net1216));
 sg13g2_buf_2 fanout1217 (.A(net1218),
    .X(net1217));
 sg13g2_buf_1 fanout1218 (.A(net1219),
    .X(net1218));
 sg13g2_buf_4 fanout1219 (.X(net1219),
    .A(net1220));
 sg13g2_buf_4 fanout1220 (.X(net1220),
    .A(\dtop.player_inst.program_addr[1] ));
 sg13g2_buf_4 fanout1221 (.X(net1221),
    .A(net1223));
 sg13g2_buf_2 fanout1222 (.A(net1223),
    .X(net1222));
 sg13g2_buf_2 fanout1223 (.A(net1224),
    .X(net1223));
 sg13g2_buf_2 fanout1224 (.A(net1225),
    .X(net1224));
 sg13g2_buf_2 fanout1225 (.A(\dtop.player_inst.program_addr[0] ),
    .X(net1225));
 sg13g2_buf_4 fanout1226 (.X(net1226),
    .A(\dtop.vtop.rs.saturated ));
 sg13g2_buf_2 fanout1227 (.A(\dtop.detune_counter[16] ),
    .X(net1227));
 sg13g2_buf_2 fanout1228 (.A(net1229),
    .X(net1228));
 sg13g2_buf_2 fanout1229 (.A(net631),
    .X(net1229));
 sg13g2_buf_2 fanout1230 (.A(net632),
    .X(net1230));
 sg13g2_buf_4 fanout1231 (.X(net1231),
    .A(net1232));
 sg13g2_buf_4 fanout1232 (.X(net1232),
    .A(\dtop.detune_counter[11] ));
 sg13g2_buf_2 fanout1233 (.A(_0073_),
    .X(net1233));
 sg13g2_buf_2 fanout1234 (.A(net1235),
    .X(net1234));
 sg13g2_buf_4 fanout1235 (.X(net1235),
    .A(net590));
 sg13g2_buf_2 fanout1236 (.A(net648),
    .X(net1236));
 sg13g2_buf_1 fanout1237 (.A(\dtop.detune_counter[7] ),
    .X(net1237));
 sg13g2_buf_2 fanout1238 (.A(net1239),
    .X(net1238));
 sg13g2_buf_2 fanout1239 (.A(net1242),
    .X(net1239));
 sg13g2_buf_1 fanout1240 (.A(net1242),
    .X(net1240));
 sg13g2_buf_2 fanout1241 (.A(net1242),
    .X(net1241));
 sg13g2_buf_2 fanout1242 (.A(net1243),
    .X(net1242));
 sg13g2_buf_2 fanout1243 (.A(rst_n),
    .X(net1243));
 sg13g2_buf_2 fanout1244 (.A(net1245),
    .X(net1244));
 sg13g2_buf_2 fanout1245 (.A(net1246),
    .X(net1245));
 sg13g2_buf_2 fanout1246 (.A(net1247),
    .X(net1246));
 sg13g2_buf_2 fanout1247 (.A(rst_n),
    .X(net1247));
 sg13g2_buf_2 fanout1248 (.A(net1249),
    .X(net1248));
 sg13g2_buf_2 fanout1249 (.A(net1252),
    .X(net1249));
 sg13g2_buf_2 fanout1250 (.A(net1251),
    .X(net1250));
 sg13g2_buf_4 fanout1251 (.X(net1251),
    .A(net1252));
 sg13g2_buf_4 fanout1252 (.X(net1252),
    .A(rst_n));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ui_in[0]));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[2]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[3]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[7]));
 sg13g2_tielo tt_um_toivoh_demo_tt08_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_36_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_38_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_1_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_24_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_33_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_10_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_16_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_17_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_23_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_34_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_20_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_21_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\dtop.vtop.pipeline.next_nstep_counter[0] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0270_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold3 (.A(\dtop.vtop.dphases[0][10] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold4 (.A(\dtop.vtop.dphases[0][1] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold5 (.A(\dtop.vtop.dphases[0][8] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold6 (.A(\dtop.vtop.dphases[0][2] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold7 (.A(\dtop.vtop.dphases[0][6] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold8 (.A(\dtop.player_inst.synth.alu.registers[4][8] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0356_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold10 (.A(\dtop.vtop.dphases[0][0] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold11 (.A(\dtop.vtop.dphases[0][9] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold12 (.A(\dtop.player_inst.synth.alu.registers[4][6] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0354_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold14 (.A(\dtop.player_inst.synth.alu.registers[4][9] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold15 (.A(\dtop.vtop.dphases[1][6] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold16 (.A(\dtop.vtop.dphases[2][10] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold17 (.A(\dtop.vtop.dphases[0][3] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold18 (.A(\dtop.vtop.dphases[2][6] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold19 (.A(\dtop.player_inst.synth.alu.registers[4][7] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0355_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold21 (.A(\dtop.player_inst.synth.alu.registers[5][5] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold22 (.A(\dtop.player_inst.synth.alu.registers[2][2] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold23 (.A(\dtop.vtop.pipeline.cosappr_acc[2] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold24 (.A(\dtop.vtop.dphases[1][0] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold25 (.A(\dtop.vtop.pipeline.zg_acc[1] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold26 (.A(\dtop.player_inst.synth.alu.registers[2][1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0341_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold28 (.A(\dtop.vtop.pipeline.cosappr_acc[1] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold29 (.A(\dtop.vtop.dphases[1][8] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold30 (.A(\dtop.vtop.dphases[2][2] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold31 (.A(\dtop.player_inst.synth.alu.registers[5][1] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0368_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold33 (.A(\dtop.player_inst.synth.alu.registers[4][3] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold34 (.A(\dtop.player_inst.synth.alu.registers[4][10] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0358_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold36 (.A(\dtop.vtop.dphases[1][9] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold37 (.A(\dtop.player_inst.synth.alu.registers[2][5] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold38 (.A(\dtop.vtop.dphases[2][8] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold39 (.A(\dtop.player_inst.synth.alu.registers[1][1] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0329_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold41 (.A(\dtop.player_inst.synth.alu.registers[1][6] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold42 (.A(\dtop.player_inst.synth.alu.registers[5][6] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold43 (.A(\dtop.player_inst.synth.alu.registers[1][3] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold44 (.A(\dtop.player_inst.synth.alu.registers[4][1] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0349_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold46 (.A(\dtop.vtop.pipeline.zg_acc[7] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold47 (.A(\dtop.player_inst.synth.alu.registers[2][4] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold48 (.A(\dtop.player_inst.synth.alu.registers[1][9] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold49 (.A(\dtop.player_inst.synth.alu.registers[4][5] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0353_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold51 (.A(\dtop.player_inst.synth.alu.registers[5][4] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0371_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold53 (.A(\dtop.vtop.dphases[2][9] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold54 (.A(\dtop.vtop.pipeline.cosappr_acc[4] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold55 (.A(\dtop.player_inst.synth.alu.registers[3][5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold56 (.A(\dtop.player_inst.synth.alu.registers[3][7] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0366_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold58 (.A(\dtop.vtop.pipeline.zg_acc[6] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold59 (.A(\dtop.player_inst.synth.alu.registers[3][1] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0360_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold61 (.A(\dtop.vtop.dphases[1][1] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold62 (.A(\dtop.vtop.dphases[1][2] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold63 (.A(\dtop.player_inst.synth.alu.registers[2][0] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0340_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold65 (.A(\dtop.vtop.dphases[2][0] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold66 (.A(\dtop.player_inst.synth.alu.registers[2][6] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold67 (.A(\dtop.player_inst.synth.alu.registers[2][3] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold68 (.A(\dtop.out_sample[0] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0310_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold70 (.A(\dtop.player_inst.synth.alu.registers[3][4] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0363_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold72 (.A(\dtop.player_inst.synth.alu.registers[1][7] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0335_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold74 (.A(\dtop.player_inst.synth.alu.registers[3][0] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold75 (.A(\dtop.player_inst.synth.alu.registers[1][4] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold76 (.A(\dtop.player_inst.synth.alu.registers[1][2] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold77 (.A(\dtop.player_inst.synth.alu.registers[1][0] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold78 (.A(\dtop.player_inst.synth.alu.registers[2][7] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0347_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold80 (.A(\dtop.vtop.dphases[1][3] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold81 (.A(\dtop.player_inst.synth.alu.registers[1][5] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold82 (.A(\dtop.vtop.pipeline.z[0] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold83 (.A(\dtop.vtop.dphases[2][1] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold84 (.A(\dtop.vtop.pipeline.phases[1][7] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold85 (.A(\dtop.vsync ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0139_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold87 (.A(\dtop.player_inst.synth.alu.registers[1][8] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0336_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold89 (.A(\dtop.vtop.pipeline.cosappr_acc[0] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold90 (.A(\dtop.out_sample[4] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0314_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold92 (.A(\dtop.player_inst.synth.alu.registers[5][3] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold93 (.A(\dtop.player_inst.synth.alu.registers[5][2] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold94 (.A(\dtop.vtop.pipeline.phases[1][5] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold95 (.A(\dtop.vtop.pipeline.cosappr_acc[5] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold96 (.A(\dtop.vtop.pipeline.phases[1][1] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold97 (.A(\dtop.vtop.pipeline.phases[1][4] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold98 (.A(\dtop.vtop.pipeline.phases[1][10] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold99 (.A(\dtop.vtop.pipeline.phases[0][7] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold100 (.A(\dtop.vtop.pipeline.phases[1][0] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0187_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold102 (.A(\dtop.vtop.dphases[0][4] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold103 (.A(\dtop.vtop.pipeline.cosappr_acc[6] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold104 (.A(\dtop.vtop.pipeline.phases[1][13] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold105 (.A(\dtop.player_inst.synth.alu.registers[3][6] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold106 (.A(\dtop.player_inst.synth.alu.registers[4][2] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold107 (.A(\dtop.vtop.pipeline.phases[0][5] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold108 (.A(\dtop.vtop.dphases[0][7] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold109 (.A(\dtop.vtop.pipeline.cosappr_acc[7] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold110 (.A(\dtop.vtop.pipeline.phases[0][9] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold111 (.A(\dtop.vtop.pipeline.phases[1][2] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold112 (.A(\dtop.out_sample[6] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold113 (.A(\dtop.player_inst.synth.alu.registers[1][10] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0338_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold115 (.A(\dtop.player_inst.synth.alu.registers[5][0] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold116 (.A(\dtop.vtop.dphases[0][5] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold117 (.A(\dtop.vtop.pipeline.phases[0][12] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold118 (.A(\dtop.vtop.pipeline.phases[0][6] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold119 (.A(\dtop.vtop.pipeline.phases[0][0] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0220_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold121 (.A(\dtop.vtop.pipeline.phases[0][4] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold122 (.A(\dtop.vtop.pipeline.phases[1][12] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold123 (.A(\dtop.vtop.pipeline.phases[1][3] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold124 (.A(uo_out[1]),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0279_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold126 (.A(\dtop.vtop.pipeline.phases[0][1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold127 (.A(\dtop.vtop.pipeline.phases[0][2] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold128 (.A(\dtop.vtop.pipeline.phases[1][6] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold129 (.A(\dtop.vtop.pipeline.phases[0][13] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold130 (.A(\dtop.vtop.pipeline.phases[0][15] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold131 (.A(\dtop.vtop.pipeline.phases[1][8] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold132 (.A(\dtop.vtop.pipeline.phases[1][11] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold133 (.A(\dtop.vtop.pipeline.phases[0][8] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold134 (.A(\dtop.player_inst.synth.alu.registers[3][3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold135 (.A(\dtop.vtop.pipeline.phases[0][3] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold136 (.A(\dtop.player_inst.synth.alu.registers[3][2] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold137 (.A(\dtop.out_sample[2] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold138 (.A(\dtop.vtop.color[5] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold139 (.A(\dtop.player_inst.synth.alu.oct_en ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold140 (.A(\dtop.out_sample[5] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0315_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold142 (.A(\dtop.player_inst.synth.alu.registers[4][0] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0348_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold144 (.A(\dtop.out_sample[3] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold145 (.A(\dtop.player_inst.synth.alu.registers[4][4] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0352_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold147 (.A(\dtop.vtop.pipeline.zg_acc[9] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold148 (.A(\dtop.vtop.dphases[2][3] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold149 (.A(\dtop.vtop.pipeline.dz[3] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold150 (.A(\dtop.vtop.pipeline.phases[0][11] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold151 (.A(\dtop.vtop.pipeline.phases[0][14] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold152 (.A(\dtop.vtop.pipeline.cosappr_acc[3] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold153 (.A(\dtop.vtop.dphases[2][7] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold154 (.A(\dtop.vtop.pipeline.phases[2][12] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold155 (.A(\dtop.vtop.dphases[1][4] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold156 (.A(uo_out[2]),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0280_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold158 (.A(\dtop.vtop.dphases[1][10] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold159 (.A(\dtop.vtop.pipeline.phases[0][10] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold160 (.A(\dtop.vtop.pipeline.phases[2][8] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold161 (.A(\dtop.vtop.pipeline.phases[1][15] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold162 (.A(\dtop.vtop.pipeline.zg[0] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold163 (.A(\dtop.vtop.pipeline.phases[1][9] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold164 (.A(uo_out[6]),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0282_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold166 (.A(uo_out[3]),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0288_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold168 (.A(uo_out[5]),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0281_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold170 (.A(\dtop.vtop.pipeline.cosappr_acc[8] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold171 (.A(\dtop.vtop.dphases[1][5] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold172 (.A(\dtop.vtop.pipeline.phases[2][4] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold173 (.A(\dtop.vtop.pipeline.zg[3] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold174 (.A(\dtop.vtop.pipeline.phases[2][9] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold175 (.A(\dtop.vtop.pipeline.phases[2][1] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold176 (.A(\dtop.vtop.pipeline.phases[2][10] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold177 (.A(\dtop.vtop.pipeline.phases[2][11] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold178 (.A(\dtop.vtop.pipeline.phases[2][14] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold179 (.A(\dtop.vtop.pipeline.nstep_counter[3] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold180 (.A(_2184_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0273_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold182 (.A(\dtop.vtop.dphases[2][5] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold183 (.A(\dtop.vtop.dphases[2][4] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold184 (.A(\dtop.vtop.pipeline.phases[2][5] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold185 (.A(\dtop.vtop.pipeline.z[2] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold186 (.A(\dtop.vtop.pipeline.z[4] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0176_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold188 (.A(\dtop.vtop.dphases[1][7] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold189 (.A(\dtop.vtop.pipeline.phases[2][0] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0203_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold191 (.A(\dtop.vtop.pipeline.phases[2][7] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold192 (.A(\dtop.vtop.pipeline.phases[1][14] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold193 (.A(\dtop.vtop.pipeline.phases[2][13] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold194 (.A(\dtop.vtop.pipeline.z[14] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold195 (.A(\dtop.out_sample[1] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0311_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold197 (.A(\dtop.vtop.pipeline.phases[2][3] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold198 (.A(\dtop.vtop.pipeline.zg_acc[0] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold199 (.A(\dtop.vtop.pipeline.zg_acc[2] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold200 (.A(\dtop.vtop.pipeline.zg_acc[5] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold201 (.A(uo_out[7]),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold202 (.A(\dtop.player_inst.synth.alu.registers[0][0] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0317_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold204 (.A(\dtop.vtop.pipeline.phases[2][2] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold205 (.A(\dtop.vtop.pipeline.zg_acc[4] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold206 (.A(\dtop.player_inst.synth.alu.registers[0][3] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold207 (.A(\dtop.vtop.pipeline.neg_t[6] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold208 (.A(\dtop.vtop.pipeline.phases[2][6] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold209 (.A(\dtop.player_inst.synth.alu.registers[0][8] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0325_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold211 (.A(\dtop.vtop.pipeline.zg_acc[8] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold212 (.A(\dtop.vtop.pipeline.neg_t[8] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold213 (.A(\dtop.vtop.pipeline.neg_t[4] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold214 (.A(_1520_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0157_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold216 (.A(\dtop.player_inst.synth.alu.registers[0][6] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold217 (.A(\dtop.vtop.pipeline.dz[2] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold218 (.A(\dtop.vtop.pipeline.zg[1] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold219 (.A(\dtop.player_inst.synth.alu.registers[0][2] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold220 (.A(\dtop.player_inst.synth.alu.registers[0][10] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0327_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold222 (.A(\dtop.vtop.pipeline.nstep_counter[2] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold223 (.A(\dtop.vtop.pipeline.nstep_counter[4] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold224 (.A(\dtop.player_inst.synth.alu.registers[0][1] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0318_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold226 (.A(uio_out[7]),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold227 (.A(\dtop.vtop.pipeline.phases[2][15] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold228 (.A(\dtop.vtop.pipeline.zg[4] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold229 (.A(\dtop.player_inst.synth.alu.registers[0][7] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0324_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold231 (.A(\dtop.vtop.pipeline.dz[7] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold232 (.A(\dtop.vtop.pipeline.nstep_counter[1] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold233 (.A(_2182_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0271_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold235 (.A(\dtop.vtop.pipeline.zg[2] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold236 (.A(\dtop.vtop.color[4] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold237 (.A(\dtop.vtop.pipeline.dz[1] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold238 (.A(\dtop.vtop.pipeline.dz[5] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold239 (.A(\dtop.vtop.pipeline.dz[6] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold240 (.A(\dtop.vtop.pipeline.zg_acc[3] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold241 (.A(\dtop.vtop.pipeline.z[11] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold242 (.A(\dtop.vtop.pipeline.z[8] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0180_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold244 (.A(\dtop.vtop.pipeline.neg_t[2] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0085_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold246 (.A(_2519_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold247 (.A(\dtop.player_inst.synth.alu.registers[0][4] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold248 (.A(\dtop.player_inst.synth.alu.registers[0][9] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold249 (.A(\dtop.vtop.pipeline.dz[0] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0163_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold251 (.A(\dtop.vtop.pipeline.dz[8] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold252 (.A(_2962_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold253 (.A(\dtop.vtop.pipeline.neg_t[0] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold254 (.A(\dtop.player_inst.synth.alu.registers[0][5] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold255 (.A(\dtop.vtop.pipeline.neg_t[1] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold256 (.A(\dtop.vtop.pipeline.z[3] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold257 (.A(\dtop.vtop.pipeline.z[6] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0178_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold259 (.A(\dtop.vtop.pipeline.neg_t[5] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold260 (.A(\dtop.vtop.color[6] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold261 (.A(\dtop.vtop.pipeline.neg_t[9] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold262 (.A(_1540_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold263 (.A(\dtop.vtop.pipeline.z[1] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold264 (.A(\dtop.detune_counter[14] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold265 (.A(\dtop.vtop.rs.scan_y.phase[1] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold266 (.A(\dtop.vtop.pipeline.zg[5] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold267 (.A(\dtop.vtop.pipeline.z[9] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold268 (.A(\dtop.detune_counter[5] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold269 (.A(\dtop.vtop.pipeline.z[10] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0053_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold271 (.A(_2512_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold272 (.A(\dtop.detune_counter[6] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold273 (.A(\dtop.vtop.pipeline.dz[4] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold274 (.A(\dtop.oct_counter[0] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold275 (.A(\dtop.vtop.logo.addr[7] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold276 (.A(\dtop.vtop.rs.x_scan.phase[0] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold277 (.A(_1438_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold278 (.A(\dtop.vtop.pipeline.z[12] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold279 (.A(\dtop.vtop.rs.x_scan.phase[1] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold280 (.A(\dtop.vtop.pipeline.neg_t[3] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold281 (.A(\dtop.player_inst.synth.alu.acc[8] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold282 (.A(\dtop.vtop.pipeline.nstep[0] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold283 (.A(\dtop.vtop.pipeline.neg_t[7] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0160_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold285 (.A(\dtop.detune_counter[8] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0962_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold287 (.A(\dtop.vtop.pipeline.z[5] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0177_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold289 (.A(uo_out[4]),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold290 (.A(\dtop.vtop.color[7] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold291 (.A(\dtop.player_inst.synth.alu.carry ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold292 (.A(\dtop.vtop.pipeline.z[7] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold293 (.A(\dtop.vtop.pipeline.nstep[1] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold294 (.A(\dtop.player_inst.synth.alu.acc[5] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold295 (.A(\dtop.vtop.pipeline.z[13] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold296 (.A(\dtop.oct_counter[4] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold297 (.A(_2511_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold298 (.A(\dtop.vtop.pipeline.nstep_zg[1] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0055_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0924_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0285_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0003_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold303 (.A(_2166_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold304 (.A(uo_out[0]),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold305 (.A(\dtop.vtop.pipeline.wave_index[0] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold306 (.A(_1756_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold307 (.A(\dtop.vtop.logo.addr[5] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0086_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold309 (.A(_2516_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0052_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold311 (.A(\dtop.vtop.logo.addr[8] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0056_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold313 (.A(_2479_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0284_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold315 (.A(\dtop.player_inst.synth.alu.acc[6] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0058_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0953_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold318 (.A(\dtop.oct_counter[6] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold319 (.A(\dtop.vtop.pipeline.zg[7] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold320 (.A(\dtop.vtop.pipeline.zg[6] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold321 (.A(\dtop.player_inst.program_addr[3] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold322 (.A(_1449_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold323 (.A(\dtop.detune_counter[10] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0965_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold325 (.A(\dtop.player_inst.synth.alu.acc[0] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold326 (.A(\dtop.detune_counter[15] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold327 (.A(\dtop.detune_counter[13] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0080_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0961_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold330 (.A(\dtop.player_inst.synth.alu.acc[4] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold331 (.A(\dtop.player_inst.synth.alu.acc[7] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0083_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold333 (.A(\dtop.player_inst.synth.alu.acc[1] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold334 (.A(\dtop.vtop.pipeline.zg_valid ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold335 (.A(\dtop.player_inst.synth.alu.acc[10] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold336 (.A(\dtop.vtop.pipeline.zg[8] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold337 (.A(\dtop.player_inst.synth.alu.acc[3] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold338 (.A(\dtop.player_inst.program_addr[5] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0070_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold340 (.A(\dtop.vtop.pipeline.zg[9] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold341 (.A(\dtop.player_inst.synth.alu.acc[2] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold342 (.A(\dtop.detune_counter[9] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold343 (.A(\dtop.detune_counter[7] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold344 (.A(\dtop.player_inst.synth.alu.acc[4] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold345 (.A(\dtop.player_inst.synth.alu.acc[0] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold346 (.A(\dtop.vtop.pipeline.zg_valid ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold347 (.A(\dtop.player_inst.synth.alu.acc[5] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold348 (.A(\dtop.vtop.rs.x_scan.phase[0] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold349 (.A(\dtop.player_inst.synth.alu.acc[6] ),
    .X(net654));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_61 ();
 sg13g2_fill_1 FILLER_0_90 ();
 sg13g2_fill_2 FILLER_0_95 ();
 sg13g2_fill_1 FILLER_0_140 ();
 sg13g2_fill_2 FILLER_0_167 ();
 sg13g2_fill_1 FILLER_0_169 ();
 sg13g2_fill_2 FILLER_0_178 ();
 sg13g2_fill_1 FILLER_0_188 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_4 FILLER_0_222 ();
 sg13g2_fill_2 FILLER_0_226 ();
 sg13g2_fill_1 FILLER_0_287 ();
 sg13g2_fill_2 FILLER_0_340 ();
 sg13g2_fill_1 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_fill_2 FILLER_1_28 ();
 sg13g2_fill_1 FILLER_1_30 ();
 sg13g2_fill_2 FILLER_1_79 ();
 sg13g2_fill_2 FILLER_1_113 ();
 sg13g2_fill_1 FILLER_1_115 ();
 sg13g2_fill_2 FILLER_1_156 ();
 sg13g2_fill_1 FILLER_1_168 ();
 sg13g2_fill_1 FILLER_1_195 ();
 sg13g2_decap_8 FILLER_1_207 ();
 sg13g2_fill_1 FILLER_1_214 ();
 sg13g2_fill_1 FILLER_1_223 ();
 sg13g2_fill_2 FILLER_1_259 ();
 sg13g2_fill_1 FILLER_1_261 ();
 sg13g2_fill_1 FILLER_1_270 ();
 sg13g2_fill_2 FILLER_1_283 ();
 sg13g2_fill_1 FILLER_1_285 ();
 sg13g2_fill_1 FILLER_1_300 ();
 sg13g2_fill_2 FILLER_1_306 ();
 sg13g2_fill_1 FILLER_1_308 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_fill_2 FILLER_2_28 ();
 sg13g2_fill_1 FILLER_2_35 ();
 sg13g2_fill_1 FILLER_2_201 ();
 sg13g2_fill_1 FILLER_2_269 ();
 sg13g2_fill_2 FILLER_2_402 ();
 sg13g2_fill_1 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_16 ();
 sg13g2_fill_1 FILLER_3_51 ();
 sg13g2_fill_2 FILLER_3_174 ();
 sg13g2_fill_1 FILLER_3_176 ();
 sg13g2_fill_2 FILLER_3_195 ();
 sg13g2_fill_2 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_4 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_11 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_fill_2 FILLER_4_145 ();
 sg13g2_fill_1 FILLER_4_147 ();
 sg13g2_fill_2 FILLER_4_266 ();
 sg13g2_fill_1 FILLER_4_276 ();
 sg13g2_fill_2 FILLER_4_304 ();
 sg13g2_fill_1 FILLER_4_316 ();
 sg13g2_fill_1 FILLER_4_396 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_9 ();
 sg13g2_fill_2 FILLER_5_83 ();
 sg13g2_fill_1 FILLER_5_136 ();
 sg13g2_fill_2 FILLER_5_198 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_fill_1 FILLER_5_227 ();
 sg13g2_fill_2 FILLER_5_235 ();
 sg13g2_fill_1 FILLER_5_237 ();
 sg13g2_fill_2 FILLER_5_244 ();
 sg13g2_fill_2 FILLER_5_266 ();
 sg13g2_fill_1 FILLER_5_268 ();
 sg13g2_fill_2 FILLER_5_284 ();
 sg13g2_fill_1 FILLER_5_286 ();
 sg13g2_fill_1 FILLER_5_323 ();
 sg13g2_fill_2 FILLER_5_335 ();
 sg13g2_fill_1 FILLER_5_337 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_47 ();
 sg13g2_fill_1 FILLER_6_90 ();
 sg13g2_fill_2 FILLER_6_192 ();
 sg13g2_fill_1 FILLER_6_194 ();
 sg13g2_fill_1 FILLER_6_231 ();
 sg13g2_fill_1 FILLER_6_242 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_27 ();
 sg13g2_fill_2 FILLER_7_85 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_157 ();
 sg13g2_fill_2 FILLER_7_210 ();
 sg13g2_fill_2 FILLER_7_224 ();
 sg13g2_fill_2 FILLER_7_261 ();
 sg13g2_fill_1 FILLER_7_263 ();
 sg13g2_fill_2 FILLER_7_312 ();
 sg13g2_fill_2 FILLER_7_329 ();
 sg13g2_fill_1 FILLER_7_331 ();
 sg13g2_fill_2 FILLER_7_358 ();
 sg13g2_fill_1 FILLER_7_360 ();
 sg13g2_fill_2 FILLER_7_396 ();
 sg13g2_fill_1 FILLER_7_398 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_4 ();
 sg13g2_fill_2 FILLER_8_36 ();
 sg13g2_fill_1 FILLER_8_38 ();
 sg13g2_fill_1 FILLER_8_89 ();
 sg13g2_fill_1 FILLER_8_124 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_193 ();
 sg13g2_fill_2 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_205 ();
 sg13g2_fill_2 FILLER_8_244 ();
 sg13g2_fill_2 FILLER_8_264 ();
 sg13g2_fill_1 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_fill_1 FILLER_8_316 ();
 sg13g2_fill_1 FILLER_8_337 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_68 ();
 sg13g2_fill_1 FILLER_9_88 ();
 sg13g2_fill_1 FILLER_9_134 ();
 sg13g2_fill_2 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_236 ();
 sg13g2_fill_2 FILLER_9_253 ();
 sg13g2_fill_1 FILLER_9_255 ();
 sg13g2_fill_2 FILLER_9_266 ();
 sg13g2_fill_1 FILLER_9_268 ();
 sg13g2_fill_1 FILLER_9_295 ();
 sg13g2_fill_2 FILLER_9_372 ();
 sg13g2_fill_1 FILLER_9_379 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_fill_1 FILLER_10_107 ();
 sg13g2_fill_2 FILLER_10_114 ();
 sg13g2_fill_1 FILLER_10_116 ();
 sg13g2_fill_2 FILLER_10_155 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_fill_2 FILLER_10_174 ();
 sg13g2_fill_1 FILLER_10_176 ();
 sg13g2_fill_2 FILLER_10_201 ();
 sg13g2_fill_1 FILLER_10_203 ();
 sg13g2_fill_2 FILLER_10_216 ();
 sg13g2_fill_2 FILLER_10_277 ();
 sg13g2_fill_1 FILLER_10_318 ();
 sg13g2_fill_1 FILLER_10_339 ();
 sg13g2_fill_1 FILLER_10_351 ();
 sg13g2_fill_2 FILLER_10_358 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_22 ();
 sg13g2_fill_2 FILLER_11_28 ();
 sg13g2_fill_2 FILLER_11_40 ();
 sg13g2_fill_2 FILLER_11_73 ();
 sg13g2_fill_1 FILLER_11_93 ();
 sg13g2_fill_2 FILLER_11_109 ();
 sg13g2_fill_1 FILLER_11_111 ();
 sg13g2_fill_1 FILLER_11_126 ();
 sg13g2_fill_2 FILLER_11_207 ();
 sg13g2_fill_1 FILLER_11_209 ();
 sg13g2_fill_1 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_273 ();
 sg13g2_fill_1 FILLER_11_338 ();
 sg13g2_fill_2 FILLER_11_348 ();
 sg13g2_fill_1 FILLER_11_350 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_59 ();
 sg13g2_fill_2 FILLER_12_78 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_2 FILLER_12_86 ();
 sg13g2_fill_1 FILLER_12_88 ();
 sg13g2_fill_2 FILLER_12_126 ();
 sg13g2_fill_2 FILLER_12_199 ();
 sg13g2_fill_1 FILLER_12_201 ();
 sg13g2_fill_2 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_fill_2 FILLER_12_280 ();
 sg13g2_fill_1 FILLER_12_308 ();
 sg13g2_fill_2 FILLER_12_387 ();
 sg13g2_fill_1 FILLER_12_389 ();
 sg13g2_fill_1 FILLER_13_69 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_183 ();
 sg13g2_fill_1 FILLER_13_185 ();
 sg13g2_fill_2 FILLER_13_191 ();
 sg13g2_fill_1 FILLER_13_193 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_2 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_261 ();
 sg13g2_fill_2 FILLER_13_274 ();
 sg13g2_fill_1 FILLER_13_276 ();
 sg13g2_fill_2 FILLER_13_301 ();
 sg13g2_fill_1 FILLER_13_317 ();
 sg13g2_fill_2 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_346 ();
 sg13g2_fill_2 FILLER_13_374 ();
 sg13g2_fill_1 FILLER_13_376 ();
 sg13g2_fill_1 FILLER_14_36 ();
 sg13g2_fill_1 FILLER_14_86 ();
 sg13g2_fill_1 FILLER_14_97 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_decap_4 FILLER_14_121 ();
 sg13g2_fill_1 FILLER_14_125 ();
 sg13g2_fill_1 FILLER_14_171 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_decap_4 FILLER_14_194 ();
 sg13g2_fill_2 FILLER_14_198 ();
 sg13g2_decap_8 FILLER_14_219 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_fill_1 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_282 ();
 sg13g2_fill_1 FILLER_14_284 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_338 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_78 ();
 sg13g2_fill_1 FILLER_15_80 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_fill_1 FILLER_15_103 ();
 sg13g2_fill_2 FILLER_15_109 ();
 sg13g2_fill_1 FILLER_15_111 ();
 sg13g2_decap_4 FILLER_15_129 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_decap_4 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_4 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_fill_1 FILLER_15_226 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_fill_2 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_1 FILLER_16_11 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_fill_1 FILLER_16_51 ();
 sg13g2_fill_2 FILLER_16_78 ();
 sg13g2_fill_2 FILLER_16_100 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_fill_2 FILLER_16_130 ();
 sg13g2_fill_1 FILLER_16_132 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_fill_2 FILLER_16_144 ();
 sg13g2_fill_1 FILLER_16_146 ();
 sg13g2_decap_4 FILLER_16_175 ();
 sg13g2_decap_4 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_209 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_237 ();
 sg13g2_fill_1 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_17_59 ();
 sg13g2_fill_2 FILLER_17_69 ();
 sg13g2_fill_1 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_143 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_decap_8 FILLER_17_158 ();
 sg13g2_decap_8 FILLER_17_165 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_174 ();
 sg13g2_fill_1 FILLER_17_201 ();
 sg13g2_decap_4 FILLER_17_224 ();
 sg13g2_fill_2 FILLER_17_233 ();
 sg13g2_fill_1 FILLER_17_235 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_fill_2 FILLER_17_282 ();
 sg13g2_fill_1 FILLER_17_299 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_336 ();
 sg13g2_fill_2 FILLER_17_352 ();
 sg13g2_fill_2 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_75 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_fill_1 FILLER_18_151 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_227 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_238 ();
 sg13g2_fill_1 FILLER_18_240 ();
 sg13g2_fill_2 FILLER_18_253 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_19_79 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_104 ();
 sg13g2_fill_2 FILLER_19_130 ();
 sg13g2_fill_1 FILLER_19_132 ();
 sg13g2_fill_1 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_283 ();
 sg13g2_fill_1 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_fill_1 FILLER_19_390 ();
 sg13g2_fill_2 FILLER_20_25 ();
 sg13g2_fill_1 FILLER_20_27 ();
 sg13g2_fill_2 FILLER_20_48 ();
 sg13g2_fill_1 FILLER_20_71 ();
 sg13g2_fill_2 FILLER_20_130 ();
 sg13g2_fill_2 FILLER_20_193 ();
 sg13g2_fill_1 FILLER_20_195 ();
 sg13g2_decap_4 FILLER_20_206 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_fill_1 FILLER_20_309 ();
 sg13g2_fill_1 FILLER_20_360 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_198 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_246 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_22_26 ();
 sg13g2_fill_1 FILLER_22_33 ();
 sg13g2_fill_2 FILLER_22_56 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_158 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_decap_8 FILLER_22_219 ();
 sg13g2_decap_4 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_256 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_fill_2 FILLER_22_339 ();
 sg13g2_fill_2 FILLER_22_354 ();
 sg13g2_fill_2 FILLER_22_384 ();
 sg13g2_fill_2 FILLER_22_395 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_fill_1 FILLER_23_96 ();
 sg13g2_fill_2 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_fill_1 FILLER_23_228 ();
 sg13g2_fill_1 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_262 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_333 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_fill_1 FILLER_24_69 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_fill_2 FILLER_24_161 ();
 sg13g2_decap_4 FILLER_24_220 ();
 sg13g2_fill_2 FILLER_24_238 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_11 ();
 sg13g2_fill_2 FILLER_25_188 ();
 sg13g2_decap_4 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_231 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_314 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_2 FILLER_25_353 ();
 sg13g2_fill_2 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_25 ();
 sg13g2_fill_1 FILLER_26_30 ();
 sg13g2_fill_2 FILLER_26_97 ();
 sg13g2_fill_1 FILLER_26_99 ();
 sg13g2_decap_4 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_decap_4 FILLER_26_210 ();
 sg13g2_fill_2 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_fill_1 FILLER_26_334 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_fill_2 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_2 FILLER_27_177 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_fill_2 FILLER_27_193 ();
 sg13g2_fill_2 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_218 ();
 sg13g2_fill_2 FILLER_27_226 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_fill_2 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_333 ();
 sg13g2_fill_1 FILLER_27_340 ();
 sg13g2_fill_1 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_9 ();
 sg13g2_decap_4 FILLER_28_176 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_fill_2 FILLER_28_398 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_48 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_fill_2 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_230 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_fill_1 FILLER_29_370 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_31 ();
 sg13g2_fill_2 FILLER_30_45 ();
 sg13g2_fill_1 FILLER_30_47 ();
 sg13g2_fill_2 FILLER_30_69 ();
 sg13g2_fill_1 FILLER_30_71 ();
 sg13g2_fill_1 FILLER_30_81 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_2 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_190 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_fill_2 FILLER_30_215 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_fill_1 FILLER_30_240 ();
 sg13g2_fill_1 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_fill_1 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_61 ();
 sg13g2_decap_4 FILLER_31_68 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_51 ();
 sg13g2_decap_4 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_fill_1 FILLER_32_139 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_189 ();
 sg13g2_decap_4 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_294 ();
 sg13g2_fill_2 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_327 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_fill_2 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_352 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_fill_1 FILLER_32_373 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_86 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_192 ();
 sg13g2_fill_1 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_243 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_258 ();
 sg13g2_fill_2 FILLER_33_317 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_fill_1 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_394 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_94 ();
 sg13g2_fill_2 FILLER_34_167 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_258 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_303 ();
 sg13g2_fill_2 FILLER_34_309 ();
 sg13g2_fill_1 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_73 ();
 sg13g2_fill_2 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_93 ();
 sg13g2_fill_2 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_fill_2 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_195 ();
 sg13g2_fill_2 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_26 ();
 sg13g2_fill_1 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_61 ();
 sg13g2_fill_2 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_2 FILLER_36_140 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_decap_8 FILLER_36_177 ();
 sg13g2_fill_2 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_190 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_decap_4 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_26 ();
 sg13g2_decap_8 FILLER_37_44 ();
 sg13g2_decap_4 FILLER_37_51 ();
 sg13g2_decap_4 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_199 ();
 sg13g2_fill_1 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_270 ();
 sg13g2_decap_8 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_fill_2 FILLER_37_309 ();
 sg13g2_fill_2 FILLER_37_324 ();
 sg13g2_fill_1 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_fill_2 FILLER_37_369 ();
 sg13g2_fill_1 FILLER_37_371 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_4 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_18 ();
 sg13g2_decap_8 FILLER_38_23 ();
 sg13g2_fill_2 FILLER_38_30 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_fill_2 FILLER_38_57 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_fill_2 FILLER_38_235 ();
 sg13g2_fill_2 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_259 ();
 sg13g2_fill_1 FILLER_38_261 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_2 FILLER_38_300 ();
 sg13g2_decap_4 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_4 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_339 ();
 sg13g2_fill_2 FILLER_38_361 ();
 sg13g2_fill_1 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_fill_1 FILLER_39_11 ();
 sg13g2_fill_2 FILLER_39_85 ();
 sg13g2_fill_2 FILLER_39_189 ();
 sg13g2_fill_1 FILLER_39_191 ();
 sg13g2_fill_1 FILLER_39_200 ();
 sg13g2_decap_4 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_243 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_fill_1 FILLER_39_284 ();
 sg13g2_fill_1 FILLER_39_290 ();
 sg13g2_decap_8 FILLER_39_316 ();
 sg13g2_decap_4 FILLER_39_323 ();
 sg13g2_fill_1 FILLER_39_332 ();
 sg13g2_fill_2 FILLER_39_373 ();
 sg13g2_fill_2 FILLER_39_380 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_51 ();
 sg13g2_fill_2 FILLER_40_87 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_fill_2 FILLER_40_151 ();
 sg13g2_fill_2 FILLER_40_227 ();
 sg13g2_decap_8 FILLER_40_272 ();
 sg13g2_decap_4 FILLER_40_279 ();
 sg13g2_fill_1 FILLER_40_317 ();
 sg13g2_fill_1 FILLER_40_344 ();
 sg13g2_fill_1 FILLER_40_355 ();
 sg13g2_fill_2 FILLER_40_377 ();
 sg13g2_fill_1 FILLER_40_379 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_29 ();
 sg13g2_fill_1 FILLER_41_31 ();
 sg13g2_fill_1 FILLER_41_45 ();
 sg13g2_fill_1 FILLER_41_127 ();
 sg13g2_fill_2 FILLER_41_133 ();
 sg13g2_fill_1 FILLER_41_135 ();
 sg13g2_fill_1 FILLER_41_157 ();
 sg13g2_fill_1 FILLER_41_173 ();
 sg13g2_fill_2 FILLER_41_192 ();
 sg13g2_fill_1 FILLER_41_194 ();
 sg13g2_fill_2 FILLER_41_218 ();
 sg13g2_fill_2 FILLER_41_282 ();
 sg13g2_fill_1 FILLER_41_298 ();
 sg13g2_fill_2 FILLER_41_303 ();
 sg13g2_fill_2 FILLER_41_321 ();
 sg13g2_fill_1 FILLER_41_323 ();
 sg13g2_fill_2 FILLER_41_395 ();
 sg13g2_fill_1 FILLER_41_397 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_4 ();
 sg13g2_decap_8 FILLER_42_24 ();
 sg13g2_decap_4 FILLER_42_31 ();
 sg13g2_fill_2 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_fill_2 FILLER_42_93 ();
 sg13g2_fill_1 FILLER_42_126 ();
 sg13g2_fill_2 FILLER_42_142 ();
 sg13g2_fill_1 FILLER_42_144 ();
 sg13g2_fill_1 FILLER_42_165 ();
 sg13g2_fill_2 FILLER_42_171 ();
 sg13g2_fill_2 FILLER_42_178 ();
 sg13g2_fill_1 FILLER_42_180 ();
 sg13g2_decap_4 FILLER_42_235 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_fill_1 FILLER_42_260 ();
 sg13g2_fill_1 FILLER_42_270 ();
 sg13g2_fill_2 FILLER_42_276 ();
 sg13g2_fill_1 FILLER_42_278 ();
 sg13g2_fill_2 FILLER_42_288 ();
 sg13g2_fill_2 FILLER_42_296 ();
 sg13g2_fill_1 FILLER_42_298 ();
 sg13g2_fill_1 FILLER_42_340 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_fill_2 FILLER_42_376 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_43_22 ();
 sg13g2_fill_1 FILLER_43_33 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_fill_2 FILLER_43_114 ();
 sg13g2_fill_1 FILLER_43_185 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_decap_4 FILLER_43_233 ();
 sg13g2_decap_4 FILLER_43_245 ();
 sg13g2_fill_2 FILLER_43_249 ();
 sg13g2_fill_1 FILLER_43_288 ();
 sg13g2_fill_2 FILLER_43_308 ();
 sg13g2_fill_1 FILLER_43_310 ();
 sg13g2_fill_2 FILLER_43_361 ();
 sg13g2_fill_1 FILLER_43_381 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_2 ();
 sg13g2_fill_1 FILLER_44_14 ();
 sg13g2_fill_2 FILLER_44_20 ();
 sg13g2_fill_1 FILLER_44_22 ();
 sg13g2_fill_1 FILLER_44_40 ();
 sg13g2_fill_2 FILLER_44_69 ();
 sg13g2_fill_1 FILLER_44_71 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_fill_2 FILLER_44_174 ();
 sg13g2_decap_8 FILLER_44_179 ();
 sg13g2_decap_8 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_193 ();
 sg13g2_decap_8 FILLER_44_200 ();
 sg13g2_decap_8 FILLER_44_207 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_fill_1 FILLER_44_229 ();
 sg13g2_decap_8 FILLER_44_242 ();
 sg13g2_fill_1 FILLER_44_335 ();
 sg13g2_fill_2 FILLER_44_344 ();
 sg13g2_fill_2 FILLER_44_358 ();
 sg13g2_fill_1 FILLER_44_380 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_27 ();
 sg13g2_fill_2 FILLER_45_36 ();
 sg13g2_fill_1 FILLER_45_61 ();
 sg13g2_fill_1 FILLER_45_75 ();
 sg13g2_fill_1 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_182 ();
 sg13g2_fill_1 FILLER_45_192 ();
 sg13g2_fill_2 FILLER_45_264 ();
 sg13g2_fill_2 FILLER_45_292 ();
 sg13g2_fill_2 FILLER_45_325 ();
 sg13g2_fill_2 FILLER_45_332 ();
 sg13g2_fill_1 FILLER_45_334 ();
 sg13g2_fill_2 FILLER_45_340 ();
 sg13g2_fill_1 FILLER_45_342 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_2 FILLER_46_12 ();
 sg13g2_fill_1 FILLER_46_22 ();
 sg13g2_fill_2 FILLER_46_38 ();
 sg13g2_fill_1 FILLER_46_40 ();
 sg13g2_fill_2 FILLER_46_49 ();
 sg13g2_fill_1 FILLER_46_51 ();
 sg13g2_fill_2 FILLER_46_66 ();
 sg13g2_fill_1 FILLER_46_68 ();
 sg13g2_fill_1 FILLER_46_74 ();
 sg13g2_fill_2 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_93 ();
 sg13g2_fill_1 FILLER_46_139 ();
 sg13g2_fill_1 FILLER_46_161 ();
 sg13g2_fill_1 FILLER_46_172 ();
 sg13g2_fill_2 FILLER_46_186 ();
 sg13g2_decap_4 FILLER_46_206 ();
 sg13g2_fill_2 FILLER_46_210 ();
 sg13g2_fill_2 FILLER_46_224 ();
 sg13g2_fill_1 FILLER_46_226 ();
 sg13g2_fill_1 FILLER_46_236 ();
 sg13g2_decap_4 FILLER_46_262 ();
 sg13g2_fill_1 FILLER_46_279 ();
 sg13g2_fill_1 FILLER_46_285 ();
 sg13g2_fill_2 FILLER_46_299 ();
 sg13g2_decap_4 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_318 ();
 sg13g2_fill_2 FILLER_46_336 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_fill_1 FILLER_46_382 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_43 ();
 sg13g2_fill_2 FILLER_47_49 ();
 sg13g2_fill_1 FILLER_47_51 ();
 sg13g2_fill_1 FILLER_47_150 ();
 sg13g2_fill_1 FILLER_47_201 ();
 sg13g2_fill_1 FILLER_47_207 ();
 sg13g2_decap_8 FILLER_47_233 ();
 sg13g2_fill_1 FILLER_47_240 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_263 ();
 sg13g2_decap_4 FILLER_47_283 ();
 sg13g2_fill_1 FILLER_47_287 ();
 sg13g2_fill_1 FILLER_47_294 ();
 sg13g2_fill_1 FILLER_47_303 ();
 sg13g2_decap_4 FILLER_47_308 ();
 sg13g2_fill_2 FILLER_47_317 ();
 sg13g2_fill_1 FILLER_47_330 ();
 sg13g2_fill_2 FILLER_47_365 ();
 sg13g2_fill_1 FILLER_47_367 ();
 sg13g2_fill_2 FILLER_47_376 ();
 sg13g2_fill_2 FILLER_47_388 ();
 sg13g2_fill_1 FILLER_47_390 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_12 ();
 sg13g2_fill_2 FILLER_48_28 ();
 sg13g2_fill_1 FILLER_48_30 ();
 sg13g2_fill_1 FILLER_48_36 ();
 sg13g2_fill_2 FILLER_48_56 ();
 sg13g2_fill_1 FILLER_48_58 ();
 sg13g2_fill_2 FILLER_48_65 ();
 sg13g2_fill_1 FILLER_48_105 ();
 sg13g2_fill_1 FILLER_48_120 ();
 sg13g2_fill_1 FILLER_48_184 ();
 sg13g2_fill_1 FILLER_48_214 ();
 sg13g2_decap_8 FILLER_48_240 ();
 sg13g2_decap_8 FILLER_48_247 ();
 sg13g2_decap_8 FILLER_48_254 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_fill_2 FILLER_48_269 ();
 sg13g2_fill_1 FILLER_48_271 ();
 sg13g2_decap_8 FILLER_48_276 ();
 sg13g2_fill_2 FILLER_48_288 ();
 sg13g2_fill_1 FILLER_48_290 ();
 sg13g2_fill_2 FILLER_48_300 ();
 sg13g2_fill_1 FILLER_48_302 ();
 sg13g2_fill_2 FILLER_48_328 ();
 sg13g2_fill_1 FILLER_48_330 ();
 sg13g2_fill_1 FILLER_48_336 ();
 sg13g2_fill_2 FILLER_48_362 ();
 sg13g2_fill_2 FILLER_48_376 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_2 ();
 sg13g2_fill_2 FILLER_49_19 ();
 sg13g2_fill_1 FILLER_49_26 ();
 sg13g2_fill_2 FILLER_49_65 ();
 sg13g2_fill_1 FILLER_49_75 ();
 sg13g2_fill_2 FILLER_49_102 ();
 sg13g2_fill_2 FILLER_49_140 ();
 sg13g2_fill_1 FILLER_49_142 ();
 sg13g2_fill_1 FILLER_49_202 ();
 sg13g2_fill_2 FILLER_49_212 ();
 sg13g2_decap_4 FILLER_49_242 ();
 sg13g2_fill_2 FILLER_49_246 ();
 sg13g2_fill_2 FILLER_49_262 ();
 sg13g2_fill_1 FILLER_49_264 ();
 sg13g2_decap_4 FILLER_49_284 ();
 sg13g2_fill_1 FILLER_49_288 ();
 sg13g2_fill_2 FILLER_49_309 ();
 sg13g2_fill_1 FILLER_49_311 ();
 sg13g2_fill_2 FILLER_49_319 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_fill_2 FILLER_49_350 ();
 sg13g2_fill_1 FILLER_49_352 ();
 sg13g2_fill_1 FILLER_49_362 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_57 ();
 sg13g2_fill_1 FILLER_50_59 ();
 sg13g2_fill_2 FILLER_50_125 ();
 sg13g2_fill_2 FILLER_50_163 ();
 sg13g2_fill_2 FILLER_50_179 ();
 sg13g2_fill_2 FILLER_50_219 ();
 sg13g2_fill_1 FILLER_50_221 ();
 sg13g2_fill_2 FILLER_50_265 ();
 sg13g2_fill_1 FILLER_50_319 ();
 sg13g2_fill_2 FILLER_50_326 ();
 sg13g2_fill_2 FILLER_50_335 ();
 sg13g2_fill_2 FILLER_50_363 ();
 sg13g2_fill_1 FILLER_50_365 ();
 sg13g2_fill_1 FILLER_50_377 ();
 sg13g2_fill_2 FILLER_50_383 ();
 sg13g2_fill_2 FILLER_50_390 ();
 sg13g2_fill_1 FILLER_50_392 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_fill_2 FILLER_51_25 ();
 sg13g2_fill_1 FILLER_51_27 ();
 sg13g2_fill_2 FILLER_51_65 ();
 sg13g2_fill_2 FILLER_51_72 ();
 sg13g2_fill_2 FILLER_51_133 ();
 sg13g2_fill_1 FILLER_51_144 ();
 sg13g2_fill_2 FILLER_51_172 ();
 sg13g2_fill_1 FILLER_51_174 ();
 sg13g2_fill_2 FILLER_51_180 ();
 sg13g2_fill_1 FILLER_51_182 ();
 sg13g2_fill_2 FILLER_51_232 ();
 sg13g2_fill_2 FILLER_51_283 ();
 sg13g2_fill_1 FILLER_51_285 ();
 sg13g2_fill_1 FILLER_51_314 ();
 sg13g2_fill_2 FILLER_51_328 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_33 ();
 sg13g2_fill_2 FILLER_52_53 ();
 sg13g2_fill_1 FILLER_52_55 ();
 sg13g2_fill_2 FILLER_52_65 ();
 sg13g2_fill_2 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_173 ();
 sg13g2_fill_2 FILLER_52_187 ();
 sg13g2_fill_1 FILLER_52_198 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_decap_8 FILLER_52_210 ();
 sg13g2_fill_2 FILLER_52_217 ();
 sg13g2_fill_1 FILLER_52_219 ();
 sg13g2_decap_4 FILLER_52_233 ();
 sg13g2_fill_2 FILLER_52_237 ();
 sg13g2_fill_1 FILLER_52_283 ();
 sg13g2_fill_2 FILLER_52_317 ();
 sg13g2_fill_1 FILLER_52_319 ();
 sg13g2_fill_2 FILLER_52_330 ();
 sg13g2_fill_1 FILLER_52_362 ();
 sg13g2_fill_1 FILLER_53_44 ();
 sg13g2_fill_1 FILLER_53_66 ();
 sg13g2_fill_1 FILLER_53_82 ();
 sg13g2_fill_2 FILLER_53_160 ();
 sg13g2_fill_1 FILLER_53_162 ();
 sg13g2_decap_4 FILLER_53_206 ();
 sg13g2_fill_2 FILLER_53_210 ();
 sg13g2_fill_1 FILLER_53_243 ();
 sg13g2_fill_1 FILLER_53_262 ();
 sg13g2_fill_1 FILLER_53_326 ();
 sg13g2_fill_1 FILLER_53_339 ();
 sg13g2_fill_2 FILLER_53_351 ();
 sg13g2_fill_1 FILLER_53_353 ();
 sg13g2_fill_2 FILLER_53_395 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_25 ();
 sg13g2_fill_1 FILLER_54_40 ();
 sg13g2_fill_1 FILLER_54_50 ();
 sg13g2_fill_1 FILLER_54_103 ();
 sg13g2_fill_2 FILLER_54_146 ();
 sg13g2_fill_2 FILLER_54_163 ();
 sg13g2_fill_1 FILLER_54_165 ();
 sg13g2_fill_2 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_260 ();
 sg13g2_fill_2 FILLER_54_335 ();
 sg13g2_fill_1 FILLER_54_337 ();
 sg13g2_fill_1 FILLER_54_385 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_24 ();
 sg13g2_fill_1 FILLER_55_26 ();
 sg13g2_fill_2 FILLER_55_43 ();
 sg13g2_fill_1 FILLER_55_45 ();
 sg13g2_fill_1 FILLER_55_54 ();
 sg13g2_fill_1 FILLER_55_76 ();
 sg13g2_fill_1 FILLER_55_94 ();
 sg13g2_fill_2 FILLER_55_135 ();
 sg13g2_fill_1 FILLER_55_137 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_2 FILLER_55_200 ();
 sg13g2_fill_1 FILLER_55_301 ();
 sg13g2_fill_1 FILLER_55_320 ();
 sg13g2_fill_2 FILLER_55_343 ();
 sg13g2_fill_1 FILLER_55_345 ();
 sg13g2_fill_1 FILLER_55_359 ();
 sg13g2_fill_2 FILLER_55_370 ();
 sg13g2_fill_1 FILLER_55_372 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_fill_2 FILLER_56_25 ();
 sg13g2_fill_1 FILLER_56_27 ();
 sg13g2_fill_1 FILLER_56_37 ();
 sg13g2_fill_1 FILLER_56_43 ();
 sg13g2_fill_1 FILLER_56_80 ();
 sg13g2_fill_1 FILLER_56_144 ();
 sg13g2_fill_1 FILLER_56_154 ();
 sg13g2_fill_2 FILLER_56_163 ();
 sg13g2_fill_2 FILLER_56_170 ();
 sg13g2_fill_1 FILLER_56_182 ();
 sg13g2_fill_2 FILLER_56_196 ();
 sg13g2_fill_1 FILLER_56_227 ();
 sg13g2_fill_2 FILLER_56_275 ();
 sg13g2_fill_1 FILLER_56_277 ();
 sg13g2_fill_2 FILLER_56_304 ();
 sg13g2_fill_2 FILLER_56_314 ();
 sg13g2_fill_1 FILLER_56_316 ();
 sg13g2_fill_1 FILLER_56_329 ();
 sg13g2_fill_1 FILLER_56_344 ();
 sg13g2_fill_1 FILLER_56_357 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_1 FILLER_57_21 ();
 sg13g2_fill_2 FILLER_57_28 ();
 sg13g2_fill_1 FILLER_57_30 ();
 sg13g2_fill_2 FILLER_57_93 ();
 sg13g2_fill_1 FILLER_57_95 ();
 sg13g2_fill_2 FILLER_57_130 ();
 sg13g2_fill_1 FILLER_57_132 ();
 sg13g2_fill_2 FILLER_57_200 ();
 sg13g2_fill_1 FILLER_57_202 ();
 sg13g2_fill_2 FILLER_57_220 ();
 sg13g2_fill_1 FILLER_57_226 ();
 sg13g2_fill_2 FILLER_57_245 ();
 sg13g2_fill_1 FILLER_57_259 ();
 sg13g2_fill_2 FILLER_57_349 ();
 sg13g2_fill_1 FILLER_57_368 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_fill_1 FILLER_58_36 ();
 sg13g2_fill_2 FILLER_58_70 ();
 sg13g2_fill_2 FILLER_58_117 ();
 sg13g2_fill_2 FILLER_58_123 ();
 sg13g2_fill_1 FILLER_58_148 ();
 sg13g2_fill_1 FILLER_58_216 ();
 sg13g2_fill_1 FILLER_58_222 ();
 sg13g2_fill_2 FILLER_58_247 ();
 sg13g2_fill_1 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_267 ();
 sg13g2_fill_2 FILLER_58_354 ();
 sg13g2_fill_1 FILLER_58_383 ();
 sg13g2_fill_2 FILLER_58_391 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_2 FILLER_59_135 ();
 sg13g2_fill_2 FILLER_59_142 ();
 sg13g2_fill_1 FILLER_59_167 ();
 sg13g2_fill_1 FILLER_59_178 ();
 sg13g2_fill_2 FILLER_59_183 ();
 sg13g2_decap_8 FILLER_59_201 ();
 sg13g2_fill_2 FILLER_59_208 ();
 sg13g2_fill_2 FILLER_59_234 ();
 sg13g2_fill_2 FILLER_59_244 ();
 sg13g2_fill_2 FILLER_59_324 ();
 sg13g2_fill_2 FILLER_59_358 ();
 sg13g2_fill_1 FILLER_59_360 ();
 sg13g2_fill_1 FILLER_59_373 ();
 sg13g2_fill_2 FILLER_60_53 ();
 sg13g2_fill_2 FILLER_60_137 ();
 sg13g2_fill_1 FILLER_60_249 ();
 sg13g2_fill_2 FILLER_60_289 ();
 sg13g2_fill_1 FILLER_60_291 ();
 sg13g2_fill_1 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_371 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_fill_1 FILLER_61_33 ();
 sg13g2_fill_2 FILLER_61_39 ();
 sg13g2_fill_2 FILLER_61_53 ();
 sg13g2_fill_2 FILLER_61_80 ();
 sg13g2_fill_2 FILLER_61_102 ();
 sg13g2_fill_2 FILLER_61_126 ();
 sg13g2_fill_2 FILLER_61_143 ();
 sg13g2_fill_2 FILLER_61_155 ();
 sg13g2_fill_1 FILLER_61_157 ();
 sg13g2_fill_2 FILLER_61_303 ();
 sg13g2_fill_1 FILLER_61_305 ();
 sg13g2_fill_2 FILLER_61_359 ();
 sg13g2_fill_1 FILLER_61_373 ();
 sg13g2_fill_2 FILLER_61_390 ();
 sg13g2_fill_1 FILLER_61_392 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_5 ();
 sg13g2_fill_1 FILLER_62_17 ();
 sg13g2_fill_1 FILLER_62_32 ();
 sg13g2_fill_2 FILLER_62_74 ();
 sg13g2_fill_2 FILLER_62_167 ();
 sg13g2_fill_2 FILLER_62_178 ();
 sg13g2_fill_1 FILLER_62_180 ();
 sg13g2_fill_1 FILLER_62_191 ();
 sg13g2_fill_1 FILLER_62_220 ();
 sg13g2_fill_2 FILLER_62_234 ();
 sg13g2_fill_2 FILLER_62_259 ();
 sg13g2_fill_1 FILLER_62_261 ();
 sg13g2_fill_2 FILLER_62_266 ();
 sg13g2_fill_2 FILLER_62_272 ();
 sg13g2_fill_2 FILLER_62_294 ();
 sg13g2_fill_2 FILLER_62_317 ();
 sg13g2_fill_1 FILLER_62_319 ();
 sg13g2_fill_1 FILLER_62_331 ();
 sg13g2_fill_2 FILLER_62_347 ();
 sg13g2_fill_1 FILLER_62_349 ();
 sg13g2_fill_2 FILLER_62_371 ();
 sg13g2_fill_1 FILLER_62_373 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_11 ();
 sg13g2_decap_8 FILLER_63_18 ();
 sg13g2_fill_1 FILLER_63_25 ();
 sg13g2_fill_1 FILLER_63_41 ();
 sg13g2_fill_1 FILLER_63_99 ();
 sg13g2_fill_2 FILLER_63_110 ();
 sg13g2_fill_1 FILLER_63_205 ();
 sg13g2_fill_1 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_237 ();
 sg13g2_fill_1 FILLER_63_246 ();
 sg13g2_fill_2 FILLER_63_261 ();
 sg13g2_fill_1 FILLER_63_263 ();
 sg13g2_fill_1 FILLER_63_269 ();
 sg13g2_fill_2 FILLER_63_288 ();
 sg13g2_fill_2 FILLER_63_319 ();
 sg13g2_fill_2 FILLER_63_340 ();
 sg13g2_fill_1 FILLER_63_342 ();
 sg13g2_fill_1 FILLER_63_351 ();
 sg13g2_fill_1 FILLER_63_370 ();
 sg13g2_fill_1 FILLER_63_379 ();
 sg13g2_fill_1 FILLER_64_26 ();
 sg13g2_fill_2 FILLER_64_71 ();
 sg13g2_fill_1 FILLER_64_163 ();
 sg13g2_fill_1 FILLER_64_174 ();
 sg13g2_fill_2 FILLER_64_245 ();
 sg13g2_fill_2 FILLER_64_259 ();
 sg13g2_fill_2 FILLER_64_272 ();
 sg13g2_fill_2 FILLER_64_402 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_28 ();
 sg13g2_fill_2 FILLER_65_37 ();
 sg13g2_fill_2 FILLER_65_94 ();
 sg13g2_fill_1 FILLER_65_129 ();
 sg13g2_fill_2 FILLER_65_135 ();
 sg13g2_fill_1 FILLER_65_152 ();
 sg13g2_fill_2 FILLER_65_207 ();
 sg13g2_fill_1 FILLER_65_209 ();
 sg13g2_fill_2 FILLER_65_218 ();
 sg13g2_fill_2 FILLER_65_266 ();
 sg13g2_fill_1 FILLER_65_268 ();
 sg13g2_fill_1 FILLER_65_292 ();
 sg13g2_fill_2 FILLER_65_303 ();
 sg13g2_fill_2 FILLER_65_326 ();
 sg13g2_fill_1 FILLER_65_328 ();
 sg13g2_fill_1 FILLER_65_361 ();
 sg13g2_fill_2 FILLER_65_373 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_29 ();
 sg13g2_fill_2 FILLER_66_73 ();
 sg13g2_fill_2 FILLER_66_83 ();
 sg13g2_fill_1 FILLER_66_85 ();
 sg13g2_fill_2 FILLER_66_96 ();
 sg13g2_fill_1 FILLER_66_103 ();
 sg13g2_fill_2 FILLER_66_123 ();
 sg13g2_fill_2 FILLER_66_138 ();
 sg13g2_fill_2 FILLER_66_159 ();
 sg13g2_fill_1 FILLER_66_202 ();
 sg13g2_fill_1 FILLER_66_214 ();
 sg13g2_fill_2 FILLER_66_246 ();
 sg13g2_fill_1 FILLER_66_248 ();
 sg13g2_fill_2 FILLER_66_272 ();
 sg13g2_fill_1 FILLER_66_274 ();
 sg13g2_fill_2 FILLER_66_295 ();
 sg13g2_fill_1 FILLER_66_297 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_363 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_fill_2 FILLER_67_116 ();
 sg13g2_fill_1 FILLER_67_145 ();
 sg13g2_fill_2 FILLER_67_165 ();
 sg13g2_fill_1 FILLER_67_186 ();
 sg13g2_fill_2 FILLER_67_192 ();
 sg13g2_fill_2 FILLER_67_202 ();
 sg13g2_fill_2 FILLER_67_213 ();
 sg13g2_fill_1 FILLER_67_215 ();
 sg13g2_fill_1 FILLER_67_236 ();
 sg13g2_fill_1 FILLER_67_247 ();
 sg13g2_fill_1 FILLER_67_263 ();
 sg13g2_fill_2 FILLER_67_273 ();
 sg13g2_fill_1 FILLER_67_275 ();
 sg13g2_fill_2 FILLER_67_304 ();
 sg13g2_fill_2 FILLER_67_318 ();
 sg13g2_fill_1 FILLER_67_320 ();
 sg13g2_fill_1 FILLER_67_332 ();
 sg13g2_fill_2 FILLER_67_346 ();
 sg13g2_fill_1 FILLER_67_348 ();
 sg13g2_fill_1 FILLER_67_362 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_fill_1 FILLER_68_78 ();
 sg13g2_fill_1 FILLER_68_100 ();
 sg13g2_fill_1 FILLER_68_127 ();
 sg13g2_fill_1 FILLER_68_137 ();
 sg13g2_fill_2 FILLER_68_143 ();
 sg13g2_fill_1 FILLER_68_219 ();
 sg13g2_fill_2 FILLER_68_315 ();
 sg13g2_fill_1 FILLER_68_348 ();
 sg13g2_fill_1 FILLER_68_357 ();
 sg13g2_fill_1 FILLER_68_375 ();
 sg13g2_fill_2 FILLER_68_381 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_19 ();
 sg13g2_fill_2 FILLER_69_37 ();
 sg13g2_fill_1 FILLER_69_39 ();
 sg13g2_fill_2 FILLER_69_44 ();
 sg13g2_fill_1 FILLER_69_46 ();
 sg13g2_fill_2 FILLER_69_105 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_fill_2 FILLER_69_231 ();
 sg13g2_fill_1 FILLER_69_233 ();
 sg13g2_fill_1 FILLER_69_247 ();
 sg13g2_fill_1 FILLER_69_308 ();
 sg13g2_fill_2 FILLER_69_314 ();
 sg13g2_fill_1 FILLER_69_354 ();
 sg13g2_fill_2 FILLER_69_380 ();
 sg13g2_fill_2 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_38 ();
 sg13g2_fill_2 FILLER_70_70 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_214 ();
 sg13g2_fill_1 FILLER_70_247 ();
 sg13g2_fill_2 FILLER_70_282 ();
 sg13g2_fill_1 FILLER_70_310 ();
 sg13g2_fill_2 FILLER_70_364 ();
 sg13g2_fill_2 FILLER_70_380 ();
 sg13g2_fill_1 FILLER_71_31 ();
 sg13g2_fill_2 FILLER_71_125 ();
 sg13g2_fill_1 FILLER_71_142 ();
 sg13g2_fill_1 FILLER_71_158 ();
 sg13g2_fill_2 FILLER_71_172 ();
 sg13g2_fill_1 FILLER_71_232 ();
 sg13g2_fill_2 FILLER_71_238 ();
 sg13g2_fill_1 FILLER_71_264 ();
 sg13g2_fill_2 FILLER_71_296 ();
 sg13g2_fill_1 FILLER_71_298 ();
 sg13g2_fill_1 FILLER_71_368 ();
 sg13g2_fill_2 FILLER_71_384 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_fill_2 FILLER_72_89 ();
 sg13g2_fill_2 FILLER_72_112 ();
 sg13g2_fill_2 FILLER_72_142 ();
 sg13g2_fill_1 FILLER_72_164 ();
 sg13g2_fill_1 FILLER_72_209 ();
 sg13g2_fill_2 FILLER_72_223 ();
 sg13g2_fill_1 FILLER_72_225 ();
 sg13g2_fill_2 FILLER_72_293 ();
 sg13g2_fill_2 FILLER_72_336 ();
 sg13g2_fill_2 FILLER_72_363 ();
 sg13g2_fill_2 FILLER_72_373 ();
 sg13g2_fill_1 FILLER_72_375 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_2 ();
 sg13g2_fill_2 FILLER_73_78 ();
 sg13g2_fill_1 FILLER_73_98 ();
 sg13g2_fill_2 FILLER_73_130 ();
 sg13g2_fill_1 FILLER_73_194 ();
 sg13g2_fill_2 FILLER_73_208 ();
 sg13g2_fill_1 FILLER_73_210 ();
 sg13g2_fill_2 FILLER_73_245 ();
 sg13g2_fill_1 FILLER_73_283 ();
 sg13g2_fill_2 FILLER_73_312 ();
 sg13g2_fill_2 FILLER_73_335 ();
 sg13g2_fill_1 FILLER_73_337 ();
 sg13g2_fill_2 FILLER_73_365 ();
 sg13g2_fill_2 FILLER_73_398 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_44 ();
 sg13g2_fill_2 FILLER_74_105 ();
 sg13g2_fill_2 FILLER_74_133 ();
 sg13g2_fill_2 FILLER_74_148 ();
 sg13g2_fill_1 FILLER_74_170 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_fill_2 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_236 ();
 sg13g2_fill_2 FILLER_74_277 ();
 sg13g2_fill_1 FILLER_74_279 ();
 sg13g2_fill_1 FILLER_74_319 ();
 sg13g2_fill_1 FILLER_74_336 ();
 sg13g2_fill_1 FILLER_74_366 ();
 sg13g2_fill_1 FILLER_74_371 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_79 ();
 sg13g2_fill_2 FILLER_75_96 ();
 sg13g2_fill_2 FILLER_75_113 ();
 sg13g2_fill_2 FILLER_75_138 ();
 sg13g2_fill_1 FILLER_75_144 ();
 sg13g2_fill_2 FILLER_75_162 ();
 sg13g2_fill_1 FILLER_75_190 ();
 sg13g2_fill_1 FILLER_75_231 ();
 sg13g2_fill_2 FILLER_75_294 ();
 sg13g2_fill_2 FILLER_75_309 ();
 sg13g2_fill_1 FILLER_75_311 ();
 sg13g2_fill_2 FILLER_75_318 ();
 sg13g2_fill_1 FILLER_75_366 ();
 sg13g2_fill_2 FILLER_75_380 ();
 sg13g2_fill_1 FILLER_75_382 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_40 ();
 sg13g2_fill_1 FILLER_76_82 ();
 sg13g2_fill_1 FILLER_76_128 ();
 sg13g2_fill_1 FILLER_76_139 ();
 sg13g2_fill_2 FILLER_76_155 ();
 sg13g2_fill_1 FILLER_76_157 ();
 sg13g2_fill_1 FILLER_76_166 ();
 sg13g2_fill_2 FILLER_76_178 ();
 sg13g2_fill_2 FILLER_76_197 ();
 sg13g2_fill_1 FILLER_76_199 ();
 sg13g2_fill_1 FILLER_76_326 ();
 sg13g2_fill_2 FILLER_76_339 ();
 sg13g2_fill_1 FILLER_76_341 ();
 sg13g2_fill_2 FILLER_76_365 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_79 ();
 sg13g2_fill_1 FILLER_77_111 ();
 sg13g2_fill_2 FILLER_77_154 ();
 sg13g2_fill_1 FILLER_77_156 ();
 sg13g2_fill_2 FILLER_77_169 ();
 sg13g2_fill_1 FILLER_77_181 ();
 sg13g2_fill_1 FILLER_77_243 ();
 sg13g2_fill_1 FILLER_77_280 ();
 sg13g2_fill_2 FILLER_77_293 ();
 sg13g2_fill_1 FILLER_77_295 ();
 sg13g2_fill_1 FILLER_77_320 ();
 sg13g2_fill_2 FILLER_77_345 ();
 sg13g2_fill_1 FILLER_77_347 ();
 sg13g2_fill_1 FILLER_77_366 ();
 sg13g2_fill_2 FILLER_77_375 ();
 sg13g2_fill_1 FILLER_77_377 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_70 ();
 sg13g2_fill_1 FILLER_78_98 ();
 sg13g2_fill_2 FILLER_78_135 ();
 sg13g2_fill_1 FILLER_78_143 ();
 sg13g2_fill_1 FILLER_78_153 ();
 sg13g2_fill_1 FILLER_78_202 ();
 sg13g2_fill_2 FILLER_78_234 ();
 sg13g2_fill_2 FILLER_78_294 ();
 sg13g2_fill_2 FILLER_78_336 ();
 sg13g2_fill_2 FILLER_78_361 ();
 sg13g2_fill_1 FILLER_78_363 ();
 sg13g2_fill_2 FILLER_78_370 ();
 sg13g2_fill_1 FILLER_78_372 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_132 ();
 sg13g2_fill_1 FILLER_79_341 ();
 sg13g2_fill_2 FILLER_79_354 ();
 sg13g2_fill_1 FILLER_79_382 ();
 sg13g2_fill_1 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_44 ();
 sg13g2_fill_1 FILLER_80_46 ();
 sg13g2_fill_2 FILLER_80_99 ();
 sg13g2_fill_2 FILLER_80_110 ();
 sg13g2_fill_1 FILLER_80_112 ();
 sg13g2_fill_2 FILLER_80_121 ();
 sg13g2_fill_2 FILLER_80_158 ();
 sg13g2_fill_2 FILLER_80_164 ();
 sg13g2_fill_1 FILLER_80_275 ();
 sg13g2_fill_1 FILLER_80_328 ();
 sg13g2_fill_1 FILLER_80_343 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_fill_2 FILLER_80_376 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net305;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
endmodule

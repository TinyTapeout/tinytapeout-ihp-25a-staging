module tt_um_cattuto_sr_latch (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire ntrig;
 wire shift;
 wire \shift_reg[0].genblk1.latch.clk ;
 wire \shift_reg[0].genblk1.latch.q ;
 wire \shift_reg[100].genblk1.genblk1.latch.clk ;
 wire \shift_reg[100].genblk1.genblk1.latch.clkout ;
 wire \shift_reg[100].genblk1.genblk1.latch.d ;
 wire \shift_reg[100].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[100].genblk1.genblk1.latch.q ;
 wire \shift_reg[101].genblk1.genblk1.latch.clk ;
 wire \shift_reg[101].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[101].genblk1.genblk1.latch.q ;
 wire \shift_reg[102].genblk1.genblk1.latch.clk ;
 wire \shift_reg[102].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[102].genblk1.genblk1.latch.q ;
 wire \shift_reg[103].genblk1.genblk1.latch.clk ;
 wire \shift_reg[103].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[103].genblk1.genblk1.latch.q ;
 wire \shift_reg[104].genblk1.genblk1.latch.clk ;
 wire \shift_reg[104].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[104].genblk1.genblk1.latch.q ;
 wire \shift_reg[105].genblk1.genblk1.latch.clk ;
 wire \shift_reg[105].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[105].genblk1.genblk1.latch.q ;
 wire \shift_reg[106].genblk1.genblk1.latch.clk ;
 wire \shift_reg[106].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[106].genblk1.genblk1.latch.q ;
 wire \shift_reg[107].genblk1.genblk1.latch.clk ;
 wire \shift_reg[107].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[107].genblk1.genblk1.latch.q ;
 wire \shift_reg[108].genblk1.genblk1.latch.clk ;
 wire \shift_reg[108].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[108].genblk1.genblk1.latch.q ;
 wire \shift_reg[109].genblk1.genblk1.latch.clk ;
 wire \shift_reg[109].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[109].genblk1.genblk1.latch.q ;
 wire \shift_reg[10].genblk1.genblk1.latch.clk ;
 wire \shift_reg[10].genblk1.genblk1.latch.clkout ;
 wire \shift_reg[10].genblk1.genblk1.latch.d ;
 wire \shift_reg[10].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[10].genblk1.genblk1.latch.q ;
 wire \shift_reg[110].genblk1.genblk1.latch.clk ;
 wire \shift_reg[110].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[110].genblk1.genblk1.latch.q ;
 wire \shift_reg[111].genblk1.genblk1.latch.clk ;
 wire \shift_reg[111].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[111].genblk1.genblk1.latch.q ;
 wire \shift_reg[112].genblk1.genblk1.latch.clk ;
 wire \shift_reg[112].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[112].genblk1.genblk1.latch.q ;
 wire \shift_reg[113].genblk1.genblk1.latch.clk ;
 wire \shift_reg[113].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[113].genblk1.genblk1.latch.q ;
 wire \shift_reg[114].genblk1.genblk1.latch.clk ;
 wire \shift_reg[114].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[114].genblk1.genblk1.latch.q ;
 wire \shift_reg[115].genblk1.genblk1.latch.clk ;
 wire \shift_reg[115].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[115].genblk1.genblk1.latch.q ;
 wire \shift_reg[116].genblk1.genblk1.latch.clk ;
 wire \shift_reg[116].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[116].genblk1.genblk1.latch.q ;
 wire \shift_reg[117].genblk1.genblk1.latch.clk ;
 wire \shift_reg[117].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[117].genblk1.genblk1.latch.q ;
 wire \shift_reg[118].genblk1.genblk1.latch.clk ;
 wire \shift_reg[118].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[118].genblk1.genblk1.latch.q ;
 wire \shift_reg[119].genblk1.genblk1.latch.clk ;
 wire \shift_reg[119].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[119].genblk1.genblk1.latch.q ;
 wire \shift_reg[11].genblk1.genblk1.latch.clk ;
 wire \shift_reg[11].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[11].genblk1.genblk1.latch.q ;
 wire \shift_reg[120].genblk1.genblk1.latch.clk ;
 wire \shift_reg[120].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[120].genblk1.genblk1.latch.q ;
 wire \shift_reg[121].genblk1.genblk1.latch.clk ;
 wire \shift_reg[121].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[121].genblk1.genblk1.latch.q ;
 wire \shift_reg[122].genblk1.genblk1.latch.clk ;
 wire \shift_reg[122].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[122].genblk1.genblk1.latch.q ;
 wire \shift_reg[123].genblk1.genblk1.latch.clk ;
 wire \shift_reg[123].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[123].genblk1.genblk1.latch.q ;
 wire \shift_reg[124].genblk1.genblk1.latch.clk ;
 wire \shift_reg[124].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[124].genblk1.genblk1.latch.q ;
 wire \shift_reg[125].genblk1.genblk1.latch.clk ;
 wire \shift_reg[125].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[125].genblk1.genblk1.latch.q ;
 wire \shift_reg[126].genblk1.genblk1.latch.clk ;
 wire \shift_reg[126].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[126].genblk1.genblk1.latch.q ;
 wire \shift_reg[127].genblk1.genblk1.latch.clk ;
 wire \shift_reg[127].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[127].genblk1.genblk1.latch.q ;
 wire \shift_reg[128].genblk1.genblk1.latch.clk ;
 wire \shift_reg[128].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[128].genblk1.genblk1.latch.q ;
 wire \shift_reg[129].genblk1.genblk1.latch.clk ;
 wire \shift_reg[129].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[129].genblk1.genblk1.latch.q ;
 wire \shift_reg[12].genblk1.genblk1.latch.clk ;
 wire \shift_reg[12].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[12].genblk1.genblk1.latch.q ;
 wire \shift_reg[130].genblk1.genblk1.latch.clk ;
 wire \shift_reg[130].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[130].genblk1.genblk1.latch.q ;
 wire \shift_reg[131].genblk1.genblk1.latch.clk ;
 wire \shift_reg[131].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[131].genblk1.genblk1.latch.q ;
 wire \shift_reg[132].genblk1.genblk1.latch.clk ;
 wire \shift_reg[132].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[132].genblk1.genblk1.latch.q ;
 wire \shift_reg[133].genblk1.genblk1.latch.clk ;
 wire \shift_reg[133].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[133].genblk1.genblk1.latch.q ;
 wire \shift_reg[134].genblk1.genblk1.latch.clk ;
 wire \shift_reg[134].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[134].genblk1.genblk1.latch.q ;
 wire \shift_reg[135].genblk1.genblk1.latch.clk ;
 wire \shift_reg[135].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[135].genblk1.genblk1.latch.q ;
 wire \shift_reg[136].genblk1.genblk1.latch.clk ;
 wire \shift_reg[136].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[136].genblk1.genblk1.latch.q ;
 wire \shift_reg[137].genblk1.genblk1.latch.clk ;
 wire \shift_reg[137].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[137].genblk1.genblk1.latch.q ;
 wire \shift_reg[138].genblk1.genblk1.latch.clk ;
 wire \shift_reg[138].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[138].genblk1.genblk1.latch.q ;
 wire \shift_reg[139].genblk1.genblk1.latch.clk ;
 wire \shift_reg[139].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[139].genblk1.genblk1.latch.q ;
 wire \shift_reg[13].genblk1.genblk1.latch.clk ;
 wire \shift_reg[13].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[13].genblk1.genblk1.latch.q ;
 wire \shift_reg[140].genblk1.genblk1.latch.clk ;
 wire \shift_reg[140].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[140].genblk1.genblk1.latch.q ;
 wire \shift_reg[141].genblk1.genblk1.latch.clk ;
 wire \shift_reg[141].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[141].genblk1.genblk1.latch.q ;
 wire \shift_reg[142].genblk1.genblk1.latch.clk ;
 wire \shift_reg[142].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[142].genblk1.genblk1.latch.q ;
 wire \shift_reg[143].genblk1.genblk1.latch.clk ;
 wire \shift_reg[143].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[143].genblk1.genblk1.latch.q ;
 wire \shift_reg[144].genblk1.genblk1.latch.clk ;
 wire \shift_reg[144].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[144].genblk1.genblk1.latch.q ;
 wire \shift_reg[145].genblk1.genblk1.latch.clk ;
 wire \shift_reg[145].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[145].genblk1.genblk1.latch.q ;
 wire \shift_reg[146].genblk1.genblk1.latch.clk ;
 wire \shift_reg[146].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[146].genblk1.genblk1.latch.q ;
 wire \shift_reg[147].genblk1.genblk1.latch.clk ;
 wire \shift_reg[147].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[147].genblk1.genblk1.latch.q ;
 wire \shift_reg[148].genblk1.genblk1.latch.clk ;
 wire \shift_reg[148].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[148].genblk1.genblk1.latch.q ;
 wire \shift_reg[149].genblk1.genblk1.latch.clk ;
 wire \shift_reg[149].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[149].genblk1.genblk1.latch.q ;
 wire \shift_reg[14].genblk1.genblk1.latch.clk ;
 wire \shift_reg[14].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[14].genblk1.genblk1.latch.q ;
 wire \shift_reg[150].genblk1.genblk1.latch.clk ;
 wire \shift_reg[150].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[150].genblk1.genblk1.latch.q ;
 wire \shift_reg[151].genblk1.genblk1.latch.clk ;
 wire \shift_reg[151].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[151].genblk1.genblk1.latch.q ;
 wire \shift_reg[152].genblk1.genblk1.latch.clk ;
 wire \shift_reg[152].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[152].genblk1.genblk1.latch.q ;
 wire \shift_reg[153].genblk1.genblk1.latch.clk ;
 wire \shift_reg[153].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[153].genblk1.genblk1.latch.q ;
 wire \shift_reg[154].genblk1.genblk1.latch.clk ;
 wire \shift_reg[154].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[154].genblk1.genblk1.latch.q ;
 wire \shift_reg[155].genblk1.genblk1.latch.clk ;
 wire \shift_reg[155].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[155].genblk1.genblk1.latch.q ;
 wire \shift_reg[156].genblk1.genblk1.latch.clk ;
 wire \shift_reg[156].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[156].genblk1.genblk1.latch.q ;
 wire \shift_reg[157].genblk1.genblk1.latch.clk ;
 wire \shift_reg[157].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[157].genblk1.genblk1.latch.q ;
 wire \shift_reg[158].genblk1.genblk1.latch.clk ;
 wire \shift_reg[158].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[158].genblk1.genblk1.latch.q ;
 wire \shift_reg[159].genblk1.genblk1.latch.clk ;
 wire \shift_reg[159].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[159].genblk1.genblk1.latch.q ;
 wire \shift_reg[15].genblk1.genblk1.latch.clk ;
 wire \shift_reg[15].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[15].genblk1.genblk1.latch.q ;
 wire \shift_reg[160].genblk1.genblk1.latch.clk ;
 wire \shift_reg[160].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[160].genblk1.genblk1.latch.q ;
 wire \shift_reg[161].genblk1.genblk1.latch.clk ;
 wire \shift_reg[161].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[161].genblk1.genblk1.latch.q ;
 wire \shift_reg[162].genblk1.genblk1.latch.clk ;
 wire \shift_reg[162].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[162].genblk1.genblk1.latch.q ;
 wire \shift_reg[163].genblk1.genblk1.latch.clk ;
 wire \shift_reg[163].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[163].genblk1.genblk1.latch.q ;
 wire \shift_reg[164].genblk1.genblk1.latch.clk ;
 wire \shift_reg[164].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[164].genblk1.genblk1.latch.q ;
 wire \shift_reg[165].genblk1.genblk1.latch.clk ;
 wire \shift_reg[165].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[165].genblk1.genblk1.latch.q ;
 wire \shift_reg[166].genblk1.genblk1.latch.clk ;
 wire \shift_reg[166].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[166].genblk1.genblk1.latch.q ;
 wire \shift_reg[167].genblk1.genblk1.latch.clk ;
 wire \shift_reg[167].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[167].genblk1.genblk1.latch.q ;
 wire \shift_reg[168].genblk1.genblk1.latch.clk ;
 wire \shift_reg[168].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[168].genblk1.genblk1.latch.q ;
 wire \shift_reg[169].genblk1.genblk1.latch.clk ;
 wire \shift_reg[169].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[169].genblk1.genblk1.latch.q ;
 wire \shift_reg[16].genblk1.genblk1.latch.clk ;
 wire \shift_reg[16].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[16].genblk1.genblk1.latch.q ;
 wire \shift_reg[170].genblk1.genblk1.latch.clk ;
 wire \shift_reg[170].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[170].genblk1.genblk1.latch.q ;
 wire \shift_reg[171].genblk1.genblk1.latch.clk ;
 wire \shift_reg[171].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[171].genblk1.genblk1.latch.q ;
 wire \shift_reg[172].genblk1.genblk1.latch.clk ;
 wire \shift_reg[172].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[172].genblk1.genblk1.latch.q ;
 wire \shift_reg[173].genblk1.genblk1.latch.clk ;
 wire \shift_reg[173].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[173].genblk1.genblk1.latch.q ;
 wire \shift_reg[174].genblk1.genblk1.latch.clk ;
 wire \shift_reg[174].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[174].genblk1.genblk1.latch.q ;
 wire \shift_reg[175].genblk1.genblk1.latch.clk ;
 wire \shift_reg[175].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[175].genblk1.genblk1.latch.q ;
 wire \shift_reg[176].genblk1.genblk1.latch.clk ;
 wire \shift_reg[176].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[176].genblk1.genblk1.latch.q ;
 wire \shift_reg[177].genblk1.genblk1.latch.clk ;
 wire \shift_reg[177].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[177].genblk1.genblk1.latch.q ;
 wire \shift_reg[178].genblk1.genblk1.latch.clk ;
 wire \shift_reg[178].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[178].genblk1.genblk1.latch.q ;
 wire \shift_reg[179].genblk1.genblk1.latch.clk ;
 wire \shift_reg[179].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[179].genblk1.genblk1.latch.q ;
 wire \shift_reg[17].genblk1.genblk1.latch.clk ;
 wire \shift_reg[17].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[17].genblk1.genblk1.latch.q ;
 wire \shift_reg[180].genblk1.genblk1.latch.clk ;
 wire \shift_reg[180].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[180].genblk1.genblk1.latch.q ;
 wire \shift_reg[181].genblk1.genblk1.latch.clk ;
 wire \shift_reg[181].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[181].genblk1.genblk1.latch.q ;
 wire \shift_reg[182].genblk1.genblk1.latch.clk ;
 wire \shift_reg[182].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[182].genblk1.genblk1.latch.q ;
 wire \shift_reg[183].genblk1.genblk1.latch.clk ;
 wire \shift_reg[183].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[183].genblk1.genblk1.latch.q ;
 wire \shift_reg[184].genblk1.genblk1.latch.clk ;
 wire \shift_reg[184].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[184].genblk1.genblk1.latch.q ;
 wire \shift_reg[185].genblk1.genblk1.latch.clk ;
 wire \shift_reg[185].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[185].genblk1.genblk1.latch.q ;
 wire \shift_reg[186].genblk1.genblk1.latch.clk ;
 wire \shift_reg[186].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[186].genblk1.genblk1.latch.q ;
 wire \shift_reg[187].genblk1.genblk1.latch.clk ;
 wire \shift_reg[187].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[187].genblk1.genblk1.latch.q ;
 wire \shift_reg[188].genblk1.genblk1.latch.clk ;
 wire \shift_reg[188].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[188].genblk1.genblk1.latch.q ;
 wire \shift_reg[189].genblk1.genblk1.latch.clk ;
 wire \shift_reg[189].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[189].genblk1.genblk1.latch.q ;
 wire \shift_reg[18].genblk1.genblk1.latch.clk ;
 wire \shift_reg[18].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[18].genblk1.genblk1.latch.q ;
 wire \shift_reg[190].genblk1.genblk1.latch.clk ;
 wire \shift_reg[190].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[190].genblk1.genblk1.latch.q ;
 wire \shift_reg[191].genblk1.genblk1.latch.clk ;
 wire \shift_reg[191].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[191].genblk1.genblk1.latch.q ;
 wire \shift_reg[192].genblk1.genblk1.latch.clk ;
 wire \shift_reg[192].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[192].genblk1.genblk1.latch.q ;
 wire \shift_reg[193].genblk1.genblk1.latch.clk ;
 wire \shift_reg[193].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[193].genblk1.genblk1.latch.q ;
 wire \shift_reg[194].genblk1.genblk1.latch.clk ;
 wire \shift_reg[194].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[194].genblk1.genblk1.latch.q ;
 wire \shift_reg[195].genblk1.genblk1.latch.clk ;
 wire \shift_reg[195].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[195].genblk1.genblk1.latch.q ;
 wire \shift_reg[196].genblk1.genblk1.latch.clk ;
 wire \shift_reg[196].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[196].genblk1.genblk1.latch.q ;
 wire \shift_reg[197].genblk1.genblk1.latch.clk ;
 wire \shift_reg[197].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[197].genblk1.genblk1.latch.q ;
 wire \shift_reg[198].genblk1.genblk1.latch.clk ;
 wire \shift_reg[198].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[198].genblk1.genblk1.latch.q ;
 wire \shift_reg[199].genblk1.genblk1.latch.clk ;
 wire \shift_reg[199].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[199].genblk1.genblk1.latch.q ;
 wire \shift_reg[19].genblk1.genblk1.latch.clk ;
 wire \shift_reg[19].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[19].genblk1.genblk1.latch.q ;
 wire \shift_reg[1].genblk1.genblk1.latch.clk ;
 wire \shift_reg[1].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[1].genblk1.genblk1.latch.q ;
 wire \shift_reg[200].genblk1.genblk1.latch.clk ;
 wire \shift_reg[200].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[200].genblk1.genblk1.latch.q ;
 wire \shift_reg[201].genblk1.genblk1.latch.clk ;
 wire \shift_reg[201].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[201].genblk1.genblk1.latch.q ;
 wire \shift_reg[202].genblk1.genblk1.latch.clk ;
 wire \shift_reg[202].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[202].genblk1.genblk1.latch.q ;
 wire \shift_reg[203].genblk1.genblk1.latch.clk ;
 wire \shift_reg[203].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[203].genblk1.genblk1.latch.q ;
 wire \shift_reg[204].genblk1.genblk1.latch.clk ;
 wire \shift_reg[204].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[204].genblk1.genblk1.latch.q ;
 wire \shift_reg[205].genblk1.genblk1.latch.clk ;
 wire \shift_reg[205].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[205].genblk1.genblk1.latch.q ;
 wire \shift_reg[206].genblk1.genblk1.latch.clk ;
 wire \shift_reg[206].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[206].genblk1.genblk1.latch.q ;
 wire \shift_reg[207].genblk1.genblk1.latch.clk ;
 wire \shift_reg[207].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[207].genblk1.genblk1.latch.q ;
 wire \shift_reg[208].genblk1.genblk1.latch.clk ;
 wire \shift_reg[208].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[208].genblk1.genblk1.latch.q ;
 wire \shift_reg[209].genblk1.genblk1.latch.clk ;
 wire \shift_reg[209].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[209].genblk1.genblk1.latch.q ;
 wire \shift_reg[20].genblk1.genblk1.latch.clk ;
 wire \shift_reg[20].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[20].genblk1.genblk1.latch.q ;
 wire \shift_reg[210].genblk1.genblk1.latch.clk ;
 wire \shift_reg[210].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[210].genblk1.genblk1.latch.q ;
 wire \shift_reg[211].genblk1.genblk1.latch.clk ;
 wire \shift_reg[211].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[211].genblk1.genblk1.latch.q ;
 wire \shift_reg[212].genblk1.genblk1.latch.clk ;
 wire \shift_reg[212].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[212].genblk1.genblk1.latch.q ;
 wire \shift_reg[213].genblk1.genblk1.latch.clk ;
 wire \shift_reg[213].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[213].genblk1.genblk1.latch.q ;
 wire \shift_reg[214].genblk1.genblk1.latch.clk ;
 wire \shift_reg[214].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[214].genblk1.genblk1.latch.q ;
 wire \shift_reg[215].genblk1.genblk1.latch.clk ;
 wire \shift_reg[215].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[215].genblk1.genblk1.latch.q ;
 wire \shift_reg[216].genblk1.genblk1.latch.clk ;
 wire \shift_reg[216].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[216].genblk1.genblk1.latch.q ;
 wire \shift_reg[217].genblk1.genblk1.latch.clk ;
 wire \shift_reg[217].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[217].genblk1.genblk1.latch.q ;
 wire \shift_reg[218].genblk1.genblk1.latch.clk ;
 wire \shift_reg[218].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[218].genblk1.genblk1.latch.q ;
 wire \shift_reg[219].genblk1.genblk1.latch.clk ;
 wire \shift_reg[219].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[219].genblk1.genblk1.latch.q ;
 wire \shift_reg[21].genblk1.genblk1.latch.clk ;
 wire \shift_reg[21].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[21].genblk1.genblk1.latch.q ;
 wire \shift_reg[220].genblk1.genblk1.latch.clk ;
 wire \shift_reg[220].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[220].genblk1.genblk1.latch.q ;
 wire \shift_reg[221].genblk1.genblk1.latch.clk ;
 wire \shift_reg[221].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[221].genblk1.genblk1.latch.q ;
 wire \shift_reg[222].genblk1.genblk1.latch.clk ;
 wire \shift_reg[222].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[222].genblk1.genblk1.latch.q ;
 wire \shift_reg[223].genblk1.genblk1.latch.clk ;
 wire \shift_reg[223].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[223].genblk1.genblk1.latch.q ;
 wire \shift_reg[224].genblk1.genblk1.latch.clk ;
 wire \shift_reg[224].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[224].genblk1.genblk1.latch.q ;
 wire \shift_reg[225].genblk1.genblk1.latch.clk ;
 wire \shift_reg[225].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[225].genblk1.genblk1.latch.q ;
 wire \shift_reg[226].genblk1.genblk1.latch.clk ;
 wire \shift_reg[226].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[226].genblk1.genblk1.latch.q ;
 wire \shift_reg[227].genblk1.genblk1.latch.clk ;
 wire \shift_reg[227].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[227].genblk1.genblk1.latch.q ;
 wire \shift_reg[228].genblk1.genblk1.latch.clk ;
 wire \shift_reg[228].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[228].genblk1.genblk1.latch.q ;
 wire \shift_reg[229].genblk1.genblk1.latch.clk ;
 wire \shift_reg[229].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[229].genblk1.genblk1.latch.q ;
 wire \shift_reg[22].genblk1.genblk1.latch.clk ;
 wire \shift_reg[22].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[22].genblk1.genblk1.latch.q ;
 wire \shift_reg[230].genblk1.genblk1.latch.clk ;
 wire \shift_reg[230].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[230].genblk1.genblk1.latch.q ;
 wire \shift_reg[231].genblk1.genblk1.latch.clk ;
 wire \shift_reg[231].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[231].genblk1.genblk1.latch.q ;
 wire \shift_reg[232].genblk1.genblk1.latch.clk ;
 wire \shift_reg[232].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[232].genblk1.genblk1.latch.q ;
 wire \shift_reg[233].genblk1.genblk1.latch.clk ;
 wire \shift_reg[233].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[233].genblk1.genblk1.latch.q ;
 wire \shift_reg[234].genblk1.genblk1.latch.clk ;
 wire \shift_reg[234].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[234].genblk1.genblk1.latch.q ;
 wire \shift_reg[235].genblk1.genblk1.latch.clk ;
 wire \shift_reg[235].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[235].genblk1.genblk1.latch.q ;
 wire \shift_reg[236].genblk1.genblk1.latch.clk ;
 wire \shift_reg[236].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[236].genblk1.genblk1.latch.q ;
 wire \shift_reg[237].genblk1.genblk1.latch.clk ;
 wire \shift_reg[237].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[237].genblk1.genblk1.latch.q ;
 wire \shift_reg[238].genblk1.genblk1.latch.clk ;
 wire \shift_reg[238].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[238].genblk1.genblk1.latch.q ;
 wire \shift_reg[239].genblk1.genblk1.latch.clk ;
 wire \shift_reg[239].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[239].genblk1.genblk1.latch.q ;
 wire \shift_reg[23].genblk1.genblk1.latch.clk ;
 wire \shift_reg[23].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[23].genblk1.genblk1.latch.q ;
 wire \shift_reg[240].genblk1.genblk1.latch.clk ;
 wire \shift_reg[240].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[240].genblk1.genblk1.latch.q ;
 wire \shift_reg[241].genblk1.genblk1.latch.clk ;
 wire \shift_reg[241].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[241].genblk1.genblk1.latch.q ;
 wire \shift_reg[242].genblk1.genblk1.latch.clk ;
 wire \shift_reg[242].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[242].genblk1.genblk1.latch.q ;
 wire \shift_reg[243].genblk1.genblk1.latch.clk ;
 wire \shift_reg[243].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[243].genblk1.genblk1.latch.q ;
 wire \shift_reg[244].genblk1.genblk1.latch.clk ;
 wire \shift_reg[244].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[244].genblk1.genblk1.latch.q ;
 wire \shift_reg[245].genblk1.genblk1.latch.clk ;
 wire \shift_reg[245].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[245].genblk1.genblk1.latch.q ;
 wire \shift_reg[246].genblk1.genblk1.latch.clk ;
 wire \shift_reg[246].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[246].genblk1.genblk1.latch.q ;
 wire \shift_reg[247].genblk1.genblk1.latch.clk ;
 wire \shift_reg[247].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[247].genblk1.genblk1.latch.q ;
 wire \shift_reg[248].genblk1.genblk1.latch.clk ;
 wire \shift_reg[248].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[248].genblk1.genblk1.latch.q ;
 wire \shift_reg[249].genblk1.genblk1.latch.clk ;
 wire \shift_reg[249].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[249].genblk1.genblk1.latch.q ;
 wire \shift_reg[24].genblk1.genblk1.latch.clk ;
 wire \shift_reg[24].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[24].genblk1.genblk1.latch.q ;
 wire \shift_reg[250].genblk1.genblk1.latch.clk ;
 wire \shift_reg[250].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[250].genblk1.genblk1.latch.q ;
 wire \shift_reg[251].genblk1.genblk1.latch.clk ;
 wire \shift_reg[251].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[251].genblk1.genblk1.latch.q ;
 wire \shift_reg[252].genblk1.genblk1.latch.clk ;
 wire \shift_reg[252].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[252].genblk1.genblk1.latch.q ;
 wire \shift_reg[253].genblk1.genblk1.latch.clk ;
 wire \shift_reg[253].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[253].genblk1.genblk1.latch.q ;
 wire \shift_reg[254].genblk1.genblk1.latch.clk ;
 wire \shift_reg[254].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[254].genblk1.genblk1.latch.q ;
 wire \shift_reg[255].genblk1.genblk1.latch.clk ;
 wire \shift_reg[255].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[255].genblk1.genblk1.latch.q ;
 wire \shift_reg[256].genblk1.genblk1.latch.clk ;
 wire \shift_reg[256].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[256].genblk1.genblk1.latch.q ;
 wire \shift_reg[257].genblk1.genblk1.latch.clk ;
 wire \shift_reg[257].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[257].genblk1.genblk1.latch.q ;
 wire \shift_reg[258].genblk1.genblk1.latch.clk ;
 wire \shift_reg[258].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[258].genblk1.genblk1.latch.q ;
 wire \shift_reg[259].genblk1.genblk1.latch.clk ;
 wire \shift_reg[259].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[259].genblk1.genblk1.latch.q ;
 wire \shift_reg[25].genblk1.genblk1.latch.clk ;
 wire \shift_reg[25].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[25].genblk1.genblk1.latch.q ;
 wire \shift_reg[260].genblk1.genblk1.latch.clk ;
 wire \shift_reg[260].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[260].genblk1.genblk1.latch.q ;
 wire \shift_reg[261].genblk1.genblk1.latch.clk ;
 wire \shift_reg[261].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[261].genblk1.genblk1.latch.q ;
 wire \shift_reg[262].genblk1.genblk1.latch.clk ;
 wire \shift_reg[262].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[262].genblk1.genblk1.latch.q ;
 wire \shift_reg[263].genblk1.genblk1.latch.clk ;
 wire \shift_reg[263].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[263].genblk1.genblk1.latch.q ;
 wire \shift_reg[264].genblk1.genblk1.latch.clk ;
 wire \shift_reg[264].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[264].genblk1.genblk1.latch.q ;
 wire \shift_reg[265].genblk1.genblk1.latch.clk ;
 wire \shift_reg[265].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[265].genblk1.genblk1.latch.q ;
 wire \shift_reg[266].genblk1.genblk1.latch.clk ;
 wire \shift_reg[266].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[266].genblk1.genblk1.latch.q ;
 wire \shift_reg[267].genblk1.genblk1.latch.clk ;
 wire \shift_reg[267].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[267].genblk1.genblk1.latch.q ;
 wire \shift_reg[268].genblk1.genblk1.latch.clk ;
 wire \shift_reg[268].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[268].genblk1.genblk1.latch.q ;
 wire \shift_reg[269].genblk1.genblk1.latch.clk ;
 wire \shift_reg[269].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[269].genblk1.genblk1.latch.q ;
 wire \shift_reg[26].genblk1.genblk1.latch.clk ;
 wire \shift_reg[26].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[26].genblk1.genblk1.latch.q ;
 wire \shift_reg[270].genblk1.genblk1.latch.clk ;
 wire \shift_reg[270].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[270].genblk1.genblk1.latch.q ;
 wire \shift_reg[271].genblk1.genblk1.latch.clk ;
 wire \shift_reg[271].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[271].genblk1.genblk1.latch.q ;
 wire \shift_reg[272].genblk1.genblk1.latch.clk ;
 wire \shift_reg[272].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[272].genblk1.genblk1.latch.q ;
 wire \shift_reg[273].genblk1.genblk1.latch.clk ;
 wire \shift_reg[273].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[273].genblk1.genblk1.latch.q ;
 wire \shift_reg[274].genblk1.genblk1.latch.clk ;
 wire \shift_reg[274].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[274].genblk1.genblk1.latch.q ;
 wire \shift_reg[275].genblk1.genblk1.latch.clk ;
 wire \shift_reg[275].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[275].genblk1.genblk1.latch.q ;
 wire \shift_reg[276].genblk1.genblk1.latch.clk ;
 wire \shift_reg[276].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[276].genblk1.genblk1.latch.q ;
 wire \shift_reg[277].genblk1.genblk1.latch.clk ;
 wire \shift_reg[277].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[277].genblk1.genblk1.latch.q ;
 wire \shift_reg[278].genblk1.genblk1.latch.clk ;
 wire \shift_reg[278].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[278].genblk1.genblk1.latch.q ;
 wire \shift_reg[279].genblk1.genblk1.latch.clk ;
 wire \shift_reg[279].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[279].genblk1.genblk1.latch.q ;
 wire \shift_reg[27].genblk1.genblk1.latch.clk ;
 wire \shift_reg[27].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[27].genblk1.genblk1.latch.q ;
 wire \shift_reg[280].genblk1.genblk1.latch.clk ;
 wire \shift_reg[280].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[280].genblk1.genblk1.latch.q ;
 wire \shift_reg[281].genblk1.genblk1.latch.clk ;
 wire \shift_reg[281].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[281].genblk1.genblk1.latch.q ;
 wire \shift_reg[282].genblk1.genblk1.latch.clk ;
 wire \shift_reg[282].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[282].genblk1.genblk1.latch.q ;
 wire \shift_reg[283].genblk1.genblk1.latch.clk ;
 wire \shift_reg[283].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[283].genblk1.genblk1.latch.q ;
 wire \shift_reg[284].genblk1.genblk1.latch.clk ;
 wire \shift_reg[284].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[284].genblk1.genblk1.latch.q ;
 wire \shift_reg[285].genblk1.genblk1.latch.clk ;
 wire \shift_reg[285].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[285].genblk1.genblk1.latch.q ;
 wire \shift_reg[286].genblk1.genblk1.latch.clk ;
 wire \shift_reg[286].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[286].genblk1.genblk1.latch.q ;
 wire \shift_reg[287].genblk1.genblk1.latch.clk ;
 wire \shift_reg[287].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[287].genblk1.genblk1.latch.q ;
 wire \shift_reg[288].genblk1.genblk1.latch.clk ;
 wire \shift_reg[288].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[288].genblk1.genblk1.latch.q ;
 wire \shift_reg[289].genblk1.genblk1.latch.clk ;
 wire \shift_reg[289].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[289].genblk1.genblk1.latch.q ;
 wire \shift_reg[28].genblk1.genblk1.latch.clk ;
 wire \shift_reg[28].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[28].genblk1.genblk1.latch.q ;
 wire \shift_reg[290].genblk1.genblk1.latch.clk ;
 wire \shift_reg[290].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[290].genblk1.genblk1.latch.q ;
 wire \shift_reg[291].genblk1.genblk1.latch.clk ;
 wire \shift_reg[291].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[291].genblk1.genblk1.latch.q ;
 wire \shift_reg[292].genblk1.genblk1.latch.clk ;
 wire \shift_reg[292].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[292].genblk1.genblk1.latch.q ;
 wire \shift_reg[293].genblk1.genblk1.latch.clk ;
 wire \shift_reg[293].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[293].genblk1.genblk1.latch.q ;
 wire \shift_reg[294].genblk1.genblk1.latch.clk ;
 wire \shift_reg[294].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[294].genblk1.genblk1.latch.q ;
 wire \shift_reg[295].genblk1.genblk1.latch.clk ;
 wire \shift_reg[295].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[295].genblk1.genblk1.latch.q ;
 wire \shift_reg[296].genblk1.genblk1.latch.clk ;
 wire \shift_reg[296].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[296].genblk1.genblk1.latch.q ;
 wire \shift_reg[297].genblk1.genblk1.latch.clk ;
 wire \shift_reg[297].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[297].genblk1.genblk1.latch.q ;
 wire \shift_reg[298].genblk1.genblk1.latch.clk ;
 wire \shift_reg[298].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[298].genblk1.genblk1.latch.q ;
 wire \shift_reg[299].genblk1.genblk1.latch.clk ;
 wire \shift_reg[299].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[299].genblk1.genblk1.latch.q ;
 wire \shift_reg[29].genblk1.genblk1.latch.clk ;
 wire \shift_reg[29].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[29].genblk1.genblk1.latch.q ;
 wire \shift_reg[2].genblk1.genblk1.latch.clk ;
 wire \shift_reg[2].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[2].genblk1.genblk1.latch.q ;
 wire \shift_reg[300].genblk1.genblk1.latch.clk ;
 wire \shift_reg[300].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[300].genblk1.genblk1.latch.q ;
 wire \shift_reg[301].genblk1.genblk1.latch.clk ;
 wire \shift_reg[301].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[301].genblk1.genblk1.latch.q ;
 wire \shift_reg[302].genblk1.genblk1.latch.clk ;
 wire \shift_reg[302].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[302].genblk1.genblk1.latch.q ;
 wire \shift_reg[303].genblk1.genblk1.latch.clk ;
 wire \shift_reg[303].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[303].genblk1.genblk1.latch.q ;
 wire \shift_reg[304].genblk1.genblk1.latch.clk ;
 wire \shift_reg[304].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[304].genblk1.genblk1.latch.q ;
 wire \shift_reg[305].genblk1.genblk1.latch.clk ;
 wire \shift_reg[305].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[305].genblk1.genblk1.latch.q ;
 wire \shift_reg[306].genblk1.genblk1.latch.clk ;
 wire \shift_reg[306].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[306].genblk1.genblk1.latch.q ;
 wire \shift_reg[307].genblk1.genblk1.latch.clk ;
 wire \shift_reg[307].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[307].genblk1.genblk1.latch.q ;
 wire \shift_reg[308].genblk1.genblk1.latch.clk ;
 wire \shift_reg[308].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[308].genblk1.genblk1.latch.q ;
 wire \shift_reg[309].genblk1.genblk1.latch.clk ;
 wire \shift_reg[309].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[309].genblk1.genblk1.latch.q ;
 wire \shift_reg[30].genblk1.genblk1.latch.clk ;
 wire \shift_reg[30].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[30].genblk1.genblk1.latch.q ;
 wire \shift_reg[310].genblk1.genblk1.latch.clk ;
 wire \shift_reg[310].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[310].genblk1.genblk1.latch.q ;
 wire \shift_reg[311].genblk1.genblk1.latch.clk ;
 wire \shift_reg[311].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[311].genblk1.genblk1.latch.q ;
 wire \shift_reg[312].genblk1.genblk1.latch.clk ;
 wire \shift_reg[312].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[312].genblk1.genblk1.latch.q ;
 wire \shift_reg[313].genblk1.genblk1.latch.clk ;
 wire \shift_reg[313].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[313].genblk1.genblk1.latch.q ;
 wire \shift_reg[314].genblk1.genblk1.latch.clk ;
 wire \shift_reg[314].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[314].genblk1.genblk1.latch.q ;
 wire \shift_reg[315].genblk1.genblk1.latch.clk ;
 wire \shift_reg[315].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[315].genblk1.genblk1.latch.q ;
 wire \shift_reg[316].genblk1.genblk1.latch.clk ;
 wire \shift_reg[316].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[316].genblk1.genblk1.latch.q ;
 wire \shift_reg[317].genblk1.genblk1.latch.clk ;
 wire \shift_reg[317].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[317].genblk1.genblk1.latch.q ;
 wire \shift_reg[318].genblk1.genblk1.latch.clk ;
 wire \shift_reg[318].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[318].genblk1.genblk1.latch.q ;
 wire \shift_reg[319].genblk1.genblk1.latch.clk ;
 wire \shift_reg[319].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[319].genblk1.genblk1.latch.q ;
 wire \shift_reg[31].genblk1.genblk1.latch.clk ;
 wire \shift_reg[31].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[31].genblk1.genblk1.latch.q ;
 wire \shift_reg[320].genblk1.genblk1.latch.clk ;
 wire \shift_reg[320].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[320].genblk1.genblk1.latch.q ;
 wire \shift_reg[321].genblk1.genblk1.latch.clk ;
 wire \shift_reg[321].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[321].genblk1.genblk1.latch.q ;
 wire \shift_reg[322].genblk1.genblk1.latch.clk ;
 wire \shift_reg[322].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[322].genblk1.genblk1.latch.q ;
 wire \shift_reg[323].genblk1.genblk1.latch.clk ;
 wire \shift_reg[323].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[323].genblk1.genblk1.latch.q ;
 wire \shift_reg[324].genblk1.genblk1.latch.clk ;
 wire \shift_reg[324].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[324].genblk1.genblk1.latch.q ;
 wire \shift_reg[325].genblk1.genblk1.latch.clk ;
 wire \shift_reg[325].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[325].genblk1.genblk1.latch.q ;
 wire \shift_reg[326].genblk1.genblk1.latch.clk ;
 wire \shift_reg[326].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[326].genblk1.genblk1.latch.q ;
 wire \shift_reg[327].genblk1.genblk1.latch.clk ;
 wire \shift_reg[327].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[327].genblk1.genblk1.latch.q ;
 wire \shift_reg[328].genblk1.genblk1.latch.clk ;
 wire \shift_reg[328].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[328].genblk1.genblk1.latch.q ;
 wire \shift_reg[329].genblk1.genblk1.latch.clk ;
 wire \shift_reg[329].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[329].genblk1.genblk1.latch.q ;
 wire \shift_reg[32].genblk1.genblk1.latch.clk ;
 wire \shift_reg[32].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[32].genblk1.genblk1.latch.q ;
 wire \shift_reg[330].genblk1.genblk1.latch.clk ;
 wire \shift_reg[330].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[330].genblk1.genblk1.latch.q ;
 wire \shift_reg[331].genblk1.genblk1.latch.clk ;
 wire \shift_reg[331].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[331].genblk1.genblk1.latch.q ;
 wire \shift_reg[332].genblk1.genblk1.latch.clk ;
 wire \shift_reg[332].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[332].genblk1.genblk1.latch.q ;
 wire \shift_reg[333].genblk1.genblk1.latch.clk ;
 wire \shift_reg[333].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[333].genblk1.genblk1.latch.q ;
 wire \shift_reg[334].genblk1.genblk1.latch.clk ;
 wire \shift_reg[334].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[334].genblk1.genblk1.latch.q ;
 wire \shift_reg[335].genblk1.genblk1.latch.clk ;
 wire \shift_reg[335].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[335].genblk1.genblk1.latch.q ;
 wire \shift_reg[336].genblk1.genblk1.latch.clk ;
 wire \shift_reg[336].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[336].genblk1.genblk1.latch.q ;
 wire \shift_reg[337].genblk1.genblk1.latch.clk ;
 wire \shift_reg[337].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[337].genblk1.genblk1.latch.q ;
 wire \shift_reg[338].genblk1.genblk1.latch.clk ;
 wire \shift_reg[338].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[338].genblk1.genblk1.latch.q ;
 wire \shift_reg[339].genblk1.genblk1.latch.clk ;
 wire \shift_reg[339].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[339].genblk1.genblk1.latch.q ;
 wire \shift_reg[33].genblk1.genblk1.latch.clk ;
 wire \shift_reg[33].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[33].genblk1.genblk1.latch.q ;
 wire \shift_reg[340].genblk1.genblk1.latch.clk ;
 wire \shift_reg[340].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[340].genblk1.genblk1.latch.q ;
 wire \shift_reg[341].genblk1.genblk1.latch.clk ;
 wire \shift_reg[341].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[341].genblk1.genblk1.latch.q ;
 wire \shift_reg[342].genblk1.genblk1.latch.clk ;
 wire \shift_reg[342].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[342].genblk1.genblk1.latch.q ;
 wire \shift_reg[343].genblk1.genblk1.latch.clk ;
 wire \shift_reg[343].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[343].genblk1.genblk1.latch.q ;
 wire \shift_reg[344].genblk1.genblk1.latch.clk ;
 wire \shift_reg[344].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[344].genblk1.genblk1.latch.q ;
 wire \shift_reg[345].genblk1.genblk1.latch.clk ;
 wire \shift_reg[345].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[345].genblk1.genblk1.latch.q ;
 wire \shift_reg[346].genblk1.genblk1.latch.clk ;
 wire \shift_reg[346].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[346].genblk1.genblk1.latch.q ;
 wire \shift_reg[347].genblk1.genblk1.latch.clk ;
 wire \shift_reg[347].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[347].genblk1.genblk1.latch.q ;
 wire \shift_reg[348].genblk1.genblk1.latch.clk ;
 wire \shift_reg[348].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[348].genblk1.genblk1.latch.q ;
 wire \shift_reg[349].genblk1.genblk1.latch.clk ;
 wire \shift_reg[349].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[349].genblk1.genblk1.latch.q ;
 wire \shift_reg[34].genblk1.genblk1.latch.clk ;
 wire \shift_reg[34].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[34].genblk1.genblk1.latch.q ;
 wire \shift_reg[350].genblk1.genblk1.latch.clk ;
 wire \shift_reg[350].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[350].genblk1.genblk1.latch.q ;
 wire \shift_reg[351].genblk1.genblk1.latch.clk ;
 wire \shift_reg[351].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[351].genblk1.genblk1.latch.q ;
 wire \shift_reg[352].genblk1.genblk1.latch.clk ;
 wire \shift_reg[352].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[352].genblk1.genblk1.latch.q ;
 wire \shift_reg[353].genblk1.genblk1.latch.clk ;
 wire \shift_reg[353].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[353].genblk1.genblk1.latch.q ;
 wire \shift_reg[354].genblk1.genblk1.latch.clk ;
 wire \shift_reg[354].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[354].genblk1.genblk1.latch.q ;
 wire \shift_reg[355].genblk1.genblk1.latch.clk ;
 wire \shift_reg[355].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[355].genblk1.genblk1.latch.q ;
 wire \shift_reg[356].genblk1.genblk1.latch.clk ;
 wire \shift_reg[356].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[356].genblk1.genblk1.latch.q ;
 wire \shift_reg[357].genblk1.genblk1.latch.clk ;
 wire \shift_reg[357].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[357].genblk1.genblk1.latch.q ;
 wire \shift_reg[358].genblk1.genblk1.latch.clk ;
 wire \shift_reg[358].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[358].genblk1.genblk1.latch.q ;
 wire \shift_reg[359].genblk1.genblk1.latch.clk ;
 wire \shift_reg[359].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[359].genblk1.genblk1.latch.q ;
 wire \shift_reg[35].genblk1.genblk1.latch.clk ;
 wire \shift_reg[35].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[35].genblk1.genblk1.latch.q ;
 wire \shift_reg[360].genblk1.genblk1.latch.clk ;
 wire \shift_reg[360].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[360].genblk1.genblk1.latch.q ;
 wire \shift_reg[361].genblk1.genblk1.latch.clk ;
 wire \shift_reg[361].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[361].genblk1.genblk1.latch.q ;
 wire \shift_reg[362].genblk1.genblk1.latch.clk ;
 wire \shift_reg[362].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[362].genblk1.genblk1.latch.q ;
 wire \shift_reg[363].genblk1.genblk1.latch.clk ;
 wire \shift_reg[363].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[363].genblk1.genblk1.latch.q ;
 wire \shift_reg[364].genblk1.genblk1.latch.clk ;
 wire \shift_reg[364].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[364].genblk1.genblk1.latch.q ;
 wire \shift_reg[365].genblk1.genblk1.latch.clk ;
 wire \shift_reg[365].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[365].genblk1.genblk1.latch.q ;
 wire \shift_reg[366].genblk1.genblk1.latch.clk ;
 wire \shift_reg[366].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[366].genblk1.genblk1.latch.q ;
 wire \shift_reg[367].genblk1.genblk1.latch.clk ;
 wire \shift_reg[367].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[367].genblk1.genblk1.latch.q ;
 wire \shift_reg[368].genblk1.genblk1.latch.clk ;
 wire \shift_reg[368].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[368].genblk1.genblk1.latch.q ;
 wire \shift_reg[369].genblk1.genblk1.latch.clk ;
 wire \shift_reg[369].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[369].genblk1.genblk1.latch.q ;
 wire \shift_reg[36].genblk1.genblk1.latch.clk ;
 wire \shift_reg[36].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[36].genblk1.genblk1.latch.q ;
 wire \shift_reg[370].genblk1.genblk1.latch.clk ;
 wire \shift_reg[370].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[370].genblk1.genblk1.latch.q ;
 wire \shift_reg[371].genblk1.genblk1.latch.clk ;
 wire \shift_reg[371].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[371].genblk1.genblk1.latch.q ;
 wire \shift_reg[372].genblk1.genblk1.latch.clk ;
 wire \shift_reg[372].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[372].genblk1.genblk1.latch.q ;
 wire \shift_reg[373].genblk1.genblk1.latch.clk ;
 wire \shift_reg[373].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[373].genblk1.genblk1.latch.q ;
 wire \shift_reg[374].genblk1.genblk1.latch.clk ;
 wire \shift_reg[374].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[374].genblk1.genblk1.latch.q ;
 wire \shift_reg[375].genblk1.genblk1.latch.clk ;
 wire \shift_reg[375].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[375].genblk1.genblk1.latch.q ;
 wire \shift_reg[376].genblk1.genblk1.latch.clk ;
 wire \shift_reg[376].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[376].genblk1.genblk1.latch.q ;
 wire \shift_reg[377].genblk1.genblk1.latch.clk ;
 wire \shift_reg[377].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[377].genblk1.genblk1.latch.q ;
 wire \shift_reg[378].genblk1.genblk1.latch.clk ;
 wire \shift_reg[378].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[378].genblk1.genblk1.latch.q ;
 wire \shift_reg[379].genblk1.genblk1.latch.clk ;
 wire \shift_reg[379].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[379].genblk1.genblk1.latch.q ;
 wire \shift_reg[37].genblk1.genblk1.latch.clk ;
 wire \shift_reg[37].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[37].genblk1.genblk1.latch.q ;
 wire \shift_reg[380].genblk1.genblk1.latch.clk ;
 wire \shift_reg[380].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[380].genblk1.genblk1.latch.q ;
 wire \shift_reg[381].genblk1.genblk1.latch.clk ;
 wire \shift_reg[381].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[381].genblk1.genblk1.latch.q ;
 wire \shift_reg[382].genblk1.genblk1.latch.clk ;
 wire \shift_reg[382].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[382].genblk1.genblk1.latch.q ;
 wire \shift_reg[383].genblk1.genblk1.latch.clk ;
 wire \shift_reg[383].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[383].genblk1.genblk1.latch.q ;
 wire \shift_reg[384].genblk1.genblk1.latch.clk ;
 wire \shift_reg[384].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[384].genblk1.genblk1.latch.q ;
 wire \shift_reg[385].genblk1.genblk1.latch.clk ;
 wire \shift_reg[385].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[385].genblk1.genblk1.latch.q ;
 wire \shift_reg[386].genblk1.genblk1.latch.clk ;
 wire \shift_reg[386].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[386].genblk1.genblk1.latch.q ;
 wire \shift_reg[387].genblk1.genblk1.latch.clk ;
 wire \shift_reg[387].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[387].genblk1.genblk1.latch.q ;
 wire \shift_reg[388].genblk1.genblk1.latch.clk ;
 wire \shift_reg[388].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[388].genblk1.genblk1.latch.q ;
 wire \shift_reg[389].genblk1.genblk1.latch.clk ;
 wire \shift_reg[389].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[389].genblk1.genblk1.latch.q ;
 wire \shift_reg[38].genblk1.genblk1.latch.clk ;
 wire \shift_reg[38].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[38].genblk1.genblk1.latch.q ;
 wire \shift_reg[390].genblk1.genblk1.latch.clk ;
 wire \shift_reg[390].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[390].genblk1.genblk1.latch.q ;
 wire \shift_reg[391].genblk1.genblk1.latch.clk ;
 wire \shift_reg[391].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[391].genblk1.genblk1.latch.q ;
 wire \shift_reg[392].genblk1.genblk1.latch.clk ;
 wire \shift_reg[392].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[392].genblk1.genblk1.latch.q ;
 wire \shift_reg[393].genblk1.genblk1.latch.clk ;
 wire \shift_reg[393].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[393].genblk1.genblk1.latch.q ;
 wire \shift_reg[394].genblk1.genblk1.latch.clk ;
 wire \shift_reg[394].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[394].genblk1.genblk1.latch.q ;
 wire \shift_reg[395].genblk1.genblk1.latch.clk ;
 wire \shift_reg[395].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[395].genblk1.genblk1.latch.q ;
 wire \shift_reg[396].genblk1.genblk1.latch.clk ;
 wire \shift_reg[396].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[396].genblk1.genblk1.latch.q ;
 wire \shift_reg[397].genblk1.genblk1.latch.clk ;
 wire \shift_reg[397].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[397].genblk1.genblk1.latch.q ;
 wire \shift_reg[398].genblk1.genblk1.latch.clk ;
 wire \shift_reg[398].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[398].genblk1.genblk1.latch.q ;
 wire \shift_reg[399].genblk1.genblk1.latch.clk ;
 wire \shift_reg[399].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[399].genblk1.genblk1.latch.q ;
 wire \shift_reg[39].genblk1.genblk1.latch.clk ;
 wire \shift_reg[39].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[39].genblk1.genblk1.latch.q ;
 wire \shift_reg[3].genblk1.genblk1.latch.clk ;
 wire \shift_reg[3].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[3].genblk1.genblk1.latch.q ;
 wire \shift_reg[400].genblk1.genblk1.latch.clk ;
 wire \shift_reg[400].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[400].genblk1.genblk1.latch.q ;
 wire \shift_reg[401].genblk1.genblk1.latch.clk ;
 wire \shift_reg[401].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[401].genblk1.genblk1.latch.q ;
 wire \shift_reg[402].genblk1.genblk1.latch.clk ;
 wire \shift_reg[402].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[402].genblk1.genblk1.latch.q ;
 wire \shift_reg[403].genblk1.genblk1.latch.clk ;
 wire \shift_reg[403].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[403].genblk1.genblk1.latch.q ;
 wire \shift_reg[404].genblk1.genblk1.latch.clk ;
 wire \shift_reg[404].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[404].genblk1.genblk1.latch.q ;
 wire \shift_reg[405].genblk1.genblk1.latch.clk ;
 wire \shift_reg[405].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[405].genblk1.genblk1.latch.q ;
 wire \shift_reg[406].genblk1.genblk1.latch.clk ;
 wire \shift_reg[406].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[406].genblk1.genblk1.latch.q ;
 wire \shift_reg[407].genblk1.genblk1.latch.clk ;
 wire \shift_reg[407].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[407].genblk1.genblk1.latch.q ;
 wire \shift_reg[408].genblk1.genblk1.latch.clk ;
 wire \shift_reg[408].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[408].genblk1.genblk1.latch.q ;
 wire \shift_reg[409].genblk1.genblk1.latch.clk ;
 wire \shift_reg[409].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[409].genblk1.genblk1.latch.q ;
 wire \shift_reg[40].genblk1.genblk1.latch.clk ;
 wire \shift_reg[40].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[40].genblk1.genblk1.latch.q ;
 wire \shift_reg[410].genblk1.genblk1.latch.clk ;
 wire \shift_reg[410].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[410].genblk1.genblk1.latch.q ;
 wire \shift_reg[411].genblk1.genblk1.latch.clk ;
 wire \shift_reg[411].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[411].genblk1.genblk1.latch.q ;
 wire \shift_reg[412].genblk1.genblk1.latch.clk ;
 wire \shift_reg[412].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[412].genblk1.genblk1.latch.q ;
 wire \shift_reg[413].genblk1.genblk1.latch.clk ;
 wire \shift_reg[413].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[413].genblk1.genblk1.latch.q ;
 wire \shift_reg[414].genblk1.genblk1.latch.clk ;
 wire \shift_reg[414].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[414].genblk1.genblk1.latch.q ;
 wire \shift_reg[415].genblk1.genblk1.latch.clk ;
 wire \shift_reg[415].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[415].genblk1.genblk1.latch.q ;
 wire \shift_reg[416].genblk1.genblk1.latch.clk ;
 wire \shift_reg[416].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[416].genblk1.genblk1.latch.q ;
 wire \shift_reg[417].genblk1.genblk1.latch.clk ;
 wire \shift_reg[417].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[417].genblk1.genblk1.latch.q ;
 wire \shift_reg[418].genblk1.genblk1.latch.clk ;
 wire \shift_reg[418].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[418].genblk1.genblk1.latch.q ;
 wire \shift_reg[419].genblk1.genblk1.latch.clk ;
 wire \shift_reg[419].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[419].genblk1.genblk1.latch.q ;
 wire \shift_reg[41].genblk1.genblk1.latch.clk ;
 wire \shift_reg[41].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[41].genblk1.genblk1.latch.q ;
 wire \shift_reg[420].genblk1.genblk1.latch.clk ;
 wire \shift_reg[420].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[420].genblk1.genblk1.latch.q ;
 wire \shift_reg[421].genblk1.genblk1.latch.clk ;
 wire \shift_reg[421].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[421].genblk1.genblk1.latch.q ;
 wire \shift_reg[422].genblk1.genblk1.latch.clk ;
 wire \shift_reg[422].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[422].genblk1.genblk1.latch.q ;
 wire \shift_reg[423].genblk1.genblk1.latch.clk ;
 wire \shift_reg[423].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[423].genblk1.genblk1.latch.q ;
 wire \shift_reg[424].genblk1.genblk1.latch.clk ;
 wire \shift_reg[424].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[424].genblk1.genblk1.latch.q ;
 wire \shift_reg[425].genblk1.genblk1.latch.clk ;
 wire \shift_reg[425].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[425].genblk1.genblk1.latch.q ;
 wire \shift_reg[426].genblk1.genblk1.latch.clk ;
 wire \shift_reg[426].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[426].genblk1.genblk1.latch.q ;
 wire \shift_reg[427].genblk1.genblk1.latch.clk ;
 wire \shift_reg[427].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[427].genblk1.genblk1.latch.q ;
 wire \shift_reg[428].genblk1.genblk1.latch.clk ;
 wire \shift_reg[428].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[428].genblk1.genblk1.latch.q ;
 wire \shift_reg[429].genblk1.genblk1.latch.clk ;
 wire \shift_reg[429].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[429].genblk1.genblk1.latch.q ;
 wire \shift_reg[42].genblk1.genblk1.latch.clk ;
 wire \shift_reg[42].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[42].genblk1.genblk1.latch.q ;
 wire \shift_reg[430].genblk1.genblk1.latch.clk ;
 wire \shift_reg[430].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[430].genblk1.genblk1.latch.q ;
 wire \shift_reg[431].genblk1.genblk1.latch.clk ;
 wire \shift_reg[431].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[431].genblk1.genblk1.latch.q ;
 wire \shift_reg[432].genblk1.genblk1.latch.clk ;
 wire \shift_reg[432].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[432].genblk1.genblk1.latch.q ;
 wire \shift_reg[433].genblk1.genblk1.latch.clk ;
 wire \shift_reg[433].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[433].genblk1.genblk1.latch.q ;
 wire \shift_reg[434].genblk1.genblk1.latch.clk ;
 wire \shift_reg[434].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[434].genblk1.genblk1.latch.q ;
 wire \shift_reg[435].genblk1.genblk1.latch.clk ;
 wire \shift_reg[435].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[435].genblk1.genblk1.latch.q ;
 wire \shift_reg[436].genblk1.genblk1.latch.clk ;
 wire \shift_reg[436].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[436].genblk1.genblk1.latch.q ;
 wire \shift_reg[437].genblk1.genblk1.latch.clk ;
 wire \shift_reg[437].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[437].genblk1.genblk1.latch.q ;
 wire \shift_reg[438].genblk1.genblk1.latch.clk ;
 wire \shift_reg[438].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[438].genblk1.genblk1.latch.q ;
 wire \shift_reg[439].genblk1.genblk1.latch.clk ;
 wire \shift_reg[439].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[439].genblk1.genblk1.latch.q ;
 wire \shift_reg[43].genblk1.genblk1.latch.clk ;
 wire \shift_reg[43].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[43].genblk1.genblk1.latch.q ;
 wire \shift_reg[440].genblk1.genblk1.latch.clk ;
 wire \shift_reg[440].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[440].genblk1.genblk1.latch.q ;
 wire \shift_reg[441].genblk1.genblk1.latch.clk ;
 wire \shift_reg[441].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[441].genblk1.genblk1.latch.q ;
 wire \shift_reg[442].genblk1.genblk1.latch.clk ;
 wire \shift_reg[442].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[442].genblk1.genblk1.latch.q ;
 wire \shift_reg[443].genblk1.genblk1.latch.clk ;
 wire \shift_reg[443].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[443].genblk1.genblk1.latch.q ;
 wire \shift_reg[444].genblk1.genblk1.latch.clk ;
 wire \shift_reg[444].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[444].genblk1.genblk1.latch.q ;
 wire \shift_reg[445].genblk1.genblk1.latch.clk ;
 wire \shift_reg[445].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[445].genblk1.genblk1.latch.q ;
 wire \shift_reg[446].genblk1.genblk1.latch.clk ;
 wire \shift_reg[446].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[446].genblk1.genblk1.latch.q ;
 wire \shift_reg[447].genblk1.genblk1.latch.clk ;
 wire \shift_reg[447].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[447].genblk1.genblk1.latch.q ;
 wire \shift_reg[448].genblk1.genblk1.latch.clk ;
 wire \shift_reg[448].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[448].genblk1.genblk1.latch.q ;
 wire \shift_reg[449].genblk1.genblk1.latch.clk ;
 wire \shift_reg[449].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[449].genblk1.genblk1.latch.q ;
 wire \shift_reg[44].genblk1.genblk1.latch.clk ;
 wire \shift_reg[44].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[44].genblk1.genblk1.latch.q ;
 wire \shift_reg[450].genblk1.genblk1.latch.clk ;
 wire \shift_reg[450].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[450].genblk1.genblk1.latch.q ;
 wire \shift_reg[451].genblk1.genblk1.latch.clk ;
 wire \shift_reg[451].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[451].genblk1.genblk1.latch.q ;
 wire \shift_reg[452].genblk1.genblk1.latch.clk ;
 wire \shift_reg[452].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[452].genblk1.genblk1.latch.q ;
 wire \shift_reg[453].genblk1.genblk1.latch.clk ;
 wire \shift_reg[453].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[453].genblk1.genblk1.latch.q ;
 wire \shift_reg[454].genblk1.genblk1.latch.clk ;
 wire \shift_reg[454].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[454].genblk1.genblk1.latch.q ;
 wire \shift_reg[455].genblk1.genblk1.latch.clk ;
 wire \shift_reg[455].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[455].genblk1.genblk1.latch.q ;
 wire \shift_reg[456].genblk1.genblk1.latch.clk ;
 wire \shift_reg[456].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[456].genblk1.genblk1.latch.q ;
 wire \shift_reg[457].genblk1.genblk1.latch.clk ;
 wire \shift_reg[457].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[457].genblk1.genblk1.latch.q ;
 wire \shift_reg[458].genblk1.genblk1.latch.clk ;
 wire \shift_reg[458].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[458].genblk1.genblk1.latch.q ;
 wire \shift_reg[459].genblk1.genblk1.latch.clk ;
 wire \shift_reg[459].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[459].genblk1.genblk1.latch.q ;
 wire \shift_reg[45].genblk1.genblk1.latch.clk ;
 wire \shift_reg[45].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[45].genblk1.genblk1.latch.q ;
 wire \shift_reg[460].genblk1.genblk1.latch.clk ;
 wire \shift_reg[460].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[460].genblk1.genblk1.latch.q ;
 wire \shift_reg[461].genblk1.genblk1.latch.clk ;
 wire \shift_reg[461].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[461].genblk1.genblk1.latch.q ;
 wire \shift_reg[462].genblk1.genblk1.latch.clk ;
 wire \shift_reg[462].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[462].genblk1.genblk1.latch.q ;
 wire \shift_reg[463].genblk1.genblk1.latch.clk ;
 wire \shift_reg[463].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[463].genblk1.genblk1.latch.q ;
 wire \shift_reg[464].genblk1.genblk1.latch.clk ;
 wire \shift_reg[464].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[464].genblk1.genblk1.latch.q ;
 wire \shift_reg[465].genblk1.genblk1.latch.clk ;
 wire \shift_reg[465].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[465].genblk1.genblk1.latch.q ;
 wire \shift_reg[466].genblk1.genblk1.latch.clk ;
 wire \shift_reg[466].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[466].genblk1.genblk1.latch.q ;
 wire \shift_reg[467].genblk1.genblk1.latch.clk ;
 wire \shift_reg[467].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[467].genblk1.genblk1.latch.q ;
 wire \shift_reg[468].genblk1.genblk1.latch.clk ;
 wire \shift_reg[468].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[468].genblk1.genblk1.latch.q ;
 wire \shift_reg[469].genblk1.genblk1.latch.clk ;
 wire \shift_reg[469].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[469].genblk1.genblk1.latch.q ;
 wire \shift_reg[46].genblk1.genblk1.latch.clk ;
 wire \shift_reg[46].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[46].genblk1.genblk1.latch.q ;
 wire \shift_reg[470].genblk1.genblk1.latch.clk ;
 wire \shift_reg[470].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[470].genblk1.genblk1.latch.q ;
 wire \shift_reg[471].genblk1.genblk1.latch.clk ;
 wire \shift_reg[471].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[471].genblk1.genblk1.latch.q ;
 wire \shift_reg[472].genblk1.genblk1.latch.clk ;
 wire \shift_reg[472].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[472].genblk1.genblk1.latch.q ;
 wire \shift_reg[473].genblk1.genblk1.latch.clk ;
 wire \shift_reg[473].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[473].genblk1.genblk1.latch.q ;
 wire \shift_reg[474].genblk1.genblk1.latch.clk ;
 wire \shift_reg[474].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[474].genblk1.genblk1.latch.q ;
 wire \shift_reg[475].genblk1.genblk1.latch.clk ;
 wire \shift_reg[475].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[475].genblk1.genblk1.latch.q ;
 wire \shift_reg[476].genblk1.genblk1.latch.clk ;
 wire \shift_reg[476].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[476].genblk1.genblk1.latch.q ;
 wire \shift_reg[477].genblk1.genblk1.latch.clk ;
 wire \shift_reg[477].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[477].genblk1.genblk1.latch.q ;
 wire \shift_reg[478].genblk1.genblk1.latch.clk ;
 wire \shift_reg[478].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[478].genblk1.genblk1.latch.q ;
 wire \shift_reg[479].genblk1.genblk1.latch.clk ;
 wire \shift_reg[479].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[479].genblk1.genblk1.latch.q ;
 wire \shift_reg[47].genblk1.genblk1.latch.clk ;
 wire \shift_reg[47].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[47].genblk1.genblk1.latch.q ;
 wire \shift_reg[480].genblk1.genblk1.latch.clk ;
 wire \shift_reg[480].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[480].genblk1.genblk1.latch.q ;
 wire \shift_reg[481].genblk1.genblk1.latch.clk ;
 wire \shift_reg[481].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[481].genblk1.genblk1.latch.q ;
 wire \shift_reg[482].genblk1.genblk1.latch.clk ;
 wire \shift_reg[482].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[482].genblk1.genblk1.latch.q ;
 wire \shift_reg[483].genblk1.genblk1.latch.clk ;
 wire \shift_reg[483].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[483].genblk1.genblk1.latch.q ;
 wire \shift_reg[484].genblk1.genblk1.latch.clk ;
 wire \shift_reg[484].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[484].genblk1.genblk1.latch.q ;
 wire \shift_reg[485].genblk1.genblk1.latch.clk ;
 wire \shift_reg[485].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[485].genblk1.genblk1.latch.q ;
 wire \shift_reg[486].genblk1.genblk1.latch.clk ;
 wire \shift_reg[486].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[486].genblk1.genblk1.latch.q ;
 wire \shift_reg[487].genblk1.genblk1.latch.clk ;
 wire \shift_reg[487].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[487].genblk1.genblk1.latch.q ;
 wire \shift_reg[488].genblk1.genblk1.latch.clk ;
 wire \shift_reg[488].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[488].genblk1.genblk1.latch.q ;
 wire \shift_reg[489].genblk1.genblk1.latch.clk ;
 wire \shift_reg[489].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[489].genblk1.genblk1.latch.q ;
 wire \shift_reg[48].genblk1.genblk1.latch.clk ;
 wire \shift_reg[48].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[48].genblk1.genblk1.latch.q ;
 wire \shift_reg[490].genblk1.genblk1.latch.clk ;
 wire \shift_reg[490].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[490].genblk1.genblk1.latch.q ;
 wire \shift_reg[491].genblk1.genblk1.latch.clk ;
 wire \shift_reg[491].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[491].genblk1.genblk1.latch.q ;
 wire \shift_reg[492].genblk1.genblk1.latch.clk ;
 wire \shift_reg[492].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[492].genblk1.genblk1.latch.q ;
 wire \shift_reg[493].genblk1.genblk1.latch.clk ;
 wire \shift_reg[493].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[493].genblk1.genblk1.latch.q ;
 wire \shift_reg[494].genblk1.genblk1.latch.clk ;
 wire \shift_reg[494].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[494].genblk1.genblk1.latch.q ;
 wire \shift_reg[495].genblk1.genblk1.latch.clk ;
 wire \shift_reg[495].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[495].genblk1.genblk1.latch.q ;
 wire \shift_reg[496].genblk1.genblk1.latch.clk ;
 wire \shift_reg[496].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[496].genblk1.genblk1.latch.q ;
 wire \shift_reg[497].genblk1.genblk1.latch.clk ;
 wire \shift_reg[497].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[497].genblk1.genblk1.latch.q ;
 wire \shift_reg[498].genblk1.genblk1.latch.clk ;
 wire \shift_reg[498].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[498].genblk1.genblk1.latch.q ;
 wire \shift_reg[499].genblk1.genblk1.latch.clk ;
 wire \shift_reg[499].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[499].genblk1.genblk1.latch.q ;
 wire \shift_reg[49].genblk1.genblk1.latch.clk ;
 wire \shift_reg[49].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[49].genblk1.genblk1.latch.q ;
 wire \shift_reg[4].genblk1.genblk1.latch.clk ;
 wire \shift_reg[4].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[4].genblk1.genblk1.latch.q ;
 wire \shift_reg[500].genblk1.genblk1.latch.clk ;
 wire \shift_reg[500].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[500].genblk1.genblk1.latch.q ;
 wire \shift_reg[501].genblk1.genblk1.latch.clk ;
 wire \shift_reg[501].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[501].genblk1.genblk1.latch.q ;
 wire \shift_reg[502].genblk1.genblk1.latch.clk ;
 wire \shift_reg[502].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[502].genblk1.genblk1.latch.q ;
 wire \shift_reg[503].genblk1.genblk1.latch.clk ;
 wire \shift_reg[503].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[503].genblk1.genblk1.latch.q ;
 wire \shift_reg[504].genblk1.genblk1.latch.clk ;
 wire \shift_reg[504].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[504].genblk1.genblk1.latch.q ;
 wire \shift_reg[505].genblk1.genblk1.latch.clk ;
 wire \shift_reg[505].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[505].genblk1.genblk1.latch.q ;
 wire \shift_reg[506].genblk1.genblk1.latch.clk ;
 wire \shift_reg[506].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[506].genblk1.genblk1.latch.q ;
 wire \shift_reg[507].genblk1.genblk1.latch.clk ;
 wire \shift_reg[507].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[507].genblk1.genblk1.latch.q ;
 wire \shift_reg[508].genblk1.genblk1.latch.clk ;
 wire \shift_reg[508].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[508].genblk1.genblk1.latch.q ;
 wire \shift_reg[509].genblk1.genblk1.latch.clk ;
 wire \shift_reg[509].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[509].genblk1.genblk1.latch.q ;
 wire \shift_reg[50].genblk1.genblk1.latch.clk ;
 wire \shift_reg[50].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[50].genblk1.genblk1.latch.q ;
 wire \shift_reg[510].genblk1.genblk1.latch.clk ;
 wire \shift_reg[510].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[510].genblk1.genblk1.latch.q ;
 wire \shift_reg[511].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[511].genblk1.genblk1.latch.q ;
 wire \shift_reg[51].genblk1.genblk1.latch.clk ;
 wire \shift_reg[51].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[51].genblk1.genblk1.latch.q ;
 wire \shift_reg[52].genblk1.genblk1.latch.clk ;
 wire \shift_reg[52].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[52].genblk1.genblk1.latch.q ;
 wire \shift_reg[53].genblk1.genblk1.latch.clk ;
 wire \shift_reg[53].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[53].genblk1.genblk1.latch.q ;
 wire \shift_reg[54].genblk1.genblk1.latch.clk ;
 wire \shift_reg[54].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[54].genblk1.genblk1.latch.q ;
 wire \shift_reg[55].genblk1.genblk1.latch.clk ;
 wire \shift_reg[55].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[55].genblk1.genblk1.latch.q ;
 wire \shift_reg[56].genblk1.genblk1.latch.clk ;
 wire \shift_reg[56].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[56].genblk1.genblk1.latch.q ;
 wire \shift_reg[57].genblk1.genblk1.latch.clk ;
 wire \shift_reg[57].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[57].genblk1.genblk1.latch.q ;
 wire \shift_reg[58].genblk1.genblk1.latch.clk ;
 wire \shift_reg[58].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[58].genblk1.genblk1.latch.q ;
 wire \shift_reg[59].genblk1.genblk1.latch.clk ;
 wire \shift_reg[59].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[59].genblk1.genblk1.latch.q ;
 wire \shift_reg[5].genblk1.genblk1.latch.clk ;
 wire \shift_reg[5].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[5].genblk1.genblk1.latch.q ;
 wire \shift_reg[60].genblk1.genblk1.latch.clk ;
 wire \shift_reg[60].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[60].genblk1.genblk1.latch.q ;
 wire \shift_reg[61].genblk1.genblk1.latch.clk ;
 wire \shift_reg[61].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[61].genblk1.genblk1.latch.q ;
 wire \shift_reg[62].genblk1.genblk1.latch.clk ;
 wire \shift_reg[62].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[62].genblk1.genblk1.latch.q ;
 wire \shift_reg[63].genblk1.genblk1.latch.clk ;
 wire \shift_reg[63].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[63].genblk1.genblk1.latch.q ;
 wire \shift_reg[64].genblk1.genblk1.latch.clk ;
 wire \shift_reg[64].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[64].genblk1.genblk1.latch.q ;
 wire \shift_reg[65].genblk1.genblk1.latch.clk ;
 wire \shift_reg[65].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[65].genblk1.genblk1.latch.q ;
 wire \shift_reg[66].genblk1.genblk1.latch.clk ;
 wire \shift_reg[66].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[66].genblk1.genblk1.latch.q ;
 wire \shift_reg[67].genblk1.genblk1.latch.clk ;
 wire \shift_reg[67].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[67].genblk1.genblk1.latch.q ;
 wire \shift_reg[68].genblk1.genblk1.latch.clk ;
 wire \shift_reg[68].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[68].genblk1.genblk1.latch.q ;
 wire \shift_reg[69].genblk1.genblk1.latch.clk ;
 wire \shift_reg[69].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[69].genblk1.genblk1.latch.q ;
 wire \shift_reg[6].genblk1.genblk1.latch.clk ;
 wire \shift_reg[6].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[6].genblk1.genblk1.latch.q ;
 wire \shift_reg[70].genblk1.genblk1.latch.clk ;
 wire \shift_reg[70].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[70].genblk1.genblk1.latch.q ;
 wire \shift_reg[71].genblk1.genblk1.latch.clk ;
 wire \shift_reg[71].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[71].genblk1.genblk1.latch.q ;
 wire \shift_reg[72].genblk1.genblk1.latch.clk ;
 wire \shift_reg[72].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[72].genblk1.genblk1.latch.q ;
 wire \shift_reg[73].genblk1.genblk1.latch.clk ;
 wire \shift_reg[73].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[73].genblk1.genblk1.latch.q ;
 wire \shift_reg[74].genblk1.genblk1.latch.clk ;
 wire \shift_reg[74].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[74].genblk1.genblk1.latch.q ;
 wire \shift_reg[75].genblk1.genblk1.latch.clk ;
 wire \shift_reg[75].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[75].genblk1.genblk1.latch.q ;
 wire \shift_reg[76].genblk1.genblk1.latch.clk ;
 wire \shift_reg[76].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[76].genblk1.genblk1.latch.q ;
 wire \shift_reg[77].genblk1.genblk1.latch.clk ;
 wire \shift_reg[77].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[77].genblk1.genblk1.latch.q ;
 wire \shift_reg[78].genblk1.genblk1.latch.clk ;
 wire \shift_reg[78].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[78].genblk1.genblk1.latch.q ;
 wire \shift_reg[79].genblk1.genblk1.latch.clk ;
 wire \shift_reg[79].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[79].genblk1.genblk1.latch.q ;
 wire \shift_reg[7].genblk1.genblk1.latch.clk ;
 wire \shift_reg[7].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[7].genblk1.genblk1.latch.q ;
 wire \shift_reg[80].genblk1.genblk1.latch.clk ;
 wire \shift_reg[80].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[80].genblk1.genblk1.latch.q ;
 wire \shift_reg[81].genblk1.genblk1.latch.clk ;
 wire \shift_reg[81].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[81].genblk1.genblk1.latch.q ;
 wire \shift_reg[82].genblk1.genblk1.latch.clk ;
 wire \shift_reg[82].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[82].genblk1.genblk1.latch.q ;
 wire \shift_reg[83].genblk1.genblk1.latch.clk ;
 wire \shift_reg[83].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[83].genblk1.genblk1.latch.q ;
 wire \shift_reg[84].genblk1.genblk1.latch.clk ;
 wire \shift_reg[84].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[84].genblk1.genblk1.latch.q ;
 wire \shift_reg[85].genblk1.genblk1.latch.clk ;
 wire \shift_reg[85].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[85].genblk1.genblk1.latch.q ;
 wire \shift_reg[86].genblk1.genblk1.latch.clk ;
 wire \shift_reg[86].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[86].genblk1.genblk1.latch.q ;
 wire \shift_reg[87].genblk1.genblk1.latch.clk ;
 wire \shift_reg[87].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[87].genblk1.genblk1.latch.q ;
 wire \shift_reg[88].genblk1.genblk1.latch.clk ;
 wire \shift_reg[88].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[88].genblk1.genblk1.latch.q ;
 wire \shift_reg[89].genblk1.genblk1.latch.clk ;
 wire \shift_reg[89].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[89].genblk1.genblk1.latch.q ;
 wire \shift_reg[8].genblk1.genblk1.latch.clk ;
 wire \shift_reg[8].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[8].genblk1.genblk1.latch.q ;
 wire \shift_reg[90].genblk1.genblk1.latch.clk ;
 wire \shift_reg[90].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[90].genblk1.genblk1.latch.q ;
 wire \shift_reg[91].genblk1.genblk1.latch.clk ;
 wire \shift_reg[91].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[91].genblk1.genblk1.latch.q ;
 wire \shift_reg[92].genblk1.genblk1.latch.clk ;
 wire \shift_reg[92].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[92].genblk1.genblk1.latch.q ;
 wire \shift_reg[93].genblk1.genblk1.latch.clk ;
 wire \shift_reg[93].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[93].genblk1.genblk1.latch.q ;
 wire \shift_reg[94].genblk1.genblk1.latch.clk ;
 wire \shift_reg[94].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[94].genblk1.genblk1.latch.q ;
 wire \shift_reg[95].genblk1.genblk1.latch.clk ;
 wire \shift_reg[95].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[95].genblk1.genblk1.latch.q ;
 wire \shift_reg[96].genblk1.genblk1.latch.clk ;
 wire \shift_reg[96].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[96].genblk1.genblk1.latch.q ;
 wire \shift_reg[97].genblk1.genblk1.latch.clk ;
 wire \shift_reg[97].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[97].genblk1.genblk1.latch.q ;
 wire \shift_reg[98].genblk1.genblk1.latch.clk ;
 wire \shift_reg[98].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[98].genblk1.genblk1.latch.q ;
 wire \shift_reg[99].genblk1.genblk1.latch.nclk ;
 wire \shift_reg[9].genblk1.genblk1.latch.nclk ;
 wire trig_delayed;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net1;
 wire net2;
 wire net3;

 sg13g2_xor2_1 _000_ (.B(net2),
    .A(trig_delayed),
    .X(shift));
 sg13g2_dlhq_1 _001_ (.D(\shift_reg[386].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[387].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[387].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _002_ (.D(\shift_reg[387].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[388].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[388].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _003_ (.D(\shift_reg[388].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[389].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[389].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _004_ (.D(\shift_reg[389].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[390].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[390].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _005_ (.D(\shift_reg[390].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[391].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[391].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _006_ (.D(\shift_reg[391].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[392].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[392].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _007_ (.D(\shift_reg[392].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[393].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[393].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _008_ (.D(\shift_reg[393].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[394].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[394].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _009_ (.D(\shift_reg[394].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[395].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[395].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _010_ (.D(\shift_reg[395].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[396].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[396].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _011_ (.D(\shift_reg[396].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[397].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[397].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _012_ (.D(\shift_reg[397].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[398].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[398].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _013_ (.D(\shift_reg[398].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[399].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[399].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _014_ (.D(\shift_reg[399].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[400].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[400].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _015_ (.D(\shift_reg[400].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[401].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[401].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _016_ (.D(\shift_reg[401].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[402].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[402].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _017_ (.D(\shift_reg[402].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[403].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[403].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _018_ (.D(\shift_reg[403].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[404].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[404].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _019_ (.D(\shift_reg[404].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[405].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[405].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _020_ (.D(\shift_reg[405].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[406].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[406].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _021_ (.D(\shift_reg[406].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[407].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[407].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _022_ (.D(\shift_reg[407].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[408].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[408].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _023_ (.D(\shift_reg[408].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[409].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[409].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _024_ (.D(\shift_reg[409].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[410].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[410].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _025_ (.D(\shift_reg[410].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[411].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[411].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _026_ (.D(\shift_reg[411].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[412].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[412].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _027_ (.D(\shift_reg[412].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[413].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[413].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _028_ (.D(\shift_reg[413].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[414].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[414].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _029_ (.D(\shift_reg[414].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[415].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[415].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _030_ (.D(\shift_reg[415].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[416].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[416].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _031_ (.D(\shift_reg[416].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[417].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[417].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _032_ (.D(\shift_reg[417].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[418].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[418].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _033_ (.D(\shift_reg[418].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[419].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[419].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _034_ (.D(\shift_reg[419].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[420].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[420].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _035_ (.D(\shift_reg[420].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[421].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[421].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _036_ (.D(\shift_reg[421].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[422].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[422].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _037_ (.D(\shift_reg[422].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[423].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[423].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _038_ (.D(\shift_reg[423].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[424].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[424].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _039_ (.D(\shift_reg[424].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[425].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[425].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _040_ (.D(\shift_reg[425].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[426].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[426].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _041_ (.D(\shift_reg[426].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[427].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[427].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _042_ (.D(\shift_reg[427].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[428].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[428].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _043_ (.D(\shift_reg[428].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[429].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[429].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _044_ (.D(\shift_reg[429].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[430].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[430].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _045_ (.D(\shift_reg[430].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[431].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[431].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _046_ (.D(\shift_reg[431].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[432].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[432].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _047_ (.D(\shift_reg[432].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[433].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[433].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _048_ (.D(\shift_reg[433].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[434].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[434].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _049_ (.D(\shift_reg[434].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[435].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[435].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _050_ (.D(\shift_reg[435].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[436].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[436].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _051_ (.D(\shift_reg[436].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[437].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[437].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _052_ (.D(\shift_reg[437].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[438].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[438].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _053_ (.D(\shift_reg[438].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[439].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[439].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _054_ (.D(\shift_reg[439].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[440].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[440].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _055_ (.D(\shift_reg[440].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[441].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[441].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _056_ (.D(\shift_reg[441].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[442].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[442].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _057_ (.D(\shift_reg[442].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[443].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[443].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _058_ (.D(\shift_reg[443].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[444].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[444].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _059_ (.D(\shift_reg[444].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[445].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[445].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _060_ (.D(\shift_reg[445].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[446].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[446].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _061_ (.D(\shift_reg[446].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[447].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[447].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _062_ (.D(\shift_reg[447].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[448].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[448].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _063_ (.D(\shift_reg[448].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[449].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[449].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _064_ (.D(\shift_reg[449].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[450].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[450].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _065_ (.D(\shift_reg[450].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[451].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[451].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _066_ (.D(\shift_reg[451].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[452].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[452].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _067_ (.D(\shift_reg[452].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[453].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[453].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _068_ (.D(\shift_reg[453].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[454].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[454].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _069_ (.D(\shift_reg[454].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[455].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[455].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _070_ (.D(\shift_reg[455].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[456].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[456].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _071_ (.D(\shift_reg[456].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[457].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[457].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _072_ (.D(\shift_reg[457].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[458].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[458].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _073_ (.D(\shift_reg[458].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[459].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[459].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _074_ (.D(\shift_reg[459].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[460].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[460].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _075_ (.D(\shift_reg[460].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[461].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[461].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _076_ (.D(\shift_reg[461].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[462].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[462].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _077_ (.D(\shift_reg[462].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[463].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[463].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _078_ (.D(\shift_reg[463].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[464].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[464].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _079_ (.D(\shift_reg[464].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[465].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[465].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _080_ (.D(\shift_reg[465].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[466].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[466].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _081_ (.D(\shift_reg[466].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[467].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[467].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _082_ (.D(\shift_reg[467].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[468].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[468].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _083_ (.D(\shift_reg[468].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[469].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[469].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _084_ (.D(\shift_reg[469].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[470].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[470].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _085_ (.D(\shift_reg[470].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[471].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[471].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _086_ (.D(\shift_reg[471].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[472].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[472].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _087_ (.D(\shift_reg[472].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[473].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[473].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _088_ (.D(\shift_reg[473].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[474].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[474].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _089_ (.D(\shift_reg[474].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[475].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[475].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _090_ (.D(\shift_reg[475].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[476].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[476].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _091_ (.D(\shift_reg[476].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[477].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[477].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _092_ (.D(\shift_reg[477].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[478].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[478].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _093_ (.D(\shift_reg[478].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[479].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[479].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _094_ (.D(\shift_reg[479].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[480].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[480].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _095_ (.D(\shift_reg[480].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[481].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[481].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _096_ (.D(\shift_reg[481].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[482].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[482].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _097_ (.D(\shift_reg[482].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[483].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[483].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _098_ (.D(\shift_reg[483].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[484].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[484].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _099_ (.D(\shift_reg[484].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[485].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[485].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _100_ (.D(\shift_reg[485].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[486].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[486].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _101_ (.D(\shift_reg[486].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[487].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[487].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _102_ (.D(\shift_reg[487].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[488].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[488].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _103_ (.D(\shift_reg[488].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[489].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[489].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _104_ (.D(\shift_reg[489].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[490].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[490].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _105_ (.D(\shift_reg[490].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[491].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[491].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _106_ (.D(\shift_reg[491].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[492].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[492].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _107_ (.D(\shift_reg[492].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[493].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[493].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _108_ (.D(\shift_reg[493].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[494].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[494].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _109_ (.D(\shift_reg[494].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[495].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[495].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _110_ (.D(\shift_reg[495].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[496].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[496].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _111_ (.D(\shift_reg[496].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[497].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[497].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _112_ (.D(\shift_reg[497].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[498].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[498].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _113_ (.D(\shift_reg[498].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[499].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[499].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _114_ (.D(\shift_reg[499].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[500].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[500].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _115_ (.D(\shift_reg[500].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[501].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[501].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _116_ (.D(\shift_reg[501].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[502].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[502].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _117_ (.D(\shift_reg[502].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[503].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[503].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _118_ (.D(\shift_reg[503].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[504].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[504].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _119_ (.D(\shift_reg[504].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[505].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[505].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _120_ (.D(\shift_reg[505].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[506].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[506].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _121_ (.D(\shift_reg[506].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[507].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[507].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _122_ (.D(\shift_reg[507].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[508].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[508].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _123_ (.D(\shift_reg[508].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[509].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[509].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _124_ (.D(\shift_reg[509].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[510].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[510].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _125_ (.D(\shift_reg[510].genblk1.genblk1.latch.q ),
    .GATE(shift),
    .Q(\shift_reg[511].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _126_ (.D(net1),
    .GATE(\shift_reg[0].genblk1.latch.clk ),
    .Q(\shift_reg[0].genblk1.latch.q ));
 sg13g2_dlhq_1 _127_ (.D(\shift_reg[0].genblk1.latch.q ),
    .GATE(\shift_reg[1].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[1].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _128_ (.D(\shift_reg[1].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[2].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[2].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _129_ (.D(\shift_reg[2].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[3].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[3].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _130_ (.D(\shift_reg[3].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[4].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[4].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _131_ (.D(\shift_reg[4].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[5].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[5].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _132_ (.D(\shift_reg[5].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[6].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[6].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _133_ (.D(\shift_reg[6].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[7].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[7].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _134_ (.D(\shift_reg[7].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[8].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[8].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _135_ (.D(\shift_reg[8].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[10].genblk1.genblk1.latch.clkout ),
    .Q(\shift_reg[10].genblk1.genblk1.latch.d ));
 sg13g2_dlhq_1 _136_ (.D(\shift_reg[10].genblk1.genblk1.latch.d ),
    .GATE(\shift_reg[10].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[10].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _137_ (.D(\shift_reg[10].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[11].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[11].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _138_ (.D(\shift_reg[11].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[12].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[12].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _139_ (.D(\shift_reg[12].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[13].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[13].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _140_ (.D(\shift_reg[13].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[14].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[14].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _141_ (.D(\shift_reg[14].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[15].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[15].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _142_ (.D(\shift_reg[15].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[16].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[16].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _143_ (.D(\shift_reg[16].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[17].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[17].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _144_ (.D(\shift_reg[17].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[18].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[18].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _145_ (.D(\shift_reg[18].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[19].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[19].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _146_ (.D(\shift_reg[19].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[20].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[20].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _147_ (.D(\shift_reg[20].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[21].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[21].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _148_ (.D(\shift_reg[21].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[22].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[22].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _149_ (.D(\shift_reg[22].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[23].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[23].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _150_ (.D(\shift_reg[23].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[24].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[24].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _151_ (.D(\shift_reg[24].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[25].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[25].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _152_ (.D(\shift_reg[25].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[26].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[26].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _153_ (.D(\shift_reg[26].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[27].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[27].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _154_ (.D(\shift_reg[27].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[28].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[28].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _155_ (.D(\shift_reg[28].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[29].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[29].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _156_ (.D(\shift_reg[29].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[30].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[30].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _157_ (.D(\shift_reg[30].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[31].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[31].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _158_ (.D(\shift_reg[31].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[32].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[32].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _159_ (.D(\shift_reg[32].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[33].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[33].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _160_ (.D(\shift_reg[33].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[34].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[34].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _161_ (.D(\shift_reg[34].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[35].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[35].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _162_ (.D(\shift_reg[35].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[36].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[36].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _163_ (.D(\shift_reg[36].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[37].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[37].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _164_ (.D(\shift_reg[37].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[38].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[38].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _165_ (.D(\shift_reg[38].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[39].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[39].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _166_ (.D(\shift_reg[39].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[40].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[40].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _167_ (.D(\shift_reg[40].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[41].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[41].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _168_ (.D(\shift_reg[41].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[42].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[42].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _169_ (.D(\shift_reg[42].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[43].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[43].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _170_ (.D(\shift_reg[43].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[44].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[44].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _171_ (.D(\shift_reg[44].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[45].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[45].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _172_ (.D(\shift_reg[45].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[46].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[46].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _173_ (.D(\shift_reg[46].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[47].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[47].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _174_ (.D(\shift_reg[47].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[48].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[48].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _175_ (.D(\shift_reg[48].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[49].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[49].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _176_ (.D(\shift_reg[49].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[50].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[50].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _177_ (.D(\shift_reg[50].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[51].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[51].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _178_ (.D(\shift_reg[51].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[52].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[52].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _179_ (.D(\shift_reg[52].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[53].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[53].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _180_ (.D(\shift_reg[53].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[54].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[54].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _181_ (.D(\shift_reg[54].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[55].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[55].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _182_ (.D(\shift_reg[55].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[56].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[56].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _183_ (.D(\shift_reg[56].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[57].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[57].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _184_ (.D(\shift_reg[57].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[58].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[58].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _185_ (.D(\shift_reg[58].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[59].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[59].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _186_ (.D(\shift_reg[59].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[60].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[60].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _187_ (.D(\shift_reg[60].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[61].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[61].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _188_ (.D(\shift_reg[61].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[62].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[62].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _189_ (.D(\shift_reg[62].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[63].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[63].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _190_ (.D(\shift_reg[63].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[64].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[64].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _191_ (.D(\shift_reg[64].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[65].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[65].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _192_ (.D(\shift_reg[65].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[66].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[66].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _193_ (.D(\shift_reg[66].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[67].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[67].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _194_ (.D(\shift_reg[67].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[68].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[68].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _195_ (.D(\shift_reg[68].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[69].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[69].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _196_ (.D(\shift_reg[69].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[70].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[70].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _197_ (.D(\shift_reg[70].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[71].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[71].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _198_ (.D(\shift_reg[71].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[72].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[72].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _199_ (.D(\shift_reg[72].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[73].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[73].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _200_ (.D(\shift_reg[73].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[74].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[74].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _201_ (.D(\shift_reg[74].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[75].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[75].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _202_ (.D(\shift_reg[75].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[76].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[76].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _203_ (.D(\shift_reg[76].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[77].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[77].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _204_ (.D(\shift_reg[77].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[78].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[78].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _205_ (.D(\shift_reg[78].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[79].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[79].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _206_ (.D(\shift_reg[79].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[80].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[80].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _207_ (.D(\shift_reg[80].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[81].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[81].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _208_ (.D(\shift_reg[81].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[82].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[82].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _209_ (.D(\shift_reg[82].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[83].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[83].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _210_ (.D(\shift_reg[83].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[84].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[84].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _211_ (.D(\shift_reg[84].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[85].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[85].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _212_ (.D(\shift_reg[85].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[86].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[86].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _213_ (.D(\shift_reg[86].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[87].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[87].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _214_ (.D(\shift_reg[87].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[88].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[88].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _215_ (.D(\shift_reg[88].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[89].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[89].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _216_ (.D(\shift_reg[89].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[90].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[90].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _217_ (.D(\shift_reg[90].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[91].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[91].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _218_ (.D(\shift_reg[91].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[92].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[92].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _219_ (.D(\shift_reg[92].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[93].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[93].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _220_ (.D(\shift_reg[93].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[94].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[94].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _221_ (.D(\shift_reg[94].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[95].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[95].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _222_ (.D(\shift_reg[95].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[96].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[96].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _223_ (.D(\shift_reg[96].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[97].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[97].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _224_ (.D(\shift_reg[97].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[98].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[98].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _225_ (.D(\shift_reg[98].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[100].genblk1.genblk1.latch.clkout ),
    .Q(\shift_reg[100].genblk1.genblk1.latch.d ));
 sg13g2_dlhq_1 _226_ (.D(\shift_reg[100].genblk1.genblk1.latch.d ),
    .GATE(\shift_reg[100].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[100].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _227_ (.D(\shift_reg[100].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[101].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[101].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _228_ (.D(\shift_reg[101].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[102].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[102].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _229_ (.D(\shift_reg[102].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[103].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[103].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _230_ (.D(\shift_reg[103].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[104].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[104].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _231_ (.D(\shift_reg[104].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[105].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[105].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _232_ (.D(\shift_reg[105].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[106].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[106].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _233_ (.D(\shift_reg[106].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[107].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[107].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _234_ (.D(\shift_reg[107].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[108].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[108].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _235_ (.D(\shift_reg[108].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[109].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[109].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _236_ (.D(\shift_reg[109].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[110].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[110].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _237_ (.D(\shift_reg[110].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[111].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[111].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _238_ (.D(\shift_reg[111].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[112].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[112].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _239_ (.D(\shift_reg[112].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[113].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[113].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _240_ (.D(\shift_reg[113].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[114].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[114].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _241_ (.D(\shift_reg[114].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[115].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[115].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _242_ (.D(\shift_reg[115].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[116].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[116].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _243_ (.D(\shift_reg[116].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[117].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[117].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _244_ (.D(\shift_reg[117].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[118].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[118].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _245_ (.D(\shift_reg[118].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[119].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[119].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _246_ (.D(\shift_reg[119].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[120].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[120].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _247_ (.D(\shift_reg[120].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[121].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[121].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _248_ (.D(\shift_reg[121].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[122].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[122].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _249_ (.D(\shift_reg[122].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[123].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[123].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _250_ (.D(\shift_reg[123].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[124].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[124].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _251_ (.D(\shift_reg[124].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[125].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[125].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _252_ (.D(\shift_reg[125].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[126].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[126].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _253_ (.D(\shift_reg[126].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[127].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[127].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _254_ (.D(\shift_reg[127].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[128].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[128].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _255_ (.D(\shift_reg[128].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[129].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[129].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _256_ (.D(\shift_reg[129].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[130].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[130].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _257_ (.D(\shift_reg[130].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[131].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[131].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _258_ (.D(\shift_reg[131].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[132].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[132].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _259_ (.D(\shift_reg[132].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[133].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[133].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _260_ (.D(\shift_reg[133].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[134].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[134].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _261_ (.D(\shift_reg[134].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[135].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[135].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _262_ (.D(\shift_reg[135].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[136].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[136].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _263_ (.D(\shift_reg[136].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[137].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[137].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _264_ (.D(\shift_reg[137].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[138].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[138].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _265_ (.D(\shift_reg[138].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[139].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[139].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _266_ (.D(\shift_reg[139].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[140].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[140].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _267_ (.D(\shift_reg[140].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[141].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[141].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _268_ (.D(\shift_reg[141].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[142].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[142].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _269_ (.D(\shift_reg[142].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[143].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[143].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _270_ (.D(\shift_reg[143].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[144].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[144].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _271_ (.D(\shift_reg[144].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[145].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[145].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _272_ (.D(\shift_reg[145].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[146].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[146].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _273_ (.D(\shift_reg[146].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[147].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[147].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _274_ (.D(\shift_reg[147].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[148].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[148].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _275_ (.D(\shift_reg[148].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[149].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[149].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _276_ (.D(\shift_reg[149].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[150].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[150].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _277_ (.D(\shift_reg[150].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[151].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[151].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _278_ (.D(\shift_reg[151].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[152].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[152].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _279_ (.D(\shift_reg[152].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[153].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[153].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _280_ (.D(\shift_reg[153].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[154].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[154].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _281_ (.D(\shift_reg[154].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[155].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[155].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _282_ (.D(\shift_reg[155].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[156].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[156].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _283_ (.D(\shift_reg[156].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[157].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[157].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _284_ (.D(\shift_reg[157].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[158].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[158].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _285_ (.D(\shift_reg[158].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[159].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[159].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _286_ (.D(\shift_reg[159].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[160].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[160].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _287_ (.D(\shift_reg[160].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[161].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[161].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _288_ (.D(\shift_reg[161].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[162].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[162].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _289_ (.D(\shift_reg[162].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[163].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[163].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _290_ (.D(\shift_reg[163].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[164].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[164].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _291_ (.D(\shift_reg[164].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[165].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[165].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _292_ (.D(\shift_reg[165].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[166].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[166].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _293_ (.D(\shift_reg[166].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[167].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[167].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _294_ (.D(\shift_reg[167].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[168].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[168].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _295_ (.D(\shift_reg[168].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[169].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[169].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _296_ (.D(\shift_reg[169].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[170].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[170].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _297_ (.D(\shift_reg[170].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[171].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[171].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _298_ (.D(\shift_reg[171].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[172].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[172].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _299_ (.D(\shift_reg[172].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[173].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[173].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _300_ (.D(\shift_reg[173].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[174].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[174].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _301_ (.D(\shift_reg[174].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[175].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[175].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _302_ (.D(\shift_reg[175].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[176].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[176].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _303_ (.D(\shift_reg[176].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[177].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[177].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _304_ (.D(\shift_reg[177].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[178].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[178].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _305_ (.D(\shift_reg[178].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[179].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[179].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _306_ (.D(\shift_reg[179].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[180].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[180].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _307_ (.D(\shift_reg[180].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[181].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[181].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _308_ (.D(\shift_reg[181].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[182].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[182].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _309_ (.D(\shift_reg[182].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[183].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[183].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _310_ (.D(\shift_reg[183].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[184].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[184].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _311_ (.D(\shift_reg[184].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[185].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[185].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _312_ (.D(\shift_reg[185].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[186].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[186].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _313_ (.D(\shift_reg[186].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[187].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[187].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _314_ (.D(\shift_reg[187].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[188].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[188].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _315_ (.D(\shift_reg[188].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[189].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[189].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _316_ (.D(\shift_reg[189].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[190].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[190].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _317_ (.D(\shift_reg[190].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[191].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[191].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _318_ (.D(\shift_reg[191].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[192].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[192].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _319_ (.D(\shift_reg[192].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[193].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[193].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _320_ (.D(\shift_reg[193].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[194].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[194].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _321_ (.D(\shift_reg[194].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[195].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[195].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _322_ (.D(\shift_reg[195].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[196].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[196].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _323_ (.D(\shift_reg[196].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[197].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[197].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _324_ (.D(\shift_reg[197].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[198].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[198].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _325_ (.D(\shift_reg[198].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[199].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[199].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _326_ (.D(\shift_reg[199].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[200].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[200].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _327_ (.D(\shift_reg[200].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[201].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[201].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _328_ (.D(\shift_reg[201].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[202].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[202].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _329_ (.D(\shift_reg[202].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[203].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[203].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _330_ (.D(\shift_reg[203].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[204].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[204].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _331_ (.D(\shift_reg[204].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[205].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[205].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _332_ (.D(\shift_reg[205].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[206].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[206].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _333_ (.D(\shift_reg[206].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[207].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[207].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _334_ (.D(\shift_reg[207].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[208].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[208].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _335_ (.D(\shift_reg[208].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[209].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[209].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _336_ (.D(\shift_reg[209].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[210].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[210].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _337_ (.D(\shift_reg[210].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[211].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[211].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _338_ (.D(\shift_reg[211].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[212].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[212].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _339_ (.D(\shift_reg[212].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[213].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[213].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _340_ (.D(\shift_reg[213].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[214].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[214].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _341_ (.D(\shift_reg[214].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[215].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[215].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _342_ (.D(\shift_reg[215].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[216].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[216].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _343_ (.D(\shift_reg[216].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[217].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[217].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _344_ (.D(\shift_reg[217].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[218].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[218].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _345_ (.D(\shift_reg[218].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[219].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[219].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _346_ (.D(\shift_reg[219].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[220].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[220].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _347_ (.D(\shift_reg[220].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[221].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[221].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _348_ (.D(\shift_reg[221].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[222].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[222].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _349_ (.D(\shift_reg[222].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[223].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[223].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _350_ (.D(\shift_reg[223].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[224].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[224].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _351_ (.D(\shift_reg[224].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[225].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[225].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _352_ (.D(\shift_reg[225].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[226].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[226].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _353_ (.D(\shift_reg[226].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[227].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[227].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _354_ (.D(\shift_reg[227].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[228].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[228].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _355_ (.D(\shift_reg[228].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[229].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[229].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _356_ (.D(\shift_reg[229].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[230].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[230].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _357_ (.D(\shift_reg[230].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[231].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[231].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _358_ (.D(\shift_reg[231].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[232].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[232].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _359_ (.D(\shift_reg[232].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[233].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[233].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _360_ (.D(\shift_reg[233].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[234].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[234].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _361_ (.D(\shift_reg[234].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[235].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[235].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _362_ (.D(\shift_reg[235].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[236].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[236].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _363_ (.D(\shift_reg[236].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[237].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[237].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _364_ (.D(\shift_reg[237].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[238].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[238].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _365_ (.D(\shift_reg[238].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[239].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[239].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _366_ (.D(\shift_reg[239].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[240].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[240].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _367_ (.D(\shift_reg[240].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[241].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[241].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _368_ (.D(\shift_reg[241].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[242].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[242].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _369_ (.D(\shift_reg[242].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[243].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[243].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _370_ (.D(\shift_reg[243].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[244].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[244].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _371_ (.D(\shift_reg[244].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[245].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[245].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _372_ (.D(\shift_reg[245].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[246].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[246].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _373_ (.D(\shift_reg[246].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[247].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[247].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _374_ (.D(\shift_reg[247].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[248].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[248].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _375_ (.D(\shift_reg[248].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[249].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[249].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _376_ (.D(\shift_reg[249].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[250].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[250].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _377_ (.D(\shift_reg[250].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[251].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[251].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _378_ (.D(\shift_reg[251].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[252].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[252].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _379_ (.D(\shift_reg[252].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[253].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[253].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _380_ (.D(\shift_reg[253].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[254].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[254].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _381_ (.D(\shift_reg[254].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[255].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[255].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _382_ (.D(\shift_reg[255].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[256].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[256].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _383_ (.D(\shift_reg[256].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[257].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[257].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _384_ (.D(\shift_reg[257].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[258].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[258].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _385_ (.D(\shift_reg[258].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[259].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[259].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _386_ (.D(\shift_reg[259].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[260].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[260].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _387_ (.D(\shift_reg[260].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[261].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[261].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _388_ (.D(\shift_reg[261].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[262].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[262].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _389_ (.D(\shift_reg[262].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[263].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[263].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _390_ (.D(\shift_reg[263].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[264].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[264].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _391_ (.D(\shift_reg[264].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[265].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[265].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _392_ (.D(\shift_reg[265].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[266].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[266].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _393_ (.D(\shift_reg[266].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[267].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[267].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _394_ (.D(\shift_reg[267].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[268].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[268].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _395_ (.D(\shift_reg[268].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[269].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[269].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _396_ (.D(\shift_reg[269].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[270].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[270].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _397_ (.D(\shift_reg[270].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[271].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[271].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _398_ (.D(\shift_reg[271].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[272].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[272].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _399_ (.D(\shift_reg[272].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[273].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[273].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _400_ (.D(\shift_reg[273].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[274].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[274].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _401_ (.D(\shift_reg[274].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[275].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[275].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _402_ (.D(\shift_reg[275].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[276].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[276].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _403_ (.D(\shift_reg[276].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[277].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[277].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _404_ (.D(\shift_reg[277].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[278].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[278].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _405_ (.D(\shift_reg[278].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[279].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[279].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _406_ (.D(\shift_reg[279].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[280].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[280].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _407_ (.D(\shift_reg[280].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[281].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[281].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _408_ (.D(\shift_reg[281].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[282].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[282].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _409_ (.D(\shift_reg[282].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[283].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[283].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _410_ (.D(\shift_reg[283].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[284].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[284].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _411_ (.D(\shift_reg[284].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[285].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[285].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _412_ (.D(\shift_reg[285].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[286].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[286].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _413_ (.D(\shift_reg[286].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[287].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[287].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _414_ (.D(\shift_reg[287].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[288].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[288].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _415_ (.D(\shift_reg[288].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[289].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[289].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _416_ (.D(\shift_reg[289].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[290].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[290].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _417_ (.D(\shift_reg[290].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[291].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[291].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _418_ (.D(\shift_reg[291].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[292].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[292].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _419_ (.D(\shift_reg[292].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[293].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[293].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _420_ (.D(\shift_reg[293].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[294].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[294].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _421_ (.D(\shift_reg[294].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[295].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[295].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _422_ (.D(\shift_reg[295].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[296].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[296].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _423_ (.D(\shift_reg[296].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[297].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[297].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _424_ (.D(\shift_reg[297].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[298].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[298].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _425_ (.D(\shift_reg[298].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[299].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[299].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _426_ (.D(\shift_reg[299].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[300].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[300].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _427_ (.D(\shift_reg[300].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[301].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[301].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _428_ (.D(\shift_reg[301].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[302].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[302].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _429_ (.D(\shift_reg[302].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[303].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[303].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _430_ (.D(\shift_reg[303].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[304].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[304].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _431_ (.D(\shift_reg[304].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[305].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[305].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _432_ (.D(\shift_reg[305].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[306].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[306].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _433_ (.D(\shift_reg[306].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[307].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[307].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _434_ (.D(\shift_reg[307].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[308].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[308].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _435_ (.D(\shift_reg[308].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[309].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[309].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _436_ (.D(\shift_reg[309].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[310].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[310].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _437_ (.D(\shift_reg[310].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[311].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[311].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _438_ (.D(\shift_reg[311].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[312].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[312].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _439_ (.D(\shift_reg[312].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[313].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[313].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _440_ (.D(\shift_reg[313].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[314].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[314].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _441_ (.D(\shift_reg[314].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[315].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[315].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _442_ (.D(\shift_reg[315].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[316].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[316].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _443_ (.D(\shift_reg[316].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[317].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[317].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _444_ (.D(\shift_reg[317].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[318].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[318].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _445_ (.D(\shift_reg[318].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[319].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[319].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _446_ (.D(\shift_reg[319].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[320].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[320].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _447_ (.D(\shift_reg[320].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[321].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[321].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _448_ (.D(\shift_reg[321].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[322].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[322].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _449_ (.D(\shift_reg[322].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[323].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[323].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _450_ (.D(\shift_reg[323].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[324].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[324].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _451_ (.D(\shift_reg[324].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[325].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[325].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _452_ (.D(\shift_reg[325].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[326].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[326].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _453_ (.D(\shift_reg[326].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[327].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[327].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _454_ (.D(\shift_reg[327].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[328].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[328].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _455_ (.D(\shift_reg[328].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[329].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[329].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _456_ (.D(\shift_reg[329].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[330].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[330].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _457_ (.D(\shift_reg[330].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[331].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[331].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _458_ (.D(\shift_reg[331].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[332].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[332].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _459_ (.D(\shift_reg[332].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[333].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[333].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _460_ (.D(\shift_reg[333].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[334].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[334].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _461_ (.D(\shift_reg[334].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[335].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[335].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _462_ (.D(\shift_reg[335].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[336].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[336].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _463_ (.D(\shift_reg[336].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[337].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[337].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _464_ (.D(\shift_reg[337].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[338].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[338].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _465_ (.D(\shift_reg[338].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[339].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[339].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _466_ (.D(\shift_reg[339].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[340].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[340].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _467_ (.D(\shift_reg[340].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[341].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[341].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _468_ (.D(\shift_reg[341].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[342].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[342].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _469_ (.D(\shift_reg[342].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[343].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[343].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _470_ (.D(\shift_reg[343].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[344].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[344].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _471_ (.D(\shift_reg[344].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[345].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[345].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _472_ (.D(\shift_reg[345].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[346].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[346].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _473_ (.D(\shift_reg[346].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[347].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[347].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _474_ (.D(\shift_reg[347].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[348].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[348].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _475_ (.D(\shift_reg[348].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[349].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[349].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _476_ (.D(\shift_reg[349].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[350].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[350].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _477_ (.D(\shift_reg[350].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[351].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[351].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _478_ (.D(\shift_reg[351].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[352].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[352].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _479_ (.D(\shift_reg[352].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[353].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[353].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _480_ (.D(\shift_reg[353].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[354].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[354].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _481_ (.D(\shift_reg[354].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[355].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[355].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _482_ (.D(\shift_reg[355].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[356].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[356].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _483_ (.D(\shift_reg[356].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[357].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[357].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _484_ (.D(\shift_reg[357].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[358].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[358].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _485_ (.D(\shift_reg[358].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[359].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[359].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _486_ (.D(\shift_reg[359].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[360].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[360].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _487_ (.D(\shift_reg[360].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[361].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[361].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _488_ (.D(\shift_reg[361].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[362].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[362].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _489_ (.D(\shift_reg[362].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[363].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[363].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _490_ (.D(\shift_reg[363].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[364].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[364].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _491_ (.D(\shift_reg[364].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[365].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[365].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _492_ (.D(\shift_reg[365].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[366].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[366].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _493_ (.D(\shift_reg[366].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[367].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[367].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _494_ (.D(\shift_reg[367].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[368].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[368].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _495_ (.D(\shift_reg[368].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[369].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[369].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _496_ (.D(\shift_reg[369].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[370].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[370].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _497_ (.D(\shift_reg[370].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[371].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[371].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _498_ (.D(\shift_reg[371].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[372].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[372].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _499_ (.D(\shift_reg[372].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[373].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[373].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _500_ (.D(\shift_reg[373].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[374].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[374].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _501_ (.D(\shift_reg[374].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[375].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[375].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _502_ (.D(\shift_reg[375].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[376].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[376].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _503_ (.D(\shift_reg[376].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[377].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[377].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _504_ (.D(\shift_reg[377].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[378].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[378].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _505_ (.D(\shift_reg[378].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[379].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[379].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _506_ (.D(\shift_reg[379].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[380].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[380].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _507_ (.D(\shift_reg[380].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[381].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[381].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _508_ (.D(\shift_reg[381].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[382].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[382].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _509_ (.D(\shift_reg[382].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[383].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[383].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _510_ (.D(\shift_reg[383].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[384].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[384].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _511_ (.D(\shift_reg[384].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[385].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[385].genblk1.genblk1.latch.q ));
 sg13g2_dlhq_1 _512_ (.D(\shift_reg[385].genblk1.genblk1.latch.q ),
    .GATE(\shift_reg[386].genblk1.genblk1.latch.clk ),
    .Q(\shift_reg[386].genblk1.genblk1.latch.q ));
 sg13g2_tielo tt_um_cattuto_sr_latch_4 (.L_LO(net4));
 sg13g2_tielo tt_um_cattuto_sr_latch_5 (.L_LO(net5));
 sg13g2_tielo tt_um_cattuto_sr_latch_6 (.L_LO(net6));
 sg13g2_tielo tt_um_cattuto_sr_latch_7 (.L_LO(net7));
 sg13g2_tielo tt_um_cattuto_sr_latch_8 (.L_LO(net8));
 sg13g2_tielo tt_um_cattuto_sr_latch_9 (.L_LO(net9));
 sg13g2_tielo tt_um_cattuto_sr_latch_10 (.L_LO(net10));
 sg13g2_tielo tt_um_cattuto_sr_latch_11 (.L_LO(net11));
 sg13g2_tielo tt_um_cattuto_sr_latch_12 (.L_LO(net12));
 sg13g2_tielo tt_um_cattuto_sr_latch_13 (.L_LO(net13));
 sg13g2_tielo tt_um_cattuto_sr_latch_14 (.L_LO(net14));
 sg13g2_tielo tt_um_cattuto_sr_latch_15 (.L_LO(net15));
 sg13g2_tielo tt_um_cattuto_sr_latch_16 (.L_LO(net16));
 sg13g2_tielo tt_um_cattuto_sr_latch_17 (.L_LO(net17));
 sg13g2_tielo tt_um_cattuto_sr_latch_18 (.L_LO(net18));
 sg13g2_tielo tt_um_cattuto_sr_latch_19 (.L_LO(net19));
 sg13g2_tielo tt_um_cattuto_sr_latch_20 (.L_LO(net20));
 sg13g2_tielo tt_um_cattuto_sr_latch_21 (.L_LO(net21));
 sg13g2_tielo tt_um_cattuto_sr_latch_22 (.L_LO(net22));
 sg13g2_tielo tt_um_cattuto_sr_latch_23 (.L_LO(net23));
 sg13g2_tielo tt_um_cattuto_sr_latch_24 (.L_LO(net24));
 sg13g2_tielo tt_um_cattuto_sr_latch_25 (.L_LO(net25));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 _536_ (.A(\shift_reg[511].genblk1.genblk1.latch.q ),
    .X(uo_out[0]));
 sg13g2_inv_1 \shift_reg[100].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[100].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[100].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[100].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[100].genblk1.genblk1.latch.clkout ),
    .A(\shift_reg[100].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[101].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[101].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[101].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[101].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[100].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[101].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[102].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[102].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[102].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[102].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[101].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[102].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[103].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[103].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[103].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[103].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[102].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[103].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[104].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[104].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[104].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[104].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[103].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[104].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[105].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[105].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[105].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[105].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[104].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[105].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[106].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[106].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[106].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[106].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[105].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[106].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[107].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[107].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[107].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[107].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[106].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[107].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[108].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[108].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[108].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[108].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[107].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[108].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[109].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[109].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[109].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[109].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[108].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[109].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[10].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[10].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[10].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[10].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[10].genblk1.genblk1.latch.clkout ),
    .A(\shift_reg[10].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[110].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[110].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[110].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[110].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[109].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[110].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[111].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[111].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[111].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[111].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[110].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[111].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[112].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[112].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[112].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[112].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[111].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[112].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[113].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[113].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[113].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[113].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[112].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[113].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[114].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[114].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[114].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[114].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[113].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[114].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[115].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[115].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[115].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[115].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[114].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[115].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[116].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[116].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[116].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[116].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[115].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[116].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[117].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[117].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[117].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[117].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[116].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[117].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[118].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[118].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[118].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[118].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[117].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[118].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[119].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[119].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[119].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[119].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[118].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[119].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[11].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[11].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[11].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[11].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[10].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[11].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[120].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[120].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[120].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[120].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[119].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[120].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[121].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[121].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[121].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[121].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[120].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[121].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[122].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[122].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[122].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[122].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[121].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[122].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[123].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[123].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[123].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[123].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[122].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[123].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[124].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[124].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[124].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[124].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[123].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[124].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[125].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[125].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[125].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[125].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[124].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[125].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[126].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[126].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[126].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[126].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[125].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[126].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[127].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[127].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[127].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[127].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[126].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[127].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[128].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[128].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[128].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[128].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[127].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[128].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[129].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[129].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[129].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[129].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[128].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[129].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[12].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[12].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[12].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[12].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[11].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[12].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[130].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[130].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[130].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[130].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[129].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[130].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[131].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[131].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[131].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[131].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[130].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[131].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[132].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[132].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[132].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[132].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[131].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[132].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[133].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[133].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[133].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[133].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[132].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[133].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[134].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[134].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[134].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[134].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[133].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[134].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[135].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[135].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[135].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[135].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[134].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[135].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[136].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[136].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[136].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[136].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[135].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[136].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[137].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[137].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[137].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[137].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[136].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[137].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[138].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[138].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[138].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[138].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[137].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[138].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[139].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[139].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[139].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[139].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[138].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[139].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[13].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[13].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[13].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[13].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[12].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[13].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[140].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[140].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[140].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[140].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[139].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[140].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[141].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[141].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[141].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[141].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[140].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[141].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[142].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[142].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[142].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[142].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[141].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[142].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[143].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[143].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[143].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[143].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[142].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[143].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[144].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[144].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[144].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[144].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[143].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[144].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[145].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[145].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[145].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[145].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[144].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[145].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[146].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[146].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[146].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[146].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[145].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[146].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[147].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[147].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[147].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[147].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[146].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[147].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[148].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[148].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[148].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[148].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[147].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[148].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[149].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[149].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[149].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[149].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[148].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[149].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[14].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[14].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[14].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[14].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[13].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[14].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[150].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[150].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[150].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[150].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[149].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[150].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[151].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[151].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[151].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[151].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[150].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[151].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[152].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[152].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[152].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[152].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[151].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[152].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[153].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[153].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[153].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[153].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[152].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[153].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[154].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[154].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[154].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[154].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[153].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[154].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[155].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[155].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[155].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[155].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[154].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[155].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[156].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[156].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[156].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[156].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[155].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[156].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[157].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[157].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[157].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[157].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[156].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[157].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[158].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[158].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[158].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[158].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[157].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[158].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[159].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[159].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[159].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[159].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[158].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[159].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[15].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[15].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[15].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[15].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[14].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[15].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[160].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[160].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[160].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[160].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[159].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[160].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[161].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[161].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[161].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[161].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[160].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[161].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[162].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[162].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[162].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[162].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[161].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[162].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[163].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[163].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[163].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[163].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[162].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[163].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[164].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[164].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[164].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[164].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[163].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[164].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[165].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[165].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[165].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[165].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[164].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[165].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[166].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[166].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[166].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[166].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[165].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[166].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[167].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[167].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[167].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[167].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[166].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[167].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[168].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[168].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[168].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[168].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[167].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[168].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[169].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[169].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[169].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[169].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[168].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[169].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[16].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[16].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[16].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[16].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[15].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[16].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[170].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[170].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[170].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[170].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[169].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[170].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[171].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[171].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[171].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[171].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[170].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[171].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[172].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[172].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[172].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[172].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[171].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[172].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[173].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[173].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[173].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[173].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[172].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[173].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[174].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[174].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[174].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[174].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[173].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[174].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[175].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[175].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[175].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[175].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[174].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[175].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[176].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[176].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[176].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[176].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[175].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[176].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[177].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[177].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[177].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[177].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[176].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[177].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[178].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[178].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[178].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[178].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[177].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[178].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[179].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[179].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[179].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[179].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[178].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[179].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[17].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[17].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[17].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[17].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[16].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[17].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[180].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[180].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[180].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[180].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[179].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[180].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[181].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[181].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[181].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[181].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[180].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[181].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[182].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[182].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[182].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[182].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[181].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[182].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[183].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[183].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[183].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[183].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[182].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[183].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[184].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[184].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[184].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[184].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[183].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[184].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[185].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[185].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[185].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[185].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[184].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[185].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[186].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[186].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[186].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[186].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[185].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[186].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[187].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[187].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[187].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[187].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[186].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[187].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[188].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[188].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[188].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[188].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[187].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[188].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[189].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[189].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[189].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[189].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[188].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[189].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[18].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[18].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[18].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[18].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[17].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[18].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[190].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[190].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[190].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[190].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[189].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[190].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[191].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[191].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[191].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[191].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[190].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[191].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[192].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[192].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[192].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[192].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[191].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[192].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[193].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[193].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[193].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[193].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[192].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[193].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[194].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[194].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[194].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[194].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[193].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[194].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[195].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[195].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[195].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[195].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[194].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[195].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[196].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[196].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[196].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[196].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[195].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[196].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[197].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[197].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[197].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[197].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[196].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[197].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[198].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[198].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[198].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[198].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[197].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[198].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[199].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[199].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[199].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[199].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[198].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[199].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[19].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[19].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[19].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[19].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[18].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[19].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[1].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[1].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[1].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[1].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[0].genblk1.latch.clk ),
    .A(\shift_reg[1].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[200].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[200].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[200].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[200].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[199].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[200].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[201].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[201].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[201].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[201].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[200].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[201].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[202].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[202].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[202].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[202].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[201].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[202].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[203].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[203].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[203].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[203].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[202].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[203].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[204].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[204].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[204].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[204].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[203].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[204].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[205].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[205].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[205].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[205].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[204].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[205].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[206].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[206].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[206].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[206].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[205].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[206].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[207].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[207].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[207].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[207].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[206].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[207].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[208].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[208].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[208].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[208].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[207].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[208].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[209].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[209].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[209].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[209].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[208].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[209].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[20].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[20].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[20].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[20].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[19].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[20].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[210].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[210].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[210].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[210].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[209].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[210].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[211].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[211].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[211].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[211].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[210].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[211].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[212].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[212].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[212].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[212].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[211].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[212].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[213].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[213].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[213].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[213].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[212].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[213].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[214].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[214].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[214].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[214].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[213].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[214].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[215].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[215].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[215].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[215].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[214].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[215].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[216].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[216].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[216].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[216].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[215].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[216].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[217].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[217].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[217].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[217].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[216].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[217].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[218].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[218].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[218].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[218].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[217].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[218].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[219].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[219].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[219].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[219].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[218].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[219].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[21].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[21].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[21].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[21].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[20].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[21].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[220].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[220].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[220].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[220].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[219].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[220].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[221].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[221].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[221].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[221].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[220].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[221].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[222].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[222].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[222].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[222].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[221].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[222].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[223].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[223].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[223].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[223].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[222].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[223].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[224].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[224].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[224].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[224].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[223].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[224].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[225].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[225].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[225].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[225].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[224].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[225].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[226].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[226].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[226].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[226].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[225].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[226].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[227].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[227].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[227].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[227].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[226].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[227].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[228].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[228].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[228].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[228].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[227].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[228].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[229].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[229].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[229].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[229].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[228].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[229].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[22].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[22].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[22].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[22].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[21].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[22].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[230].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[230].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[230].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[230].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[229].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[230].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[231].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[231].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[231].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[231].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[230].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[231].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[232].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[232].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[232].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[232].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[231].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[232].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[233].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[233].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[233].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[233].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[232].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[233].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[234].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[234].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[234].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[234].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[233].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[234].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[235].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[235].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[235].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[235].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[234].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[235].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[236].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[236].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[236].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[236].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[235].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[236].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[237].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[237].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[237].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[237].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[236].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[237].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[238].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[238].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[238].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[238].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[237].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[238].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[239].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[239].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[239].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[239].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[238].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[239].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[23].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[23].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[23].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[23].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[22].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[23].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[240].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[240].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[240].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[240].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[239].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[240].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[241].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[241].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[241].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[241].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[240].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[241].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[242].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[242].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[242].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[242].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[241].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[242].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[243].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[243].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[243].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[243].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[242].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[243].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[244].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[244].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[244].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[244].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[243].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[244].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[245].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[245].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[245].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[245].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[244].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[245].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[246].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[246].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[246].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[246].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[245].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[246].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[247].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[247].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[247].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[247].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[246].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[247].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[248].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[248].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[248].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[248].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[247].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[248].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[249].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[249].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[249].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[249].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[248].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[249].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[24].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[24].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[24].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[24].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[23].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[24].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[250].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[250].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[250].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[250].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[249].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[250].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[251].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[251].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[251].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[251].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[250].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[251].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[252].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[252].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[252].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[252].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[251].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[252].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[253].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[253].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[253].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[253].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[252].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[253].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[254].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[254].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[254].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[254].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[253].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[254].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[255].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[255].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[255].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[255].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[254].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[255].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[256].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[256].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[256].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[256].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[255].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[256].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[257].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[257].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[257].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[257].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[256].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[257].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[258].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[258].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[258].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[258].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[257].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[258].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[259].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[259].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[259].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[259].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[258].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[259].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[25].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[25].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[25].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[25].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[24].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[25].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[260].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[260].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[260].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[260].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[259].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[260].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[261].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[261].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[261].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[261].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[260].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[261].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[262].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[262].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[262].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[262].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[261].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[262].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[263].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[263].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[263].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[263].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[262].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[263].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[264].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[264].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[264].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[264].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[263].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[264].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[265].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[265].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[265].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[265].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[264].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[265].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[266].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[266].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[266].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[266].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[265].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[266].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[267].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[267].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[267].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[267].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[266].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[267].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[268].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[268].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[268].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[268].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[267].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[268].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[269].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[269].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[269].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[269].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[268].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[269].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[26].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[26].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[26].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[26].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[25].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[26].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[270].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[270].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[270].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[270].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[269].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[270].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[271].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[271].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[271].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[271].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[270].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[271].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[272].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[272].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[272].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[272].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[271].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[272].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[273].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[273].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[273].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[273].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[272].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[273].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[274].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[274].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[274].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[274].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[273].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[274].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[275].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[275].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[275].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[275].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[274].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[275].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[276].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[276].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[276].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[276].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[275].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[276].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[277].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[277].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[277].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[277].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[276].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[277].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[278].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[278].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[278].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[278].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[277].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[278].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[279].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[279].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[279].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[279].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[278].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[279].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[27].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[27].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[27].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[27].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[26].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[27].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[280].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[280].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[280].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[280].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[279].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[280].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[281].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[281].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[281].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[281].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[280].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[281].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[282].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[282].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[282].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[282].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[281].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[282].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[283].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[283].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[283].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[283].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[282].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[283].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[284].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[284].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[284].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[284].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[283].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[284].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[285].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[285].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[285].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[285].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[284].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[285].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[286].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[286].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[286].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[286].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[285].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[286].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[287].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[287].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[287].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[287].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[286].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[287].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[288].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[288].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[288].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[288].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[287].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[288].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[289].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[289].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[289].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[289].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[288].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[289].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[28].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[28].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[28].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[28].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[27].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[28].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[290].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[290].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[290].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[290].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[289].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[290].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[291].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[291].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[291].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[291].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[290].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[291].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[292].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[292].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[292].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[292].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[291].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[292].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[293].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[293].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[293].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[293].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[292].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[293].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[294].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[294].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[294].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[294].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[293].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[294].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[295].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[295].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[295].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[295].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[294].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[295].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[296].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[296].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[296].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[296].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[295].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[296].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[297].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[297].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[297].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[297].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[296].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[297].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[298].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[298].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[298].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[298].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[297].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[298].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[299].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[299].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[299].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[299].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[298].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[299].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[29].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[29].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[29].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[29].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[28].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[29].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[2].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[2].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[2].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[2].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[1].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[2].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[300].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[300].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[300].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[300].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[299].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[300].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[301].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[301].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[301].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[301].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[300].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[301].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[302].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[302].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[302].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[302].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[301].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[302].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[303].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[303].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[303].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[303].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[302].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[303].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[304].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[304].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[304].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[304].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[303].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[304].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[305].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[305].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[305].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[305].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[304].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[305].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[306].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[306].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[306].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[306].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[305].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[306].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[307].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[307].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[307].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[307].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[306].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[307].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[308].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[308].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[308].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[308].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[307].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[308].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[309].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[309].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[309].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[309].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[308].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[309].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[30].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[30].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[30].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[30].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[29].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[30].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[310].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[310].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[310].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[310].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[309].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[310].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[311].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[311].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[311].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[311].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[310].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[311].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[312].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[312].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[312].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[312].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[311].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[312].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[313].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[313].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[313].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[313].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[312].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[313].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[314].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[314].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[314].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[314].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[313].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[314].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[315].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[315].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[315].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[315].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[314].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[315].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[316].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[316].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[316].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[316].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[315].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[316].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[317].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[317].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[317].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[317].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[316].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[317].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[318].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[318].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[318].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[318].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[317].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[318].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[319].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[319].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[319].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[319].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[318].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[319].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[31].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[31].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[31].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[31].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[30].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[31].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[320].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[320].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[320].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[320].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[319].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[320].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[321].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[321].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[321].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[321].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[320].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[321].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[322].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[322].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[322].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[322].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[321].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[322].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[323].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[323].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[323].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[323].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[322].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[323].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[324].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[324].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[324].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[324].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[323].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[324].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[325].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[325].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[325].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[325].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[324].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[325].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[326].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[326].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[326].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[326].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[325].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[326].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[327].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[327].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[327].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[327].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[326].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[327].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[328].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[328].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[328].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[328].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[327].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[328].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[329].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[329].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[329].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[329].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[328].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[329].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[32].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[32].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[32].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[32].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[31].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[32].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[330].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[330].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[330].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[330].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[329].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[330].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[331].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[331].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[331].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[331].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[330].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[331].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[332].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[332].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[332].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[332].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[331].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[332].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[333].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[333].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[333].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[333].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[332].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[333].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[334].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[334].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[334].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[334].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[333].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[334].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[335].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[335].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[335].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[335].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[334].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[335].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[336].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[336].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[336].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[336].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[335].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[336].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[337].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[337].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[337].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[337].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[336].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[337].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[338].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[338].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[338].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[338].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[337].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[338].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[339].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[339].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[339].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[339].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[338].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[339].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[33].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[33].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[33].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[33].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[32].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[33].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[340].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[340].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[340].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[340].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[339].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[340].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[341].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[341].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[341].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[341].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[340].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[341].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[342].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[342].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[342].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[342].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[341].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[342].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[343].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[343].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[343].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[343].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[342].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[343].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[344].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[344].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[344].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[344].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[343].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[344].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[345].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[345].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[345].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[345].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[344].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[345].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[346].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[346].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[346].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[346].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[345].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[346].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[347].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[347].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[347].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[347].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[346].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[347].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[348].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[348].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[348].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[348].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[347].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[348].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[349].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[349].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[349].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[349].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[348].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[349].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[34].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[34].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[34].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[34].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[33].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[34].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[350].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[350].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[350].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[350].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[349].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[350].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[351].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[351].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[351].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[351].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[350].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[351].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[352].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[352].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[352].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[352].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[351].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[352].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[353].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[353].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[353].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[353].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[352].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[353].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[354].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[354].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[354].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[354].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[353].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[354].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[355].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[355].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[355].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[355].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[354].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[355].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[356].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[356].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[356].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[356].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[355].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[356].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[357].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[357].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[357].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[357].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[356].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[357].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[358].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[358].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[358].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[358].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[357].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[358].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[359].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[359].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[359].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[359].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[358].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[359].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[35].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[35].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[35].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[35].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[34].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[35].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[360].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[360].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[360].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[360].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[359].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[360].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[361].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[361].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[361].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[361].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[360].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[361].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[362].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[362].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[362].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[362].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[361].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[362].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[363].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[363].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[363].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[363].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[362].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[363].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[364].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[364].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[364].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[364].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[363].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[364].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[365].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[365].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[365].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[365].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[364].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[365].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[366].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[366].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[366].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[366].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[365].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[366].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[367].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[367].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[367].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[367].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[366].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[367].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[368].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[368].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[368].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[368].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[367].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[368].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[369].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[369].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[369].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[369].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[368].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[369].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[36].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[36].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[36].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[36].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[35].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[36].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[370].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[370].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[370].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[370].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[369].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[370].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[371].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[371].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[371].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[371].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[370].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[371].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[372].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[372].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[372].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[372].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[371].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[372].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[373].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[373].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[373].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[373].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[372].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[373].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[374].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[374].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[374].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[374].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[373].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[374].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[375].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[375].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[375].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[375].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[374].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[375].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[376].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[376].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[376].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[376].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[375].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[376].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[377].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[377].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[377].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[377].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[376].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[377].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[378].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[378].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[378].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[378].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[377].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[378].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[379].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[379].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[379].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[379].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[378].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[379].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[37].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[37].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[37].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[37].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[36].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[37].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[380].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[380].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[380].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[380].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[379].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[380].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[381].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[381].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[381].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[381].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[380].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[381].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[382].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[382].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[382].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[382].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[381].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[382].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[383].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[383].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[383].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[383].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[382].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[383].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[384].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[384].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[384].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[384].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[383].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[384].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[385].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[385].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[385].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[385].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[384].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[385].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[386].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[386].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[386].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[386].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[385].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[386].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[387].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[387].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[387].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[387].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[386].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[387].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[388].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[388].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[388].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[388].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[387].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[388].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[389].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[389].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[389].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[389].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[388].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[389].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[38].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[38].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[38].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[38].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[37].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[38].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[390].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[390].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[390].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[390].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[389].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[390].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[391].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[391].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[391].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[391].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[390].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[391].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[392].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[392].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[392].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[392].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[391].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[392].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[393].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[393].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[393].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[393].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[392].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[393].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[394].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[394].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[394].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[394].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[393].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[394].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[395].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[395].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[395].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[395].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[394].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[395].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[396].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[396].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[396].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[396].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[395].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[396].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[397].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[397].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[397].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[397].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[396].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[397].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[398].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[398].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[398].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[398].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[397].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[398].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[399].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[399].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[399].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[399].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[398].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[399].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[39].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[39].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[39].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[39].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[38].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[39].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[3].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[3].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[3].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[3].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[2].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[3].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[400].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[400].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[400].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[400].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[399].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[400].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[401].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[401].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[401].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[401].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[400].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[401].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[402].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[402].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[402].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[402].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[401].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[402].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[403].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[403].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[403].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[403].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[402].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[403].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[404].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[404].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[404].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[404].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[403].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[404].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[405].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[405].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[405].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[405].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[404].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[405].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[406].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[406].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[406].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[406].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[405].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[406].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[407].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[407].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[407].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[407].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[406].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[407].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[408].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[408].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[408].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[408].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[407].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[408].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[409].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[409].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[409].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[409].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[408].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[409].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[40].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[40].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[40].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[40].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[39].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[40].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[410].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[410].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[410].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[410].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[409].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[410].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[411].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[411].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[411].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[411].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[410].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[411].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[412].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[412].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[412].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[412].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[411].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[412].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[413].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[413].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[413].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[413].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[412].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[413].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[414].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[414].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[414].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[414].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[413].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[414].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[415].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[415].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[415].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[415].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[414].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[415].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[416].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[416].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[416].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[416].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[415].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[416].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[417].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[417].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[417].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[417].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[416].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[417].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[418].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[418].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[418].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[418].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[417].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[418].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[419].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[419].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[419].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[419].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[418].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[419].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[41].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[41].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[41].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[41].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[40].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[41].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[420].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[420].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[420].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[420].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[419].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[420].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[421].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[421].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[421].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[421].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[420].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[421].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[422].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[422].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[422].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[422].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[421].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[422].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[423].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[423].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[423].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[423].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[422].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[423].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[424].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[424].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[424].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[424].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[423].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[424].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[425].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[425].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[425].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[425].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[424].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[425].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[426].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[426].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[426].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[426].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[425].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[426].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[427].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[427].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[427].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[427].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[426].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[427].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[428].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[428].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[428].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[428].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[427].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[428].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[429].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[429].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[429].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[429].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[428].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[429].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[42].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[42].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[42].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[42].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[41].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[42].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[430].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[430].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[430].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[430].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[429].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[430].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[431].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[431].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[431].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[431].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[430].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[431].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[432].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[432].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[432].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[432].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[431].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[432].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[433].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[433].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[433].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[433].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[432].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[433].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[434].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[434].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[434].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[434].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[433].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[434].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[435].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[435].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[435].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[435].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[434].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[435].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[436].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[436].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[436].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[436].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[435].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[436].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[437].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[437].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[437].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[437].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[436].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[437].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[438].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[438].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[438].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[438].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[437].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[438].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[439].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[439].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[439].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[439].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[438].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[439].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[43].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[43].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[43].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[43].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[42].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[43].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[440].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[440].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[440].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[440].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[439].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[440].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[441].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[441].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[441].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[441].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[440].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[441].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[442].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[442].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[442].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[442].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[441].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[442].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[443].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[443].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[443].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[443].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[442].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[443].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[444].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[444].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[444].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[444].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[443].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[444].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[445].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[445].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[445].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[445].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[444].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[445].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[446].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[446].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[446].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[446].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[445].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[446].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[447].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[447].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[447].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[447].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[446].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[447].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[448].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[448].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[448].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[448].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[447].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[448].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[449].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[449].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[449].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[449].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[448].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[449].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[44].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[44].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[44].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[44].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[43].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[44].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[450].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[450].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[450].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[450].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[449].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[450].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[451].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[451].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[451].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[451].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[450].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[451].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[452].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[452].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[452].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[452].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[451].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[452].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[453].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[453].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[453].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[453].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[452].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[453].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[454].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[454].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[454].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[454].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[453].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[454].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[455].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[455].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[455].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[455].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[454].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[455].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[456].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[456].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[456].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[456].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[455].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[456].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[457].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[457].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[457].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[457].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[456].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[457].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[458].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[458].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[458].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[458].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[457].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[458].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[459].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[459].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[459].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[459].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[458].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[459].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[45].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[45].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[45].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[45].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[44].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[45].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[460].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[460].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[460].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[460].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[459].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[460].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[461].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[461].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[461].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[461].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[460].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[461].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[462].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[462].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[462].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[462].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[461].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[462].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[463].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[463].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[463].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[463].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[462].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[463].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[464].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[464].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[464].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[464].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[463].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[464].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[465].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[465].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[465].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[465].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[464].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[465].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[466].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[466].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[466].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[466].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[465].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[466].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[467].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[467].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[467].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[467].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[466].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[467].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[468].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[468].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[468].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[468].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[467].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[468].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[469].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[469].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[469].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[469].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[468].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[469].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[46].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[46].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[46].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[46].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[45].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[46].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[470].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[470].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[470].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[470].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[469].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[470].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[471].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[471].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[471].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[471].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[470].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[471].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[472].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[472].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[472].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[472].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[471].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[472].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[473].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[473].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[473].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[473].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[472].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[473].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[474].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[474].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[474].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[474].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[473].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[474].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[475].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[475].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[475].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[475].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[474].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[475].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[476].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[476].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[476].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[476].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[475].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[476].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[477].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[477].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[477].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[477].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[476].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[477].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[478].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[478].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[478].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[478].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[477].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[478].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[479].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[479].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[479].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[479].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[478].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[479].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[47].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[47].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[47].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[47].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[46].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[47].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[480].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[480].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[480].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[480].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[479].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[480].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[481].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[481].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[481].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[481].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[480].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[481].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[482].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[482].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[482].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[482].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[481].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[482].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[483].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[483].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[483].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[483].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[482].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[483].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[484].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[484].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[484].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[484].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[483].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[484].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[485].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[485].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[485].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[485].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[484].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[485].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[486].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[486].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[486].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[486].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[485].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[486].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[487].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[487].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[487].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[487].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[486].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[487].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[488].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[488].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[488].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[488].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[487].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[488].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[489].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[489].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[489].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[489].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[488].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[489].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[48].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[48].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[48].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[48].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[47].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[48].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[490].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[490].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[490].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[490].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[489].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[490].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[491].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[491].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[491].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[491].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[490].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[491].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[492].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[492].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[492].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[492].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[491].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[492].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[493].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[493].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[493].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[493].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[492].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[493].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[494].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[494].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[494].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[494].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[493].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[494].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[495].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[495].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[495].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[495].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[494].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[495].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[496].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[496].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[496].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[496].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[495].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[496].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[497].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[497].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[497].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[497].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[496].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[497].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[498].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[498].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[498].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[498].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[497].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[498].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[499].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[499].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[499].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[499].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[498].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[499].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[49].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[49].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[49].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[49].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[48].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[49].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[4].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[4].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[4].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[4].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[3].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[4].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[500].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[500].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[500].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[500].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[499].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[500].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[501].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[501].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[501].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[501].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[500].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[501].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[502].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[502].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[502].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[502].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[501].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[502].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[503].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[503].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[503].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[503].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[502].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[503].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[504].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[504].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[504].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[504].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[503].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[504].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[505].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[505].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[505].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[505].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[504].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[505].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[506].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[506].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[506].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[506].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[505].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[506].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[507].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[507].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[507].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[507].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[506].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[507].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[508].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[508].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[508].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[508].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[507].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[508].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[509].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[509].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[509].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[509].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[508].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[509].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[50].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[50].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[50].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[50].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[49].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[50].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[510].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[510].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[510].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[510].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[509].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[510].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[511].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[511].genblk1.genblk1.latch.nclk ),
    .A(shift));
 sg13g2_inv_1 \shift_reg[511].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[510].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[511].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[51].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[51].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[51].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[51].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[50].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[51].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[52].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[52].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[52].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[52].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[51].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[52].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[53].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[53].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[53].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[53].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[52].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[53].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[54].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[54].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[54].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[54].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[53].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[54].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[55].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[55].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[55].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[55].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[54].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[55].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[56].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[56].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[56].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[56].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[55].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[56].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[57].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[57].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[57].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[57].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[56].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[57].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[58].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[58].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[58].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[58].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[57].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[58].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[59].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[59].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[59].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[59].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[58].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[59].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[5].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[5].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[5].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[5].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[4].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[5].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[60].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[60].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[60].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[60].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[59].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[60].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[61].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[61].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[61].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[61].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[60].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[61].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[62].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[62].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[62].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[62].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[61].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[62].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[63].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[63].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[63].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[63].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[62].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[63].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[64].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[64].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[64].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[64].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[63].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[64].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[65].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[65].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[65].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[65].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[64].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[65].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[66].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[66].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[66].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[66].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[65].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[66].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[67].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[67].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[67].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[67].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[66].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[67].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[68].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[68].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[68].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[68].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[67].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[68].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[69].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[69].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[69].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[69].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[68].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[69].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[6].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[6].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[6].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[6].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[5].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[6].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[70].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[70].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[70].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[70].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[69].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[70].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[71].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[71].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[71].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[71].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[70].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[71].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[72].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[72].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[72].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[72].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[71].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[72].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[73].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[73].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[73].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[73].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[72].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[73].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[74].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[74].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[74].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[74].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[73].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[74].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[75].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[75].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[75].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[75].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[74].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[75].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[76].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[76].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[76].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[76].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[75].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[76].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[77].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[77].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[77].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[77].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[76].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[77].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[78].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[78].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[78].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[78].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[77].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[78].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[79].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[79].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[79].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[79].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[78].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[79].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[7].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[7].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[7].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[7].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[6].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[7].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[80].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[80].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[80].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[80].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[79].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[80].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[81].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[81].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[81].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[81].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[80].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[81].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[82].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[82].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[82].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[82].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[81].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[82].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[83].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[83].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[83].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[83].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[82].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[83].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[84].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[84].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[84].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[84].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[83].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[84].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[85].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[85].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[85].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[85].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[84].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[85].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[86].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[86].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[86].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[86].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[85].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[86].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[87].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[87].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[87].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[87].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[86].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[87].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[88].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[88].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[88].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[88].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[87].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[88].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[89].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[89].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[89].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[89].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[88].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[89].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[8].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[8].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[8].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[8].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[7].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[8].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[90].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[90].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[90].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[90].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[89].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[90].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[91].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[91].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[91].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[91].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[90].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[91].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[92].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[92].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[92].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[92].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[91].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[92].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[93].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[93].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[93].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[93].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[92].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[93].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[94].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[94].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[94].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[94].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[93].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[94].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[95].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[95].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[95].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[95].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[94].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[95].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[96].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[96].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[96].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[96].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[95].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[96].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[97].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[97].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[97].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[97].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[96].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[97].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[98].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[98].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[98].genblk1.genblk1.latch.clk ));
 sg13g2_inv_1 \shift_reg[98].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[97].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[98].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[99].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[99].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[100].genblk1.genblk1.latch.clkout ));
 sg13g2_inv_1 \shift_reg[99].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[98].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[99].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \shift_reg[9].genblk1.genblk1.latch.u_inv1.inv  (.Y(\shift_reg[9].genblk1.genblk1.latch.nclk ),
    .A(\shift_reg[10].genblk1.genblk1.latch.clkout ));
 sg13g2_inv_1 \shift_reg[9].genblk1.genblk1.latch.u_inv2.inv  (.Y(\shift_reg[8].genblk1.genblk1.latch.clk ),
    .A(\shift_reg[9].genblk1.genblk1.latch.nclk ));
 sg13g2_inv_1 \u_invA.inv  (.Y(ntrig),
    .A(net2));
 sg13g2_inv_1 \u_invB.inv  (.Y(trig_delayed),
    .A(ntrig));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_cattuto_sr_latch_3 (.L_LO(net3));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_38 ();
 sg13g2_fill_1 FILLER_0_46 ();
 sg13g2_fill_2 FILLER_0_64 ();
 sg13g2_decap_4 FILLER_0_72 ();
 sg13g2_fill_1 FILLER_0_79 ();
 sg13g2_decap_8 FILLER_0_83 ();
 sg13g2_decap_8 FILLER_0_90 ();
 sg13g2_fill_1 FILLER_0_114 ();
 sg13g2_decap_4 FILLER_0_130 ();
 sg13g2_fill_2 FILLER_0_137 ();
 sg13g2_fill_1 FILLER_0_162 ();
 sg13g2_fill_1 FILLER_0_169 ();
 sg13g2_fill_1 FILLER_0_199 ();
 sg13g2_decap_4 FILLER_0_203 ();
 sg13g2_fill_2 FILLER_0_210 ();
 sg13g2_fill_1 FILLER_0_212 ();
 sg13g2_decap_4 FILLER_0_216 ();
 sg13g2_fill_1 FILLER_0_223 ();
 sg13g2_fill_1 FILLER_0_227 ();
 sg13g2_fill_2 FILLER_0_248 ();
 sg13g2_decap_4 FILLER_0_267 ();
 sg13g2_fill_1 FILLER_0_294 ();
 sg13g2_fill_2 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_fill_1 FILLER_0_344 ();
 sg13g2_fill_2 FILLER_0_385 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_fill_1 FILLER_1_149 ();
 sg13g2_decap_4 FILLER_1_241 ();
 sg13g2_decap_4 FILLER_1_248 ();
 sg13g2_fill_1 FILLER_1_267 ();
 sg13g2_fill_2 FILLER_1_288 ();
 sg13g2_fill_1 FILLER_1_293 ();
 sg13g2_fill_2 FILLER_1_300 ();
 sg13g2_fill_1 FILLER_1_302 ();
 sg13g2_decap_4 FILLER_1_315 ();
 sg13g2_fill_1 FILLER_1_322 ();
 sg13g2_fill_2 FILLER_1_349 ();
 sg13g2_fill_2 FILLER_1_354 ();
 sg13g2_fill_1 FILLER_1_356 ();
 sg13g2_fill_1 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_4 FILLER_1_377 ();
 sg13g2_fill_1 FILLER_1_381 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_7 ();
 sg13g2_fill_1 FILLER_2_9 ();
 sg13g2_fill_1 FILLER_2_30 ();
 sg13g2_decap_8 FILLER_2_37 ();
 sg13g2_decap_8 FILLER_2_44 ();
 sg13g2_fill_2 FILLER_2_54 ();
 sg13g2_fill_1 FILLER_2_56 ();
 sg13g2_fill_2 FILLER_2_60 ();
 sg13g2_fill_1 FILLER_2_82 ();
 sg13g2_fill_1 FILLER_2_86 ();
 sg13g2_fill_1 FILLER_2_93 ();
 sg13g2_decap_4 FILLER_2_100 ();
 sg13g2_fill_2 FILLER_2_104 ();
 sg13g2_decap_4 FILLER_2_135 ();
 sg13g2_fill_1 FILLER_2_139 ();
 sg13g2_fill_1 FILLER_2_160 ();
 sg13g2_fill_1 FILLER_2_164 ();
 sg13g2_decap_4 FILLER_2_168 ();
 sg13g2_fill_2 FILLER_2_175 ();
 sg13g2_fill_1 FILLER_2_180 ();
 sg13g2_fill_2 FILLER_2_198 ();
 sg13g2_fill_1 FILLER_2_200 ();
 sg13g2_decap_4 FILLER_2_204 ();
 sg13g2_fill_2 FILLER_2_208 ();
 sg13g2_decap_8 FILLER_2_213 ();
 sg13g2_decap_8 FILLER_2_220 ();
 sg13g2_decap_4 FILLER_2_227 ();
 sg13g2_fill_1 FILLER_2_231 ();
 sg13g2_fill_1 FILLER_2_334 ();
 sg13g2_fill_1 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_11 ();
 sg13g2_fill_1 FILLER_3_36 ();
 sg13g2_decap_8 FILLER_3_108 ();
 sg13g2_fill_2 FILLER_3_132 ();
 sg13g2_fill_2 FILLER_3_185 ();
 sg13g2_fill_1 FILLER_3_227 ();
 sg13g2_decap_4 FILLER_3_231 ();
 sg13g2_fill_2 FILLER_3_235 ();
 sg13g2_fill_2 FILLER_3_240 ();
 sg13g2_decap_4 FILLER_3_245 ();
 sg13g2_fill_1 FILLER_3_249 ();
 sg13g2_fill_1 FILLER_3_253 ();
 sg13g2_fill_2 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_285 ();
 sg13g2_decap_8 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_299 ();
 sg13g2_fill_1 FILLER_3_306 ();
 sg13g2_fill_1 FILLER_3_330 ();
 sg13g2_fill_1 FILLER_3_334 ();
 sg13g2_fill_1 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_fill_1 FILLER_3_355 ();
 sg13g2_fill_2 FILLER_3_359 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_decap_4 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_57 ();
 sg13g2_decap_4 FILLER_4_64 ();
 sg13g2_fill_2 FILLER_4_68 ();
 sg13g2_decap_8 FILLER_4_73 ();
 sg13g2_decap_4 FILLER_4_80 ();
 sg13g2_fill_1 FILLER_4_84 ();
 sg13g2_decap_4 FILLER_4_88 ();
 sg13g2_fill_1 FILLER_4_92 ();
 sg13g2_fill_2 FILLER_4_96 ();
 sg13g2_fill_2 FILLER_4_101 ();
 sg13g2_fill_1 FILLER_4_103 ();
 sg13g2_decap_4 FILLER_4_121 ();
 sg13g2_decap_8 FILLER_4_131 ();
 sg13g2_decap_8 FILLER_4_138 ();
 sg13g2_fill_2 FILLER_4_145 ();
 sg13g2_decap_8 FILLER_4_162 ();
 sg13g2_decap_8 FILLER_4_169 ();
 sg13g2_decap_8 FILLER_4_176 ();
 sg13g2_fill_1 FILLER_4_183 ();
 sg13g2_decap_8 FILLER_4_187 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_fill_2 FILLER_4_214 ();
 sg13g2_fill_1 FILLER_4_216 ();
 sg13g2_fill_1 FILLER_4_271 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_11 ();
 sg13g2_fill_1 FILLER_5_29 ();
 sg13g2_fill_2 FILLER_5_47 ();
 sg13g2_decap_8 FILLER_5_58 ();
 sg13g2_decap_8 FILLER_5_65 ();
 sg13g2_fill_1 FILLER_5_72 ();
 sg13g2_fill_2 FILLER_5_107 ();
 sg13g2_fill_1 FILLER_5_163 ();
 sg13g2_fill_2 FILLER_5_167 ();
 sg13g2_fill_1 FILLER_5_169 ();
 sg13g2_decap_4 FILLER_5_173 ();
 sg13g2_fill_1 FILLER_5_180 ();
 sg13g2_fill_2 FILLER_5_184 ();
 sg13g2_fill_1 FILLER_5_186 ();
 sg13g2_decap_4 FILLER_5_210 ();
 sg13g2_fill_2 FILLER_5_217 ();
 sg13g2_fill_1 FILLER_5_219 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_8 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_decap_8 FILLER_5_251 ();
 sg13g2_decap_4 FILLER_5_258 ();
 sg13g2_fill_1 FILLER_5_262 ();
 sg13g2_fill_2 FILLER_5_266 ();
 sg13g2_decap_4 FILLER_5_271 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_282 ();
 sg13g2_decap_8 FILLER_5_289 ();
 sg13g2_fill_2 FILLER_5_299 ();
 sg13g2_fill_1 FILLER_5_301 ();
 sg13g2_fill_2 FILLER_5_308 ();
 sg13g2_fill_1 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_fill_1 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_decap_8 FILLER_5_332 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_decap_8 FILLER_5_353 ();
 sg13g2_fill_1 FILLER_5_360 ();
 sg13g2_decap_4 FILLER_5_364 ();
 sg13g2_fill_1 FILLER_5_368 ();
 sg13g2_decap_4 FILLER_5_378 ();
 sg13g2_fill_1 FILLER_5_382 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_27 ();
 sg13g2_decap_4 FILLER_6_34 ();
 sg13g2_fill_1 FILLER_6_38 ();
 sg13g2_fill_1 FILLER_6_82 ();
 sg13g2_decap_8 FILLER_6_92 ();
 sg13g2_decap_8 FILLER_6_99 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_4 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_4 FILLER_6_147 ();
 sg13g2_decap_4 FILLER_6_191 ();
 sg13g2_fill_1 FILLER_6_195 ();
 sg13g2_fill_2 FILLER_6_233 ();
 sg13g2_fill_2 FILLER_6_252 ();
 sg13g2_fill_1 FILLER_6_254 ();
 sg13g2_fill_1 FILLER_6_258 ();
 sg13g2_fill_2 FILLER_6_279 ();
 sg13g2_fill_2 FILLER_6_315 ();
 sg13g2_fill_1 FILLER_6_317 ();
 sg13g2_decap_4 FILLER_6_321 ();
 sg13g2_fill_2 FILLER_6_325 ();
 sg13g2_decap_4 FILLER_6_330 ();
 sg13g2_decap_4 FILLER_6_337 ();
 sg13g2_fill_1 FILLER_6_341 ();
 sg13g2_fill_2 FILLER_6_345 ();
 sg13g2_fill_1 FILLER_6_350 ();
 sg13g2_decap_4 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_30 ();
 sg13g2_decap_8 FILLER_7_37 ();
 sg13g2_fill_1 FILLER_7_44 ();
 sg13g2_fill_2 FILLER_7_51 ();
 sg13g2_fill_1 FILLER_7_56 ();
 sg13g2_fill_2 FILLER_7_94 ();
 sg13g2_decap_4 FILLER_7_99 ();
 sg13g2_fill_1 FILLER_7_103 ();
 sg13g2_fill_2 FILLER_7_107 ();
 sg13g2_decap_4 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_116 ();
 sg13g2_decap_4 FILLER_7_121 ();
 sg13g2_fill_1 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_decap_8 FILLER_7_153 ();
 sg13g2_decap_8 FILLER_7_160 ();
 sg13g2_decap_8 FILLER_7_167 ();
 sg13g2_decap_4 FILLER_7_174 ();
 sg13g2_fill_2 FILLER_7_178 ();
 sg13g2_fill_2 FILLER_7_183 ();
 sg13g2_fill_1 FILLER_7_185 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_194 ();
 sg13g2_decap_4 FILLER_7_201 ();
 sg13g2_fill_1 FILLER_7_225 ();
 sg13g2_fill_2 FILLER_7_229 ();
 sg13g2_fill_2 FILLER_7_254 ();
 sg13g2_fill_2 FILLER_7_279 ();
 sg13g2_fill_2 FILLER_7_284 ();
 sg13g2_fill_1 FILLER_7_286 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_4 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_fill_2 FILLER_7_395 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_18 ();
 sg13g2_fill_1 FILLER_8_25 ();
 sg13g2_fill_1 FILLER_8_29 ();
 sg13g2_decap_4 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_4 FILLER_8_135 ();
 sg13g2_fill_1 FILLER_8_139 ();
 sg13g2_fill_1 FILLER_8_163 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_decap_8 FILLER_8_205 ();
 sg13g2_fill_2 FILLER_8_212 ();
 sg13g2_fill_1 FILLER_8_234 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_fill_2 FILLER_8_278 ();
 sg13g2_decap_8 FILLER_8_283 ();
 sg13g2_fill_2 FILLER_8_293 ();
 sg13g2_decap_4 FILLER_8_298 ();
 sg13g2_fill_1 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_fill_2 FILLER_8_333 ();
 sg13g2_fill_1 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_fill_2 FILLER_8_366 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_41 ();
 sg13g2_fill_2 FILLER_9_48 ();
 sg13g2_fill_1 FILLER_9_50 ();
 sg13g2_fill_2 FILLER_9_57 ();
 sg13g2_fill_2 FILLER_9_82 ();
 sg13g2_fill_1 FILLER_9_84 ();
 sg13g2_fill_2 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_107 ();
 sg13g2_decap_4 FILLER_9_111 ();
 sg13g2_fill_1 FILLER_9_115 ();
 sg13g2_fill_2 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_decap_4 FILLER_9_125 ();
 sg13g2_fill_1 FILLER_9_129 ();
 sg13g2_fill_2 FILLER_9_133 ();
 sg13g2_fill_1 FILLER_9_135 ();
 sg13g2_fill_2 FILLER_9_139 ();
 sg13g2_fill_1 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_decap_4 FILLER_9_216 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_decap_4 FILLER_9_230 ();
 sg13g2_decap_4 FILLER_9_237 ();
 sg13g2_decap_8 FILLER_9_244 ();
 sg13g2_decap_8 FILLER_9_251 ();
 sg13g2_decap_4 FILLER_9_312 ();
 sg13g2_fill_1 FILLER_9_316 ();
 sg13g2_fill_2 FILLER_9_385 ();
 sg13g2_fill_1 FILLER_9_390 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_9 ();
 sg13g2_fill_1 FILLER_10_27 ();
 sg13g2_decap_8 FILLER_10_34 ();
 sg13g2_fill_2 FILLER_10_41 ();
 sg13g2_fill_1 FILLER_10_43 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_77 ();
 sg13g2_fill_2 FILLER_10_81 ();
 sg13g2_fill_1 FILLER_10_86 ();
 sg13g2_fill_1 FILLER_10_144 ();
 sg13g2_decap_4 FILLER_10_148 ();
 sg13g2_fill_2 FILLER_10_172 ();
 sg13g2_decap_4 FILLER_10_177 ();
 sg13g2_decap_4 FILLER_10_187 ();
 sg13g2_fill_1 FILLER_10_191 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_fill_1 FILLER_10_242 ();
 sg13g2_fill_2 FILLER_10_246 ();
 sg13g2_fill_1 FILLER_10_251 ();
 sg13g2_fill_2 FILLER_10_269 ();
 sg13g2_fill_1 FILLER_10_271 ();
 sg13g2_decap_4 FILLER_10_275 ();
 sg13g2_decap_4 FILLER_10_282 ();
 sg13g2_decap_4 FILLER_10_289 ();
 sg13g2_fill_1 FILLER_10_293 ();
 sg13g2_fill_2 FILLER_10_297 ();
 sg13g2_decap_4 FILLER_10_302 ();
 sg13g2_fill_1 FILLER_10_323 ();
 sg13g2_decap_4 FILLER_10_327 ();
 sg13g2_fill_2 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_fill_1 FILLER_10_379 ();
 sg13g2_fill_1 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_18 ();
 sg13g2_decap_4 FILLER_11_31 ();
 sg13g2_fill_1 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_59 ();
 sg13g2_fill_2 FILLER_11_94 ();
 sg13g2_fill_1 FILLER_11_99 ();
 sg13g2_decap_4 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_110 ();
 sg13g2_fill_2 FILLER_11_114 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_fill_2 FILLER_11_150 ();
 sg13g2_decap_4 FILLER_11_155 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_220 ();
 sg13g2_fill_1 FILLER_11_227 ();
 sg13g2_fill_1 FILLER_11_268 ();
 sg13g2_fill_2 FILLER_11_272 ();
 sg13g2_fill_2 FILLER_11_277 ();
 sg13g2_decap_4 FILLER_11_356 ();
 sg13g2_fill_1 FILLER_11_363 ();
 sg13g2_decap_4 FILLER_11_367 ();
 sg13g2_fill_1 FILLER_11_371 ();
 sg13g2_decap_4 FILLER_11_375 ();
 sg13g2_fill_1 FILLER_11_379 ();
 sg13g2_decap_4 FILLER_11_383 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_11 ();
 sg13g2_fill_2 FILLER_12_30 ();
 sg13g2_fill_1 FILLER_12_49 ();
 sg13g2_fill_2 FILLER_12_67 ();
 sg13g2_fill_1 FILLER_12_69 ();
 sg13g2_decap_8 FILLER_12_73 ();
 sg13g2_fill_2 FILLER_12_83 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_fill_2 FILLER_12_186 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_192 ();
 sg13g2_fill_2 FILLER_12_199 ();
 sg13g2_fill_2 FILLER_12_204 ();
 sg13g2_fill_1 FILLER_12_206 ();
 sg13g2_decap_4 FILLER_12_210 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_decap_4 FILLER_12_218 ();
 sg13g2_decap_8 FILLER_12_239 ();
 sg13g2_fill_1 FILLER_12_246 ();
 sg13g2_fill_2 FILLER_12_250 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_fill_2 FILLER_12_316 ();
 sg13g2_decap_4 FILLER_12_321 ();
 sg13g2_fill_2 FILLER_12_328 ();
 sg13g2_fill_1 FILLER_12_330 ();
 sg13g2_decap_4 FILLER_12_334 ();
 sg13g2_fill_2 FILLER_12_338 ();
 sg13g2_fill_2 FILLER_12_383 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_18 ();
 sg13g2_fill_2 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_36 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_fill_2 FILLER_13_116 ();
 sg13g2_fill_1 FILLER_13_118 ();
 sg13g2_fill_2 FILLER_13_139 ();
 sg13g2_decap_4 FILLER_13_144 ();
 sg13g2_fill_2 FILLER_13_148 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_157 ();
 sg13g2_decap_8 FILLER_13_261 ();
 sg13g2_fill_1 FILLER_13_268 ();
 sg13g2_decap_8 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_302 ();
 sg13g2_fill_2 FILLER_13_346 ();
 sg13g2_fill_1 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_41 ();
 sg13g2_decap_8 FILLER_14_48 ();
 sg13g2_decap_4 FILLER_14_58 ();
 sg13g2_fill_1 FILLER_14_65 ();
 sg13g2_decap_4 FILLER_14_69 ();
 sg13g2_fill_1 FILLER_14_90 ();
 sg13g2_decap_4 FILLER_14_100 ();
 sg13g2_fill_2 FILLER_14_104 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_167 ();
 sg13g2_decap_4 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_fill_1 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_4 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_231 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_240 ();
 sg13g2_fill_2 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_4 FILLER_14_276 ();
 sg13g2_fill_2 FILLER_14_280 ();
 sg13g2_decap_4 FILLER_14_308 ();
 sg13g2_fill_2 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_fill_2 FILLER_14_324 ();
 sg13g2_fill_1 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_4 FILLER_14_368 ();
 sg13g2_fill_2 FILLER_14_372 ();
 sg13g2_fill_1 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_31 ();
 sg13g2_fill_2 FILLER_15_36 ();
 sg13g2_fill_1 FILLER_15_38 ();
 sg13g2_decap_4 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_46 ();
 sg13g2_decap_4 FILLER_15_51 ();
 sg13g2_fill_1 FILLER_15_55 ();
 sg13g2_fill_1 FILLER_15_73 ();
 sg13g2_decap_4 FILLER_15_77 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_fill_2 FILLER_15_116 ();
 sg13g2_fill_1 FILLER_15_118 ();
 sg13g2_fill_1 FILLER_15_122 ();
 sg13g2_decap_8 FILLER_15_129 ();
 sg13g2_decap_8 FILLER_15_136 ();
 sg13g2_decap_8 FILLER_15_143 ();
 sg13g2_fill_2 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_2 FILLER_15_170 ();
 sg13g2_fill_1 FILLER_15_178 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_decap_4 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_190 ();
 sg13g2_fill_2 FILLER_15_218 ();
 sg13g2_fill_1 FILLER_15_220 ();
 sg13g2_decap_8 FILLER_15_258 ();
 sg13g2_decap_4 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_309 ();
 sg13g2_fill_2 FILLER_15_313 ();
 sg13g2_fill_1 FILLER_15_318 ();
 sg13g2_fill_2 FILLER_15_356 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_64 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_decap_4 FILLER_16_83 ();
 sg13g2_decap_4 FILLER_16_90 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_113 ();
 sg13g2_fill_1 FILLER_16_115 ();
 sg13g2_decap_4 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_123 ();
 sg13g2_fill_1 FILLER_16_134 ();
 sg13g2_fill_1 FILLER_16_138 ();
 sg13g2_decap_8 FILLER_16_145 ();
 sg13g2_decap_4 FILLER_16_152 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_fill_2 FILLER_16_200 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_4 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_234 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_fill_2 FILLER_16_245 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_4 FILLER_16_337 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_345 ();
 sg13g2_decap_4 FILLER_16_350 ();
 sg13g2_fill_1 FILLER_16_354 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_384 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_16 ();
 sg13g2_fill_2 FILLER_17_20 ();
 sg13g2_fill_1 FILLER_17_42 ();
 sg13g2_decap_4 FILLER_17_46 ();
 sg13g2_fill_1 FILLER_17_50 ();
 sg13g2_fill_2 FILLER_17_54 ();
 sg13g2_fill_1 FILLER_17_79 ();
 sg13g2_decap_4 FILLER_17_83 ();
 sg13g2_fill_1 FILLER_17_87 ();
 sg13g2_fill_1 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_97 ();
 sg13g2_fill_2 FILLER_17_152 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_172 ();
 sg13g2_fill_2 FILLER_17_179 ();
 sg13g2_fill_2 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_fill_2 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_246 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_decap_4 FILLER_17_300 ();
 sg13g2_fill_2 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_315 ();
 sg13g2_decap_4 FILLER_17_319 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_decap_4 FILLER_17_381 ();
 sg13g2_fill_1 FILLER_17_385 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_fill_2 FILLER_18_22 ();
 sg13g2_fill_2 FILLER_18_64 ();
 sg13g2_decap_8 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_114 ();
 sg13g2_decap_8 FILLER_18_121 ();
 sg13g2_decap_4 FILLER_18_128 ();
 sg13g2_fill_2 FILLER_18_132 ();
 sg13g2_fill_1 FILLER_18_137 ();
 sg13g2_fill_1 FILLER_18_155 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_decap_8 FILLER_18_191 ();
 sg13g2_decap_4 FILLER_18_201 ();
 sg13g2_fill_2 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_247 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_decap_8 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_4 FILLER_18_334 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_fill_2 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_395 ();
 sg13g2_fill_1 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_fill_2 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_51 ();
 sg13g2_fill_2 FILLER_19_58 ();
 sg13g2_fill_1 FILLER_19_66 ();
 sg13g2_decap_4 FILLER_19_73 ();
 sg13g2_fill_2 FILLER_19_80 ();
 sg13g2_fill_1 FILLER_19_82 ();
 sg13g2_decap_4 FILLER_19_86 ();
 sg13g2_fill_2 FILLER_19_90 ();
 sg13g2_fill_2 FILLER_19_95 ();
 sg13g2_fill_1 FILLER_19_97 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_153 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_171 ();
 sg13g2_decap_8 FILLER_19_178 ();
 sg13g2_fill_1 FILLER_19_185 ();
 sg13g2_fill_1 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_224 ();
 sg13g2_fill_2 FILLER_19_228 ();
 sg13g2_decap_4 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_237 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_4 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_fill_2 FILLER_19_396 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_37 ();
 sg13g2_fill_1 FILLER_20_41 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_fill_2 FILLER_20_130 ();
 sg13g2_fill_1 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_206 ();
 sg13g2_decap_4 FILLER_20_258 ();
 sg13g2_fill_2 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_decap_8 FILLER_20_288 ();
 sg13g2_decap_4 FILLER_20_295 ();
 sg13g2_fill_2 FILLER_20_299 ();
 sg13g2_decap_4 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_312 ();
 sg13g2_decap_4 FILLER_20_336 ();
 sg13g2_decap_4 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_347 ();
 sg13g2_fill_2 FILLER_20_351 ();
 sg13g2_fill_1 FILLER_20_353 ();
 sg13g2_decap_4 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_361 ();
 sg13g2_fill_2 FILLER_20_365 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_fill_2 FILLER_20_385 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_52 ();
 sg13g2_decap_4 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_64 ();
 sg13g2_decap_8 FILLER_21_71 ();
 sg13g2_decap_8 FILLER_21_78 ();
 sg13g2_fill_2 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_fill_2 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_136 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_183 ();
 sg13g2_fill_1 FILLER_21_185 ();
 sg13g2_decap_4 FILLER_21_192 ();
 sg13g2_fill_2 FILLER_21_196 ();
 sg13g2_decap_4 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_229 ();
 sg13g2_decap_4 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_240 ();
 sg13g2_fill_2 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_308 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_18 ();
 sg13g2_fill_2 FILLER_22_32 ();
 sg13g2_fill_2 FILLER_22_40 ();
 sg13g2_decap_8 FILLER_22_45 ();
 sg13g2_decap_8 FILLER_22_52 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_decap_4 FILLER_22_80 ();
 sg13g2_decap_8 FILLER_22_101 ();
 sg13g2_fill_2 FILLER_22_108 ();
 sg13g2_fill_1 FILLER_22_110 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_149 ();
 sg13g2_fill_1 FILLER_22_151 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_206 ();
 sg13g2_decap_4 FILLER_22_213 ();
 sg13g2_decap_8 FILLER_22_237 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_fill_2 FILLER_22_251 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_decap_4 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_271 ();
 sg13g2_decap_8 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_1 FILLER_22_308 ();
 sg13g2_decap_4 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_4 FILLER_22_343 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_fill_1 FILLER_22_352 ();
 sg13g2_decap_4 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_360 ();
 sg13g2_fill_2 FILLER_22_364 ();
 sg13g2_decap_4 FILLER_22_369 ();
 sg13g2_fill_1 FILLER_22_373 ();
 sg13g2_fill_2 FILLER_22_377 ();
 sg13g2_decap_4 FILLER_22_382 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_1 FILLER_23_80 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_2 FILLER_23_107 ();
 sg13g2_fill_2 FILLER_23_129 ();
 sg13g2_decap_4 FILLER_23_134 ();
 sg13g2_fill_2 FILLER_23_141 ();
 sg13g2_fill_2 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_168 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_2 FILLER_23_294 ();
 sg13g2_fill_2 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_23 ();
 sg13g2_decap_8 FILLER_24_30 ();
 sg13g2_fill_2 FILLER_24_37 ();
 sg13g2_fill_1 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_fill_2 FILLER_24_53 ();
 sg13g2_decap_4 FILLER_24_78 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_decap_8 FILLER_24_86 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_4 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_151 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_decap_4 FILLER_24_176 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_fill_1 FILLER_24_187 ();
 sg13g2_decap_4 FILLER_24_211 ();
 sg13g2_decap_4 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_222 ();
 sg13g2_decap_4 FILLER_24_226 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_fill_2 FILLER_24_234 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_266 ();
 sg13g2_fill_2 FILLER_24_270 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_276 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_4 FILLER_24_370 ();
 sg13g2_fill_1 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_48 ();
 sg13g2_fill_1 FILLER_25_50 ();
 sg13g2_decap_4 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_decap_8 FILLER_25_123 ();
 sg13g2_decap_4 FILLER_25_130 ();
 sg13g2_fill_1 FILLER_25_134 ();
 sg13g2_decap_4 FILLER_25_138 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_decap_4 FILLER_25_146 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_192 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_decap_4 FILLER_25_201 ();
 sg13g2_fill_2 FILLER_25_205 ();
 sg13g2_decap_4 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_214 ();
 sg13g2_fill_2 FILLER_25_250 ();
 sg13g2_decap_4 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_decap_4 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_fill_2 FILLER_25_344 ();
 sg13g2_fill_1 FILLER_25_346 ();
 sg13g2_fill_1 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_4 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_18 ();
 sg13g2_decap_8 FILLER_26_31 ();
 sg13g2_decap_4 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_59 ();
 sg13g2_decap_4 FILLER_26_66 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_78 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_decap_4 FILLER_26_89 ();
 sg13g2_fill_2 FILLER_26_93 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_decap_4 FILLER_26_103 ();
 sg13g2_decap_8 FILLER_26_113 ();
 sg13g2_fill_1 FILLER_26_120 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_fill_2 FILLER_26_193 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_4 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_decap_4 FILLER_26_251 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_decap_4 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_4 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_decap_4 FILLER_26_344 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_fill_1 FILLER_26_387 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_55 ();
 sg13g2_decap_8 FILLER_27_62 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_decap_4 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_decap_4 FILLER_27_145 ();
 sg13g2_decap_4 FILLER_27_152 ();
 sg13g2_fill_2 FILLER_27_156 ();
 sg13g2_fill_2 FILLER_27_161 ();
 sg13g2_decap_4 FILLER_27_166 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_decap_4 FILLER_27_229 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_decap_4 FILLER_27_277 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_27_354 ();
 sg13g2_decap_4 FILLER_27_358 ();
 sg13g2_fill_2 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_387 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_27 ();
 sg13g2_fill_2 FILLER_28_31 ();
 sg13g2_fill_2 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_97 ();
 sg13g2_decap_4 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_106 ();
 sg13g2_fill_2 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_199 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_decap_4 FILLER_28_335 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_9 ();
 sg13g2_decap_4 FILLER_29_30 ();
 sg13g2_fill_2 FILLER_29_34 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_60 ();
 sg13g2_fill_1 FILLER_29_62 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_156 ();
 sg13g2_fill_2 FILLER_29_174 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_fill_1 FILLER_29_186 ();
 sg13g2_decap_4 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_194 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_decap_4 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_230 ();
 sg13g2_decap_4 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_269 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_decap_4 FILLER_29_275 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_decap_4 FILLER_29_319 ();
 sg13g2_decap_4 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_334 ();
 sg13g2_decap_4 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_decap_4 FILLER_29_347 ();
 sg13g2_decap_4 FILLER_29_391 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_24 ();
 sg13g2_decap_4 FILLER_30_31 ();
 sg13g2_fill_2 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_decap_4 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_85 ();
 sg13g2_decap_8 FILLER_30_106 ();
 sg13g2_fill_2 FILLER_30_113 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_decap_4 FILLER_30_394 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_46 ();
 sg13g2_fill_2 FILLER_31_50 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_fill_2 FILLER_31_76 ();
 sg13g2_decap_4 FILLER_31_87 ();
 sg13g2_decap_4 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_fill_2 FILLER_31_150 ();
 sg13g2_decap_4 FILLER_31_155 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_decap_8 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_fill_2 FILLER_31_176 ();
 sg13g2_decap_4 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_228 ();
 sg13g2_decap_8 FILLER_31_233 ();
 sg13g2_decap_8 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_247 ();
 sg13g2_decap_4 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_261 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_decap_4 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_4 FILLER_31_329 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_fill_2 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_340 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_fill_1 FILLER_31_348 ();
 sg13g2_decap_8 FILLER_31_366 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_4 FILLER_31_380 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_24 ();
 sg13g2_fill_2 FILLER_32_31 ();
 sg13g2_fill_1 FILLER_32_33 ();
 sg13g2_decap_8 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_64 ();
 sg13g2_decap_8 FILLER_32_82 ();
 sg13g2_fill_2 FILLER_32_89 ();
 sg13g2_decap_4 FILLER_32_94 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_decap_4 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_4 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_4 FILLER_32_259 ();
 sg13g2_decap_4 FILLER_32_320 ();
 sg13g2_fill_1 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_62 ();
 sg13g2_fill_2 FILLER_33_66 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_decap_4 FILLER_33_92 ();
 sg13g2_fill_1 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_134 ();
 sg13g2_fill_2 FILLER_33_138 ();
 sg13g2_fill_1 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_144 ();
 sg13g2_fill_1 FILLER_33_146 ();
 sg13g2_decap_8 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_159 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_decap_8 FILLER_33_205 ();
 sg13g2_decap_4 FILLER_33_212 ();
 sg13g2_decap_8 FILLER_33_219 ();
 sg13g2_decap_8 FILLER_33_226 ();
 sg13g2_decap_4 FILLER_33_276 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_313 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_decap_8 FILLER_33_345 ();
 sg13g2_decap_8 FILLER_33_352 ();
 sg13g2_decap_4 FILLER_33_379 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_18 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_fill_2 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_71 ();
 sg13g2_decap_8 FILLER_34_129 ();
 sg13g2_decap_4 FILLER_34_142 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_decap_4 FILLER_34_156 ();
 sg13g2_decap_4 FILLER_34_200 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_213 ();
 sg13g2_decap_4 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_226 ();
 sg13g2_decap_4 FILLER_34_230 ();
 sg13g2_decap_4 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_341 ();
 sg13g2_decap_8 FILLER_34_348 ();
 sg13g2_decap_4 FILLER_34_355 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_decap_4 FILLER_34_383 ();
 sg13g2_fill_1 FILLER_34_387 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_32 ();
 sg13g2_fill_1 FILLER_35_51 ();
 sg13g2_fill_1 FILLER_35_55 ();
 sg13g2_decap_8 FILLER_35_82 ();
 sg13g2_decap_8 FILLER_35_89 ();
 sg13g2_decap_4 FILLER_35_96 ();
 sg13g2_decap_4 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_110 ();
 sg13g2_decap_8 FILLER_35_169 ();
 sg13g2_decap_4 FILLER_35_176 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_fill_2 FILLER_35_185 ();
 sg13g2_fill_1 FILLER_35_187 ();
 sg13g2_fill_1 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_11 ();
 sg13g2_decap_8 FILLER_36_33 ();
 sg13g2_fill_2 FILLER_36_40 ();
 sg13g2_fill_1 FILLER_36_45 ();
 sg13g2_fill_2 FILLER_36_49 ();
 sg13g2_fill_1 FILLER_36_51 ();
 sg13g2_fill_1 FILLER_36_55 ();
 sg13g2_fill_2 FILLER_36_62 ();
 sg13g2_fill_1 FILLER_36_64 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_127 ();
 sg13g2_fill_2 FILLER_36_131 ();
 sg13g2_fill_1 FILLER_36_133 ();
 sg13g2_decap_4 FILLER_36_143 ();
 sg13g2_fill_2 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_decap_8 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_fill_2 FILLER_36_208 ();
 sg13g2_decap_4 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_221 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_decap_4 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_251 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_fill_2 FILLER_36_283 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_decap_4 FILLER_36_292 ();
 sg13g2_fill_1 FILLER_36_296 ();
 sg13g2_fill_2 FILLER_36_300 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_fill_2 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_36_386 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_decap_8 FILLER_37_79 ();
 sg13g2_decap_8 FILLER_37_86 ();
 sg13g2_decap_8 FILLER_37_184 ();
 sg13g2_decap_8 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_267 ();
 sg13g2_fill_1 FILLER_37_336 ();
 sg13g2_fill_2 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_365 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_30 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_decap_8 FILLER_38_36 ();
 sg13g2_decap_8 FILLER_38_43 ();
 sg13g2_decap_4 FILLER_38_50 ();
 sg13g2_fill_2 FILLER_38_54 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_71 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_decap_4 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_fill_2 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_238 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_247 ();
 sg13g2_decap_4 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_fill_2 FILLER_38_263 ();
 sg13g2_decap_4 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_272 ();
 sg13g2_decap_8 FILLER_38_276 ();
 sg13g2_decap_8 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_decap_8 FILLER_38_297 ();
 sg13g2_decap_4 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_308 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_fill_2 FILLER_38_324 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
 assign uo_out[1] = net19;
 assign uo_out[2] = net20;
 assign uo_out[3] = net21;
 assign uo_out[4] = net22;
 assign uo_out[5] = net23;
 assign uo_out[6] = net24;
 assign uo_out[7] = net25;
endmodule

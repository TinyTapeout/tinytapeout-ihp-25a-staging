module tt_um_rebeccargb_tt09ball_screensaver (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire clknet_0_clk;
 wire \color_index[0] ;
 wire \color_index[1] ;
 wire \color_index[2] ;
 wire dir_x;
 wire dir_y;
 wire hsync;
 wire \logo_left[0] ;
 wire \logo_left[1] ;
 wire \logo_left[2] ;
 wire \logo_left[3] ;
 wire \logo_left[4] ;
 wire \logo_left[5] ;
 wire \logo_left[6] ;
 wire \logo_left[7] ;
 wire \logo_left[8] ;
 wire \logo_left[9] ;
 wire \logo_top[0] ;
 wire \logo_top[1] ;
 wire \logo_top[2] ;
 wire \logo_top[3] ;
 wire \logo_top[4] ;
 wire \logo_top[5] ;
 wire \logo_top[6] ;
 wire \logo_top[7] ;
 wire \logo_top[8] ;
 wire \logo_top[9] ;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire \prev_y[0] ;
 wire \prev_y[1] ;
 wire \prev_y[2] ;
 wire \prev_y[3] ;
 wire \prev_y[4] ;
 wire \prev_y[5] ;
 wire \prev_y[6] ;
 wire \prev_y[7] ;
 wire \prev_y[8] ;
 wire \prev_y[9] ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire \vga_sync_gen.vsync ;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;

 sg13g2_inv_1 _1192_ (.Y(_0264_),
    .A(net95));
 sg13g2_inv_1 _1193_ (.Y(_0265_),
    .A(net87));
 sg13g2_inv_2 _1194_ (.Y(_0266_),
    .A(net625));
 sg13g2_inv_2 _1195_ (.Y(_0267_),
    .A(net627));
 sg13g2_inv_1 _1196_ (.Y(_0268_),
    .A(\logo_top[5] ));
 sg13g2_inv_1 _1197_ (.Y(_0269_),
    .A(\logo_top[4] ));
 sg13g2_inv_1 _1198_ (.Y(_0270_),
    .A(net165));
 sg13g2_inv_1 _1199_ (.Y(_0271_),
    .A(net91));
 sg13g2_inv_1 _1200_ (.Y(_0272_),
    .A(\logo_left[7] ));
 sg13g2_inv_1 _1201_ (.Y(_0273_),
    .A(\logo_left[5] ));
 sg13g2_inv_1 _1202_ (.Y(_0274_),
    .A(\logo_left[4] ));
 sg13g2_inv_1 _1203_ (.Y(_0275_),
    .A(net631));
 sg13g2_inv_1 _1204_ (.Y(_0276_),
    .A(net89));
 sg13g2_inv_1 _1205_ (.Y(_0277_),
    .A(\pix_y[1] ));
 sg13g2_inv_1 _1206_ (.Y(_0278_),
    .A(\pix_y[0] ));
 sg13g2_inv_1 _1207_ (.Y(_0279_),
    .A(net622));
 sg13g2_inv_2 _1208_ (.Y(_0280_),
    .A(net175));
 sg13g2_inv_1 _1209_ (.Y(_0281_),
    .A(net621));
 sg13g2_inv_2 _1210_ (.Y(_0282_),
    .A(net633));
 sg13g2_inv_2 _1211_ (.Y(_0283_),
    .A(net146));
 sg13g2_inv_2 _1212_ (.Y(_0284_),
    .A(net168));
 sg13g2_inv_1 _1213_ (.Y(_0285_),
    .A(\prev_y[0] ));
 sg13g2_inv_1 _1214_ (.Y(_0286_),
    .A(net97));
 sg13g2_inv_1 _1215_ (.Y(_0287_),
    .A(\prev_y[4] ));
 sg13g2_inv_1 _1216_ (.Y(_0288_),
    .A(\prev_y[6] ));
 sg13g2_inv_1 _1217_ (.Y(_0289_),
    .A(\prev_y[8] ));
 sg13g2_inv_1 _1218_ (.Y(_0290_),
    .A(net81));
 sg13g2_nand3_1 _1219_ (.B(\pix_y[6] ),
    .C(\pix_y[7] ),
    .A(\pix_y[5] ),
    .Y(_0291_));
 sg13g2_nor2_1 _1220_ (.A(_0283_),
    .B(net151),
    .Y(_0292_));
 sg13g2_nand3_1 _1221_ (.B(\pix_y[3] ),
    .C(_0292_),
    .A(\pix_y[1] ),
    .Y(_0293_));
 sg13g2_nor4_2 _1222_ (.A(net624),
    .B(net85),
    .C(_0291_),
    .Y(_0001_),
    .D(_0293_));
 sg13g2_and2_1 _1223_ (.A(net173),
    .B(\pix_x[5] ),
    .X(_0294_));
 sg13g2_and2_1 _1224_ (.A(net132),
    .B(_0294_),
    .X(_0295_));
 sg13g2_nor3_1 _1225_ (.A(\pix_x[4] ),
    .B(\pix_x[5] ),
    .C(net132),
    .Y(_0296_));
 sg13g2_nand2_1 _1226_ (.Y(_0297_),
    .A(\pix_x[7] ),
    .B(net133));
 sg13g2_nor4_2 _1227_ (.A(\pix_x[8] ),
    .B(_0295_),
    .C(_0296_),
    .Y(_0000_),
    .D(net134));
 sg13g2_and3_1 _1228_ (.X(_0298_),
    .A(net127),
    .B(net129),
    .C(\pix_x[1] ));
 sg13g2_and2_2 _1229_ (.A(net139),
    .B(_0298_),
    .X(_0299_));
 sg13g2_nand2_2 _1230_ (.Y(_0300_),
    .A(net166),
    .B(_0299_));
 sg13g2_nand3b_1 _1231_ (.B(\pix_x[8] ),
    .C(net133),
    .Y(_0301_),
    .A_N(\pix_x[7] ));
 sg13g2_nor4_2 _1232_ (.A(\pix_x[5] ),
    .B(net132),
    .C(_0300_),
    .Y(_0302_),
    .D(_0301_));
 sg13g2_nand2b_2 _1233_ (.Y(_0303_),
    .B(net637),
    .A_N(_0302_));
 sg13g2_nor2_1 _1234_ (.A(_0290_),
    .B(_0303_),
    .Y(_0016_));
 sg13g2_xnor2_1 _1235_ (.Y(_0304_),
    .A(net127),
    .B(\pix_x[1] ));
 sg13g2_nor2_1 _1236_ (.A(_0303_),
    .B(net128),
    .Y(_0017_));
 sg13g2_a21oi_1 _1237_ (.A1(net127),
    .A2(\pix_x[1] ),
    .Y(_0305_),
    .B1(net129));
 sg13g2_nor3_1 _1238_ (.A(_0282_),
    .B(_0298_),
    .C(net130),
    .Y(_0018_));
 sg13g2_o21ai_1 _1239_ (.B1(net638),
    .Y(_0306_),
    .A1(net139),
    .A2(_0298_));
 sg13g2_nor2_1 _1240_ (.A(_0299_),
    .B(net140),
    .Y(_0019_));
 sg13g2_o21ai_1 _1241_ (.B1(net638),
    .Y(_0307_),
    .A1(net166),
    .A2(_0299_));
 sg13g2_nor2b_1 _1242_ (.A(_0307_),
    .B_N(_0300_),
    .Y(_0020_));
 sg13g2_xor2_1 _1243_ (.B(_0300_),
    .A(net156),
    .X(_0308_));
 sg13g2_nor2_1 _1244_ (.A(_0303_),
    .B(net157),
    .Y(_0021_));
 sg13g2_a21oi_1 _1245_ (.A1(net174),
    .A2(_0299_),
    .Y(_0309_),
    .B1(net132));
 sg13g2_and2_1 _1246_ (.A(_0295_),
    .B(_0299_),
    .X(_0310_));
 sg13g2_nor3_1 _1247_ (.A(net546),
    .B(_0309_),
    .C(_0310_),
    .Y(_0022_));
 sg13g2_xnor2_1 _1248_ (.Y(_0311_),
    .A(net144),
    .B(_0310_));
 sg13g2_nor2_1 _1249_ (.A(net546),
    .B(_0311_),
    .Y(_0023_));
 sg13g2_a21oi_1 _1250_ (.A1(\pix_x[7] ),
    .A2(_0310_),
    .Y(_0312_),
    .B1(net141));
 sg13g2_and3_1 _1251_ (.X(_0313_),
    .A(net145),
    .B(net141),
    .C(_0310_));
 sg13g2_nor3_1 _1252_ (.A(net546),
    .B(net142),
    .C(_0313_),
    .Y(_0024_));
 sg13g2_a21oi_1 _1253_ (.A1(net133),
    .A2(_0313_),
    .Y(_0314_),
    .B1(net546));
 sg13g2_o21ai_1 _1254_ (.B1(_0314_),
    .Y(_0315_),
    .A1(net133),
    .A2(_0313_));
 sg13g2_inv_1 _1255_ (.Y(_0025_),
    .A(_0315_));
 sg13g2_a21oi_1 _1256_ (.A1(_0278_),
    .A2(\prev_y[0] ),
    .Y(_0316_),
    .B1(\prev_y[3] ));
 sg13g2_a22oi_1 _1257_ (.Y(_0317_),
    .B1(\prev_y[6] ),
    .B2(_0281_),
    .A2(_0287_),
    .A1(net622));
 sg13g2_xnor2_1 _1258_ (.Y(_0318_),
    .A(\pix_y[1] ),
    .B(\prev_y[1] ));
 sg13g2_nor2_1 _1259_ (.A(_0280_),
    .B(\prev_y[5] ),
    .Y(_0319_));
 sg13g2_xnor2_1 _1260_ (.Y(_0320_),
    .A(\pix_y[9] ),
    .B(\prev_y[9] ));
 sg13g2_xnor2_1 _1261_ (.Y(_0321_),
    .A(net624),
    .B(\prev_y[2] ));
 sg13g2_and4_1 _1262_ (.A(_0316_),
    .B(_0317_),
    .C(_0320_),
    .D(_0321_),
    .X(_0322_));
 sg13g2_nor2b_1 _1263_ (.A(\pix_y[7] ),
    .B_N(\prev_y[7] ),
    .Y(_0323_));
 sg13g2_nor2_1 _1264_ (.A(_0284_),
    .B(\prev_y[7] ),
    .Y(_0324_));
 sg13g2_a22oi_1 _1265_ (.Y(_0325_),
    .B1(\prev_y[8] ),
    .B2(_0283_),
    .A2(\prev_y[5] ),
    .A1(_0280_));
 sg13g2_a22oi_1 _1266_ (.Y(_0326_),
    .B1(_0289_),
    .B2(\pix_y[8] ),
    .A2(_0288_),
    .A1(net621));
 sg13g2_a22oi_1 _1267_ (.Y(_0327_),
    .B1(\prev_y[4] ),
    .B2(_0279_),
    .A2(_0285_),
    .A1(\pix_y[0] ));
 sg13g2_nand4_1 _1268_ (.B(_0325_),
    .C(_0326_),
    .A(_0318_),
    .Y(_0328_),
    .D(_0327_));
 sg13g2_nor4_1 _1269_ (.A(_0319_),
    .B(_0323_),
    .C(_0324_),
    .D(_0328_),
    .Y(_0329_));
 sg13g2_nor3_1 _1270_ (.A(net621),
    .B(\pix_y[8] ),
    .C(\pix_y[7] ),
    .Y(_0330_));
 sg13g2_nor4_1 _1271_ (.A(\pix_y[1] ),
    .B(\pix_y[0] ),
    .C(net622),
    .D(\pix_y[5] ),
    .Y(_0331_));
 sg13g2_nor3_1 _1272_ (.A(net624),
    .B(net623),
    .C(\pix_y[9] ),
    .Y(_0332_));
 sg13g2_nand3_1 _1273_ (.B(_0331_),
    .C(_0332_),
    .A(_0330_),
    .Y(_0333_));
 sg13g2_a21oi_1 _1274_ (.A1(_0322_),
    .A2(_0329_),
    .Y(_0334_),
    .B1(_0333_));
 sg13g2_o21ai_1 _1275_ (.B1(net639),
    .Y(_0335_),
    .A1(\logo_left[0] ),
    .A2(net544));
 sg13g2_a21oi_1 _1276_ (.A1(_0276_),
    .A2(net544),
    .Y(_0026_),
    .B1(_0335_));
 sg13g2_nor2b_1 _1277_ (.A(net628),
    .B_N(\logo_left[1] ),
    .Y(_0336_));
 sg13g2_nand2b_1 _1278_ (.Y(_0337_),
    .B(net628),
    .A_N(\logo_left[1] ));
 sg13g2_nand2b_1 _1279_ (.Y(_0338_),
    .B(_0337_),
    .A_N(_0336_));
 sg13g2_xnor2_1 _1280_ (.Y(_0339_),
    .A(net89),
    .B(_0338_));
 sg13g2_o21ai_1 _1281_ (.B1(net639),
    .Y(_0340_),
    .A1(net120),
    .A2(net543));
 sg13g2_a21oi_1 _1282_ (.A1(net543),
    .A2(_0339_),
    .Y(_0027_),
    .B1(_0340_));
 sg13g2_xor2_1 _1283_ (.B(\logo_left[2] ),
    .A(net628),
    .X(_0341_));
 sg13g2_o21ai_1 _1284_ (.B1(_0337_),
    .Y(_0342_),
    .A1(\logo_left[0] ),
    .A2(_0336_));
 sg13g2_nor2_1 _1285_ (.A(_0341_),
    .B(_0342_),
    .Y(_0343_));
 sg13g2_xnor2_1 _1286_ (.Y(_0344_),
    .A(_0341_),
    .B(_0342_));
 sg13g2_o21ai_1 _1287_ (.B1(net639),
    .Y(_0345_),
    .A1(net158),
    .A2(net543));
 sg13g2_a21oi_1 _1288_ (.A1(net543),
    .A2(_0344_),
    .Y(_0028_),
    .B1(_0345_));
 sg13g2_nand2_1 _1289_ (.Y(_0346_),
    .A(net628),
    .B(_0275_));
 sg13g2_xnor2_1 _1290_ (.Y(_0347_),
    .A(net628),
    .B(net631));
 sg13g2_a21oi_1 _1291_ (.A1(_0267_),
    .A2(\logo_left[2] ),
    .Y(_0348_),
    .B1(_0343_));
 sg13g2_xnor2_1 _1292_ (.Y(_0349_),
    .A(_0347_),
    .B(_0348_));
 sg13g2_a21oi_1 _1293_ (.A1(net544),
    .A2(_0349_),
    .Y(_0350_),
    .B1(_0282_));
 sg13g2_o21ai_1 _1294_ (.B1(_0350_),
    .Y(_0029_),
    .A1(_0275_),
    .A2(net543));
 sg13g2_xnor2_1 _1295_ (.Y(_0351_),
    .A(net628),
    .B(\logo_left[4] ));
 sg13g2_or2_1 _1296_ (.X(_0352_),
    .B(\logo_left[2] ),
    .A(net631));
 sg13g2_a22oi_1 _1297_ (.Y(_0353_),
    .B1(_0352_),
    .B2(_0267_),
    .A2(_0346_),
    .A1(_0343_));
 sg13g2_nand2b_1 _1298_ (.Y(_0354_),
    .B(_0351_),
    .A_N(_0353_));
 sg13g2_xnor2_1 _1299_ (.Y(_0355_),
    .A(_0351_),
    .B(_0353_));
 sg13g2_mux2_1 _1300_ (.A0(net171),
    .A1(_0355_),
    .S(net543),
    .X(_0356_));
 sg13g2_and2_1 _1301_ (.A(net638),
    .B(_0356_),
    .X(_0030_));
 sg13g2_o21ai_1 _1302_ (.B1(net638),
    .Y(_0357_),
    .A1(net160),
    .A2(net545));
 sg13g2_xnor2_1 _1303_ (.Y(_0358_),
    .A(net627),
    .B(\logo_left[5] ));
 sg13g2_o21ai_1 _1304_ (.B1(_0354_),
    .Y(_0359_),
    .A1(net627),
    .A2(_0274_));
 sg13g2_xnor2_1 _1305_ (.Y(_0360_),
    .A(_0358_),
    .B(_0359_));
 sg13g2_a21oi_1 _1306_ (.A1(net542),
    .A2(_0360_),
    .Y(_0031_),
    .B1(_0357_));
 sg13g2_nand2_1 _1307_ (.Y(_0361_),
    .A(_0267_),
    .B(net630));
 sg13g2_xor2_1 _1308_ (.B(net630),
    .A(net627),
    .X(_0362_));
 sg13g2_o21ai_1 _1309_ (.B1(_0267_),
    .Y(_0363_),
    .A1(\logo_left[5] ),
    .A2(\logo_left[4] ));
 sg13g2_nand2b_1 _1310_ (.Y(_0364_),
    .B(_0358_),
    .A_N(_0354_));
 sg13g2_and2_1 _1311_ (.A(_0363_),
    .B(_0364_),
    .X(_0365_));
 sg13g2_nand2_1 _1312_ (.Y(_0366_),
    .A(_0362_),
    .B(_0365_));
 sg13g2_or2_1 _1313_ (.X(_0367_),
    .B(_0365_),
    .A(_0362_));
 sg13g2_nand2b_1 _1314_ (.Y(_0368_),
    .B(net630),
    .A_N(net542));
 sg13g2_nand3_1 _1315_ (.B(_0366_),
    .C(_0367_),
    .A(net542),
    .Y(_0369_));
 sg13g2_nand3_1 _1316_ (.B(_0368_),
    .C(_0369_),
    .A(net633),
    .Y(_0032_));
 sg13g2_xor2_1 _1317_ (.B(\logo_left[7] ),
    .A(net627),
    .X(_0370_));
 sg13g2_a21o_1 _1318_ (.A2(_0367_),
    .A1(_0361_),
    .B1(_0370_),
    .X(_0371_));
 sg13g2_nand3_1 _1319_ (.B(_0367_),
    .C(_0370_),
    .A(_0361_),
    .Y(_0372_));
 sg13g2_nand3_1 _1320_ (.B(_0371_),
    .C(_0372_),
    .A(net542),
    .Y(_0373_));
 sg13g2_o21ai_1 _1321_ (.B1(net638),
    .Y(_0374_),
    .A1(_0272_),
    .A2(net542));
 sg13g2_nand2b_1 _1322_ (.Y(_0033_),
    .B(_0373_),
    .A_N(_0374_));
 sg13g2_nor3_1 _1323_ (.A(_0362_),
    .B(_0364_),
    .C(_0370_),
    .Y(_0375_));
 sg13g2_o21ai_1 _1324_ (.B1(_0267_),
    .Y(_0376_),
    .A1(\logo_left[7] ),
    .A2(net630));
 sg13g2_nand2_1 _1325_ (.Y(_0377_),
    .A(_0363_),
    .B(_0376_));
 sg13g2_nor2_1 _1326_ (.A(_0375_),
    .B(_0377_),
    .Y(_0378_));
 sg13g2_xor2_1 _1327_ (.B(net629),
    .A(net627),
    .X(_0379_));
 sg13g2_xnor2_1 _1328_ (.Y(_0380_),
    .A(_0378_),
    .B(_0379_));
 sg13g2_o21ai_1 _1329_ (.B1(net638),
    .Y(_0381_),
    .A1(net629),
    .A2(net542));
 sg13g2_a21oi_1 _1330_ (.A1(net542),
    .A2(_0380_),
    .Y(_0034_),
    .B1(_0381_));
 sg13g2_a21o_1 _1331_ (.A2(net629),
    .A1(net627),
    .B1(_0378_),
    .X(_0382_));
 sg13g2_o21ai_1 _1332_ (.B1(_0378_),
    .Y(_0383_),
    .A1(net627),
    .A2(net629));
 sg13g2_and3_1 _1333_ (.X(_0384_),
    .A(net542),
    .B(_0382_),
    .C(_0383_));
 sg13g2_o21ai_1 _1334_ (.B1(net638),
    .Y(_0385_),
    .A1(net138),
    .A2(_0384_));
 sg13g2_a21oi_1 _1335_ (.A1(net138),
    .A2(_0384_),
    .Y(_0035_),
    .B1(_0385_));
 sg13g2_o21ai_1 _1336_ (.B1(net632),
    .Y(_0386_),
    .A1(\logo_top[0] ),
    .A2(net539));
 sg13g2_a21oi_1 _1337_ (.A1(_0271_),
    .A2(net539),
    .Y(_0036_),
    .B1(_0386_));
 sg13g2_nor2b_1 _1338_ (.A(net625),
    .B_N(\logo_top[1] ),
    .Y(_0387_));
 sg13g2_nand2b_1 _1339_ (.Y(_0388_),
    .B(net625),
    .A_N(\logo_top[1] ));
 sg13g2_nand2b_1 _1340_ (.Y(_0389_),
    .B(_0388_),
    .A_N(_0387_));
 sg13g2_xnor2_1 _1341_ (.Y(_0390_),
    .A(net91),
    .B(_0389_));
 sg13g2_o21ai_1 _1342_ (.B1(net632),
    .Y(_0391_),
    .A1(net126),
    .A2(net539));
 sg13g2_a21oi_1 _1343_ (.A1(net539),
    .A2(_0390_),
    .Y(_0037_),
    .B1(_0391_));
 sg13g2_xor2_1 _1344_ (.B(\logo_top[2] ),
    .A(net625),
    .X(_0392_));
 sg13g2_o21ai_1 _1345_ (.B1(_0388_),
    .Y(_0393_),
    .A1(\logo_top[0] ),
    .A2(_0387_));
 sg13g2_nor2_1 _1346_ (.A(_0392_),
    .B(_0393_),
    .Y(_0394_));
 sg13g2_xnor2_1 _1347_ (.Y(_0395_),
    .A(_0392_),
    .B(_0393_));
 sg13g2_o21ai_1 _1348_ (.B1(net632),
    .Y(_0396_),
    .A1(net167),
    .A2(net539));
 sg13g2_a21oi_1 _1349_ (.A1(net539),
    .A2(_0395_),
    .Y(_0038_),
    .B1(_0396_));
 sg13g2_a21oi_1 _1350_ (.A1(_0266_),
    .A2(\logo_top[2] ),
    .Y(_0397_),
    .B1(_0394_));
 sg13g2_nand2_1 _1351_ (.Y(_0398_),
    .A(_0266_),
    .B(\logo_top[3] ));
 sg13g2_nor2_1 _1352_ (.A(_0266_),
    .B(\logo_top[3] ),
    .Y(_0399_));
 sg13g2_xnor2_1 _1353_ (.Y(_0400_),
    .A(net625),
    .B(\logo_top[3] ));
 sg13g2_xnor2_1 _1354_ (.Y(_0401_),
    .A(_0397_),
    .B(_0400_));
 sg13g2_a21oi_1 _1355_ (.A1(net541),
    .A2(_0401_),
    .Y(_0402_),
    .B1(_0282_));
 sg13g2_o21ai_1 _1356_ (.B1(_0402_),
    .Y(_0039_),
    .A1(_0270_),
    .A2(net541));
 sg13g2_xor2_1 _1357_ (.B(\logo_top[4] ),
    .A(net625),
    .X(_0403_));
 sg13g2_a21oi_1 _1358_ (.A1(_0397_),
    .A2(_0398_),
    .Y(_0404_),
    .B1(_0399_));
 sg13g2_nor2b_1 _1359_ (.A(_0403_),
    .B_N(_0404_),
    .Y(_0405_));
 sg13g2_xor2_1 _1360_ (.B(_0404_),
    .A(_0403_),
    .X(_0406_));
 sg13g2_o21ai_1 _1361_ (.B1(net632),
    .Y(_0407_),
    .A1(net161),
    .A2(net539));
 sg13g2_a21oi_1 _1362_ (.A1(net539),
    .A2(_0406_),
    .Y(_0040_),
    .B1(_0407_));
 sg13g2_o21ai_1 _1363_ (.B1(net632),
    .Y(_0408_),
    .A1(net162),
    .A2(net540));
 sg13g2_xor2_1 _1364_ (.B(\logo_top[5] ),
    .A(net626),
    .X(_0409_));
 sg13g2_inv_1 _1365_ (.Y(_0410_),
    .A(_0409_));
 sg13g2_a21oi_1 _1366_ (.A1(_0266_),
    .A2(\logo_top[4] ),
    .Y(_0411_),
    .B1(_0405_));
 sg13g2_xnor2_1 _1367_ (.Y(_0412_),
    .A(_0409_),
    .B(_0411_));
 sg13g2_a21oi_1 _1368_ (.A1(net540),
    .A2(_0412_),
    .Y(_0041_),
    .B1(_0408_));
 sg13g2_nor2b_1 _1369_ (.A(net626),
    .B_N(\logo_top[6] ),
    .Y(_0413_));
 sg13g2_xor2_1 _1370_ (.B(\logo_top[6] ),
    .A(net625),
    .X(_0414_));
 sg13g2_a21oi_2 _1371_ (.B1(net626),
    .Y(_0415_),
    .A2(_0269_),
    .A1(_0268_));
 sg13g2_nand2_1 _1372_ (.Y(_0416_),
    .A(_0405_),
    .B(_0410_));
 sg13g2_a21oi_1 _1373_ (.A1(_0405_),
    .A2(_0410_),
    .Y(_0417_),
    .B1(_0415_));
 sg13g2_nand2_1 _1374_ (.Y(_0418_),
    .A(_0414_),
    .B(_0417_));
 sg13g2_or2_1 _1375_ (.X(_0419_),
    .B(_0417_),
    .A(_0414_));
 sg13g2_nand2b_1 _1376_ (.Y(_0420_),
    .B(net163),
    .A_N(net540));
 sg13g2_nand3_1 _1377_ (.B(_0418_),
    .C(_0419_),
    .A(net540),
    .Y(_0421_));
 sg13g2_nand3_1 _1378_ (.B(_0420_),
    .C(_0421_),
    .A(net632),
    .Y(_0042_));
 sg13g2_nand2b_1 _1379_ (.Y(_0422_),
    .B(net148),
    .A_N(net540));
 sg13g2_nor2b_1 _1380_ (.A(net625),
    .B_N(\logo_top[7] ),
    .Y(_0423_));
 sg13g2_xor2_1 _1381_ (.B(\logo_top[7] ),
    .A(net626),
    .X(_0424_));
 sg13g2_nor2b_1 _1382_ (.A(_0413_),
    .B_N(_0419_),
    .Y(_0425_));
 sg13g2_o21ai_1 _1383_ (.B1(net540),
    .Y(_0426_),
    .A1(_0424_),
    .A2(_0425_));
 sg13g2_a21oi_1 _1384_ (.A1(_0424_),
    .A2(_0425_),
    .Y(_0427_),
    .B1(_0426_));
 sg13g2_nand3b_1 _1385_ (.B(net633),
    .C(_0422_),
    .Y(_0043_),
    .A_N(_0427_));
 sg13g2_nor3_1 _1386_ (.A(_0414_),
    .B(_0416_),
    .C(_0424_),
    .Y(_0428_));
 sg13g2_nor4_2 _1387_ (.A(_0413_),
    .B(_0415_),
    .C(_0423_),
    .Y(_0429_),
    .D(_0428_));
 sg13g2_xor2_1 _1388_ (.B(\logo_top[8] ),
    .A(net626),
    .X(_0430_));
 sg13g2_xnor2_1 _1389_ (.Y(_0431_),
    .A(_0429_),
    .B(_0430_));
 sg13g2_o21ai_1 _1390_ (.B1(net633),
    .Y(_0432_),
    .A1(net149),
    .A2(net541));
 sg13g2_a21oi_1 _1391_ (.A1(net541),
    .A2(_0431_),
    .Y(_0044_),
    .B1(_0432_));
 sg13g2_a21o_1 _1392_ (.A2(\logo_top[8] ),
    .A1(net626),
    .B1(_0429_),
    .X(_0433_));
 sg13g2_o21ai_1 _1393_ (.B1(_0429_),
    .Y(_0434_),
    .A1(net626),
    .A2(\logo_top[8] ));
 sg13g2_and3_1 _1394_ (.X(_0435_),
    .A(net540),
    .B(_0433_),
    .C(_0434_));
 sg13g2_o21ai_1 _1395_ (.B1(net633),
    .Y(_0436_),
    .A1(net110),
    .A2(_0435_));
 sg13g2_a21oi_1 _1396_ (.A1(net110),
    .A2(_0435_),
    .Y(_0045_),
    .B1(_0436_));
 sg13g2_nor2_1 _1397_ (.A(\logo_left[8] ),
    .B(net631),
    .Y(_0437_));
 sg13g2_a21oi_1 _1398_ (.A1(_0009_),
    .A2(_0437_),
    .Y(_0438_),
    .B1(\logo_left[4] ));
 sg13g2_nor2b_1 _1399_ (.A(_0009_),
    .B_N(net631),
    .Y(_0439_));
 sg13g2_o21ai_1 _1400_ (.B1(_0439_),
    .Y(_0440_),
    .A1(net629),
    .A2(_0007_));
 sg13g2_a21oi_1 _1401_ (.A1(\logo_left[4] ),
    .A2(_0440_),
    .Y(_0441_),
    .B1(_0438_));
 sg13g2_nand4_1 _1402_ (.B(\logo_left[1] ),
    .C(\logo_left[0] ),
    .A(\logo_left[2] ),
    .Y(_0442_),
    .D(_0441_));
 sg13g2_nor3_1 _1403_ (.A(\logo_left[7] ),
    .B(net630),
    .C(\logo_left[5] ),
    .Y(_0443_));
 sg13g2_a21oi_1 _1404_ (.A1(\logo_left[9] ),
    .A2(_0443_),
    .Y(_0444_),
    .B1(net629));
 sg13g2_nand2_1 _1405_ (.Y(_0445_),
    .A(net630),
    .B(\logo_left[5] ));
 sg13g2_nor4_1 _1406_ (.A(\logo_left[9] ),
    .B(_0272_),
    .C(_0007_),
    .D(_0445_),
    .Y(_0446_));
 sg13g2_nor2b_1 _1407_ (.A(_0446_),
    .B_N(net629),
    .Y(_0447_));
 sg13g2_nor3_1 _1408_ (.A(_0442_),
    .B(_0444_),
    .C(_0447_),
    .Y(_0448_));
 sg13g2_o21ai_1 _1409_ (.B1(net543),
    .Y(_0449_),
    .A1(_0267_),
    .A2(_0448_));
 sg13g2_nor3_1 _1410_ (.A(\logo_left[9] ),
    .B(\logo_left[1] ),
    .C(_0352_),
    .Y(_0450_));
 sg13g2_nand4_1 _1411_ (.B(_0007_),
    .C(_0008_),
    .A(\logo_left[0] ),
    .Y(_0451_),
    .D(_0450_));
 sg13g2_nor4_2 _1412_ (.A(\logo_left[7] ),
    .B(net630),
    .C(\logo_left[5] ),
    .Y(_0452_),
    .D(_0451_));
 sg13g2_nor2_1 _1413_ (.A(net628),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_nand3_1 _1414_ (.B(net543),
    .C(_0452_),
    .A(_0267_),
    .Y(_0454_));
 sg13g2_o21ai_1 _1415_ (.B1(net628),
    .Y(_0455_),
    .A1(net99),
    .A2(_0449_));
 sg13g2_nand3_1 _1416_ (.B(_0454_),
    .C(net100),
    .A(net638),
    .Y(_0046_));
 sg13g2_nand4_1 _1417_ (.B(\logo_top[4] ),
    .C(\logo_top[2] ),
    .A(\logo_top[6] ),
    .Y(_0456_),
    .D(\logo_top[1] ));
 sg13g2_nor3_1 _1418_ (.A(_0270_),
    .B(_0003_),
    .C(_0456_),
    .Y(_0457_));
 sg13g2_nor3_1 _1419_ (.A(\logo_top[9] ),
    .B(\logo_top[7] ),
    .C(\logo_top[5] ),
    .Y(_0458_));
 sg13g2_nor2_1 _1420_ (.A(\logo_top[2] ),
    .B(\logo_top[1] ),
    .Y(_0459_));
 sg13g2_nand3_1 _1421_ (.B(_0003_),
    .C(_0459_),
    .A(_0002_),
    .Y(_0460_));
 sg13g2_nor3_1 _1422_ (.A(\logo_top[6] ),
    .B(\logo_top[3] ),
    .C(_0460_),
    .Y(_0461_));
 sg13g2_mux2_1 _1423_ (.A0(_0457_),
    .A1(_0461_),
    .S(_0266_),
    .X(_0462_));
 sg13g2_nand4_1 _1424_ (.B(net540),
    .C(_0458_),
    .A(\logo_top[0] ),
    .Y(_0463_),
    .D(_0462_));
 sg13g2_and2_1 _1425_ (.A(_0266_),
    .B(_0463_),
    .X(_0464_));
 sg13g2_nor3_1 _1426_ (.A(_0266_),
    .B(net106),
    .C(_0463_),
    .Y(_0465_));
 sg13g2_nor3_1 _1427_ (.A(_0282_),
    .B(_0464_),
    .C(_0465_),
    .Y(_0047_));
 sg13g2_o21ai_1 _1428_ (.B1(_0463_),
    .Y(_0466_),
    .A1(_0449_),
    .A2(_0453_));
 sg13g2_o21ai_1 _1429_ (.B1(net639),
    .Y(_0467_),
    .A1(\color_index[0] ),
    .A2(_0466_));
 sg13g2_a21oi_1 _1430_ (.A1(_0265_),
    .A2(_0466_),
    .Y(_0048_),
    .B1(_0467_));
 sg13g2_and2_1 _1431_ (.A(\color_index[0] ),
    .B(_0466_),
    .X(_0468_));
 sg13g2_nand2_1 _1432_ (.Y(_0469_),
    .A(net123),
    .B(_0468_));
 sg13g2_o21ai_1 _1433_ (.B1(net639),
    .Y(_0470_),
    .A1(net123),
    .A2(_0468_));
 sg13g2_nor2b_1 _1434_ (.A(net124),
    .B_N(_0469_),
    .Y(_0049_));
 sg13g2_o21ai_1 _1435_ (.B1(net639),
    .Y(_0471_),
    .A1(_0264_),
    .A2(_0469_));
 sg13g2_a21oi_1 _1436_ (.A1(_0264_),
    .A2(_0469_),
    .Y(_0050_),
    .B1(_0471_));
 sg13g2_nor2_1 _1437_ (.A(net634),
    .B(net102),
    .Y(_0472_));
 sg13g2_a21oi_1 _1438_ (.A1(_0278_),
    .A2(net634),
    .Y(_0051_),
    .B1(_0472_));
 sg13g2_nand2_1 _1439_ (.Y(_0473_),
    .A(\pix_y[1] ),
    .B(net633));
 sg13g2_o21ai_1 _1440_ (.B1(_0473_),
    .Y(_0052_),
    .A1(net632),
    .A2(_0286_));
 sg13g2_mux2_1 _1441_ (.A0(net108),
    .A1(net624),
    .S(net634),
    .X(_0053_));
 sg13g2_nor2b_1 _1442_ (.A(net623),
    .B_N(net634),
    .Y(_0474_));
 sg13g2_nor2_1 _1443_ (.A(net634),
    .B(net93),
    .Y(_0475_));
 sg13g2_nor2_1 _1444_ (.A(_0474_),
    .B(_0475_),
    .Y(_0054_));
 sg13g2_mux2_1 _1445_ (.A0(net119),
    .A1(net622),
    .S(net634),
    .X(_0055_));
 sg13g2_nor2_1 _1446_ (.A(net636),
    .B(net115),
    .Y(_0476_));
 sg13g2_a21oi_1 _1447_ (.A1(_0280_),
    .A2(net636),
    .Y(_0056_),
    .B1(_0476_));
 sg13g2_mux2_1 _1448_ (.A0(net121),
    .A1(net621),
    .S(net635),
    .X(_0057_));
 sg13g2_nor2_1 _1449_ (.A(net635),
    .B(net104),
    .Y(_0477_));
 sg13g2_a21oi_1 _1450_ (.A1(net635),
    .A2(_0284_),
    .Y(_0058_),
    .B1(_0477_));
 sg13g2_nor2_1 _1451_ (.A(net635),
    .B(net111),
    .Y(_0478_));
 sg13g2_a21oi_1 _1452_ (.A1(net635),
    .A2(_0283_),
    .Y(_0059_),
    .B1(_0478_));
 sg13g2_mux2_1 _1453_ (.A0(net113),
    .A1(\pix_y[9] ),
    .S(net635),
    .X(_0060_));
 sg13g2_nor2b_1 _1454_ (.A(\logo_left[4] ),
    .B_N(\pix_x[4] ),
    .Y(_0479_));
 sg13g2_nor2b_1 _1455_ (.A(\logo_left[1] ),
    .B_N(\pix_x[1] ),
    .Y(_0480_));
 sg13g2_nand2b_1 _1456_ (.Y(_0481_),
    .B(\logo_left[0] ),
    .A_N(\pix_x[0] ));
 sg13g2_xnor2_1 _1457_ (.Y(_0482_),
    .A(\logo_left[1] ),
    .B(\pix_x[1] ));
 sg13g2_nand2_1 _1458_ (.Y(_0483_),
    .A(_0481_),
    .B(_0482_));
 sg13g2_a21oi_2 _1459_ (.B1(_0480_),
    .Y(_0484_),
    .A2(_0482_),
    .A1(_0481_));
 sg13g2_inv_1 _1460_ (.Y(_0485_),
    .A(_0484_));
 sg13g2_nor2b_1 _1461_ (.A(\logo_left[3] ),
    .B_N(\pix_x[3] ),
    .Y(_0486_));
 sg13g2_nand2b_1 _1462_ (.Y(_0487_),
    .B(\logo_left[3] ),
    .A_N(\pix_x[3] ));
 sg13g2_xnor2_1 _1463_ (.Y(_0488_),
    .A(\logo_left[3] ),
    .B(\pix_x[3] ));
 sg13g2_nor2b_1 _1464_ (.A(\logo_left[2] ),
    .B_N(\pix_x[2] ),
    .Y(_0489_));
 sg13g2_xnor2_1 _1465_ (.Y(_0490_),
    .A(\logo_left[2] ),
    .B(\pix_x[2] ));
 sg13g2_nand2_1 _1466_ (.Y(_0491_),
    .A(_0488_),
    .B(_0490_));
 sg13g2_a21oi_1 _1467_ (.A1(_0487_),
    .A2(_0489_),
    .Y(_0492_),
    .B1(_0486_));
 sg13g2_o21ai_1 _1468_ (.B1(_0492_),
    .Y(_0493_),
    .A1(_0484_),
    .A2(_0491_));
 sg13g2_xnor2_1 _1469_ (.Y(_0494_),
    .A(\logo_left[4] ),
    .B(\pix_x[4] ));
 sg13g2_a21o_1 _1470_ (.A2(_0494_),
    .A1(_0493_),
    .B1(_0479_),
    .X(_0495_));
 sg13g2_nor2_2 _1471_ (.A(_0273_),
    .B(\pix_x[5] ),
    .Y(_0496_));
 sg13g2_inv_1 _1472_ (.Y(_0497_),
    .A(_0496_));
 sg13g2_nor2b_1 _1473_ (.A(\logo_left[5] ),
    .B_N(\pix_x[5] ),
    .Y(_0498_));
 sg13g2_nor2_1 _1474_ (.A(_0496_),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_xor2_1 _1475_ (.B(_0499_),
    .A(_0495_),
    .X(_0500_));
 sg13g2_xnor2_1 _1476_ (.Y(_0501_),
    .A(_0495_),
    .B(_0499_));
 sg13g2_xor2_1 _1477_ (.B(_0494_),
    .A(_0493_),
    .X(_0502_));
 sg13g2_xnor2_1 _1478_ (.Y(_0503_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_nor2_2 _1479_ (.A(net535),
    .B(net568),
    .Y(_0504_));
 sg13g2_nand2_1 _1480_ (.Y(_0505_),
    .A(net532),
    .B(net573));
 sg13g2_nand2b_2 _1481_ (.Y(_0506_),
    .B(\logo_top[0] ),
    .A_N(\pix_y[0] ));
 sg13g2_nor2b_1 _1482_ (.A(\logo_top[1] ),
    .B_N(\pix_y[1] ),
    .Y(_0507_));
 sg13g2_xnor2_1 _1483_ (.Y(_0508_),
    .A(\logo_top[1] ),
    .B(\pix_y[1] ));
 sg13g2_xor2_1 _1484_ (.B(_0508_),
    .A(_0506_),
    .X(_0509_));
 sg13g2_xnor2_1 _1485_ (.Y(_0510_),
    .A(_0506_),
    .B(_0508_));
 sg13g2_nand2b_1 _1486_ (.Y(_0511_),
    .B(\pix_x[6] ),
    .A_N(\logo_left[6] ));
 sg13g2_nand2b_1 _1487_ (.Y(_0512_),
    .B(net630),
    .A_N(\pix_x[6] ));
 sg13g2_and2_1 _1488_ (.A(_0511_),
    .B(_0512_),
    .X(_0513_));
 sg13g2_nand2_1 _1489_ (.Y(_0514_),
    .A(_0511_),
    .B(_0512_));
 sg13g2_a221oi_1 _1490_ (.B2(_0494_),
    .C1(_0479_),
    .B1(_0493_),
    .A1(_0273_),
    .Y(_0515_),
    .A2(\pix_x[5] ));
 sg13g2_nor3_2 _1491_ (.A(_0496_),
    .B(_0514_),
    .C(_0515_),
    .Y(_0516_));
 sg13g2_or3_1 _1492_ (.A(_0496_),
    .B(_0514_),
    .C(_0515_),
    .X(_0517_));
 sg13g2_a221oi_1 _1493_ (.B2(_0512_),
    .C1(_0498_),
    .B1(_0511_),
    .A1(_0495_),
    .Y(_0518_),
    .A2(_0497_));
 sg13g2_o21ai_1 _1494_ (.B1(_0514_),
    .Y(_0519_),
    .A1(_0496_),
    .A2(_0515_));
 sg13g2_or3_1 _1495_ (.A(_0496_),
    .B(_0513_),
    .C(_0515_),
    .X(_0520_));
 sg13g2_o21ai_1 _1496_ (.B1(_0513_),
    .Y(_0521_),
    .A1(_0496_),
    .A2(_0515_));
 sg13g2_nor2_1 _1497_ (.A(net530),
    .B(net527),
    .Y(_0522_));
 sg13g2_nand2_2 _1498_ (.Y(_0523_),
    .A(net528),
    .B(net525));
 sg13g2_nand2_2 _1499_ (.Y(_0524_),
    .A(net537),
    .B(net570));
 sg13g2_nor3_2 _1500_ (.A(net572),
    .B(net530),
    .C(net527),
    .Y(_0525_));
 sg13g2_nand3_1 _1501_ (.B(net528),
    .C(net525),
    .A(net569),
    .Y(_0526_));
 sg13g2_nor4_2 _1502_ (.A(net531),
    .B(net571),
    .C(net530),
    .Y(_0527_),
    .D(net527));
 sg13g2_nand4_1 _1503_ (.B(net568),
    .C(net529),
    .A(net535),
    .Y(_0528_),
    .D(net526));
 sg13g2_nor2_2 _1504_ (.A(net610),
    .B(_0527_),
    .Y(_0529_));
 sg13g2_nor2_1 _1505_ (.A(net538),
    .B(_0502_),
    .Y(_0530_));
 sg13g2_nand2_2 _1506_ (.Y(_0531_),
    .A(net533),
    .B(net570));
 sg13g2_nor2_2 _1507_ (.A(net531),
    .B(net568),
    .Y(_0532_));
 sg13g2_nand2_2 _1508_ (.Y(_0533_),
    .A(net537),
    .B(net572));
 sg13g2_a21oi_2 _1509_ (.B1(net573),
    .Y(_0534_),
    .A2(net526),
    .A1(net529));
 sg13g2_o21ai_1 _1510_ (.B1(net569),
    .Y(_0535_),
    .A1(net530),
    .A2(net527));
 sg13g2_nor2_1 _1511_ (.A(_0504_),
    .B(_0527_),
    .Y(_0536_));
 sg13g2_nand2_1 _1512_ (.Y(_0537_),
    .A(net537),
    .B(net605));
 sg13g2_a21oi_2 _1513_ (.B1(net610),
    .Y(_0538_),
    .A2(net572),
    .A1(net531));
 sg13g2_nand2_1 _1514_ (.Y(_0539_),
    .A(net505),
    .B(net504));
 sg13g2_a21oi_2 _1515_ (.B1(_0507_),
    .Y(_0540_),
    .A2(_0508_),
    .A1(_0506_));
 sg13g2_nand2b_1 _1516_ (.Y(_0541_),
    .B(\pix_y[2] ),
    .A_N(\logo_top[2] ));
 sg13g2_nor2b_1 _1517_ (.A(\pix_y[2] ),
    .B_N(\logo_top[2] ),
    .Y(_0542_));
 sg13g2_xnor2_1 _1518_ (.Y(_0543_),
    .A(\logo_top[2] ),
    .B(net624));
 sg13g2_xnor2_1 _1519_ (.Y(_0544_),
    .A(_0540_),
    .B(_0543_));
 sg13g2_xor2_1 _1520_ (.B(_0543_),
    .A(_0540_),
    .X(_0545_));
 sg13g2_nor2_2 _1521_ (.A(net609),
    .B(net591),
    .Y(_0546_));
 sg13g2_nand2_2 _1522_ (.Y(_0547_),
    .A(net602),
    .B(net579));
 sg13g2_xnor2_1 _1523_ (.Y(_0548_),
    .A(net533),
    .B(net572));
 sg13g2_xnor2_1 _1524_ (.Y(_0549_),
    .A(net535),
    .B(net571));
 sg13g2_nor3_2 _1525_ (.A(net531),
    .B(net530),
    .C(net527),
    .Y(_0550_));
 sg13g2_nand3_1 _1526_ (.B(net528),
    .C(net525),
    .A(net535),
    .Y(_0551_));
 sg13g2_nor2_2 _1527_ (.A(_0532_),
    .B(_0550_),
    .Y(_0552_));
 sg13g2_a21oi_2 _1528_ (.B1(net532),
    .Y(_0553_),
    .A2(net525),
    .A1(net528));
 sg13g2_o21ai_1 _1529_ (.B1(net536),
    .Y(_0554_),
    .A1(_0516_),
    .A2(_0518_));
 sg13g2_and4_2 _1530_ (.A(net535),
    .B(net569),
    .C(net524),
    .D(net523),
    .X(_0555_));
 sg13g2_nand4_1 _1531_ (.B(net568),
    .C(_0520_),
    .A(net536),
    .Y(_0556_),
    .D(_0521_));
 sg13g2_nand2_1 _1532_ (.Y(_0557_),
    .A(net512),
    .B(net501));
 sg13g2_a21o_1 _1533_ (.A2(_0557_),
    .A1(net587),
    .B1(_0546_),
    .X(_0558_));
 sg13g2_nor2b_1 _1534_ (.A(\logo_top[3] ),
    .B_N(net623),
    .Y(_0559_));
 sg13g2_xnor2_1 _1535_ (.Y(_0560_),
    .A(\logo_top[3] ),
    .B(net623));
 sg13g2_o21ai_1 _1536_ (.B1(_0541_),
    .Y(_0561_),
    .A1(_0540_),
    .A2(_0542_));
 sg13g2_xor2_1 _1537_ (.B(_0561_),
    .A(_0560_),
    .X(_0562_));
 sg13g2_xnor2_1 _1538_ (.Y(_0563_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_nor3_2 _1539_ (.A(net536),
    .B(_0516_),
    .C(_0518_),
    .Y(_0564_));
 sg13g2_nand3_1 _1540_ (.B(net529),
    .C(net525),
    .A(net531),
    .Y(_0565_));
 sg13g2_nand2_2 _1541_ (.Y(_0566_),
    .A(net503),
    .B(net500));
 sg13g2_nand3_1 _1542_ (.B(net502),
    .C(net499),
    .A(net571),
    .Y(_0567_));
 sg13g2_nand2_1 _1543_ (.Y(_0568_),
    .A(net613),
    .B(_0567_));
 sg13g2_nand2_2 _1544_ (.Y(_0569_),
    .A(net571),
    .B(net589));
 sg13g2_nor2_1 _1545_ (.A(_0564_),
    .B(_0569_),
    .Y(_0570_));
 sg13g2_a221oi_1 _1546_ (.B2(_0570_),
    .C1(net552),
    .B1(_0568_),
    .A1(_0539_),
    .Y(_0571_),
    .A2(_0558_));
 sg13g2_nand2_1 _1547_ (.Y(_0572_),
    .A(_0269_),
    .B(net622));
 sg13g2_a21oi_2 _1548_ (.B1(_0559_),
    .Y(_0573_),
    .A2(_0561_),
    .A1(_0560_));
 sg13g2_xor2_1 _1549_ (.B(net622),
    .A(\logo_top[4] ),
    .X(_0574_));
 sg13g2_o21ai_1 _1550_ (.B1(_0572_),
    .Y(_0575_),
    .A1(_0573_),
    .A2(_0574_));
 sg13g2_xnor2_1 _1551_ (.Y(_0576_),
    .A(\logo_top[5] ),
    .B(\pix_y[5] ));
 sg13g2_xnor2_1 _1552_ (.Y(_0577_),
    .A(_0575_),
    .B(_0576_));
 sg13g2_xor2_1 _1553_ (.B(_0576_),
    .A(_0575_),
    .X(_0578_));
 sg13g2_nand2_2 _1554_ (.Y(_0579_),
    .A(_0526_),
    .B(net500));
 sg13g2_nor2_1 _1555_ (.A(_0525_),
    .B(_0564_),
    .Y(_0580_));
 sg13g2_a221oi_1 _1556_ (.B2(net523),
    .C1(net594),
    .B1(net524),
    .A1(net536),
    .Y(_0581_),
    .A2(net573));
 sg13g2_nor2_1 _1557_ (.A(net603),
    .B(net594),
    .Y(_0582_));
 sg13g2_nand2_1 _1558_ (.Y(_0583_),
    .A(net616),
    .B(net587));
 sg13g2_nand2b_1 _1559_ (.Y(_0584_),
    .B(_0583_),
    .A_N(_0581_));
 sg13g2_a21oi_1 _1560_ (.A1(net528),
    .A2(net525),
    .Y(_0585_),
    .B1(net569));
 sg13g2_o21ai_1 _1561_ (.B1(net571),
    .Y(_0586_),
    .A1(net530),
    .A2(net527));
 sg13g2_nor2_2 _1562_ (.A(net605),
    .B(_0564_),
    .Y(_0587_));
 sg13g2_nand2_1 _1563_ (.Y(_0588_),
    .A(net614),
    .B(net500));
 sg13g2_nand3_1 _1564_ (.B(net528),
    .C(net525),
    .A(net610),
    .Y(_0589_));
 sg13g2_nand2_2 _1565_ (.Y(_0590_),
    .A(net570),
    .B(net611));
 sg13g2_nor2_2 _1566_ (.A(net602),
    .B(net493),
    .Y(_0591_));
 sg13g2_a221oi_1 _1567_ (.B2(_0587_),
    .C1(net595),
    .B1(_0586_),
    .A1(net605),
    .Y(_0592_),
    .A2(_0580_));
 sg13g2_nor2_2 _1568_ (.A(net589),
    .B(net559),
    .Y(_0593_));
 sg13g2_nand2_2 _1569_ (.Y(_0594_),
    .A(net574),
    .B(net547));
 sg13g2_and2_1 _1570_ (.A(net534),
    .B(_0589_),
    .X(_0595_));
 sg13g2_nand2_1 _1571_ (.Y(_0596_),
    .A(_0504_),
    .B(_0589_));
 sg13g2_a21oi_1 _1572_ (.A1(_0504_),
    .A2(_0589_),
    .Y(_0597_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1573_ (.B1(net555),
    .Y(_0598_),
    .A1(net584),
    .A2(_0597_));
 sg13g2_xor2_1 _1574_ (.B(_0574_),
    .A(_0573_),
    .X(_0599_));
 sg13g2_xnor2_1 _1575_ (.Y(_0600_),
    .A(_0573_),
    .B(_0574_));
 sg13g2_and4_2 _1576_ (.A(net535),
    .B(net571),
    .C(net524),
    .D(net523),
    .X(_0601_));
 sg13g2_nand4_1 _1577_ (.B(net571),
    .C(net524),
    .A(net535),
    .Y(_0602_),
    .D(net523));
 sg13g2_a21oi_2 _1578_ (.B1(net609),
    .Y(_0603_),
    .A2(net526),
    .A1(net529));
 sg13g2_o21ai_1 _1579_ (.B1(net602),
    .Y(_0604_),
    .A1(net530),
    .A2(net527));
 sg13g2_nor2_1 _1580_ (.A(net597),
    .B(_0601_),
    .Y(_0605_));
 sg13g2_a21oi_1 _1581_ (.A1(net604),
    .A2(_0601_),
    .Y(_0606_),
    .B1(net592));
 sg13g2_o21ai_1 _1582_ (.B1(net586),
    .Y(_0607_),
    .A1(net617),
    .A2(net491));
 sg13g2_nor2_1 _1583_ (.A(net534),
    .B(net603),
    .Y(_0608_));
 sg13g2_nand2_1 _1584_ (.Y(_0609_),
    .A(net538),
    .B(net609));
 sg13g2_nand2_1 _1585_ (.Y(_0610_),
    .A(net573),
    .B(net510));
 sg13g2_nor2_1 _1586_ (.A(_0525_),
    .B(net493),
    .Y(_0611_));
 sg13g2_nand2_1 _1587_ (.Y(_0612_),
    .A(net506),
    .B(_0586_));
 sg13g2_a21oi_2 _1588_ (.B1(net536),
    .Y(_0613_),
    .A2(net526),
    .A1(net529));
 sg13g2_o21ai_1 _1589_ (.B1(net531),
    .Y(_0614_),
    .A1(_0516_),
    .A2(_0518_));
 sg13g2_a22oi_1 _1590_ (.Y(_0615_),
    .B1(net529),
    .B2(net526),
    .A2(net569),
    .A1(net535));
 sg13g2_nand2_1 _1591_ (.Y(_0616_),
    .A(_0591_),
    .B(net490));
 sg13g2_nor2_2 _1592_ (.A(net618),
    .B(_0530_),
    .Y(_0617_));
 sg13g2_nand2_1 _1593_ (.Y(_0618_),
    .A(net509),
    .B(_0531_));
 sg13g2_nand2_2 _1594_ (.Y(_0619_),
    .A(net510),
    .B(_0548_));
 sg13g2_a22oi_1 _1595_ (.Y(_0620_),
    .B1(_0617_),
    .B2(_0579_),
    .A2(_0611_),
    .A1(_0608_));
 sg13g2_a221oi_1 _1596_ (.B2(net592),
    .C1(net550),
    .B1(_0620_),
    .A1(net499),
    .Y(_0621_),
    .A2(_0606_));
 sg13g2_nand4_1 _1597_ (.B(net568),
    .C(net524),
    .A(net532),
    .Y(_0622_),
    .D(net523));
 sg13g2_nand2_2 _1598_ (.Y(_0623_),
    .A(net615),
    .B(_0622_));
 sg13g2_a21oi_2 _1599_ (.B1(net595),
    .Y(_0624_),
    .A2(net505),
    .A1(net600));
 sg13g2_nor2_1 _1600_ (.A(net583),
    .B(_0550_),
    .Y(_0625_));
 sg13g2_a22oi_1 _1601_ (.Y(_0626_),
    .B1(_0625_),
    .B2(_0616_),
    .A2(_0624_),
    .A1(_0623_));
 sg13g2_nor2b_1 _1602_ (.A(\logo_top[6] ),
    .B_N(net621),
    .Y(_0627_));
 sg13g2_nand2b_1 _1603_ (.Y(_0628_),
    .B(\logo_top[6] ),
    .A_N(net621));
 sg13g2_nand2b_1 _1604_ (.Y(_0629_),
    .B(_0628_),
    .A_N(_0627_));
 sg13g2_a21oi_1 _1605_ (.A1(_0268_),
    .A2(\pix_y[5] ),
    .Y(_0630_),
    .B1(_0575_));
 sg13g2_a21oi_2 _1606_ (.B1(_0630_),
    .Y(_0631_),
    .A2(_0280_),
    .A1(\logo_top[5] ));
 sg13g2_xnor2_1 _1607_ (.Y(_0632_),
    .A(_0629_),
    .B(_0631_));
 sg13g2_xor2_1 _1608_ (.B(_0631_),
    .A(_0629_),
    .X(_0633_));
 sg13g2_nand2_1 _1609_ (.Y(_0634_),
    .A(_0504_),
    .B(net509));
 sg13g2_nor2_1 _1610_ (.A(_0538_),
    .B(_0603_),
    .Y(_0635_));
 sg13g2_nand2_1 _1611_ (.Y(_0636_),
    .A(net534),
    .B(net614));
 sg13g2_a21oi_2 _1612_ (.B1(net587),
    .Y(_0637_),
    .A2(_0602_),
    .A1(net616));
 sg13g2_a221oi_1 _1613_ (.B2(_0637_),
    .C1(net554),
    .B1(_0635_),
    .A1(net587),
    .Y(_0638_),
    .A2(_0557_));
 sg13g2_nand3_1 _1614_ (.B(net581),
    .C(net503),
    .A(net512),
    .Y(_0639_));
 sg13g2_nand4_1 _1615_ (.B(net573),
    .C(net524),
    .A(net534),
    .Y(_0640_),
    .D(net523));
 sg13g2_nor2_2 _1616_ (.A(net608),
    .B(net493),
    .Y(_0641_));
 sg13g2_and2_1 _1617_ (.A(net606),
    .B(net488),
    .X(_0642_));
 sg13g2_nand2_2 _1618_ (.Y(_0643_),
    .A(net604),
    .B(net487));
 sg13g2_a21oi_2 _1619_ (.B1(net592),
    .Y(_0644_),
    .A2(net487),
    .A1(net604));
 sg13g2_a22oi_1 _1620_ (.Y(_0645_),
    .B1(net524),
    .B2(net523),
    .A2(net568),
    .A1(net538));
 sg13g2_nand2_1 _1621_ (.Y(_0646_),
    .A(net509),
    .B(_0524_));
 sg13g2_nor2_2 _1622_ (.A(_0523_),
    .B(_0548_),
    .Y(_0647_));
 sg13g2_nand2_2 _1623_ (.Y(_0648_),
    .A(net512),
    .B(_0645_));
 sg13g2_nor2_1 _1624_ (.A(_0534_),
    .B(net581),
    .Y(_0649_));
 sg13g2_a21o_1 _1625_ (.A2(_0649_),
    .A1(_0648_),
    .B1(_0644_),
    .X(_0650_));
 sg13g2_a21oi_1 _1626_ (.A1(_0639_),
    .A2(_0650_),
    .Y(_0651_),
    .B1(net563));
 sg13g2_nand2_1 _1627_ (.Y(_0652_),
    .A(net504),
    .B(_0645_));
 sg13g2_a21oi_1 _1628_ (.A1(net507),
    .A2(net489),
    .Y(_0653_),
    .B1(net597));
 sg13g2_nor2_2 _1629_ (.A(net600),
    .B(_0525_),
    .Y(_0654_));
 sg13g2_nand2_2 _1630_ (.Y(_0655_),
    .A(net608),
    .B(net506));
 sg13g2_or2_1 _1631_ (.X(_0656_),
    .B(_0653_),
    .A(_0546_));
 sg13g2_nand3_1 _1632_ (.B(net499),
    .C(_0622_),
    .A(net602),
    .Y(_0657_));
 sg13g2_and2_1 _1633_ (.A(net596),
    .B(_0657_),
    .X(_0658_));
 sg13g2_o21ai_1 _1634_ (.B1(net616),
    .Y(_0659_),
    .A1(net512),
    .A2(_0523_));
 sg13g2_nand2_1 _1635_ (.Y(_0660_),
    .A(net612),
    .B(_0619_));
 sg13g2_nand2b_1 _1636_ (.Y(_0661_),
    .B(net503),
    .A_N(_0659_));
 sg13g2_nand2_1 _1637_ (.Y(_0662_),
    .A(net606),
    .B(net501));
 sg13g2_a21oi_2 _1638_ (.B1(net584),
    .Y(_0663_),
    .A2(net501),
    .A1(net605));
 sg13g2_nand4_1 _1639_ (.B(net569),
    .C(net528),
    .A(net532),
    .Y(_0664_),
    .D(net525));
 sg13g2_nor4_2 _1640_ (.A(net537),
    .B(net530),
    .C(net527),
    .Y(_0665_),
    .D(_0590_));
 sg13g2_nor2_1 _1641_ (.A(net604),
    .B(net501),
    .Y(_0666_));
 sg13g2_a21oi_1 _1642_ (.A1(net501),
    .A2(net486),
    .Y(_0667_),
    .B1(net606));
 sg13g2_o21ai_1 _1643_ (.B1(net514),
    .Y(_0668_),
    .A1(_0638_),
    .A2(_0651_));
 sg13g2_o21ai_1 _1644_ (.B1(net521),
    .Y(_0669_),
    .A1(net565),
    .A2(_0626_));
 sg13g2_o21ai_1 _1645_ (.B1(_0668_),
    .Y(_0670_),
    .A1(_0621_),
    .A2(_0669_));
 sg13g2_a221oi_1 _1646_ (.B2(net585),
    .C1(net565),
    .B1(_0667_),
    .A1(_0661_),
    .Y(_0671_),
    .A2(_0663_));
 sg13g2_a221oi_1 _1647_ (.B2(_0660_),
    .C1(net553),
    .B1(_0658_),
    .A1(_0652_),
    .Y(_0672_),
    .A2(_0656_));
 sg13g2_nor3_1 _1648_ (.A(net521),
    .B(_0671_),
    .C(_0672_),
    .Y(_0673_));
 sg13g2_o21ai_1 _1649_ (.B1(net519),
    .Y(_0674_),
    .A1(_0592_),
    .A2(_0598_));
 sg13g2_o21ai_1 _1650_ (.B1(net497),
    .Y(_0675_),
    .A1(_0571_),
    .A2(_0674_));
 sg13g2_o21ai_1 _1651_ (.B1(net484),
    .Y(_0676_),
    .A1(_0673_),
    .A2(_0675_));
 sg13g2_a21o_1 _1652_ (.A2(_0670_),
    .A1(net494),
    .B1(_0676_),
    .X(_0677_));
 sg13g2_or2_1 _1653_ (.X(_0678_),
    .B(_0482_),
    .A(_0481_));
 sg13g2_and2_2 _1654_ (.A(_0483_),
    .B(_0678_),
    .X(_0679_));
 sg13g2_nand2_2 _1655_ (.Y(_0680_),
    .A(_0483_),
    .B(_0678_));
 sg13g2_nand3_1 _1656_ (.B(net491),
    .C(_0619_),
    .A(net617),
    .Y(_0681_));
 sg13g2_nor2_1 _1657_ (.A(net585),
    .B(_0617_),
    .Y(_0682_));
 sg13g2_nand2_1 _1658_ (.Y(_0683_),
    .A(_0531_),
    .B(net490));
 sg13g2_a221oi_1 _1659_ (.B2(net585),
    .C1(net553),
    .B1(_0683_),
    .A1(_0681_),
    .Y(_0684_),
    .A2(_0682_));
 sg13g2_a21oi_2 _1660_ (.B1(net578),
    .Y(_0685_),
    .A2(net505),
    .A1(net603));
 sg13g2_a221oi_1 _1661_ (.B2(_0685_),
    .C1(net566),
    .B1(_0659_),
    .A1(net585),
    .Y(_0686_),
    .A2(_0601_));
 sg13g2_o21ai_1 _1662_ (.B1(net515),
    .Y(_0687_),
    .A1(_0684_),
    .A2(_0686_));
 sg13g2_a21oi_1 _1663_ (.A1(_0537_),
    .A2(_0590_),
    .Y(_0688_),
    .B1(_0594_));
 sg13g2_a21oi_1 _1664_ (.A1(_0646_),
    .A2(_0688_),
    .Y(_0689_),
    .B1(net516));
 sg13g2_nand2_1 _1665_ (.Y(_0690_),
    .A(net618),
    .B(_0535_));
 sg13g2_nor2_2 _1666_ (.A(net602),
    .B(net577),
    .Y(_0691_));
 sg13g2_nand2_2 _1667_ (.Y(_0692_),
    .A(net608),
    .B(net591));
 sg13g2_o21ai_1 _1668_ (.B1(net591),
    .Y(_0693_),
    .A1(net531),
    .A2(net568));
 sg13g2_nor2_1 _1669_ (.A(_0566_),
    .B(_0693_),
    .Y(_0694_));
 sg13g2_nor3_1 _1670_ (.A(net573),
    .B(net580),
    .C(_0566_),
    .Y(_0695_));
 sg13g2_nand2_1 _1671_ (.Y(_0696_),
    .A(net512),
    .B(net614));
 sg13g2_nand2_1 _1672_ (.Y(_0697_),
    .A(net614),
    .B(net487));
 sg13g2_and2_2 _1673_ (.A(net616),
    .B(net488),
    .X(_0698_));
 sg13g2_nand3_1 _1674_ (.B(_0524_),
    .C(net488),
    .A(net616),
    .Y(_0699_));
 sg13g2_a21oi_1 _1675_ (.A1(net613),
    .A2(_0535_),
    .Y(_0700_),
    .B1(net560));
 sg13g2_o21ai_1 _1676_ (.B1(_0700_),
    .Y(_0701_),
    .A1(_0691_),
    .A2(_0695_));
 sg13g2_nor2_1 _1677_ (.A(net574),
    .B(_0698_),
    .Y(_0702_));
 sg13g2_a21oi_2 _1678_ (.B1(net578),
    .Y(_0703_),
    .A2(net568),
    .A1(net536));
 sg13g2_nand4_1 _1679_ (.B(_0583_),
    .C(_0662_),
    .A(net566),
    .Y(_0704_),
    .D(_0699_));
 sg13g2_nand3_1 _1680_ (.B(_0701_),
    .C(_0704_),
    .A(_0689_),
    .Y(_0705_));
 sg13g2_a21o_1 _1681_ (.A2(_0705_),
    .A1(_0687_),
    .B1(net495),
    .X(_0706_));
 sg13g2_nor4_1 _1682_ (.A(_0546_),
    .B(net501),
    .C(net550),
    .D(_0691_),
    .Y(_0707_));
 sg13g2_nor2_2 _1683_ (.A(net509),
    .B(_0549_),
    .Y(_0708_));
 sg13g2_nand2_2 _1684_ (.Y(_0709_),
    .A(net508),
    .B(_0548_));
 sg13g2_o21ai_1 _1685_ (.B1(net602),
    .Y(_0710_),
    .A1(net510),
    .A2(_0549_));
 sg13g2_nand3_1 _1686_ (.B(_0535_),
    .C(net489),
    .A(net613),
    .Y(_0711_));
 sg13g2_nand3_1 _1687_ (.B(_0710_),
    .C(_0711_),
    .A(net578),
    .Y(_0712_));
 sg13g2_o21ai_1 _1688_ (.B1(_0692_),
    .Y(_0713_),
    .A1(net509),
    .A2(_0693_));
 sg13g2_nand2_2 _1689_ (.Y(_0714_),
    .A(net614),
    .B(net489));
 sg13g2_nand2_1 _1690_ (.Y(_0715_),
    .A(_0713_),
    .B(_0714_));
 sg13g2_a21oi_1 _1691_ (.A1(_0712_),
    .A2(_0715_),
    .Y(_0716_),
    .B1(net560));
 sg13g2_o21ai_1 _1692_ (.B1(net520),
    .Y(_0717_),
    .A1(_0707_),
    .A2(_0716_));
 sg13g2_a21oi_2 _1693_ (.B1(net606),
    .Y(_0718_),
    .A2(_0548_),
    .A1(net508));
 sg13g2_o21ai_1 _1694_ (.B1(net614),
    .Y(_0719_),
    .A1(net509),
    .A2(_0549_));
 sg13g2_o21ai_1 _1695_ (.B1(net587),
    .Y(_0720_),
    .A1(_0642_),
    .A2(_0718_));
 sg13g2_o21ai_1 _1696_ (.B1(_0708_),
    .Y(_0721_),
    .A1(net593),
    .A2(_0643_));
 sg13g2_nand2_2 _1697_ (.Y(_0722_),
    .A(net604),
    .B(_0527_));
 sg13g2_nor4_1 _1698_ (.A(_0553_),
    .B(_0564_),
    .C(_0585_),
    .D(_0594_),
    .Y(_0723_));
 sg13g2_nor2_2 _1699_ (.A(net577),
    .B(net559),
    .Y(_0724_));
 sg13g2_nand2_2 _1700_ (.Y(_0725_),
    .A(net590),
    .B(net548));
 sg13g2_a21oi_1 _1701_ (.A1(net512),
    .A2(_0586_),
    .Y(_0726_),
    .B1(_0608_));
 sg13g2_o21ai_1 _1702_ (.B1(net515),
    .Y(_0727_),
    .A1(_0725_),
    .A2(_0726_));
 sg13g2_a221oi_1 _1703_ (.B2(_0723_),
    .C1(_0727_),
    .B1(_0722_),
    .A1(net561),
    .Y(_0728_),
    .A2(_0721_));
 sg13g2_nor2_1 _1704_ (.A(net496),
    .B(_0728_),
    .Y(_0729_));
 sg13g2_a21oi_1 _1705_ (.A1(_0717_),
    .A2(_0729_),
    .Y(_0730_),
    .B1(net484));
 sg13g2_a21oi_1 _1706_ (.A1(_0706_),
    .A2(_0730_),
    .Y(_0731_),
    .B1(_0680_));
 sg13g2_xnor2_1 _1707_ (.Y(_0732_),
    .A(_0484_),
    .B(_0490_));
 sg13g2_xor2_1 _1708_ (.B(_0490_),
    .A(_0484_),
    .X(_0733_));
 sg13g2_a221oi_1 _1709_ (.B2(net490),
    .C1(net595),
    .B1(_0654_),
    .A1(_0619_),
    .Y(_0734_),
    .A2(_0641_));
 sg13g2_a21oi_1 _1710_ (.A1(net611),
    .A2(net499),
    .Y(_0735_),
    .B1(net583));
 sg13g2_nand3_1 _1711_ (.B(net577),
    .C(_0548_),
    .A(net508),
    .Y(_0736_));
 sg13g2_nand2_1 _1712_ (.Y(_0737_),
    .A(net608),
    .B(net505));
 sg13g2_nand3_1 _1713_ (.B(net505),
    .C(net502),
    .A(net609),
    .Y(_0738_));
 sg13g2_a22oi_1 _1714_ (.Y(_0739_),
    .B1(_0738_),
    .B2(_0663_),
    .A2(_0708_),
    .A1(net583));
 sg13g2_nor2_1 _1715_ (.A(net618),
    .B(_0553_),
    .Y(_0740_));
 sg13g2_nand2_1 _1716_ (.Y(_0741_),
    .A(net603),
    .B(net502));
 sg13g2_nand3_1 _1717_ (.B(_0524_),
    .C(_0586_),
    .A(net612),
    .Y(_0742_));
 sg13g2_a21oi_1 _1718_ (.A1(_0529_),
    .A2(net502),
    .Y(_0743_),
    .B1(net583));
 sg13g2_nor2_1 _1719_ (.A(net573),
    .B(_0613_),
    .Y(_0744_));
 sg13g2_nand3b_1 _1720_ (.B(_0699_),
    .C(net598),
    .Y(_0745_),
    .A_N(_0641_));
 sg13g2_or2_1 _1721_ (.X(_0746_),
    .B(_0720_),
    .A(_0665_));
 sg13g2_nor2_1 _1722_ (.A(net579),
    .B(_0553_),
    .Y(_0747_));
 sg13g2_a221oi_1 _1723_ (.B2(_0596_),
    .C1(net496),
    .B1(_0747_),
    .A1(net561),
    .Y(_0748_),
    .A2(_0721_));
 sg13g2_nand3_1 _1724_ (.B(_0657_),
    .C(_0659_),
    .A(net598),
    .Y(_0749_));
 sg13g2_nor2_2 _1725_ (.A(_0534_),
    .B(net594),
    .Y(_0750_));
 sg13g2_o21ai_1 _1726_ (.B1(_0595_),
    .Y(_0751_),
    .A1(_0582_),
    .A2(_0750_));
 sg13g2_nand3_1 _1727_ (.B(_0749_),
    .C(_0751_),
    .A(net563),
    .Y(_0752_));
 sg13g2_o21ai_1 _1728_ (.B1(net551),
    .Y(_0753_),
    .A1(_0547_),
    .A2(net491));
 sg13g2_a21oi_1 _1729_ (.A1(_0685_),
    .A2(_0696_),
    .Y(_0754_),
    .B1(_0753_));
 sg13g2_nor2_1 _1730_ (.A(net494),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_a22oi_1 _1731_ (.Y(_0756_),
    .B1(_0752_),
    .B2(_0755_),
    .A2(_0748_),
    .A1(_0746_));
 sg13g2_a21oi_1 _1732_ (.A1(net605),
    .A2(_0619_),
    .Y(_0757_),
    .B1(net595));
 sg13g2_o21ai_1 _1733_ (.B1(net503),
    .Y(_0758_),
    .A1(net570),
    .A2(_0603_));
 sg13g2_a21oi_1 _1734_ (.A1(net618),
    .A2(_0553_),
    .Y(_0759_),
    .B1(net584));
 sg13g2_nor2_2 _1735_ (.A(net606),
    .B(_0555_),
    .Y(_0760_));
 sg13g2_nand2_1 _1736_ (.Y(_0761_),
    .A(net613),
    .B(net501));
 sg13g2_nand2_1 _1737_ (.Y(_0762_),
    .A(_0610_),
    .B(_0760_));
 sg13g2_a221oi_1 _1738_ (.B2(_0610_),
    .C1(net585),
    .B1(_0760_),
    .A1(net605),
    .Y(_0763_),
    .A2(_0618_));
 sg13g2_nor4_1 _1739_ (.A(_0534_),
    .B(net595),
    .C(_0550_),
    .D(_0587_),
    .Y(_0764_));
 sg13g2_nor2_2 _1740_ (.A(net618),
    .B(_0525_),
    .Y(_0765_));
 sg13g2_a21oi_1 _1741_ (.A1(_0580_),
    .A2(_0740_),
    .Y(_0766_),
    .B1(net595));
 sg13g2_nand3_1 _1742_ (.B(net618),
    .C(net503),
    .A(net511),
    .Y(_0767_));
 sg13g2_nand2_1 _1743_ (.Y(_0768_),
    .A(_0587_),
    .B(_0709_));
 sg13g2_a21oi_1 _1744_ (.A1(net604),
    .A2(net489),
    .Y(_0769_),
    .B1(net580));
 sg13g2_o21ai_1 _1745_ (.B1(net591),
    .Y(_0770_),
    .A1(net613),
    .A2(_0613_));
 sg13g2_a21oi_1 _1746_ (.A1(_0587_),
    .A2(_0709_),
    .Y(_0771_),
    .B1(_0770_));
 sg13g2_nor2_1 _1747_ (.A(net597),
    .B(net489),
    .Y(_0772_));
 sg13g2_and2_1 _1748_ (.A(_0718_),
    .B(_0772_),
    .X(_0773_));
 sg13g2_a21oi_2 _1749_ (.B1(net591),
    .Y(_0774_),
    .A2(net608),
    .A1(net532));
 sg13g2_o21ai_1 _1750_ (.B1(net578),
    .Y(_0775_),
    .A1(net536),
    .A2(net603));
 sg13g2_a21oi_1 _1751_ (.A1(net603),
    .A2(net501),
    .Y(_0776_),
    .B1(_0775_));
 sg13g2_a22oi_1 _1752_ (.Y(_0777_),
    .B1(_0776_),
    .B2(_0655_),
    .A2(_0697_),
    .A1(_0685_));
 sg13g2_a21oi_1 _1753_ (.A1(_0710_),
    .A2(_0761_),
    .Y(_0778_),
    .B1(net592));
 sg13g2_a22oi_1 _1754_ (.Y(_0779_),
    .B1(_0719_),
    .B2(_0713_),
    .A2(_0714_),
    .A1(_0644_));
 sg13g2_nand4_1 _1755_ (.B(net505),
    .C(net580),
    .A(net613),
    .Y(_0780_),
    .D(net489));
 sg13g2_nor2_2 _1756_ (.A(net617),
    .B(_0601_),
    .Y(_0781_));
 sg13g2_a221oi_1 _1757_ (.B2(_0703_),
    .C1(net562),
    .B1(net489),
    .A1(_0546_),
    .Y(_0782_),
    .A2(net491));
 sg13g2_a21oi_1 _1758_ (.A1(_0780_),
    .A2(_0782_),
    .Y(_0783_),
    .B1(net494));
 sg13g2_o21ai_1 _1759_ (.B1(_0783_),
    .Y(_0784_),
    .A1(net551),
    .A2(_0777_));
 sg13g2_nor2_1 _1760_ (.A(net560),
    .B(_0779_),
    .Y(_0785_));
 sg13g2_nand2b_1 _1761_ (.Y(_0786_),
    .B(net562),
    .A_N(_0703_));
 sg13g2_o21ai_1 _1762_ (.B1(net494),
    .Y(_0787_),
    .A1(_0778_),
    .A2(_0786_));
 sg13g2_o21ai_1 _1763_ (.B1(_0784_),
    .Y(_0788_),
    .A1(_0785_),
    .A2(_0787_));
 sg13g2_a21oi_1 _1764_ (.A1(_0657_),
    .A2(_0735_),
    .Y(_0789_),
    .B1(net552));
 sg13g2_nand2b_1 _1765_ (.Y(_0790_),
    .B(_0789_),
    .A_N(_0734_));
 sg13g2_a221oi_1 _1766_ (.B2(_0624_),
    .C1(net557),
    .B1(_0744_),
    .A1(_0742_),
    .Y(_0791_),
    .A2(_0743_));
 sg13g2_nand3b_1 _1767_ (.B(net498),
    .C(_0790_),
    .Y(_0792_),
    .A_N(_0791_));
 sg13g2_a21oi_1 _1768_ (.A1(net587),
    .A2(_0557_),
    .Y(_0793_),
    .B1(net565));
 sg13g2_a221oi_1 _1769_ (.B2(_0793_),
    .C1(net497),
    .B1(_0745_),
    .A1(net565),
    .Y(_0794_),
    .A2(_0739_));
 sg13g2_nor2_1 _1770_ (.A(net521),
    .B(_0794_),
    .Y(_0795_));
 sg13g2_nor3_1 _1771_ (.A(net552),
    .B(_0763_),
    .C(_0764_),
    .Y(_0796_));
 sg13g2_nor3_1 _1772_ (.A(net565),
    .B(_0771_),
    .C(_0773_),
    .Y(_0797_));
 sg13g2_nor3_1 _1773_ (.A(net497),
    .B(_0796_),
    .C(_0797_),
    .Y(_0798_));
 sg13g2_a221oi_1 _1774_ (.B2(_0759_),
    .C1(net552),
    .B1(_0758_),
    .A1(_0661_),
    .Y(_0799_),
    .A2(_0757_));
 sg13g2_a221oi_1 _1775_ (.B2(_0767_),
    .C1(net566),
    .B1(_0766_),
    .A1(_0548_),
    .Y(_0800_),
    .A2(_0625_));
 sg13g2_nor3_1 _1776_ (.A(_0578_),
    .B(_0799_),
    .C(_0800_),
    .Y(_0801_));
 sg13g2_nor3_1 _1777_ (.A(net516),
    .B(_0798_),
    .C(_0801_),
    .Y(_0802_));
 sg13g2_a21oi_1 _1778_ (.A1(_0792_),
    .A2(_0795_),
    .Y(_0803_),
    .B1(net482));
 sg13g2_nand2b_1 _1779_ (.Y(_0804_),
    .B(_0803_),
    .A_N(_0802_));
 sg13g2_nand2_1 _1780_ (.Y(_0805_),
    .A(net515),
    .B(_0756_));
 sg13g2_a21oi_1 _1781_ (.A1(net520),
    .A2(_0788_),
    .Y(_0806_),
    .B1(net484));
 sg13g2_a21oi_1 _1782_ (.A1(_0805_),
    .A2(_0806_),
    .Y(_0807_),
    .B1(_0679_));
 sg13g2_a221oi_1 _1783_ (.B2(_0807_),
    .C1(_0733_),
    .B1(_0804_),
    .A1(_0677_),
    .Y(_0808_),
    .A2(_0731_));
 sg13g2_nand3_1 _1784_ (.B(net499),
    .C(net492),
    .A(net602),
    .Y(_0809_));
 sg13g2_a221oi_1 _1785_ (.B2(_0580_),
    .C1(net585),
    .B1(_0781_),
    .A1(_0610_),
    .Y(_0810_),
    .A2(_0760_));
 sg13g2_nand2_1 _1786_ (.Y(_0811_),
    .A(_0524_),
    .B(_0587_));
 sg13g2_a21oi_1 _1787_ (.A1(net504),
    .A2(_0646_),
    .Y(_0812_),
    .B1(net596));
 sg13g2_a21oi_1 _1788_ (.A1(_0811_),
    .A2(_0812_),
    .Y(_0813_),
    .B1(_0810_));
 sg13g2_nor2_1 _1789_ (.A(_0534_),
    .B(_0564_),
    .Y(_0814_));
 sg13g2_nand2_1 _1790_ (.Y(_0815_),
    .A(_0535_),
    .B(net500));
 sg13g2_nand3_1 _1791_ (.B(net507),
    .C(net589),
    .A(net611),
    .Y(_0816_));
 sg13g2_o21ai_1 _1792_ (.B1(_0814_),
    .Y(_0817_),
    .A1(_0655_),
    .A2(_0693_));
 sg13g2_nor3_1 _1793_ (.A(net583),
    .B(_0550_),
    .C(net493),
    .Y(_0818_));
 sg13g2_nor2_1 _1794_ (.A(net564),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_a21oi_1 _1795_ (.A1(_0817_),
    .A2(_0819_),
    .Y(_0820_),
    .B1(net497));
 sg13g2_o21ai_1 _1796_ (.B1(_0820_),
    .Y(_0821_),
    .A1(net552),
    .A2(_0813_));
 sg13g2_nor3_2 _1797_ (.A(net537),
    .B(net570),
    .C(net600),
    .Y(_0822_));
 sg13g2_o21ai_1 _1798_ (.B1(net508),
    .Y(_0823_),
    .A1(net504),
    .A2(_0822_));
 sg13g2_a21oi_1 _1799_ (.A1(net507),
    .A2(_0823_),
    .Y(_0824_),
    .B1(net598));
 sg13g2_a21oi_2 _1800_ (.B1(net574),
    .Y(_0825_),
    .A2(net600),
    .A1(net537));
 sg13g2_a21oi_1 _1801_ (.A1(net616),
    .A2(net486),
    .Y(_0826_),
    .B1(net587));
 sg13g2_and2_1 _1802_ (.A(_0643_),
    .B(_0826_),
    .X(_0827_));
 sg13g2_o21ai_1 _1803_ (.B1(net554),
    .Y(_0828_),
    .A1(_0824_),
    .A2(_0827_));
 sg13g2_nand2_1 _1804_ (.Y(_0829_),
    .A(_0525_),
    .B(_0537_));
 sg13g2_nor2_1 _1805_ (.A(net585),
    .B(_0555_),
    .Y(_0830_));
 sg13g2_a221oi_1 _1806_ (.B2(_0652_),
    .C1(net553),
    .B1(_0830_),
    .A1(_0605_),
    .Y(_0831_),
    .A2(_0829_));
 sg13g2_nor2_1 _1807_ (.A(_0578_),
    .B(_0831_),
    .Y(_0832_));
 sg13g2_a21oi_1 _1808_ (.A1(_0828_),
    .A2(_0832_),
    .Y(_0833_),
    .B1(net516));
 sg13g2_nor3_1 _1809_ (.A(net601),
    .B(_0532_),
    .C(_0550_),
    .Y(_0834_));
 sg13g2_nor2_1 _1810_ (.A(net595),
    .B(_0834_),
    .Y(_0835_));
 sg13g2_a21oi_1 _1811_ (.A1(net511),
    .A2(_0645_),
    .Y(_0836_),
    .B1(net611));
 sg13g2_nor3_1 _1812_ (.A(net595),
    .B(_0834_),
    .C(_0836_),
    .Y(_0837_));
 sg13g2_nor2_1 _1813_ (.A(_0527_),
    .B(net493),
    .Y(_0838_));
 sg13g2_nor3_1 _1814_ (.A(net600),
    .B(_0527_),
    .C(net493),
    .Y(_0839_));
 sg13g2_a21oi_1 _1815_ (.A1(net601),
    .A2(_0552_),
    .Y(_0840_),
    .B1(net584));
 sg13g2_a221oi_1 _1816_ (.B2(net505),
    .C1(net583),
    .B1(_0591_),
    .A1(net600),
    .Y(_0841_),
    .A2(_0552_));
 sg13g2_o21ai_1 _1817_ (.B1(net552),
    .Y(_0842_),
    .A1(_0837_),
    .A2(_0841_));
 sg13g2_nor2_2 _1818_ (.A(_0546_),
    .B(_0581_),
    .Y(_0843_));
 sg13g2_a21oi_1 _1819_ (.A1(_0619_),
    .A2(_0641_),
    .Y(_0844_),
    .B1(_0843_));
 sg13g2_o21ai_1 _1820_ (.B1(net566),
    .Y(_0845_),
    .A1(_0818_),
    .A2(_0844_));
 sg13g2_nand3_1 _1821_ (.B(_0842_),
    .C(_0845_),
    .A(net496),
    .Y(_0846_));
 sg13g2_nor2_1 _1822_ (.A(net598),
    .B(net487),
    .Y(_0847_));
 sg13g2_nor2_1 _1823_ (.A(net579),
    .B(_0822_),
    .Y(_0848_));
 sg13g2_nand2b_1 _1824_ (.Y(_0849_),
    .B(net598),
    .A_N(_0822_));
 sg13g2_a21oi_1 _1825_ (.A1(net616),
    .A2(_0645_),
    .Y(_0850_),
    .B1(_0849_));
 sg13g2_nor2_1 _1826_ (.A(net554),
    .B(_0642_),
    .Y(_0851_));
 sg13g2_o21ai_1 _1827_ (.B1(_0851_),
    .Y(_0852_),
    .A1(_0847_),
    .A2(_0850_));
 sg13g2_nand2_2 _1828_ (.Y(_0853_),
    .A(net509),
    .B(_0532_));
 sg13g2_mux2_1 _1829_ (.A0(_0533_),
    .A1(_0549_),
    .S(net508),
    .X(_0854_));
 sg13g2_nor2_1 _1830_ (.A(_0698_),
    .B(_0854_),
    .Y(_0855_));
 sg13g2_nor3_1 _1831_ (.A(net534),
    .B(_0603_),
    .C(_0611_),
    .Y(_0856_));
 sg13g2_a221oi_1 _1832_ (.B2(_0724_),
    .C1(net498),
    .B1(_0856_),
    .A1(_0593_),
    .Y(_0857_),
    .A2(_0855_));
 sg13g2_a21oi_1 _1833_ (.A1(_0852_),
    .A2(_0857_),
    .Y(_0858_),
    .B1(net521));
 sg13g2_a221oi_1 _1834_ (.B2(_0858_),
    .C1(net482),
    .B1(_0846_),
    .A1(_0821_),
    .Y(_0859_),
    .A2(_0833_));
 sg13g2_and2_1 _1835_ (.A(_0625_),
    .B(net488),
    .X(_0860_));
 sg13g2_a22oi_1 _1836_ (.Y(_0861_),
    .B1(_0602_),
    .B2(net618),
    .A2(_0586_),
    .A1(net511));
 sg13g2_a221oi_1 _1837_ (.B2(net583),
    .C1(net552),
    .B1(_0861_),
    .A1(_0690_),
    .Y(_0862_),
    .A2(_0860_));
 sg13g2_nand2_1 _1838_ (.Y(_0863_),
    .A(_0591_),
    .B(net485));
 sg13g2_a221oi_1 _1839_ (.B2(_0863_),
    .C1(net562),
    .B1(_0685_),
    .A1(_0523_),
    .Y(_0864_),
    .A2(_0532_));
 sg13g2_o21ai_1 _1840_ (.B1(net496),
    .Y(_0865_),
    .A1(_0862_),
    .A2(_0864_));
 sg13g2_nand2_1 _1841_ (.Y(_0866_),
    .A(net507),
    .B(_0606_));
 sg13g2_nand3_1 _1842_ (.B(_0586_),
    .C(_0604_),
    .A(net502),
    .Y(_0867_));
 sg13g2_o21ai_1 _1843_ (.B1(net593),
    .Y(_0868_),
    .A1(_0647_),
    .A2(_0867_));
 sg13g2_nand3_1 _1844_ (.B(_0866_),
    .C(_0868_),
    .A(net561),
    .Y(_0869_));
 sg13g2_nand3b_1 _1845_ (.B(net593),
    .C(net491),
    .Y(_0870_),
    .A_N(_0665_));
 sg13g2_and3_1 _1846_ (.X(_0871_),
    .A(net550),
    .B(_0639_),
    .C(_0870_));
 sg13g2_nor2_1 _1847_ (.A(net496),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_a21oi_1 _1848_ (.A1(_0869_),
    .A2(_0872_),
    .Y(_0873_),
    .B1(net520));
 sg13g2_o21ai_1 _1849_ (.B1(net578),
    .Y(_0874_),
    .A1(net603),
    .A2(_0615_));
 sg13g2_a21oi_1 _1850_ (.A1(net603),
    .A2(_0535_),
    .Y(_0875_),
    .B1(_0874_));
 sg13g2_o21ai_1 _1851_ (.B1(net551),
    .Y(_0876_),
    .A1(_0694_),
    .A2(_0875_));
 sg13g2_nand3_1 _1852_ (.B(_0691_),
    .C(_0708_),
    .A(net560),
    .Y(_0877_));
 sg13g2_nand3_1 _1853_ (.B(_0876_),
    .C(_0877_),
    .A(net496),
    .Y(_0878_));
 sg13g2_a21oi_1 _1854_ (.A1(net614),
    .A2(net508),
    .Y(_0879_),
    .B1(net511));
 sg13g2_nand3_1 _1855_ (.B(_0770_),
    .C(_0879_),
    .A(net560),
    .Y(_0880_));
 sg13g2_o21ai_1 _1856_ (.B1(net551),
    .Y(_0881_),
    .A1(net579),
    .A2(_0822_));
 sg13g2_a21oi_1 _1857_ (.A1(_0722_),
    .A2(_0750_),
    .Y(_0882_),
    .B1(_0881_));
 sg13g2_o21ai_1 _1858_ (.B1(net494),
    .Y(_0883_),
    .A1(net560),
    .A2(_0634_));
 sg13g2_nor2_1 _1859_ (.A(_0882_),
    .B(_0883_),
    .Y(_0884_));
 sg13g2_a21oi_1 _1860_ (.A1(_0880_),
    .A2(_0884_),
    .Y(_0885_),
    .B1(net514));
 sg13g2_a221oi_1 _1861_ (.B2(_0885_),
    .C1(net484),
    .B1(_0878_),
    .A1(_0865_),
    .Y(_0886_),
    .A2(_0873_));
 sg13g2_or3_1 _1862_ (.A(_0679_),
    .B(_0859_),
    .C(_0886_),
    .X(_0887_));
 sg13g2_nand2b_1 _1863_ (.Y(_0888_),
    .B(net499),
    .A_N(_0710_));
 sg13g2_a21oi_1 _1864_ (.A1(_0533_),
    .A2(_0587_),
    .Y(_0889_),
    .B1(net599));
 sg13g2_a221oi_1 _1865_ (.B2(_0889_),
    .C1(net555),
    .B1(_0888_),
    .A1(_0685_),
    .Y(_0890_),
    .A2(_0762_));
 sg13g2_o21ai_1 _1866_ (.B1(net574),
    .Y(_0891_),
    .A1(net533),
    .A2(net600));
 sg13g2_o21ai_1 _1867_ (.B1(net548),
    .Y(_0892_),
    .A1(_0535_),
    .A2(_0891_));
 sg13g2_a21oi_1 _1868_ (.A1(_0657_),
    .A2(_0702_),
    .Y(_0893_),
    .B1(_0892_));
 sg13g2_o21ai_1 _1869_ (.B1(net519),
    .Y(_0894_),
    .A1(_0890_),
    .A2(_0893_));
 sg13g2_a21o_1 _1870_ (.A2(_0738_),
    .A1(_0710_),
    .B1(net583),
    .X(_0895_));
 sg13g2_nand3_1 _1871_ (.B(_0720_),
    .C(_0895_),
    .A(net557),
    .Y(_0896_));
 sg13g2_o21ai_1 _1872_ (.B1(net547),
    .Y(_0897_),
    .A1(net611),
    .A2(_0601_));
 sg13g2_o21ai_1 _1873_ (.B1(_0594_),
    .Y(_0898_),
    .A1(_0839_),
    .A2(_0897_));
 sg13g2_o21ai_1 _1874_ (.B1(net574),
    .Y(_0899_),
    .A1(_0698_),
    .A2(_0854_));
 sg13g2_a21oi_1 _1875_ (.A1(_0898_),
    .A2(_0899_),
    .Y(_0900_),
    .B1(net519));
 sg13g2_a21oi_1 _1876_ (.A1(_0896_),
    .A2(_0900_),
    .Y(_0901_),
    .B1(net498));
 sg13g2_and2_1 _1877_ (.A(_0815_),
    .B(_0825_),
    .X(_0902_));
 sg13g2_or3_1 _1878_ (.A(_0773_),
    .B(_0844_),
    .C(_0902_),
    .X(_0903_));
 sg13g2_nor2_1 _1879_ (.A(net590),
    .B(_0555_),
    .Y(_0904_));
 sg13g2_nand2_1 _1880_ (.Y(_0905_),
    .A(net584),
    .B(_0556_));
 sg13g2_nor2_1 _1881_ (.A(_0548_),
    .B(_0589_),
    .Y(_0906_));
 sg13g2_nand2b_1 _1882_ (.Y(_0907_),
    .B(_0904_),
    .A_N(_0906_));
 sg13g2_a221oi_1 _1883_ (.B2(_0898_),
    .C1(net519),
    .B1(_0907_),
    .A1(net558),
    .Y(_0908_),
    .A2(_0903_));
 sg13g2_nand2_1 _1884_ (.Y(_0909_),
    .A(net511),
    .B(_0615_));
 sg13g2_a221oi_1 _1885_ (.B2(_0735_),
    .C1(net564),
    .B1(_0888_),
    .A1(_0766_),
    .Y(_0910_),
    .A2(_0768_));
 sg13g2_o21ai_1 _1886_ (.B1(_0619_),
    .Y(_0911_),
    .A1(net600),
    .A2(net492));
 sg13g2_a21oi_2 _1887_ (.B1(net574),
    .Y(_0912_),
    .A2(net611),
    .A1(_0503_));
 sg13g2_nor2_1 _1888_ (.A(net533),
    .B(_0612_),
    .Y(_0913_));
 sg13g2_a221oi_1 _1889_ (.B2(_0913_),
    .C1(net548),
    .B1(_0912_),
    .A1(net584),
    .Y(_0914_),
    .A2(_0911_));
 sg13g2_o21ai_1 _1890_ (.B1(net518),
    .Y(_0915_),
    .A1(_0910_),
    .A2(_0914_));
 sg13g2_nand3b_1 _1891_ (.B(_0915_),
    .C(net498),
    .Y(_0916_),
    .A_N(_0908_));
 sg13g2_a21oi_1 _1892_ (.A1(_0894_),
    .A2(_0901_),
    .Y(_0917_),
    .B1(net482));
 sg13g2_nand3_1 _1893_ (.B(net487),
    .C(net486),
    .A(net617),
    .Y(_0918_));
 sg13g2_a21oi_1 _1894_ (.A1(_0685_),
    .A2(_0918_),
    .Y(_0919_),
    .B1(_0753_));
 sg13g2_nor2_1 _1895_ (.A(_0538_),
    .B(net591),
    .Y(_0920_));
 sg13g2_nand3_1 _1896_ (.B(_0657_),
    .C(_0848_),
    .A(_0589_),
    .Y(_0921_));
 sg13g2_a21oi_1 _1897_ (.A1(_0623_),
    .A2(_0920_),
    .Y(_0922_),
    .B1(net551));
 sg13g2_a21o_1 _1898_ (.A2(_0922_),
    .A1(_0921_),
    .B1(_0919_),
    .X(_0923_));
 sg13g2_o21ai_1 _1899_ (.B1(_0713_),
    .Y(_0924_),
    .A1(_0527_),
    .A2(_0714_));
 sg13g2_nand3_1 _1900_ (.B(_0711_),
    .C(_0741_),
    .A(net578),
    .Y(_0925_));
 sg13g2_a21o_1 _1901_ (.A2(_0925_),
    .A1(_0924_),
    .B1(net562),
    .X(_0926_));
 sg13g2_o21ai_1 _1902_ (.B1(net562),
    .Y(_0927_),
    .A1(_0546_),
    .A2(_0691_));
 sg13g2_nor3_1 _1903_ (.A(_0529_),
    .B(_0591_),
    .C(_0927_),
    .Y(_0928_));
 sg13g2_nor2_1 _1904_ (.A(net514),
    .B(_0928_),
    .Y(_0929_));
 sg13g2_a221oi_1 _1905_ (.B2(_0929_),
    .C1(net495),
    .B1(_0926_),
    .A1(net514),
    .Y(_0930_),
    .A2(_0923_));
 sg13g2_nand3_1 _1906_ (.B(net502),
    .C(net485),
    .A(net608),
    .Y(_0931_));
 sg13g2_and3_1 _1907_ (.X(_0932_),
    .A(_0724_),
    .B(_0809_),
    .C(_0931_));
 sg13g2_nand2_1 _1908_ (.Y(_0933_),
    .A(_0504_),
    .B(_0593_));
 sg13g2_a21oi_1 _1909_ (.A1(_0809_),
    .A2(_0931_),
    .Y(_0934_),
    .B1(_0933_));
 sg13g2_nor2_1 _1910_ (.A(net493),
    .B(_0692_),
    .Y(_0935_));
 sg13g2_nor3_1 _1911_ (.A(net502),
    .B(net549),
    .C(_0935_),
    .Y(_0936_));
 sg13g2_nor4_1 _1912_ (.A(net518),
    .B(_0932_),
    .C(_0934_),
    .D(_0936_),
    .Y(_0937_));
 sg13g2_a221oi_1 _1913_ (.B2(_0909_),
    .C1(net562),
    .B1(_0692_),
    .A1(net591),
    .Y(_0938_),
    .A2(_0591_));
 sg13g2_nand3_1 _1914_ (.B(net559),
    .C(_0691_),
    .A(_0555_),
    .Y(_0939_));
 sg13g2_nand3_1 _1915_ (.B(net493),
    .C(_0774_),
    .A(net559),
    .Y(_0940_));
 sg13g2_nand3_1 _1916_ (.B(_0939_),
    .C(_0940_),
    .A(net518),
    .Y(_0941_));
 sg13g2_o21ai_1 _1917_ (.B1(net495),
    .Y(_0942_),
    .A1(_0938_),
    .A2(_0941_));
 sg13g2_o21ai_1 _1918_ (.B1(net482),
    .Y(_0943_),
    .A1(_0937_),
    .A2(_0942_));
 sg13g2_o21ai_1 _1919_ (.B1(_0679_),
    .Y(_0944_),
    .A1(_0930_),
    .A2(_0943_));
 sg13g2_a21o_1 _1920_ (.A2(_0917_),
    .A1(_0916_),
    .B1(_0944_),
    .X(_0945_));
 sg13g2_nand3_1 _1921_ (.B(net506),
    .C(_0533_),
    .A(net612),
    .Y(_0946_));
 sg13g2_a21oi_1 _1922_ (.A1(_0887_),
    .A2(_0945_),
    .Y(_0947_),
    .B1(_0732_));
 sg13g2_a21oi_1 _1923_ (.A1(_0485_),
    .A2(_0490_),
    .Y(_0948_),
    .B1(_0489_));
 sg13g2_xor2_1 _1924_ (.B(_0948_),
    .A(_0488_),
    .X(_0949_));
 sg13g2_nor3_2 _1925_ (.A(_0808_),
    .B(_0947_),
    .C(_0949_),
    .Y(_0950_));
 sg13g2_nand3_1 _1926_ (.B(net506),
    .C(net492),
    .A(net601),
    .Y(_0951_));
 sg13g2_nand3_1 _1927_ (.B(_0946_),
    .C(_0951_),
    .A(net589),
    .Y(_0952_));
 sg13g2_nand3_1 _1928_ (.B(net491),
    .C(net485),
    .A(net604),
    .Y(_0953_));
 sg13g2_nand4_1 _1929_ (.B(net506),
    .C(net499),
    .A(net609),
    .Y(_0954_),
    .D(net492));
 sg13g2_nand3_1 _1930_ (.B(_0953_),
    .C(_0954_),
    .A(net577),
    .Y(_0955_));
 sg13g2_a21oi_1 _1931_ (.A1(_0952_),
    .A2(_0955_),
    .Y(_0956_),
    .B1(net557));
 sg13g2_o21ai_1 _1932_ (.B1(_0825_),
    .Y(_0957_),
    .A1(net511),
    .A2(net508));
 sg13g2_o21ai_1 _1933_ (.B1(_0957_),
    .Y(_0958_),
    .A1(net589),
    .A2(_0622_));
 sg13g2_o21ai_1 _1934_ (.B1(net513),
    .Y(_0959_),
    .A1(net549),
    .A2(_0958_));
 sg13g2_nor4_1 _1935_ (.A(net504),
    .B(net559),
    .C(_0603_),
    .D(_0843_),
    .Y(_0960_));
 sg13g2_nand2_1 _1936_ (.Y(_0961_),
    .A(_0569_),
    .B(_0692_));
 sg13g2_and3_1 _1937_ (.X(_0962_),
    .A(net506),
    .B(net490),
    .C(_0961_));
 sg13g2_a221oi_1 _1938_ (.B2(net610),
    .C1(net589),
    .B1(_0549_),
    .A1(net524),
    .Y(_0963_),
    .A2(net523));
 sg13g2_nor3_1 _1939_ (.A(net549),
    .B(_0962_),
    .C(_0963_),
    .Y(_0964_));
 sg13g2_a22oi_1 _1940_ (.Y(_0965_),
    .B1(_0604_),
    .B2(net569),
    .A2(_0589_),
    .A1(net531));
 sg13g2_o21ai_1 _1941_ (.B1(net518),
    .Y(_0966_),
    .A1(_0725_),
    .A2(_0965_));
 sg13g2_or3_1 _1942_ (.A(_0960_),
    .B(_0964_),
    .C(_0966_),
    .X(_0967_));
 sg13g2_o21ai_1 _1943_ (.B1(_0770_),
    .Y(_0968_),
    .A1(net578),
    .A2(_0853_));
 sg13g2_o21ai_1 _1944_ (.B1(net562),
    .Y(_0969_),
    .A1(_0641_),
    .A2(_0874_));
 sg13g2_a21o_1 _1945_ (.A2(_0968_),
    .A1(_0711_),
    .B1(_0969_),
    .X(_0970_));
 sg13g2_nor2_1 _1946_ (.A(_0613_),
    .B(_0693_),
    .Y(_0971_));
 sg13g2_or2_1 _1947_ (.X(_0972_),
    .B(_0615_),
    .A(net613));
 sg13g2_nor3_1 _1948_ (.A(net608),
    .B(net577),
    .C(_0615_),
    .Y(_0973_));
 sg13g2_o21ai_1 _1949_ (.B1(net549),
    .Y(_0974_),
    .A1(_0971_),
    .A2(_0973_));
 sg13g2_o21ai_1 _1950_ (.B1(_0593_),
    .Y(_0975_),
    .A1(_0529_),
    .A2(_0591_));
 sg13g2_and3_1 _1951_ (.X(_0976_),
    .A(net518),
    .B(_0974_),
    .C(_0975_));
 sg13g2_a22oi_1 _1952_ (.Y(_0977_),
    .B1(_0724_),
    .B2(_0550_),
    .A2(_0665_),
    .A1(_0593_));
 sg13g2_nor2_1 _1953_ (.A(_0912_),
    .B(_0977_),
    .Y(_0978_));
 sg13g2_o21ai_1 _1954_ (.B1(_0556_),
    .Y(_0979_),
    .A1(net504),
    .A2(_0603_));
 sg13g2_nand3_1 _1955_ (.B(net492),
    .C(net485),
    .A(net612),
    .Y(_0980_));
 sg13g2_a21oi_1 _1956_ (.A1(_0979_),
    .A2(_0980_),
    .Y(_0981_),
    .B1(net575));
 sg13g2_and2_1 _1957_ (.A(net575),
    .B(_0597_),
    .X(_0982_));
 sg13g2_nor3_1 _1958_ (.A(net547),
    .B(_0981_),
    .C(_0982_),
    .Y(_0983_));
 sg13g2_o21ai_1 _1959_ (.B1(net517),
    .Y(_0984_),
    .A1(_0978_),
    .A2(_0983_));
 sg13g2_a21oi_1 _1960_ (.A1(_0970_),
    .A2(_0976_),
    .Y(_0985_),
    .B1(net483));
 sg13g2_o21ai_1 _1961_ (.B1(_0967_),
    .Y(_0986_),
    .A1(_0956_),
    .A2(_0959_));
 sg13g2_a221oi_1 _1962_ (.B2(net483),
    .C1(net495),
    .B1(_0986_),
    .A1(_0984_),
    .Y(_0987_),
    .A2(_0985_));
 sg13g2_nand3_1 _1963_ (.B(_0531_),
    .C(net489),
    .A(net617),
    .Y(_0988_));
 sg13g2_o21ai_1 _1964_ (.B1(_0988_),
    .Y(_0989_),
    .A1(_0624_),
    .A2(_0772_));
 sg13g2_a221oi_1 _1965_ (.B2(net486),
    .C1(net586),
    .B1(_0642_),
    .A1(net617),
    .Y(_0990_),
    .A2(net507));
 sg13g2_nand3b_1 _1966_ (.B(net565),
    .C(_0989_),
    .Y(_0991_),
    .A_N(_0990_));
 sg13g2_nand3_1 _1967_ (.B(net605),
    .C(net490),
    .A(net573),
    .Y(_0992_));
 sg13g2_o21ai_1 _1968_ (.B1(_0992_),
    .Y(_0993_),
    .A1(_0550_),
    .A2(_0690_));
 sg13g2_o21ai_1 _1969_ (.B1(net511),
    .Y(_0994_),
    .A1(_0613_),
    .A2(_0655_));
 sg13g2_a221oi_1 _1970_ (.B2(_0724_),
    .C1(net518),
    .B1(_0994_),
    .A1(_0593_),
    .Y(_0995_),
    .A2(_0993_));
 sg13g2_o21ai_1 _1971_ (.B1(_0953_),
    .Y(_0996_),
    .A1(net604),
    .A2(_0647_));
 sg13g2_a21oi_1 _1972_ (.A1(_0584_),
    .A2(_0588_),
    .Y(_0997_),
    .B1(net550));
 sg13g2_o21ai_1 _1973_ (.B1(_0997_),
    .Y(_0998_),
    .A1(net581),
    .A2(_0996_));
 sg13g2_o21ai_1 _1974_ (.B1(_0953_),
    .Y(_0999_),
    .A1(_0647_),
    .A2(_0761_));
 sg13g2_and2_1 _1975_ (.A(_0596_),
    .B(_0703_),
    .X(_1000_));
 sg13g2_a221oi_1 _1976_ (.B2(net551),
    .C1(net514),
    .B1(_1000_),
    .A1(_0593_),
    .Y(_1001_),
    .A2(_0999_));
 sg13g2_a221oi_1 _1977_ (.B2(_1001_),
    .C1(net482),
    .B1(_0998_),
    .A1(_0991_),
    .Y(_1002_),
    .A2(_0995_));
 sg13g2_o21ai_1 _1978_ (.B1(_0551_),
    .Y(_1003_),
    .A1(net611),
    .A2(net492));
 sg13g2_nand2_1 _1979_ (.Y(_1004_),
    .A(net590),
    .B(_1003_));
 sg13g2_nor2_1 _1980_ (.A(_0564_),
    .B(_0822_),
    .Y(_1005_));
 sg13g2_mux2_1 _1981_ (.A0(_0531_),
    .A1(net533),
    .S(_0589_),
    .X(_1006_));
 sg13g2_o21ai_1 _1982_ (.B1(_0774_),
    .Y(_1007_),
    .A1(_0525_),
    .A2(_0532_));
 sg13g2_o21ai_1 _1983_ (.B1(net574),
    .Y(_1008_),
    .A1(_0552_),
    .A2(net557));
 sg13g2_a221oi_1 _1984_ (.B2(_0838_),
    .C1(net513),
    .B1(_0724_),
    .A1(_0533_),
    .Y(_1009_),
    .A2(net557));
 sg13g2_o21ai_1 _1985_ (.B1(_1007_),
    .Y(_1010_),
    .A1(net575),
    .A2(_1006_));
 sg13g2_a21oi_1 _1986_ (.A1(_0904_),
    .A2(_1005_),
    .Y(_1011_),
    .B1(net547));
 sg13g2_a221oi_1 _1987_ (.B2(_1004_),
    .C1(net518),
    .B1(_1011_),
    .A1(net547),
    .Y(_1012_),
    .A2(_1010_));
 sg13g2_a21o_1 _1988_ (.A2(_1009_),
    .A1(_1008_),
    .B1(net483),
    .X(_1013_));
 sg13g2_o21ai_1 _1989_ (.B1(net495),
    .Y(_1014_),
    .A1(_1012_),
    .A2(_1013_));
 sg13g2_o21ai_1 _1990_ (.B1(_0679_),
    .Y(_1015_),
    .A1(_1002_),
    .A2(_1014_));
 sg13g2_o21ai_1 _1991_ (.B1(net564),
    .Y(_1016_),
    .A1(_0524_),
    .A2(_0547_));
 sg13g2_a21o_1 _1992_ (.A2(_0685_),
    .A1(_0655_),
    .B1(_1016_),
    .X(_1017_));
 sg13g2_a21oi_1 _1993_ (.A1(net612),
    .A2(_0553_),
    .Y(_1018_),
    .B1(_0530_));
 sg13g2_a22oi_1 _1994_ (.Y(_1019_),
    .B1(_1018_),
    .B2(_0750_),
    .A2(_0912_),
    .A1(_0539_));
 sg13g2_o21ai_1 _1995_ (.B1(_1017_),
    .Y(_1020_),
    .A1(net564),
    .A2(_1019_));
 sg13g2_nor2b_1 _1996_ (.A(_0836_),
    .B_N(_0637_),
    .Y(_1021_));
 sg13g2_o21ai_1 _1997_ (.B1(net564),
    .Y(_1022_),
    .A1(_0581_),
    .A2(_1021_));
 sg13g2_nor2_1 _1998_ (.A(_0594_),
    .B(_0603_),
    .Y(_1023_));
 sg13g2_o21ai_1 _1999_ (.B1(net506),
    .Y(_1024_),
    .A1(net510),
    .A2(_0549_));
 sg13g2_a221oi_1 _2000_ (.B2(_0724_),
    .C1(net513),
    .B1(_1024_),
    .A1(_0954_),
    .Y(_1025_),
    .A2(_1023_));
 sg13g2_a221oi_1 _2001_ (.B2(_1025_),
    .C1(net498),
    .B1(_1022_),
    .A1(net513),
    .Y(_1026_),
    .A2(_1020_));
 sg13g2_a221oi_1 _2002_ (.B2(_0946_),
    .C1(net557),
    .B1(_0840_),
    .A1(_0624_),
    .Y(_1027_),
    .A2(_0660_));
 sg13g2_and4_1 _2003_ (.A(net533),
    .B(net506),
    .C(_0586_),
    .D(_0589_),
    .X(_1028_));
 sg13g2_o21ai_1 _2004_ (.B1(net575),
    .Y(_1029_),
    .A1(_0906_),
    .A2(_1028_));
 sg13g2_a22oi_1 _2005_ (.Y(_1030_),
    .B1(_0825_),
    .B2(net570),
    .A2(net590),
    .A1(net508));
 sg13g2_a21oi_1 _2006_ (.A1(_1029_),
    .A2(_1030_),
    .Y(_1031_),
    .B1(net547));
 sg13g2_o21ai_1 _2007_ (.B1(net513),
    .Y(_1032_),
    .A1(_1027_),
    .A2(_1031_));
 sg13g2_nor4_1 _2008_ (.A(net504),
    .B(net557),
    .C(_0603_),
    .D(_0654_),
    .Y(_1033_));
 sg13g2_o21ai_1 _2009_ (.B1(_0703_),
    .Y(_1034_),
    .A1(_0596_),
    .A2(_0603_));
 sg13g2_o21ai_1 _2010_ (.B1(_1034_),
    .Y(_1035_),
    .A1(_0724_),
    .A2(_1033_));
 sg13g2_o21ai_1 _2011_ (.B1(_0569_),
    .Y(_1036_),
    .A1(_0550_),
    .A2(_0891_));
 sg13g2_nand3_1 _2012_ (.B(net490),
    .C(_1036_),
    .A(_0535_),
    .Y(_1037_));
 sg13g2_a21oi_1 _2013_ (.A1(net557),
    .A2(_1037_),
    .Y(_1038_),
    .B1(net517));
 sg13g2_a21oi_1 _2014_ (.A1(_1035_),
    .A2(_1038_),
    .Y(_1039_),
    .B1(net495));
 sg13g2_a21o_1 _2015_ (.A2(_1039_),
    .A1(_1032_),
    .B1(_1026_),
    .X(_1040_));
 sg13g2_nor3_1 _2016_ (.A(net577),
    .B(_0567_),
    .C(_0698_),
    .Y(_1041_));
 sg13g2_a221oi_1 _2017_ (.B2(_0529_),
    .C1(net589),
    .B1(net492),
    .A1(net610),
    .Y(_1042_),
    .A2(_0586_));
 sg13g2_o21ai_1 _2018_ (.B1(net549),
    .Y(_1043_),
    .A1(_1041_),
    .A2(_1042_));
 sg13g2_nand2b_1 _2019_ (.Y(_1044_),
    .B(_0615_),
    .A_N(net504));
 sg13g2_a221oi_1 _2020_ (.B2(net577),
    .C1(net549),
    .B1(_1044_),
    .A1(_0737_),
    .Y(_1045_),
    .A2(_0971_));
 sg13g2_nor2_1 _2021_ (.A(net513),
    .B(_1045_),
    .Y(_1046_));
 sg13g2_nor3_1 _2022_ (.A(net572),
    .B(net611),
    .C(net574),
    .Y(_1047_));
 sg13g2_a21oi_1 _2023_ (.A1(net571),
    .A2(net510),
    .Y(_1048_),
    .B1(_0691_));
 sg13g2_a221oi_1 _2024_ (.B2(_1048_),
    .C1(net549),
    .B1(_0736_),
    .A1(net589),
    .Y(_1049_),
    .A2(_0654_));
 sg13g2_o21ai_1 _2025_ (.B1(net513),
    .Y(_1050_),
    .A1(_0977_),
    .A2(_1047_));
 sg13g2_o21ai_1 _2026_ (.B1(net498),
    .Y(_1051_),
    .A1(_1049_),
    .A2(_1050_));
 sg13g2_a21o_1 _2027_ (.A2(_1046_),
    .A1(_1043_),
    .B1(_1051_),
    .X(_1052_));
 sg13g2_nand4_1 _2028_ (.B(_0710_),
    .C(_0742_),
    .A(net547),
    .Y(_1053_),
    .D(_0905_));
 sg13g2_nand4_1 _2029_ (.B(net558),
    .C(_0612_),
    .A(net537),
    .Y(_1054_),
    .D(_0816_));
 sg13g2_nand3_1 _2030_ (.B(_1053_),
    .C(_1054_),
    .A(net519),
    .Y(_1055_));
 sg13g2_a21oi_2 _2031_ (.B1(net578),
    .Y(_1056_),
    .A2(_0535_),
    .A1(net608));
 sg13g2_nand2_1 _2032_ (.Y(_1057_),
    .A(net502),
    .B(_0609_));
 sg13g2_a22oi_1 _2033_ (.Y(_1058_),
    .B1(_1056_),
    .B2(_1057_),
    .A2(_0738_),
    .A1(net579));
 sg13g2_o21ai_1 _2034_ (.B1(net559),
    .Y(_1059_),
    .A1(_0547_),
    .A2(_1024_));
 sg13g2_nor2_1 _2035_ (.A(net570),
    .B(_0546_),
    .Y(_1060_));
 sg13g2_o21ai_1 _2036_ (.B1(_1060_),
    .Y(_1061_),
    .A1(_0553_),
    .A2(_0564_));
 sg13g2_a21oi_1 _2037_ (.A1(_0527_),
    .A2(net579),
    .Y(_1062_),
    .B1(net559));
 sg13g2_a21oi_1 _2038_ (.A1(_1061_),
    .A2(_1062_),
    .Y(_1063_),
    .B1(net518));
 sg13g2_o21ai_1 _2039_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_1058_),
    .A2(_1059_));
 sg13g2_nand3_1 _2040_ (.B(_1055_),
    .C(_1064_),
    .A(net495),
    .Y(_1065_));
 sg13g2_a21oi_1 _2041_ (.A1(_1052_),
    .A2(_1065_),
    .Y(_1066_),
    .B1(net483));
 sg13g2_a221oi_1 _2042_ (.B2(net483),
    .C1(_1066_),
    .B1(_1040_),
    .A1(_0483_),
    .Y(_1067_),
    .A2(_0678_));
 sg13g2_o21ai_1 _2043_ (.B1(_0733_),
    .Y(_1068_),
    .A1(_0987_),
    .A2(_1015_));
 sg13g2_nand2_1 _2044_ (.Y(_1069_),
    .A(net507),
    .B(_0551_));
 sg13g2_a21oi_1 _2045_ (.A1(_0765_),
    .A2(_0815_),
    .Y(_1070_),
    .B1(net596));
 sg13g2_a221oi_1 _2046_ (.B2(_0815_),
    .C1(net598),
    .B1(_0765_),
    .A1(_0646_),
    .Y(_1071_),
    .A2(_0718_));
 sg13g2_o21ai_1 _2047_ (.B1(_0637_),
    .Y(_1072_),
    .A1(net618),
    .A2(_0566_));
 sg13g2_nand3b_1 _2048_ (.B(_1072_),
    .C(net565),
    .Y(_1073_),
    .A_N(_1071_));
 sg13g2_a21oi_1 _2049_ (.A1(net509),
    .A2(_0531_),
    .Y(_1074_),
    .B1(net564));
 sg13g2_o21ai_1 _2050_ (.B1(_1074_),
    .Y(_1075_),
    .A1(_0582_),
    .A2(_1056_));
 sg13g2_nand3_1 _2051_ (.B(_0533_),
    .C(net485),
    .A(net601),
    .Y(_1076_));
 sg13g2_or2_1 _2052_ (.X(_1077_),
    .B(_1076_),
    .A(_0594_));
 sg13g2_nand4_1 _2053_ (.B(_1073_),
    .C(_1075_),
    .A(net483),
    .Y(_1078_),
    .D(_1077_));
 sg13g2_a21oi_1 _2054_ (.A1(_0547_),
    .A2(_0905_),
    .Y(_1079_),
    .B1(_0504_));
 sg13g2_nor3_1 _2055_ (.A(net548),
    .B(_0981_),
    .C(_1079_),
    .Y(_1080_));
 sg13g2_a221oi_1 _2056_ (.B2(net505),
    .C1(_0725_),
    .B1(_0698_),
    .A1(net601),
    .Y(_1081_),
    .A2(net485));
 sg13g2_o21ai_1 _2057_ (.B1(net482),
    .Y(_0076_),
    .A1(_1080_),
    .A2(_1081_));
 sg13g2_a21oi_1 _2058_ (.A1(_1078_),
    .A2(_0076_),
    .Y(_0077_),
    .B1(net521));
 sg13g2_and2_1 _2059_ (.A(_0825_),
    .B(_0988_),
    .X(_0078_));
 sg13g2_and2_1 _2060_ (.A(_0546_),
    .B(_0622_),
    .X(_0079_));
 sg13g2_a21oi_1 _2061_ (.A1(_0634_),
    .A2(_0079_),
    .Y(_0080_),
    .B1(net560));
 sg13g2_o21ai_1 _2062_ (.B1(_0080_),
    .Y(_0081_),
    .A1(_0656_),
    .A2(_0078_));
 sg13g2_a22oi_1 _2063_ (.Y(_0082_),
    .B1(_0648_),
    .B2(_0698_),
    .A2(_0641_),
    .A1(_0531_));
 sg13g2_or2_1 _2064_ (.X(_0083_),
    .B(_0082_),
    .A(net593));
 sg13g2_a21oi_1 _2065_ (.A1(_0643_),
    .A2(_0719_),
    .Y(_0084_),
    .B1(net580));
 sg13g2_a21oi_1 _2066_ (.A1(_0722_),
    .A2(_0084_),
    .Y(_0085_),
    .B1(net550));
 sg13g2_a21oi_1 _2067_ (.A1(_0083_),
    .A2(_0085_),
    .Y(_0086_),
    .B1(_0633_));
 sg13g2_a21oi_1 _2068_ (.A1(net581),
    .A2(_0567_),
    .Y(_0087_),
    .B1(net556));
 sg13g2_nand2b_1 _2069_ (.Y(_0088_),
    .B(_0087_),
    .A_N(_0084_));
 sg13g2_o21ai_1 _2070_ (.B1(net550),
    .Y(_0089_),
    .A1(net580),
    .A2(_0615_));
 sg13g2_nor2_1 _2071_ (.A(_0079_),
    .B(_0089_),
    .Y(_0090_));
 sg13g2_a21oi_1 _2072_ (.A1(_0780_),
    .A2(_0090_),
    .Y(_0091_),
    .B1(net483));
 sg13g2_a221oi_1 _2073_ (.B2(_0091_),
    .C1(net514),
    .B1(_0088_),
    .A1(_0081_),
    .Y(_0092_),
    .A2(_0086_));
 sg13g2_o21ai_1 _2074_ (.B1(net497),
    .Y(_0093_),
    .A1(_0077_),
    .A2(_0092_));
 sg13g2_nand4_1 _2075_ (.B(_0528_),
    .C(net491),
    .A(net613),
    .Y(_0094_),
    .D(_0622_));
 sg13g2_a21oi_1 _2076_ (.A1(_0972_),
    .A2(_0094_),
    .Y(_0095_),
    .B1(net592));
 sg13g2_and3_1 _2077_ (.X(_0096_),
    .A(net592),
    .B(_0722_),
    .C(_0909_));
 sg13g2_o21ai_1 _2078_ (.B1(net561),
    .Y(_0097_),
    .A1(_0095_),
    .A2(_0096_));
 sg13g2_o21ai_1 _2079_ (.B1(net551),
    .Y(_0098_),
    .A1(net591),
    .A2(net485));
 sg13g2_a221oi_1 _2080_ (.B2(_0595_),
    .C1(_0098_),
    .B1(_0961_),
    .A1(net579),
    .Y(_0099_),
    .A2(_0708_));
 sg13g2_nor2_1 _2081_ (.A(net520),
    .B(_0099_),
    .Y(_0100_));
 sg13g2_a221oi_1 _2082_ (.B2(_0853_),
    .C1(net581),
    .B1(_0709_),
    .A1(net615),
    .Y(_0101_),
    .A2(_0567_));
 sg13g2_nor4_1 _2083_ (.A(net534),
    .B(_0525_),
    .C(net596),
    .D(_0781_),
    .Y(_0102_));
 sg13g2_or3_1 _2084_ (.A(net565),
    .B(_0101_),
    .C(_0102_),
    .X(_0103_));
 sg13g2_o21ai_1 _2085_ (.B1(net562),
    .Y(_0104_),
    .A1(_0547_),
    .A2(net487));
 sg13g2_a21oi_1 _2086_ (.A1(_0532_),
    .A2(_0691_),
    .Y(_0105_),
    .B1(_0104_));
 sg13g2_nor2_1 _2087_ (.A(net515),
    .B(_0105_),
    .Y(_0106_));
 sg13g2_a221oi_1 _2088_ (.B2(_0106_),
    .C1(net483),
    .B1(_0103_),
    .A1(_0097_),
    .Y(_0107_),
    .A2(_0100_));
 sg13g2_a221oi_1 _2089_ (.B2(_0760_),
    .C1(net586),
    .B1(_0648_),
    .A1(net605),
    .Y(_0108_),
    .A2(net491));
 sg13g2_nor4_1 _2090_ (.A(_0532_),
    .B(_0534_),
    .C(net596),
    .D(_0587_),
    .Y(_0109_));
 sg13g2_nor3_1 _2091_ (.A(net553),
    .B(_0108_),
    .C(_0109_),
    .Y(_0110_));
 sg13g2_nor2_1 _2092_ (.A(_0607_),
    .B(_0667_),
    .Y(_0111_));
 sg13g2_a21oi_1 _2093_ (.A1(net553),
    .A2(_0111_),
    .Y(_0112_),
    .B1(net516));
 sg13g2_a22oi_1 _2094_ (.Y(_0113_),
    .B1(_0972_),
    .B2(_0536_),
    .A2(_0617_),
    .A1(_0579_));
 sg13g2_o21ai_1 _2095_ (.B1(_0112_),
    .Y(_0114_),
    .A1(_0725_),
    .A2(_0113_));
 sg13g2_nand4_1 _2096_ (.B(_0610_),
    .C(_0709_),
    .A(net596),
    .Y(_0115_),
    .D(_0951_));
 sg13g2_o21ai_1 _2097_ (.B1(net553),
    .Y(_0116_),
    .A1(net597),
    .A2(net487));
 sg13g2_a21oi_1 _2098_ (.A1(_0624_),
    .A2(_1069_),
    .Y(_0117_),
    .B1(_0116_));
 sg13g2_o21ai_1 _2099_ (.B1(_0769_),
    .Y(_0118_),
    .A1(_0527_),
    .A2(_0623_));
 sg13g2_a21oi_1 _2100_ (.A1(_0653_),
    .A2(_0988_),
    .Y(_0119_),
    .B1(net553));
 sg13g2_a22oi_1 _2101_ (.Y(_0120_),
    .B1(_0118_),
    .B2(_0119_),
    .A2(_0117_),
    .A1(_0115_));
 sg13g2_a21oi_1 _2102_ (.A1(net515),
    .A2(_0120_),
    .Y(_0121_),
    .B1(net482));
 sg13g2_o21ai_1 _2103_ (.B1(_0121_),
    .Y(_0122_),
    .A1(_0110_),
    .A2(_0114_));
 sg13g2_nor2_1 _2104_ (.A(net496),
    .B(_0107_),
    .Y(_0123_));
 sg13g2_a21oi_1 _2105_ (.A1(_0122_),
    .A2(_0123_),
    .Y(_0124_),
    .B1(_0679_));
 sg13g2_o21ai_1 _2106_ (.B1(net580),
    .Y(_0125_),
    .A1(_0666_),
    .A2(_0879_));
 sg13g2_o21ai_1 _2107_ (.B1(_1056_),
    .Y(_0126_),
    .A1(net614),
    .A2(_0566_));
 sg13g2_nand3_1 _2108_ (.B(_0125_),
    .C(_0126_),
    .A(net561),
    .Y(_0127_));
 sg13g2_nand3b_1 _2109_ (.B(_0697_),
    .C(net592),
    .Y(_0128_),
    .A_N(_0765_));
 sg13g2_a21oi_1 _2110_ (.A1(net550),
    .A2(_0128_),
    .Y(_0129_),
    .B1(net520));
 sg13g2_nor2_1 _2111_ (.A(_0613_),
    .B(_0692_),
    .Y(_0130_));
 sg13g2_nor4_1 _2112_ (.A(_0555_),
    .B(_0645_),
    .C(_0079_),
    .D(_0130_),
    .Y(_0131_));
 sg13g2_nor2_1 _2113_ (.A(net560),
    .B(_0131_),
    .Y(_0132_));
 sg13g2_a221oi_1 _2114_ (.B2(_0587_),
    .C1(net587),
    .B1(_0709_),
    .A1(net606),
    .Y(_0133_),
    .A2(net486));
 sg13g2_o21ai_1 _2115_ (.B1(net563),
    .Y(_0134_),
    .A1(_0583_),
    .A2(_0853_));
 sg13g2_o21ai_1 _2116_ (.B1(net520),
    .Y(_0135_),
    .A1(_0133_),
    .A2(_0134_));
 sg13g2_a21oi_1 _2117_ (.A1(_0127_),
    .A2(_0129_),
    .Y(_0136_),
    .B1(net494));
 sg13g2_o21ai_1 _2118_ (.B1(_0136_),
    .Y(_0137_),
    .A1(_0132_),
    .A2(_0135_));
 sg13g2_a221oi_1 _2119_ (.B2(_0534_),
    .C1(net564),
    .B1(_0774_),
    .A1(_0568_),
    .Y(_0138_),
    .A2(_0663_));
 sg13g2_nand2b_1 _2120_ (.Y(_0139_),
    .B(_0853_),
    .A_N(_0104_));
 sg13g2_nand3b_1 _2121_ (.B(_0139_),
    .C(net520),
    .Y(_0140_),
    .A_N(_0138_));
 sg13g2_nand3_1 _2122_ (.B(_0623_),
    .C(_0953_),
    .A(net580),
    .Y(_0141_));
 sg13g2_nand3b_1 _2123_ (.B(_0141_),
    .C(net561),
    .Y(_0142_),
    .A_N(_0695_));
 sg13g2_o21ai_1 _2124_ (.B1(net579),
    .Y(_0143_),
    .A1(_0564_),
    .A2(_0708_));
 sg13g2_o21ai_1 _2125_ (.B1(_0848_),
    .Y(_0144_),
    .A1(_0579_),
    .A2(_0601_));
 sg13g2_nand3_1 _2126_ (.B(_0143_),
    .C(_0144_),
    .A(net550),
    .Y(_0145_));
 sg13g2_nand3_1 _2127_ (.B(_0142_),
    .C(_0145_),
    .A(net514),
    .Y(_0146_));
 sg13g2_nand3_1 _2128_ (.B(_0140_),
    .C(_0146_),
    .A(net494),
    .Y(_0147_));
 sg13g2_nand3_1 _2129_ (.B(_0137_),
    .C(_0147_),
    .A(_0633_),
    .Y(_0148_));
 sg13g2_a221oi_1 _2130_ (.B2(_0835_),
    .C1(net564),
    .B1(_1076_),
    .A1(_0814_),
    .Y(_0149_),
    .A2(_0840_));
 sg13g2_a221oi_1 _2131_ (.B2(_0811_),
    .C1(net552),
    .B1(_1070_),
    .A1(_0860_),
    .Y(_0150_),
    .A2(_0979_));
 sg13g2_nor3_1 _2132_ (.A(net521),
    .B(_0149_),
    .C(_0150_),
    .Y(_0151_));
 sg13g2_o21ai_1 _2133_ (.B1(net596),
    .Y(_0152_),
    .A1(_0662_),
    .A2(_1069_));
 sg13g2_a21o_1 _2134_ (.A2(_0718_),
    .A1(net485),
    .B1(_0152_),
    .X(_0153_));
 sg13g2_a221oi_1 _2135_ (.B2(_0781_),
    .C1(net596),
    .B1(net486),
    .A1(net617),
    .Y(_0154_),
    .A2(_0551_));
 sg13g2_nor2_1 _2136_ (.A(net554),
    .B(_0154_),
    .Y(_0155_));
 sg13g2_a22oi_1 _2137_ (.Y(_0156_),
    .B1(_0612_),
    .B2(_0617_),
    .A2(_0526_),
    .A1(net537));
 sg13g2_a21o_1 _2138_ (.A2(_0918_),
    .A1(_0683_),
    .B1(net586),
    .X(_0157_));
 sg13g2_o21ai_1 _2139_ (.B1(_0157_),
    .Y(_0158_),
    .A1(_0607_),
    .A2(_0156_));
 sg13g2_a221oi_1 _2140_ (.B2(net553),
    .C1(net515),
    .B1(_0158_),
    .A1(_0153_),
    .Y(_0159_),
    .A2(_0155_));
 sg13g2_or3_1 _2141_ (.A(net494),
    .B(_0151_),
    .C(_0159_),
    .X(_0160_));
 sg13g2_a221oi_1 _2142_ (.B2(_0094_),
    .C1(net520),
    .B1(_0769_),
    .A1(_0644_),
    .Y(_0161_),
    .A2(_0714_));
 sg13g2_a221oi_1 _2143_ (.B2(_0648_),
    .C1(net585),
    .B1(_0760_),
    .A1(net499),
    .Y(_0162_),
    .A2(_0740_));
 sg13g2_a21oi_1 _2144_ (.A1(net511),
    .A2(net507),
    .Y(_0163_),
    .B1(_0843_));
 sg13g2_nor3_1 _2145_ (.A(net515),
    .B(_0162_),
    .C(_0163_),
    .Y(_0164_));
 sg13g2_or3_1 _2146_ (.A(net554),
    .B(_0161_),
    .C(_0164_),
    .X(_0165_));
 sg13g2_a221oi_1 _2147_ (.B2(net616),
    .C1(_0849_),
    .B1(_0645_),
    .A1(_0566_),
    .Y(_0166_),
    .A2(_0641_));
 sg13g2_a21oi_1 _2148_ (.A1(_0534_),
    .A2(_0636_),
    .Y(_0167_),
    .B1(net592));
 sg13g2_o21ai_1 _2149_ (.B1(net521),
    .Y(_0168_),
    .A1(_0166_),
    .A2(_0167_));
 sg13g2_nand2b_1 _2150_ (.Y(_0169_),
    .B(_0637_),
    .A_N(_0529_));
 sg13g2_o21ai_1 _2151_ (.B1(net514),
    .Y(_0170_),
    .A1(net593),
    .A2(net487));
 sg13g2_a21oi_1 _2152_ (.A1(net580),
    .A2(_0647_),
    .Y(_0171_),
    .B1(_0170_));
 sg13g2_a21oi_1 _2153_ (.A1(_0169_),
    .A2(_0171_),
    .Y(_0172_),
    .B1(net561));
 sg13g2_a21oi_1 _2154_ (.A1(_0168_),
    .A2(_0172_),
    .Y(_0173_),
    .B1(net496));
 sg13g2_a21oi_1 _2155_ (.A1(_0165_),
    .A2(_0173_),
    .Y(_0174_),
    .B1(net482));
 sg13g2_a21oi_1 _2156_ (.A1(_0160_),
    .A2(_0174_),
    .Y(_0175_),
    .B1(_0680_));
 sg13g2_a221oi_1 _2157_ (.B2(_0175_),
    .C1(_0733_),
    .B1(_0148_),
    .A1(_0093_),
    .Y(_0176_),
    .A2(_0124_));
 sg13g2_o21ai_1 _2158_ (.B1(_0949_),
    .Y(_0177_),
    .A1(_1067_),
    .A2(_1068_));
 sg13g2_a21oi_2 _2159_ (.B1(_0627_),
    .Y(_0178_),
    .A2(_0631_),
    .A1(_0628_));
 sg13g2_xor2_1 _2160_ (.B(\pix_y[9] ),
    .A(\logo_top[9] ),
    .X(_0179_));
 sg13g2_nor2_1 _2161_ (.A(\logo_top[8] ),
    .B(_0283_),
    .Y(_0180_));
 sg13g2_nor2b_1 _2162_ (.A(\pix_y[7] ),
    .B_N(\logo_top[7] ),
    .Y(_0181_));
 sg13g2_nor2_1 _2163_ (.A(\logo_top[7] ),
    .B(_0284_),
    .Y(_0182_));
 sg13g2_nor2b_1 _2164_ (.A(_0178_),
    .B_N(_0182_),
    .Y(_0183_));
 sg13g2_nor2b_1 _2165_ (.A(\pix_x[8] ),
    .B_N(\logo_left[8] ),
    .Y(_0184_));
 sg13g2_xor2_1 _2166_ (.B(\pix_x[8] ),
    .A(net629),
    .X(_0185_));
 sg13g2_nor2b_1 _2167_ (.A(\logo_left[7] ),
    .B_N(\pix_x[7] ),
    .Y(_0186_));
 sg13g2_and2_1 _2168_ (.A(_0511_),
    .B(net528),
    .X(_0187_));
 sg13g2_nor2b_1 _2169_ (.A(\pix_x[7] ),
    .B_N(\logo_left[7] ),
    .Y(_0188_));
 sg13g2_nor3_1 _2170_ (.A(_0186_),
    .B(_0187_),
    .C(_0188_),
    .Y(_0189_));
 sg13g2_o21ai_1 _2171_ (.B1(_0185_),
    .Y(_0190_),
    .A1(_0186_),
    .A2(_0189_));
 sg13g2_a21o_1 _2172_ (.A2(_0188_),
    .A1(_0185_),
    .B1(_0186_),
    .X(_0191_));
 sg13g2_a21oi_1 _2173_ (.A1(_0187_),
    .A2(_0191_),
    .Y(_0192_),
    .B1(_0189_));
 sg13g2_nand2_1 _2174_ (.Y(_0193_),
    .A(\logo_top[8] ),
    .B(_0283_));
 sg13g2_xnor2_1 _2175_ (.Y(_0194_),
    .A(_0179_),
    .B(_0193_));
 sg13g2_xnor2_1 _2176_ (.Y(_0195_),
    .A(\logo_left[9] ),
    .B(\pix_x[9] ));
 sg13g2_xnor2_1 _2177_ (.Y(_0196_),
    .A(_0184_),
    .B(_0195_));
 sg13g2_nor4_1 _2178_ (.A(_0183_),
    .B(_0192_),
    .C(_0194_),
    .D(_0196_),
    .Y(_0197_));
 sg13g2_nand2_1 _2179_ (.Y(_0198_),
    .A(_0178_),
    .B(_0181_));
 sg13g2_o21ai_1 _2180_ (.B1(_0198_),
    .Y(_0199_),
    .A1(_0179_),
    .A2(_0180_));
 sg13g2_nor3_1 _2181_ (.A(_0179_),
    .B(_0180_),
    .C(_0182_),
    .Y(_0200_));
 sg13g2_o21ai_1 _2182_ (.B1(_0200_),
    .Y(_0201_),
    .A1(_0178_),
    .A2(_0181_));
 sg13g2_nand4_1 _2183_ (.B(_0197_),
    .C(_0199_),
    .A(_0190_),
    .Y(_0202_),
    .D(_0201_));
 sg13g2_nor2b_1 _2184_ (.A(net1),
    .B_N(_0202_),
    .Y(_0203_));
 sg13g2_nor2_2 _2185_ (.A(_0283_),
    .B(_0291_),
    .Y(_0204_));
 sg13g2_o21ai_1 _2186_ (.B1(\pix_x[9] ),
    .Y(_0205_),
    .A1(\pix_x[7] ),
    .A2(\pix_x[8] ));
 sg13g2_nand3b_1 _2187_ (.B(_0205_),
    .C(net637),
    .Y(_0206_),
    .A_N(\pix_y[9] ));
 sg13g2_nor3_2 _2188_ (.A(_0203_),
    .B(_0204_),
    .C(_0206_),
    .Y(_0207_));
 sg13g2_o21ai_1 _2189_ (.B1(_0207_),
    .Y(_0208_),
    .A1(_0176_),
    .A2(_0177_));
 sg13g2_nor2_1 _2190_ (.A(_0950_),
    .B(_0208_),
    .Y(_0061_));
 sg13g2_and2_1 _2191_ (.A(net623),
    .B(\pix_y[9] ),
    .X(_0209_));
 sg13g2_nand4_1 _2192_ (.B(_0330_),
    .C(_0331_),
    .A(net624),
    .Y(_0210_),
    .D(_0209_));
 sg13g2_nand2_1 _2193_ (.Y(_0211_),
    .A(net636),
    .B(_0210_));
 sg13g2_nand4_1 _2194_ (.B(net634),
    .C(_0302_),
    .A(net82),
    .Y(_0212_),
    .D(_0210_));
 sg13g2_o21ai_1 _2195_ (.B1(net83),
    .Y(_0062_),
    .A1(_0278_),
    .A2(net546));
 sg13g2_nand3_1 _2196_ (.B(net632),
    .C(_0302_),
    .A(net136),
    .Y(_0213_));
 sg13g2_nor2_1 _2197_ (.A(_0277_),
    .B(_0278_),
    .Y(_0214_));
 sg13g2_a22oi_1 _2198_ (.Y(_0063_),
    .B1(_0214_),
    .B2(_0302_),
    .A2(_0213_),
    .A1(_0473_));
 sg13g2_and3_1 _2199_ (.X(_0215_),
    .A(net624),
    .B(net546),
    .C(_0214_));
 sg13g2_and2_2 _2200_ (.A(net546),
    .B(_0211_),
    .X(_0216_));
 sg13g2_nor2_1 _2201_ (.A(_0215_),
    .B(_0216_),
    .Y(_0217_));
 sg13g2_a21oi_1 _2202_ (.A1(net546),
    .A2(_0214_),
    .Y(_0218_),
    .B1(net624));
 sg13g2_nor3_1 _2203_ (.A(_0215_),
    .B(_0216_),
    .C(_0218_),
    .Y(_0064_));
 sg13g2_a22oi_1 _2204_ (.Y(_0219_),
    .B1(_0217_),
    .B2(net623),
    .A2(_0215_),
    .A1(_0474_));
 sg13g2_inv_1 _2205_ (.Y(_0065_),
    .A(_0219_));
 sg13g2_and3_2 _2206_ (.X(_0220_),
    .A(net623),
    .B(net622),
    .C(_0215_));
 sg13g2_a21oi_1 _2207_ (.A1(net623),
    .A2(_0215_),
    .Y(_0221_),
    .B1(net622));
 sg13g2_nor3_1 _2208_ (.A(_0216_),
    .B(_0220_),
    .C(_0221_),
    .Y(_0066_));
 sg13g2_nor3_1 _2209_ (.A(_0280_),
    .B(_0216_),
    .C(_0220_),
    .Y(_0222_));
 sg13g2_nand4_1 _2210_ (.B(net635),
    .C(_0210_),
    .A(_0280_),
    .Y(_0223_),
    .D(_0220_));
 sg13g2_nand2b_1 _2211_ (.Y(_0067_),
    .B(_0223_),
    .A_N(_0222_));
 sg13g2_and3_1 _2212_ (.X(_0224_),
    .A(net176),
    .B(net621),
    .C(_0220_));
 sg13g2_a21oi_1 _2213_ (.A1(net153),
    .A2(_0220_),
    .Y(_0225_),
    .B1(net621));
 sg13g2_nor3_1 _2214_ (.A(_0216_),
    .B(_0224_),
    .C(net154),
    .Y(_0068_));
 sg13g2_nor3_1 _2215_ (.A(_0284_),
    .B(_0216_),
    .C(_0224_),
    .Y(_0226_));
 sg13g2_nand4_1 _2216_ (.B(_0284_),
    .C(_0210_),
    .A(net635),
    .Y(_0227_),
    .D(_0224_));
 sg13g2_nand2b_1 _2217_ (.Y(_0069_),
    .B(_0227_),
    .A_N(_0226_));
 sg13g2_nand2b_1 _2218_ (.Y(_0228_),
    .B(_0220_),
    .A_N(_0291_));
 sg13g2_a21oi_1 _2219_ (.A1(_0204_),
    .A2(_0220_),
    .Y(_0229_),
    .B1(_0216_));
 sg13g2_a221oi_1 _2220_ (.B2(_0283_),
    .C1(_0216_),
    .B1(_0228_),
    .A1(_0204_),
    .Y(_0070_),
    .A2(_0220_));
 sg13g2_nand2_1 _2221_ (.Y(_0230_),
    .A(net151),
    .B(_0229_));
 sg13g2_nand2_1 _2222_ (.Y(_0231_),
    .A(net634),
    .B(_0292_));
 sg13g2_o21ai_1 _2223_ (.B1(_0230_),
    .Y(_0071_),
    .A1(_0228_),
    .A2(_0231_));
 sg13g2_xnor2_1 _2224_ (.Y(_0232_),
    .A(\pix_x[2] ),
    .B(_0484_));
 sg13g2_xnor2_1 _2225_ (.Y(_0233_),
    .A(net590),
    .B(_0232_));
 sg13g2_nand2_1 _2226_ (.Y(_0234_),
    .A(net117),
    .B(net2));
 sg13g2_o21ai_1 _2227_ (.B1(_0234_),
    .Y(_0235_),
    .A1(net2),
    .A2(_0233_));
 sg13g2_nand2_1 _2228_ (.Y(_0236_),
    .A(_0009_),
    .B(_0732_));
 sg13g2_and2_1 _2229_ (.A(net631),
    .B(net558),
    .X(_0237_));
 sg13g2_nand2b_1 _2230_ (.Y(_0238_),
    .B(net547),
    .A_N(net631));
 sg13g2_xnor2_1 _2231_ (.Y(_0239_),
    .A(net631),
    .B(net558));
 sg13g2_xnor2_1 _2232_ (.Y(_0240_),
    .A(_0949_),
    .B(_0239_));
 sg13g2_xnor2_1 _2233_ (.Y(_0241_),
    .A(_0236_),
    .B(_0240_));
 sg13g2_nor3_1 _2234_ (.A(net576),
    .B(_0232_),
    .C(_0241_),
    .Y(_0242_));
 sg13g2_o21ai_1 _2235_ (.B1(_0241_),
    .Y(_0243_),
    .A1(net576),
    .A2(_0232_));
 sg13g2_nor2b_1 _2236_ (.A(_0242_),
    .B_N(_0243_),
    .Y(_0244_));
 sg13g2_nand2_1 _2237_ (.Y(_0245_),
    .A(net2),
    .B(net164));
 sg13g2_o21ai_1 _2238_ (.B1(_0245_),
    .Y(_0246_),
    .A1(net2),
    .A2(_0244_));
 sg13g2_nand2_1 _2239_ (.Y(_0247_),
    .A(_0235_),
    .B(_0246_));
 sg13g2_or2_1 _2240_ (.X(_0248_),
    .B(_0246_),
    .A(_0235_));
 sg13g2_a21oi_1 _2241_ (.A1(_0236_),
    .A2(_0240_),
    .Y(_0249_),
    .B1(_0242_));
 sg13g2_a21oi_1 _2242_ (.A1(_0949_),
    .A2(_0238_),
    .Y(_0250_),
    .B1(_0237_));
 sg13g2_xor2_1 _2243_ (.B(_0493_),
    .A(\pix_x[4] ),
    .X(_0251_));
 sg13g2_xnor2_1 _2244_ (.Y(_0252_),
    .A(net513),
    .B(_0251_));
 sg13g2_xnor2_1 _2245_ (.Y(_0253_),
    .A(_0250_),
    .B(_0252_));
 sg13g2_xnor2_1 _2246_ (.Y(_0254_),
    .A(_0249_),
    .B(_0253_));
 sg13g2_nand2_1 _2247_ (.Y(_0255_),
    .A(net87),
    .B(net2));
 sg13g2_o21ai_1 _2248_ (.B1(_0255_),
    .Y(_0256_),
    .A1(net2),
    .A2(_0254_));
 sg13g2_inv_1 _2249_ (.Y(_0257_),
    .A(_0256_));
 sg13g2_o21ai_1 _2250_ (.B1(_0247_),
    .Y(_0258_),
    .A1(_0248_),
    .A2(_0257_));
 sg13g2_nor3_1 _2251_ (.A(_0950_),
    .B(_0208_),
    .C(_0258_),
    .Y(_0072_));
 sg13g2_nand2_1 _2252_ (.Y(_0259_),
    .A(_0247_),
    .B(_0256_));
 sg13g2_nor2b_1 _2253_ (.A(_0259_),
    .B_N(_0248_),
    .Y(_0260_));
 sg13g2_nor3_1 _2254_ (.A(_0950_),
    .B(_0208_),
    .C(_0260_),
    .Y(_0073_));
 sg13g2_nand2_1 _2255_ (.Y(_0261_),
    .A(_0246_),
    .B(_0257_));
 sg13g2_inv_1 _2256_ (.Y(_0262_),
    .A(_0261_));
 sg13g2_nor4_1 _2257_ (.A(_0950_),
    .B(_0208_),
    .C(_0235_),
    .D(_0262_),
    .Y(_0074_));
 sg13g2_nand2_1 _2258_ (.Y(_0263_),
    .A(_0259_),
    .B(_0261_));
 sg13g2_nor3_1 _2259_ (.A(_0950_),
    .B(_0208_),
    .C(_0263_),
    .Y(_0075_));
 sg13g2_dfrbp_1 _2260_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net65),
    .D(_0016_),
    .Q_N(_0015_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _2261_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net24),
    .D(_0017_),
    .Q_N(_1127_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _2262_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net23),
    .D(net131),
    .Q_N(_1126_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _2263_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net22),
    .D(_0019_),
    .Q_N(_1125_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _2264_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net21),
    .D(_0020_),
    .Q_N(_1124_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _2265_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net20),
    .D(_0021_),
    .Q_N(_1123_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net19),
    .D(_0022_),
    .Q_N(_1122_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _2267_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net80),
    .D(_0023_),
    .Q_N(_1121_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net79),
    .D(net143),
    .Q_N(_1120_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net78),
    .D(_0025_),
    .Q_N(_1119_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _2270_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net77),
    .D(net90),
    .Q_N(_0014_),
    .Q(\logo_left[0] ));
 sg13g2_dfrbp_1 _2271_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net74),
    .D(_0027_),
    .Q_N(_1118_),
    .Q(\logo_left[1] ));
 sg13g2_dfrbp_1 _2272_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net72),
    .D(_0028_),
    .Q_N(_0009_),
    .Q(\logo_left[2] ));
 sg13g2_dfrbp_1 _2273_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net70),
    .D(_0029_),
    .Q_N(_1117_),
    .Q(\logo_left[3] ));
 sg13g2_dfrbp_1 _2274_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net68),
    .D(_0030_),
    .Q_N(_0007_),
    .Q(\logo_left[4] ));
 sg13g2_dfrbp_1 _2275_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net66),
    .D(_0031_),
    .Q_N(_1116_),
    .Q(\logo_left[5] ));
 sg13g2_dfrbp_1 _2276_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net63),
    .D(_0032_),
    .Q_N(_1115_),
    .Q(\logo_left[6] ));
 sg13g2_dfrbp_1 _2277_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net61),
    .D(_0033_),
    .Q_N(_1114_),
    .Q(\logo_left[7] ));
 sg13g2_dfrbp_1 _2278_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net59),
    .D(_0034_),
    .Q_N(_0008_),
    .Q(\logo_left[8] ));
 sg13g2_dfrbp_1 _2279_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net57),
    .D(_0035_),
    .Q_N(_1113_),
    .Q(\logo_left[9] ));
 sg13g2_dfrbp_1 _2280_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net55),
    .D(net92),
    .Q_N(_0013_),
    .Q(\logo_top[0] ));
 sg13g2_dfrbp_1 _2281_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net53),
    .D(_0037_),
    .Q_N(_1112_),
    .Q(\logo_top[1] ));
 sg13g2_dfrbp_1 _2282_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net51),
    .D(_0038_),
    .Q_N(_1111_),
    .Q(\logo_top[2] ));
 sg13g2_dfrbp_1 _2283_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net49),
    .D(_0039_),
    .Q_N(_1110_),
    .Q(\logo_top[3] ));
 sg13g2_dfrbp_1 _2284_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net47),
    .D(_0040_),
    .Q_N(_0002_),
    .Q(\logo_top[4] ));
 sg13g2_dfrbp_1 _2285_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net45),
    .D(_0041_),
    .Q_N(_1109_),
    .Q(\logo_top[5] ));
 sg13g2_dfrbp_1 _2286_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net43),
    .D(_0042_),
    .Q_N(_1108_),
    .Q(\logo_top[6] ));
 sg13g2_dfrbp_1 _2287_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net41),
    .D(_0043_),
    .Q_N(_1107_),
    .Q(\logo_top[7] ));
 sg13g2_dfrbp_1 _2288_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net39),
    .D(net150),
    .Q_N(_0003_),
    .Q(\logo_top[8] ));
 sg13g2_dfrbp_1 _2289_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net37),
    .D(_0045_),
    .Q_N(_1106_),
    .Q(\logo_top[9] ));
 sg13g2_dfrbp_1 _2290_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net35),
    .D(net101),
    .Q_N(_0006_),
    .Q(dir_x));
 sg13g2_dfrbp_1 _2291_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net33),
    .D(net107),
    .Q_N(_0010_),
    .Q(dir_y));
 sg13g2_dfrbp_1 _2292_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net31),
    .D(net88),
    .Q_N(_0012_),
    .Q(\color_index[0] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net29),
    .D(net125),
    .Q_N(_0005_),
    .Q(\color_index[1] ));
 sg13g2_dfrbp_1 _2294_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net27),
    .D(net96),
    .Q_N(_0004_),
    .Q(\color_index[2] ));
 sg13g2_dfrbp_1 _2295_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net25),
    .D(net103),
    .Q_N(_1105_),
    .Q(\prev_y[0] ));
 sg13g2_dfrbp_1 _2296_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net75),
    .D(net98),
    .Q_N(_1104_),
    .Q(\prev_y[1] ));
 sg13g2_dfrbp_1 _2297_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net73),
    .D(net109),
    .Q_N(_1103_),
    .Q(\prev_y[2] ));
 sg13g2_dfrbp_1 _2298_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net71),
    .D(net94),
    .Q_N(_1102_),
    .Q(\prev_y[3] ));
 sg13g2_dfrbp_1 _2299_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net69),
    .D(_0055_),
    .Q_N(_1101_),
    .Q(\prev_y[4] ));
 sg13g2_dfrbp_1 _2300_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net67),
    .D(net116),
    .Q_N(_1100_),
    .Q(\prev_y[5] ));
 sg13g2_dfrbp_1 _2301_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net64),
    .D(net122),
    .Q_N(_1099_),
    .Q(\prev_y[6] ));
 sg13g2_dfrbp_1 _2302_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net62),
    .D(net105),
    .Q_N(_1098_),
    .Q(\prev_y[7] ));
 sg13g2_dfrbp_1 _2303_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net60),
    .D(net112),
    .Q_N(_1097_),
    .Q(\prev_y[8] ));
 sg13g2_dfrbp_1 _2304_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net58),
    .D(net114),
    .Q_N(_1096_),
    .Q(\prev_y[9] ));
 sg13g2_dfrbp_1 _2305_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net76),
    .D(_0061_),
    .Q_N(_1128_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2306_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net56),
    .D(net135),
    .Q_N(_1095_),
    .Q(hsync));
 sg13g2_dfrbp_1 _2307_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net54),
    .D(net84),
    .Q_N(_0011_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _2308_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net50),
    .D(net137),
    .Q_N(_1094_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _2309_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net46),
    .D(_0064_),
    .Q_N(_1093_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _2310_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net42),
    .D(_0065_),
    .Q_N(_1092_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _2311_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net38),
    .D(_0066_),
    .Q_N(_1091_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _2312_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net34),
    .D(_0067_),
    .Q_N(_1090_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _2313_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net30),
    .D(_0068_),
    .Q_N(_1089_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _2314_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net26),
    .D(net169),
    .Q_N(_1088_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _2315_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(net147),
    .Q_N(_1087_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _2316_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net36),
    .D(net152),
    .Q_N(_1129_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 _2317_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net40),
    .D(net86),
    .Q_N(_1086_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _2318_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net32),
    .D(_0072_),
    .Q_N(_1085_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2319_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net28),
    .D(_0073_),
    .Q_N(_1084_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2320_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net52),
    .D(net118),
    .Q_N(_1083_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2321_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net44),
    .D(_0075_),
    .Q_N(_1082_),
    .Q(uo_out[0]));
 sg13g2_tiehi _2265__20 (.L_HI(net20));
 sg13g2_tiehi _2264__21 (.L_HI(net21));
 sg13g2_tiehi _2263__22 (.L_HI(net22));
 sg13g2_tiehi _2262__23 (.L_HI(net23));
 sg13g2_tiehi _2261__24 (.L_HI(net24));
 sg13g2_tiehi _2295__25 (.L_HI(net25));
 sg13g2_tiehi _2314__26 (.L_HI(net26));
 sg13g2_tiehi _2294__27 (.L_HI(net27));
 sg13g2_tiehi _2319__28 (.L_HI(net28));
 sg13g2_tiehi _2293__29 (.L_HI(net29));
 sg13g2_tiehi _2313__30 (.L_HI(net30));
 sg13g2_tiehi _2292__31 (.L_HI(net31));
 sg13g2_tiehi _2318__32 (.L_HI(net32));
 sg13g2_tiehi _2291__33 (.L_HI(net33));
 sg13g2_tiehi _2312__34 (.L_HI(net34));
 sg13g2_tiehi _2290__35 (.L_HI(net35));
 sg13g2_tiehi _2316__36 (.L_HI(net36));
 sg13g2_tiehi _2289__37 (.L_HI(net37));
 sg13g2_tiehi _2311__38 (.L_HI(net38));
 sg13g2_tiehi _2288__39 (.L_HI(net39));
 sg13g2_tiehi _2317__40 (.L_HI(net40));
 sg13g2_tiehi _2287__41 (.L_HI(net41));
 sg13g2_tiehi _2310__42 (.L_HI(net42));
 sg13g2_tiehi _2286__43 (.L_HI(net43));
 sg13g2_tiehi _2321__44 (.L_HI(net44));
 sg13g2_tiehi _2285__45 (.L_HI(net45));
 sg13g2_tiehi _2309__46 (.L_HI(net46));
 sg13g2_tiehi _2284__47 (.L_HI(net47));
 sg13g2_tiehi _2315__48 (.L_HI(net48));
 sg13g2_tiehi _2283__49 (.L_HI(net49));
 sg13g2_tiehi _2308__50 (.L_HI(net50));
 sg13g2_tiehi _2282__51 (.L_HI(net51));
 sg13g2_tiehi _2320__52 (.L_HI(net52));
 sg13g2_tiehi _2281__53 (.L_HI(net53));
 sg13g2_tiehi _2307__54 (.L_HI(net54));
 sg13g2_tiehi _2280__55 (.L_HI(net55));
 sg13g2_tiehi _2306__56 (.L_HI(net56));
 sg13g2_tiehi _2279__57 (.L_HI(net57));
 sg13g2_tiehi _2304__58 (.L_HI(net58));
 sg13g2_tiehi _2278__59 (.L_HI(net59));
 sg13g2_tiehi _2303__60 (.L_HI(net60));
 sg13g2_tiehi _2277__61 (.L_HI(net61));
 sg13g2_tiehi _2302__62 (.L_HI(net62));
 sg13g2_tiehi _2276__63 (.L_HI(net63));
 sg13g2_tiehi _2301__64 (.L_HI(net64));
 sg13g2_tiehi _2260__65 (.L_HI(net65));
 sg13g2_tiehi _2275__66 (.L_HI(net66));
 sg13g2_tiehi _2300__67 (.L_HI(net67));
 sg13g2_tiehi _2274__68 (.L_HI(net68));
 sg13g2_tiehi _2299__69 (.L_HI(net69));
 sg13g2_tiehi _2273__70 (.L_HI(net70));
 sg13g2_tiehi _2298__71 (.L_HI(net71));
 sg13g2_tiehi _2272__72 (.L_HI(net72));
 sg13g2_tiehi _2297__73 (.L_HI(net73));
 sg13g2_tiehi _2271__74 (.L_HI(net74));
 sg13g2_tiehi _2296__75 (.L_HI(net75));
 sg13g2_tiehi _2305__76 (.L_HI(net76));
 sg13g2_tiehi _2270__77 (.L_HI(net77));
 sg13g2_tiehi _2269__78 (.L_HI(net78));
 sg13g2_tiehi _2268__79 (.L_HI(net79));
 sg13g2_tiehi _2267__80 (.L_HI(net80));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_4 (.L_LO(net4));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_5 (.L_LO(net5));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_6 (.L_LO(net6));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_7 (.L_LO(net7));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_8 (.L_LO(net8));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_9 (.L_LO(net9));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_10 (.L_LO(net10));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_18 (.L_LO(net18));
 sg13g2_tiehi _2266__19 (.L_HI(net19));
 sg13g2_buf_1 _2400_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _2401_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2402_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(_0633_));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(_0632_));
 sg13g2_buf_2 fanout484 (.A(_0632_),
    .X(net484));
 sg13g2_buf_4 fanout485 (.X(net485),
    .A(_0664_));
 sg13g2_buf_2 fanout486 (.A(_0664_),
    .X(net486));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(_0640_));
 sg13g2_buf_1 fanout488 (.A(_0640_),
    .X(net488));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(net490));
 sg13g2_buf_4 fanout490 (.X(net490),
    .A(_0614_));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net492));
 sg13g2_buf_2 fanout492 (.A(_0602_),
    .X(net492));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(_0585_));
 sg13g2_buf_2 fanout494 (.A(net495),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(_0578_));
 sg13g2_buf_4 fanout496 (.X(net496),
    .A(net498));
 sg13g2_buf_2 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(_0577_));
 sg13g2_buf_4 fanout499 (.X(net499),
    .A(_0565_));
 sg13g2_buf_2 fanout500 (.A(_0565_),
    .X(net500));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(_0556_));
 sg13g2_buf_2 fanout502 (.A(_0554_),
    .X(net502));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(_0554_));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(_0538_));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(_0528_));
 sg13g2_buf_2 fanout506 (.A(net507),
    .X(net506));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(_0526_));
 sg13g2_buf_4 fanout508 (.X(net508),
    .A(_0523_));
 sg13g2_buf_4 fanout509 (.X(net509),
    .A(net510));
 sg13g2_buf_2 fanout510 (.A(_0522_),
    .X(net510));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(_0505_));
 sg13g2_buf_2 fanout512 (.A(_0505_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net517),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(net515),
    .X(net514));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(net517));
 sg13g2_buf_1 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_0600_),
    .X(net517));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net522));
 sg13g2_buf_1 fanout519 (.A(net522),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(net522),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_0599_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_0521_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_0520_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_0519_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_0519_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_0518_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_0517_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_0517_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_0516_),
    .X(net530));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(net533));
 sg13g2_buf_2 fanout532 (.A(net533),
    .X(net532));
 sg13g2_buf_4 fanout533 (.X(net533),
    .A(net534));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(_0501_));
 sg13g2_buf_2 fanout535 (.A(net536),
    .X(net535));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net538));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(net538));
 sg13g2_buf_2 fanout538 (.A(_0500_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(net541),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net541),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net545),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net545),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_1 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_0334_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_0303_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net556),
    .X(net547));
 sg13g2_buf_1 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(net556),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net556),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net555),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_1 fanout555 (.A(net556),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_0563_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(net567));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net563),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net567),
    .X(net562));
 sg13g2_buf_1 fanout563 (.A(net567),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net566),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_0562_),
    .X(net567));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(net569));
 sg13g2_buf_2 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_0503_));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_0502_),
    .X(net572));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(_0502_));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(net576));
 sg13g2_buf_1 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_1 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_4 fanout577 (.X(net577),
    .A(_0545_));
 sg13g2_buf_2 fanout578 (.A(net582),
    .X(net578));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(net582));
 sg13g2_buf_2 fanout580 (.A(net582),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_0545_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(net588),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net588),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net588),
    .X(net585));
 sg13g2_buf_1 fanout586 (.A(net588),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_0545_),
    .X(net588));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(_0544_));
 sg13g2_buf_2 fanout590 (.A(_0544_),
    .X(net590));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(net594));
 sg13g2_buf_2 fanout592 (.A(net594),
    .X(net592));
 sg13g2_buf_1 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net599),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(net599),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(net598),
    .X(net596));
 sg13g2_buf_1 fanout597 (.A(net598),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_0544_),
    .X(net599));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(_0510_));
 sg13g2_buf_1 fanout601 (.A(net602),
    .X(net601));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(_0510_));
 sg13g2_buf_2 fanout603 (.A(net607),
    .X(net603));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(net607));
 sg13g2_buf_2 fanout605 (.A(net607),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_0510_),
    .X(net607));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(net609));
 sg13g2_buf_2 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(net620),
    .X(net610));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(net620));
 sg13g2_buf_1 fanout612 (.A(net620),
    .X(net612));
 sg13g2_buf_4 fanout613 (.X(net613),
    .A(net615));
 sg13g2_buf_2 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net619),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(net619),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(net619),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_0509_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(\pix_y[6] ),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(net85),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(net155),
    .X(net623));
 sg13g2_buf_4 fanout624 (.X(net624),
    .A(net159));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(dir_y));
 sg13g2_buf_2 fanout626 (.A(dir_y),
    .X(net626));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(dir_x));
 sg13g2_buf_2 fanout628 (.A(dir_x),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(\logo_left[8] ),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(net170),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(net172),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(net637),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net636),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net637),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(rst_n),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(rst_n),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(rst_n),
    .X(net639));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_rebeccargb_tt09ball_screensaver_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0015_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0011_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0212_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0062_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold5 (.A(\pix_y[4] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0001_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0012_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0048_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0014_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0026_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0013_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0036_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold13 (.A(\prev_y[3] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0054_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold15 (.A(\color_index[2] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0050_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold17 (.A(\prev_y[1] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0052_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0006_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0455_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0046_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold22 (.A(\prev_y[0] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0051_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold24 (.A(\prev_y[7] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0058_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0010_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0047_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold28 (.A(\prev_y[2] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0053_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold30 (.A(\logo_top[9] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold31 (.A(\prev_y[8] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0059_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold33 (.A(\prev_y[9] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0060_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold35 (.A(\prev_y[5] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0056_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0004_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0074_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold39 (.A(\prev_y[4] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold40 (.A(\logo_left[1] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold41 (.A(\prev_y[6] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0057_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold43 (.A(\color_index[1] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0470_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0049_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold46 (.A(\logo_top[1] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold47 (.A(\pix_x[0] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0304_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold49 (.A(\pix_x[2] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0305_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0018_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold52 (.A(\pix_x[6] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold53 (.A(\pix_x[9] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0297_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0000_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold56 (.A(\pix_y[0] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0063_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold58 (.A(\logo_left[9] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold59 (.A(\pix_x[3] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0306_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold61 (.A(\pix_x[8] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0312_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0024_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold64 (.A(\pix_x[7] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold65 (.A(\pix_x[7] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold66 (.A(\pix_y[8] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0070_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold68 (.A(\logo_top[7] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold69 (.A(\logo_top[8] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0044_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold71 (.A(\pix_y[9] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0071_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold73 (.A(\pix_y[5] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0225_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold75 (.A(\pix_y[3] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold76 (.A(\pix_x[5] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0308_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold78 (.A(\logo_left[2] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold79 (.A(\pix_y[2] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold80 (.A(\logo_left[5] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold81 (.A(\logo_top[4] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold82 (.A(\logo_top[5] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold83 (.A(\logo_top[6] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0005_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold85 (.A(\logo_top[3] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold86 (.A(\pix_x[4] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold87 (.A(\logo_top[2] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold88 (.A(\pix_y[7] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0069_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold90 (.A(\logo_left[6] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold91 (.A(\logo_left[4] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold92 (.A(\logo_left[3] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold93 (.A(\pix_x[4] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0294_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold95 (.A(\pix_y[5] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold96 (.A(\pix_y[5] ),
    .X(net176));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_fill_2 FILLER_4_182 ();
 sg13g2_fill_1 FILLER_4_184 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_4 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_fill_2 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_171 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_4 FILLER_5_237 ();
 sg13g2_fill_2 FILLER_5_241 ();
 sg13g2_decap_8 FILLER_5_247 ();
 sg13g2_decap_8 FILLER_5_254 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_decap_8 FILLER_5_268 ();
 sg13g2_decap_8 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_282 ();
 sg13g2_decap_8 FILLER_5_289 ();
 sg13g2_decap_8 FILLER_5_296 ();
 sg13g2_decap_8 FILLER_5_303 ();
 sg13g2_decap_8 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_317 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_331 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_fill_2 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_30 ();
 sg13g2_decap_4 FILLER_6_35 ();
 sg13g2_fill_1 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_45 ();
 sg13g2_decap_8 FILLER_6_52 ();
 sg13g2_decap_8 FILLER_6_59 ();
 sg13g2_decap_8 FILLER_6_66 ();
 sg13g2_decap_8 FILLER_6_73 ();
 sg13g2_decap_8 FILLER_6_80 ();
 sg13g2_decap_8 FILLER_6_87 ();
 sg13g2_decap_8 FILLER_6_94 ();
 sg13g2_decap_8 FILLER_6_101 ();
 sg13g2_decap_8 FILLER_6_108 ();
 sg13g2_decap_8 FILLER_6_115 ();
 sg13g2_fill_2 FILLER_6_122 ();
 sg13g2_fill_1 FILLER_6_124 ();
 sg13g2_fill_1 FILLER_6_134 ();
 sg13g2_fill_2 FILLER_6_143 ();
 sg13g2_decap_4 FILLER_6_228 ();
 sg13g2_fill_1 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_50 ();
 sg13g2_fill_1 FILLER_7_52 ();
 sg13g2_fill_2 FILLER_7_66 ();
 sg13g2_fill_1 FILLER_7_68 ();
 sg13g2_fill_1 FILLER_7_79 ();
 sg13g2_decap_8 FILLER_7_100 ();
 sg13g2_decap_8 FILLER_7_107 ();
 sg13g2_decap_4 FILLER_7_114 ();
 sg13g2_fill_1 FILLER_7_118 ();
 sg13g2_fill_1 FILLER_7_150 ();
 sg13g2_fill_2 FILLER_7_190 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_fill_2 FILLER_7_201 ();
 sg13g2_fill_1 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_281 ();
 sg13g2_decap_8 FILLER_7_288 ();
 sg13g2_decap_8 FILLER_7_295 ();
 sg13g2_decap_8 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_309 ();
 sg13g2_decap_8 FILLER_7_316 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_8 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_34 ();
 sg13g2_fill_2 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_1 FILLER_8_215 ();
 sg13g2_fill_1 FILLER_8_219 ();
 sg13g2_decap_8 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_288 ();
 sg13g2_decap_8 FILLER_8_295 ();
 sg13g2_decap_8 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_309 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_decap_8 FILLER_8_323 ();
 sg13g2_decap_8 FILLER_8_330 ();
 sg13g2_decap_8 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_51 ();
 sg13g2_decap_4 FILLER_9_58 ();
 sg13g2_fill_2 FILLER_9_67 ();
 sg13g2_fill_2 FILLER_9_79 ();
 sg13g2_fill_2 FILLER_9_96 ();
 sg13g2_fill_1 FILLER_9_98 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_fill_2 FILLER_9_187 ();
 sg13g2_decap_4 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_295 ();
 sg13g2_decap_8 FILLER_9_302 ();
 sg13g2_decap_8 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_351 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_15 ();
 sg13g2_fill_1 FILLER_10_42 ();
 sg13g2_fill_1 FILLER_10_60 ();
 sg13g2_fill_2 FILLER_10_132 ();
 sg13g2_fill_2 FILLER_10_225 ();
 sg13g2_fill_1 FILLER_10_227 ();
 sg13g2_decap_8 FILLER_10_288 ();
 sg13g2_decap_8 FILLER_10_295 ();
 sg13g2_decap_8 FILLER_10_302 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_10_337 ();
 sg13g2_decap_8 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_14 ();
 sg13g2_decap_4 FILLER_11_30 ();
 sg13g2_fill_1 FILLER_11_42 ();
 sg13g2_fill_2 FILLER_11_78 ();
 sg13g2_fill_2 FILLER_11_92 ();
 sg13g2_fill_2 FILLER_11_114 ();
 sg13g2_fill_2 FILLER_11_143 ();
 sg13g2_fill_2 FILLER_11_170 ();
 sg13g2_fill_1 FILLER_11_172 ();
 sg13g2_fill_2 FILLER_11_179 ();
 sg13g2_fill_2 FILLER_11_199 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_fill_2 FILLER_12_54 ();
 sg13g2_fill_1 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_66 ();
 sg13g2_fill_2 FILLER_12_80 ();
 sg13g2_fill_1 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_115 ();
 sg13g2_fill_1 FILLER_12_142 ();
 sg13g2_fill_2 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_decap_8 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_fill_1 FILLER_13_48 ();
 sg13g2_fill_1 FILLER_13_68 ();
 sg13g2_fill_1 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_118 ();
 sg13g2_fill_2 FILLER_13_146 ();
 sg13g2_fill_1 FILLER_13_233 ();
 sg13g2_fill_1 FILLER_13_244 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_11 ();
 sg13g2_fill_1 FILLER_14_52 ();
 sg13g2_fill_2 FILLER_14_58 ();
 sg13g2_fill_2 FILLER_14_84 ();
 sg13g2_fill_1 FILLER_14_86 ();
 sg13g2_fill_2 FILLER_14_118 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_fill_2 FILLER_14_129 ();
 sg13g2_fill_1 FILLER_14_148 ();
 sg13g2_fill_2 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_165 ();
 sg13g2_fill_2 FILLER_14_192 ();
 sg13g2_fill_1 FILLER_14_209 ();
 sg13g2_fill_2 FILLER_14_248 ();
 sg13g2_fill_1 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_15 ();
 sg13g2_fill_1 FILLER_15_22 ();
 sg13g2_fill_2 FILLER_15_27 ();
 sg13g2_fill_1 FILLER_15_29 ();
 sg13g2_fill_2 FILLER_15_39 ();
 sg13g2_fill_1 FILLER_15_49 ();
 sg13g2_fill_2 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_fill_2 FILLER_15_155 ();
 sg13g2_fill_1 FILLER_15_188 ();
 sg13g2_fill_2 FILLER_15_213 ();
 sg13g2_fill_2 FILLER_15_241 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_decap_8 FILLER_15_279 ();
 sg13g2_decap_8 FILLER_15_286 ();
 sg13g2_decap_8 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_307 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_fill_2 FILLER_16_40 ();
 sg13g2_decap_4 FILLER_16_47 ();
 sg13g2_fill_1 FILLER_16_64 ();
 sg13g2_fill_1 FILLER_16_74 ();
 sg13g2_fill_1 FILLER_16_107 ();
 sg13g2_fill_2 FILLER_16_132 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_fill_1 FILLER_16_172 ();
 sg13g2_fill_2 FILLER_16_177 ();
 sg13g2_fill_1 FILLER_16_179 ();
 sg13g2_decap_8 FILLER_16_197 ();
 sg13g2_fill_1 FILLER_16_204 ();
 sg13g2_fill_1 FILLER_16_218 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_283 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_fill_2 FILLER_17_76 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_decap_4 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_fill_1 FILLER_17_278 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_4 FILLER_18_31 ();
 sg13g2_fill_1 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_50 ();
 sg13g2_fill_1 FILLER_18_52 ();
 sg13g2_fill_2 FILLER_18_58 ();
 sg13g2_fill_2 FILLER_18_65 ();
 sg13g2_fill_1 FILLER_18_67 ();
 sg13g2_fill_1 FILLER_18_94 ();
 sg13g2_fill_2 FILLER_18_118 ();
 sg13g2_fill_1 FILLER_18_137 ();
 sg13g2_fill_2 FILLER_18_153 ();
 sg13g2_decap_8 FILLER_18_171 ();
 sg13g2_decap_8 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_201 ();
 sg13g2_decap_8 FILLER_18_208 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_decap_4 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_240 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_decap_8 FILLER_18_261 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_4 FILLER_18_319 ();
 sg13g2_fill_2 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_17 ();
 sg13g2_fill_2 FILLER_19_65 ();
 sg13g2_fill_1 FILLER_19_125 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_208 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_fill_2 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_223 ();
 sg13g2_fill_2 FILLER_19_272 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_fill_2 FILLER_19_297 ();
 sg13g2_fill_1 FILLER_19_327 ();
 sg13g2_fill_1 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_19 ();
 sg13g2_fill_1 FILLER_20_24 ();
 sg13g2_fill_2 FILLER_20_35 ();
 sg13g2_fill_1 FILLER_20_42 ();
 sg13g2_decap_4 FILLER_20_48 ();
 sg13g2_fill_1 FILLER_20_52 ();
 sg13g2_decap_4 FILLER_20_60 ();
 sg13g2_fill_1 FILLER_20_64 ();
 sg13g2_fill_2 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_decap_4 FILLER_20_160 ();
 sg13g2_fill_2 FILLER_20_169 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_decap_4 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_228 ();
 sg13g2_fill_1 FILLER_20_230 ();
 sg13g2_decap_4 FILLER_20_243 ();
 sg13g2_decap_4 FILLER_20_282 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_4 FILLER_20_346 ();
 sg13g2_fill_2 FILLER_20_355 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_fill_2 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_1 FILLER_21_31 ();
 sg13g2_fill_2 FILLER_21_68 ();
 sg13g2_fill_1 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_86 ();
 sg13g2_fill_2 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_146 ();
 sg13g2_fill_2 FILLER_21_153 ();
 sg13g2_fill_1 FILLER_21_155 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_decap_4 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_fill_1 FILLER_21_190 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_284 ();
 sg13g2_fill_2 FILLER_21_291 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_2 FILLER_21_299 ();
 sg13g2_fill_2 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_21_341 ();
 sg13g2_fill_1 FILLER_21_366 ();
 sg13g2_fill_1 FILLER_21_372 ();
 sg13g2_decap_4 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_9 ();
 sg13g2_fill_1 FILLER_22_13 ();
 sg13g2_decap_4 FILLER_22_19 ();
 sg13g2_fill_2 FILLER_22_47 ();
 sg13g2_fill_1 FILLER_22_49 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_fill_2 FILLER_22_142 ();
 sg13g2_fill_1 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_150 ();
 sg13g2_decap_4 FILLER_22_157 ();
 sg13g2_fill_2 FILLER_22_171 ();
 sg13g2_fill_2 FILLER_22_183 ();
 sg13g2_fill_1 FILLER_22_185 ();
 sg13g2_fill_2 FILLER_22_204 ();
 sg13g2_fill_1 FILLER_22_206 ();
 sg13g2_decap_4 FILLER_22_212 ();
 sg13g2_decap_4 FILLER_22_220 ();
 sg13g2_decap_8 FILLER_22_230 ();
 sg13g2_decap_4 FILLER_22_237 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_decap_4 FILLER_22_302 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_338 ();
 sg13g2_decap_4 FILLER_22_345 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_fill_2 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_38 ();
 sg13g2_fill_2 FILLER_23_45 ();
 sg13g2_fill_1 FILLER_23_47 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_189 ();
 sg13g2_decap_4 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_209 ();
 sg13g2_fill_2 FILLER_23_232 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_2 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_decap_4 FILLER_23_292 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_333 ();
 sg13g2_fill_2 FILLER_23_366 ();
 sg13g2_fill_1 FILLER_23_368 ();
 sg13g2_fill_2 FILLER_23_374 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_fill_2 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_387 ();
 sg13g2_fill_1 FILLER_23_393 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_fill_2 FILLER_24_52 ();
 sg13g2_fill_2 FILLER_24_70 ();
 sg13g2_fill_1 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_decap_4 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_141 ();
 sg13g2_decap_4 FILLER_24_151 ();
 sg13g2_fill_2 FILLER_24_155 ();
 sg13g2_fill_2 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_fill_2 FILLER_24_183 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_208 ();
 sg13g2_fill_1 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_fill_2 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_fill_2 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_fill_2 FILLER_24_338 ();
 sg13g2_fill_2 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_fill_1 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_32 ();
 sg13g2_fill_2 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_85 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_decap_8 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_266 ();
 sg13g2_fill_2 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_301 ();
 sg13g2_decap_4 FILLER_25_307 ();
 sg13g2_fill_1 FILLER_25_311 ();
 sg13g2_fill_1 FILLER_25_335 ();
 sg13g2_fill_2 FILLER_25_341 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_4 FILLER_25_372 ();
 sg13g2_fill_2 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_48 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_123 ();
 sg13g2_decap_4 FILLER_26_133 ();
 sg13g2_decap_4 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_204 ();
 sg13g2_decap_4 FILLER_26_221 ();
 sg13g2_fill_2 FILLER_26_230 ();
 sg13g2_decap_8 FILLER_26_240 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_300 ();
 sg13g2_decap_4 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_fill_2 FILLER_26_347 ();
 sg13g2_fill_1 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_55 ();
 sg13g2_fill_1 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_85 ();
 sg13g2_decap_4 FILLER_27_122 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_decap_4 FILLER_27_172 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_fill_2 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_decap_4 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_307 ();
 sg13g2_decap_4 FILLER_27_332 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_decap_4 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_28_86 ();
 sg13g2_fill_1 FILLER_28_101 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_4 FILLER_28_134 ();
 sg13g2_fill_2 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_171 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_decap_4 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_212 ();
 sg13g2_decap_4 FILLER_28_229 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_decap_8 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_340 ();
 sg13g2_fill_2 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_fill_1 FILLER_28_386 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_31 ();
 sg13g2_fill_2 FILLER_29_66 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_decap_8 FILLER_29_135 ();
 sg13g2_decap_4 FILLER_29_155 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_187 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_decap_4 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_fill_2 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_decap_4 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_decap_4 FILLER_29_284 ();
 sg13g2_fill_1 FILLER_29_294 ();
 sg13g2_decap_4 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_decap_4 FILLER_29_315 ();
 sg13g2_fill_2 FILLER_29_319 ();
 sg13g2_decap_4 FILLER_29_351 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_363 ();
 sg13g2_fill_2 FILLER_29_379 ();
 sg13g2_fill_1 FILLER_29_381 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_23 ();
 sg13g2_fill_1 FILLER_30_38 ();
 sg13g2_fill_2 FILLER_30_76 ();
 sg13g2_fill_2 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_98 ();
 sg13g2_decap_4 FILLER_30_139 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_164 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_decap_8 FILLER_30_208 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_decap_4 FILLER_30_276 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_4 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_decap_4 FILLER_30_364 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_30 ();
 sg13g2_fill_2 FILLER_31_115 ();
 sg13g2_fill_1 FILLER_31_117 ();
 sg13g2_decap_4 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_130 ();
 sg13g2_decap_4 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_decap_4 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_decap_8 FILLER_31_234 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_243 ();
 sg13g2_fill_1 FILLER_31_256 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_decap_4 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_293 ();
 sg13g2_decap_4 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_4 FILLER_31_379 ();
 sg13g2_fill_2 FILLER_31_383 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_26 ();
 sg13g2_fill_1 FILLER_32_41 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_decap_8 FILLER_32_113 ();
 sg13g2_decap_4 FILLER_32_120 ();
 sg13g2_decap_4 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_146 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_173 ();
 sg13g2_fill_2 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_208 ();
 sg13g2_fill_2 FILLER_32_227 ();
 sg13g2_decap_8 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_fill_1 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_283 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_decap_4 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_347 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_decap_4 FILLER_32_362 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_fill_1 FILLER_32_373 ();
 sg13g2_fill_1 FILLER_32_379 ();
 sg13g2_fill_1 FILLER_32_390 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_55 ();
 sg13g2_fill_2 FILLER_33_64 ();
 sg13g2_fill_1 FILLER_33_66 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_136 ();
 sg13g2_fill_1 FILLER_33_143 ();
 sg13g2_fill_2 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_183 ();
 sg13g2_decap_4 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_241 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_fill_2 FILLER_33_291 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_321 ();
 sg13g2_fill_1 FILLER_33_323 ();
 sg13g2_fill_2 FILLER_33_333 ();
 sg13g2_decap_4 FILLER_33_340 ();
 sg13g2_decap_4 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_fill_1 FILLER_33_380 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_46 ();
 sg13g2_fill_2 FILLER_34_73 ();
 sg13g2_fill_1 FILLER_34_75 ();
 sg13g2_decap_8 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_113 ();
 sg13g2_decap_8 FILLER_34_118 ();
 sg13g2_decap_8 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_decap_4 FILLER_34_137 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_173 ();
 sg13g2_decap_4 FILLER_34_200 ();
 sg13g2_decap_4 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_decap_8 FILLER_34_265 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_fill_2 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_decap_4 FILLER_34_304 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_323 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_decap_4 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_379 ();
 sg13g2_fill_2 FILLER_34_386 ();
 sg13g2_fill_1 FILLER_34_388 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_4 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_80 ();
 sg13g2_fill_2 FILLER_35_87 ();
 sg13g2_decap_4 FILLER_35_130 ();
 sg13g2_fill_2 FILLER_35_134 ();
 sg13g2_fill_2 FILLER_35_151 ();
 sg13g2_fill_1 FILLER_35_163 ();
 sg13g2_fill_2 FILLER_35_169 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_4 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_decap_4 FILLER_35_230 ();
 sg13g2_decap_4 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_fill_2 FILLER_35_320 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_decap_4 FILLER_35_357 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_35 ();
 sg13g2_fill_1 FILLER_36_113 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_fill_2 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_fill_2 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_236 ();
 sg13g2_fill_2 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_decap_4 FILLER_36_319 ();
 sg13g2_decap_4 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_4 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_fill_1 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_61 ();
 sg13g2_fill_1 FILLER_37_68 ();
 sg13g2_fill_1 FILLER_37_76 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_fill_2 FILLER_37_118 ();
 sg13g2_fill_1 FILLER_37_120 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_fill_2 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_156 ();
 sg13g2_fill_2 FILLER_37_173 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_decap_4 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_fill_2 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_320 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_fill_2 FILLER_38_233 ();
 sg13g2_decap_4 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_256 ();
 sg13g2_decap_4 FILLER_38_263 ();
 sg13g2_decap_4 FILLER_38_272 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_304 ();
 sg13g2_decap_4 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_fill_2 FILLER_38_331 ();
 sg13g2_fill_1 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_339 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_decap_4 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule

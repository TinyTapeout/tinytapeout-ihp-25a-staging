module tt_um_toivoh_pio_ram_emu_example (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire \rx_pins[0] ;
 wire \rx_pins[1] ;
 wire \top.buttons_stable ;
 wire \top.c_x[0] ;
 wire \top.c_x[10] ;
 wire \top.c_x[11] ;
 wire \top.c_x[1] ;
 wire \top.c_x[2] ;
 wire \top.c_x[3] ;
 wire \top.c_x[4] ;
 wire \top.c_x[5] ;
 wire \top.c_x[6] ;
 wire \top.c_x[7] ;
 wire \top.c_x[8] ;
 wire \top.c_x[9] ;
 wire \top.c_y[0] ;
 wire \top.c_y[10] ;
 wire \top.c_y[11] ;
 wire \top.c_y[1] ;
 wire \top.c_y[2] ;
 wire \top.c_y[3] ;
 wire \top.c_y[4] ;
 wire \top.c_y[5] ;
 wire \top.c_y[6] ;
 wire \top.c_y[7] ;
 wire \top.c_y[8] ;
 wire \top.c_y[9] ;
 wire \top.debouncer_inst.last_data[0] ;
 wire \top.debouncer_inst.last_data[1] ;
 wire \top.debouncer_inst.last_data[2] ;
 wire \top.debouncer_inst.last_data[3] ;
 wire \top.debouncer_inst.last_data[4] ;
 wire \top.debouncer_inst.last_data[5] ;
 wire \top.debouncer_inst.timer[0] ;
 wire \top.debouncer_inst.timer[10] ;
 wire \top.debouncer_inst.timer[11] ;
 wire \top.debouncer_inst.timer[12] ;
 wire \top.debouncer_inst.timer[13] ;
 wire \top.debouncer_inst.timer[14] ;
 wire \top.debouncer_inst.timer[15] ;
 wire \top.debouncer_inst.timer[16] ;
 wire \top.debouncer_inst.timer[17] ;
 wire \top.debouncer_inst.timer[18] ;
 wire \top.debouncer_inst.timer[1] ;
 wire \top.debouncer_inst.timer[2] ;
 wire \top.debouncer_inst.timer[3] ;
 wire \top.debouncer_inst.timer[4] ;
 wire \top.debouncer_inst.timer[5] ;
 wire \top.debouncer_inst.timer[6] ;
 wire \top.debouncer_inst.timer[7] ;
 wire \top.debouncer_inst.timer[8] ;
 wire \top.debouncer_inst.timer[9] ;
 wire \top.early_x[0] ;
 wire \top.early_x[1] ;
 wire \top.early_x[2] ;
 wire \top.early_x[3] ;
 wire \top.julia_calc.dest_x[0] ;
 wire \top.julia_calc.dest_x[1] ;
 wire \top.julia_calc.dest_x[2] ;
 wire \top.julia_calc.dest_x[3] ;
 wire \top.julia_calc.dest_x[4] ;
 wire \top.julia_calc.dest_x[5] ;
 wire \top.julia_calc.dest_x[6] ;
 wire \top.julia_calc.dest_x[7] ;
 wire \top.julia_calc.dest_x[8] ;
 wire \top.julia_calc.dest_y[0] ;
 wire \top.julia_calc.dest_y[1] ;
 wire \top.julia_calc.dest_y[2] ;
 wire \top.julia_calc.dest_y[3] ;
 wire \top.julia_calc.dest_y[4] ;
 wire \top.julia_calc.dest_y[5] ;
 wire \top.julia_calc.dest_y[6] ;
 wire \top.julia_calc.dest_y[7] ;
 wire \top.julia_calc.dest_y[8] ;
 wire \top.julia_calc.far_outside_reg ;
 wire \top.julia_calc.iter[0] ;
 wire \top.julia_calc.iter[1] ;
 wire \top.julia_calc.iter[2] ;
 wire \top.julia_calc.iter[3] ;
 wire \top.julia_calc.iter[4] ;
 wire \top.julia_calc.iter[5] ;
 wire \top.julia_calc.iter[6] ;
 wire \top.julia_calc.iter[7] ;
 wire \top.julia_calc.iter[8] ;
 wire \top.julia_calc.iter_done_reg ;
 wire \top.julia_calc.new_pixel_group ;
 wire \top.julia_calc.new_pixel_group1 ;
 wire \top.julia_calc.phase[0] ;
 wire \top.julia_calc.phase[1] ;
 wire \top.julia_calc.pixel_sreg[0] ;
 wire \top.julia_calc.pixel_sreg[10] ;
 wire \top.julia_calc.pixel_sreg[11] ;
 wire \top.julia_calc.pixel_sreg[12] ;
 wire \top.julia_calc.pixel_sreg[13] ;
 wire \top.julia_calc.pixel_sreg[14] ;
 wire \top.julia_calc.pixel_sreg[15] ;
 wire \top.julia_calc.pixel_sreg[1] ;
 wire \top.julia_calc.pixel_sreg[2] ;
 wire \top.julia_calc.pixel_sreg[3] ;
 wire \top.julia_calc.pixel_sreg[4] ;
 wire \top.julia_calc.pixel_sreg[5] ;
 wire \top.julia_calc.pixel_sreg[6] ;
 wire \top.julia_calc.pixel_sreg[7] ;
 wire \top.julia_calc.pixel_sreg[8] ;
 wire \top.julia_calc.pixel_sreg[9] ;
 wire \top.julia_calc.w_addr[0] ;
 wire \top.julia_calc.w_addr[10] ;
 wire \top.julia_calc.w_addr[11] ;
 wire \top.julia_calc.w_addr[12] ;
 wire \top.julia_calc.w_addr[13] ;
 wire \top.julia_calc.w_addr[14] ;
 wire \top.julia_calc.w_addr[1] ;
 wire \top.julia_calc.w_addr[2] ;
 wire \top.julia_calc.w_addr[3] ;
 wire \top.julia_calc.w_addr[4] ;
 wire \top.julia_calc.w_addr[5] ;
 wire \top.julia_calc.w_addr[6] ;
 wire \top.julia_calc.w_addr[7] ;
 wire \top.julia_calc.w_addr[8] ;
 wire \top.julia_calc.w_addr[9] ;
 wire \top.julia_calc.write_addr_available ;
 wire \top.julia_calc.write_data_available ;
 wire \top.julia_calc.write_mode_data ;
 wire \top.julia_calc.z_x2[0] ;
 wire \top.julia_calc.z_x2[10] ;
 wire \top.julia_calc.z_x2[11] ;
 wire \top.julia_calc.z_x2[12] ;
 wire \top.julia_calc.z_x2[1] ;
 wire \top.julia_calc.z_x2[2] ;
 wire \top.julia_calc.z_x2[3] ;
 wire \top.julia_calc.z_x2[4] ;
 wire \top.julia_calc.z_x2[5] ;
 wire \top.julia_calc.z_x2[6] ;
 wire \top.julia_calc.z_x2[7] ;
 wire \top.julia_calc.z_x2[8] ;
 wire \top.julia_calc.z_x2[9] ;
 wire \top.julia_calc.z_x[0] ;
 wire \top.julia_calc.z_x[10] ;
 wire \top.julia_calc.z_x[11] ;
 wire \top.julia_calc.z_x[1] ;
 wire \top.julia_calc.z_x[2] ;
 wire \top.julia_calc.z_x[3] ;
 wire \top.julia_calc.z_x[4] ;
 wire \top.julia_calc.z_x[5] ;
 wire \top.julia_calc.z_x[6] ;
 wire \top.julia_calc.z_x[7] ;
 wire \top.julia_calc.z_x[8] ;
 wire \top.julia_calc.z_x[9] ;
 wire \top.julia_calc.z_xy[0] ;
 wire \top.julia_calc.z_xy[10] ;
 wire \top.julia_calc.z_xy[11] ;
 wire \top.julia_calc.z_xy[1] ;
 wire \top.julia_calc.z_xy[2] ;
 wire \top.julia_calc.z_xy[3] ;
 wire \top.julia_calc.z_xy[4] ;
 wire \top.julia_calc.z_xy[5] ;
 wire \top.julia_calc.z_xy[6] ;
 wire \top.julia_calc.z_xy[7] ;
 wire \top.julia_calc.z_xy[8] ;
 wire \top.julia_calc.z_xy[9] ;
 wire \top.julia_calc.z_y2[0] ;
 wire \top.julia_calc.z_y2[10] ;
 wire \top.julia_calc.z_y2[11] ;
 wire \top.julia_calc.z_y2[12] ;
 wire \top.julia_calc.z_y2[1] ;
 wire \top.julia_calc.z_y2[2] ;
 wire \top.julia_calc.z_y2[3] ;
 wire \top.julia_calc.z_y2[4] ;
 wire \top.julia_calc.z_y2[5] ;
 wire \top.julia_calc.z_y2[6] ;
 wire \top.julia_calc.z_y2[7] ;
 wire \top.julia_calc.z_y2[8] ;
 wire \top.julia_calc.z_y2[9] ;
 wire \top.julia_calc.z_y[0] ;
 wire \top.julia_calc.z_y[10] ;
 wire \top.julia_calc.z_y[11] ;
 wire \top.julia_calc.z_y[1] ;
 wire \top.julia_calc.z_y[2] ;
 wire \top.julia_calc.z_y[3] ;
 wire \top.julia_calc.z_y[4] ;
 wire \top.julia_calc.z_y[5] ;
 wire \top.julia_calc.z_y[6] ;
 wire \top.julia_calc.z_y[7] ;
 wire \top.julia_calc.z_y[8] ;
 wire \top.julia_calc.z_y[9] ;
 wire \top.last_stable_buttons[0] ;
 wire \top.last_stable_buttons[1] ;
 wire \top.last_stable_buttons[2] ;
 wire \top.last_stable_buttons[3] ;
 wire \top.last_stable_buttons[4] ;
 wire \top.last_stable_buttons[5] ;
 wire \top.next_read_addr[10] ;
 wire \top.next_read_addr[11] ;
 wire \top.next_read_addr[12] ;
 wire \top.next_read_addr[13] ;
 wire \top.next_read_addr[14] ;
 wire \top.next_read_addr[6] ;
 wire \top.next_read_addr[7] ;
 wire \top.next_read_addr[8] ;
 wire \top.next_read_addr[9] ;
 wire \top.pixel_buffer[0][0] ;
 wire \top.pixel_buffer[0][1] ;
 wire \top.pixel_buffer[10][0] ;
 wire \top.pixel_buffer[10][1] ;
 wire \top.pixel_buffer[11][0] ;
 wire \top.pixel_buffer[11][1] ;
 wire \top.pixel_buffer[12][0] ;
 wire \top.pixel_buffer[12][1] ;
 wire \top.pixel_buffer[13][0] ;
 wire \top.pixel_buffer[13][1] ;
 wire \top.pixel_buffer[14][0] ;
 wire \top.pixel_buffer[14][1] ;
 wire \top.pixel_buffer[15][0] ;
 wire \top.pixel_buffer[15][1] ;
 wire \top.pixel_buffer[1][0] ;
 wire \top.pixel_buffer[1][1] ;
 wire \top.pixel_buffer[2][0] ;
 wire \top.pixel_buffer[2][1] ;
 wire \top.pixel_buffer[3][0] ;
 wire \top.pixel_buffer[3][1] ;
 wire \top.pixel_buffer[4][0] ;
 wire \top.pixel_buffer[4][1] ;
 wire \top.pixel_buffer[5][0] ;
 wire \top.pixel_buffer[5][1] ;
 wire \top.pixel_buffer[6][0] ;
 wire \top.pixel_buffer[6][1] ;
 wire \top.pixel_buffer[7][0] ;
 wire \top.pixel_buffer[7][1] ;
 wire \top.pixel_buffer[8][0] ;
 wire \top.pixel_buffer[8][1] ;
 wire \top.pixel_buffer[9][0] ;
 wire \top.pixel_buffer[9][1] ;
 wire \top.receiver.data[0] ;
 wire \top.receiver.data[10] ;
 wire \top.receiver.data[11] ;
 wire \top.receiver.data[12] ;
 wire \top.receiver.data[13] ;
 wire \top.receiver.data[1] ;
 wire \top.receiver.data[2] ;
 wire \top.receiver.data[3] ;
 wire \top.receiver.data[4] ;
 wire \top.receiver.data[5] ;
 wire \top.receiver.data[6] ;
 wire \top.receiver.data[7] ;
 wire \top.receiver.data[8] ;
 wire \top.receiver.data[9] ;
 wire \top.receiver.receiver.counter[0] ;
 wire \top.receiver.receiver.counter[1] ;
 wire \top.receiver.receiver.counter[2] ;
 wire \top.receiver.receiver.counter[3] ;
 wire \top.rs.x[10] ;
 wire \top.rs.x[11] ;
 wire \top.rs.x[4] ;
 wire \top.rs.x[5] ;
 wire \top.rs.x[6] ;
 wire \top.rs.x[7] ;
 wire \top.rs.x[8] ;
 wire \top.rs.x[9] ;
 wire \top.rs.y[9] ;
 wire \top.step_size[0] ;
 wire \top.step_size[1] ;
 wire \top.step_size[2] ;
 wire \top.step_size[3] ;
 wire \top.transmitter.message_accepted ;
 wire \top.transmitter.transmitter.counter[0] ;
 wire \top.transmitter.transmitter.counter[1] ;
 wire \top.transmitter.transmitter.counter[2] ;
 wire \top.transmitter.transmitter.counter[3] ;
 wire \top.transmitter.transmitter.tx_sreg[0] ;
 wire \top.transmitter.transmitter.tx_sreg[10] ;
 wire \top.transmitter.transmitter.tx_sreg[11] ;
 wire \top.transmitter.transmitter.tx_sreg[12] ;
 wire \top.transmitter.transmitter.tx_sreg[13] ;
 wire \top.transmitter.transmitter.tx_sreg[14] ;
 wire \top.transmitter.transmitter.tx_sreg[15] ;
 wire \top.transmitter.transmitter.tx_sreg[16] ;
 wire \top.transmitter.transmitter.tx_sreg[17] ;
 wire \top.transmitter.transmitter.tx_sreg[18] ;
 wire \top.transmitter.transmitter.tx_sreg[19] ;
 wire \top.transmitter.transmitter.tx_sreg[1] ;
 wire \top.transmitter.transmitter.tx_sreg[20] ;
 wire \top.transmitter.transmitter.tx_sreg[2] ;
 wire \top.transmitter.transmitter.tx_sreg[3] ;
 wire \top.transmitter.transmitter.tx_sreg[4] ;
 wire \top.transmitter.transmitter.tx_sreg[5] ;
 wire \top.transmitter.transmitter.tx_sreg[6] ;
 wire \top.transmitter.transmitter.tx_sreg[7] ;
 wire \top.transmitter.transmitter.tx_sreg[8] ;
 wire \top.transmitter.transmitter.tx_sreg[9] ;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net320;
 wire clknet_leaf_0_clk;
 wire net15;
 wire net16;
 wire \uio_out0[4] ;
 wire \uio_out0[5] ;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire \uo_out0[3] ;
 wire \uo_out0[7] ;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;

 sg13g2_and2_1 _2724_ (.A(net557),
    .B(_1880_),
    .X(_1881_));
 sg13g2_nand2_1 _2725_ (.Y(_1882_),
    .A(net557),
    .B(_1880_));
 sg13g2_nor2b_1 _2726_ (.A(net557),
    .B_N(_1880_),
    .Y(_1883_));
 sg13g2_nand2_1 _2727_ (.Y(_1884_),
    .A(net631),
    .B(_1883_));
 sg13g2_nor2_1 _2728_ (.A(net564),
    .B(_1884_),
    .Y(_1885_));
 sg13g2_nand3_1 _2729_ (.B(\top.julia_calc.write_data_available ),
    .C(_1883_),
    .A(net564),
    .Y(_1886_));
 sg13g2_nor2b_1 _2730_ (.A(_1885_),
    .B_N(_1886_),
    .Y(_1887_));
 sg13g2_nand3_1 _2731_ (.B(net817),
    .C(net836),
    .A(\top.transmitter.transmitter.counter[0] ),
    .Y(_1888_));
 sg13g2_nand4_1 _2732_ (.B(\top.transmitter.transmitter.counter[1] ),
    .C(\top.transmitter.transmitter.counter[2] ),
    .A(\top.transmitter.transmitter.counter[0] ),
    .Y(_1889_),
    .D(\top.transmitter.transmitter.counter[3] ));
 sg13g2_a21o_2 _2733_ (.A2(_1887_),
    .A1(net462),
    .B1(net576),
    .X(_1890_));
 sg13g2_nor2_2 _2734_ (.A(_1889_),
    .B(_1890_),
    .Y(\top.transmitter.message_accepted ));
 sg13g2_and3_1 _2735_ (.X(_1891_),
    .A(\top.next_read_addr[13] ),
    .B(\top.next_read_addr[12] ),
    .C(\top.next_read_addr[11] ));
 sg13g2_nand3_1 _2736_ (.B(\top.next_read_addr[12] ),
    .C(\top.next_read_addr[11] ),
    .A(net720),
    .Y(_1892_));
 sg13g2_a21oi_2 _2737_ (.B1(\top.rs.y[9] ),
    .Y(_1893_),
    .A2(_1891_),
    .A1(\top.next_read_addr[14] ));
 sg13g2_o21ai_1 _2738_ (.B1(_1893_),
    .Y(_1894_),
    .A1(\top.next_read_addr[6] ),
    .A2(_1892_));
 sg13g2_nor2b_1 _2739_ (.A(\top.next_read_addr[10] ),
    .B_N(\top.next_read_addr[7] ),
    .Y(_1895_));
 sg13g2_a21oi_1 _2740_ (.A1(\top.next_read_addr[9] ),
    .A2(_1895_),
    .Y(_1896_),
    .B1(_1892_));
 sg13g2_nor3_1 _2741_ (.A(\top.rs.y[9] ),
    .B(\top.next_read_addr[8] ),
    .C(_1896_),
    .Y(_1897_));
 sg13g2_nand3_1 _2742_ (.B(_1894_),
    .C(_1897_),
    .A(net783),
    .Y(\uo_out0[3] ));
 sg13g2_or2_1 _2743_ (.X(_1898_),
    .B(\top.rs.x[6] ),
    .A(\top.rs.x[7] ));
 sg13g2_nor3_1 _2744_ (.A(\top.early_x[0] ),
    .B(\top.rs.x[11] ),
    .C(_1898_),
    .Y(_1899_));
 sg13g2_a21oi_1 _2745_ (.A1(_1883_),
    .A2(_1899_),
    .Y(_1900_),
    .B1(net791));
 sg13g2_nand3_1 _2746_ (.B(\top.rs.x[8] ),
    .C(_1842_),
    .A(\top.rs.x[10] ),
    .Y(_1901_));
 sg13g2_nand2_2 _2747_ (.Y(_1902_),
    .A(\top.rs.x[7] ),
    .B(\top.rs.x[6] ));
 sg13g2_nand3_1 _2748_ (.B(\top.rs.x[7] ),
    .C(\top.rs.x[6] ),
    .A(net556),
    .Y(_1903_));
 sg13g2_o21ai_1 _2749_ (.B1(_1903_),
    .Y(_1904_),
    .A1(net556),
    .A2(_1898_));
 sg13g2_or3_1 _2750_ (.A(net792),
    .B(_1901_),
    .C(_1904_),
    .X(\uo_out0[7] ));
 sg13g2_nor2b_1 _2751_ (.A(\top.julia_calc.phase[0] ),
    .B_N(\top.julia_calc.phase[1] ),
    .Y(_1905_));
 sg13g2_nand2_1 _2752_ (.Y(_1906_),
    .A(\top.julia_calc.phase[1] ),
    .B(_1835_));
 sg13g2_nor2b_1 _2753_ (.A(\top.julia_calc.far_outside_reg ),
    .B_N(_0056_),
    .Y(_1907_));
 sg13g2_nor2_1 _2754_ (.A(\top.julia_calc.z_x2[6] ),
    .B(\top.julia_calc.z_y2[6] ),
    .Y(_1908_));
 sg13g2_and2_1 _2755_ (.A(\top.julia_calc.z_x2[3] ),
    .B(\top.julia_calc.z_y2[3] ),
    .X(_1909_));
 sg13g2_a22oi_1 _2756_ (.Y(_1910_),
    .B1(\top.julia_calc.z_x2[1] ),
    .B2(\top.julia_calc.z_y2[1] ),
    .A2(\top.julia_calc.z_y2[2] ),
    .A1(\top.julia_calc.z_x2[2] ));
 sg13g2_nand2_1 _2757_ (.Y(_1911_),
    .A(\top.julia_calc.z_x2[0] ),
    .B(\top.julia_calc.z_y2[0] ));
 sg13g2_xnor2_1 _2758_ (.Y(_1912_),
    .A(\top.julia_calc.z_x2[1] ),
    .B(\top.julia_calc.z_y2[1] ));
 sg13g2_o21ai_1 _2759_ (.B1(_1910_),
    .Y(_1913_),
    .A1(_1911_),
    .A2(_1912_));
 sg13g2_nor2_1 _2760_ (.A(\top.julia_calc.z_x2[2] ),
    .B(\top.julia_calc.z_y2[2] ),
    .Y(_1914_));
 sg13g2_xnor2_1 _2761_ (.Y(_1915_),
    .A(\top.julia_calc.z_x2[3] ),
    .B(\top.julia_calc.z_y2[3] ));
 sg13g2_nor2_1 _2762_ (.A(_1914_),
    .B(_1915_),
    .Y(_1916_));
 sg13g2_a221oi_1 _2763_ (.B2(_1916_),
    .C1(_1909_),
    .B1(_1913_),
    .A1(\top.julia_calc.z_x2[4] ),
    .Y(_1917_),
    .A2(\top.julia_calc.z_y2[4] ));
 sg13g2_or2_1 _2764_ (.X(_1918_),
    .B(\top.julia_calc.z_y2[4] ),
    .A(\top.julia_calc.z_x2[4] ));
 sg13g2_o21ai_1 _2765_ (.B1(_1918_),
    .Y(_1919_),
    .A1(\top.julia_calc.z_x2[5] ),
    .A2(\top.julia_calc.z_y2[5] ));
 sg13g2_a22oi_1 _2766_ (.Y(_1920_),
    .B1(\top.julia_calc.z_x2[5] ),
    .B2(\top.julia_calc.z_y2[5] ),
    .A2(\top.julia_calc.z_y2[6] ),
    .A1(\top.julia_calc.z_x2[6] ));
 sg13g2_o21ai_1 _2767_ (.B1(_1920_),
    .Y(_1921_),
    .A1(_1917_),
    .A2(_1919_));
 sg13g2_nor2_1 _2768_ (.A(\top.julia_calc.z_x2[8] ),
    .B(\top.julia_calc.z_y2[8] ),
    .Y(_1922_));
 sg13g2_xnor2_1 _2769_ (.Y(_1923_),
    .A(\top.julia_calc.z_x2[7] ),
    .B(\top.julia_calc.z_y2[7] ));
 sg13g2_nor2_1 _2770_ (.A(_1908_),
    .B(_1923_),
    .Y(_1924_));
 sg13g2_a22oi_1 _2771_ (.Y(_1925_),
    .B1(_1921_),
    .B2(_1924_),
    .A2(\top.julia_calc.z_y2[7] ),
    .A1(\top.julia_calc.z_x2[7] ));
 sg13g2_nor2_1 _2772_ (.A(\top.julia_calc.z_x2[9] ),
    .B(\top.julia_calc.z_y2[9] ),
    .Y(_1926_));
 sg13g2_nand2_1 _2773_ (.Y(_1927_),
    .A(\top.julia_calc.z_x2[10] ),
    .B(\top.julia_calc.z_y2[10] ));
 sg13g2_xnor2_1 _2774_ (.Y(_1928_),
    .A(\top.julia_calc.z_x2[11] ),
    .B(\top.julia_calc.z_y2[11] ));
 sg13g2_nor2_1 _2775_ (.A(_1927_),
    .B(_1928_),
    .Y(_1929_));
 sg13g2_a22oi_1 _2776_ (.Y(_1930_),
    .B1(\top.julia_calc.z_x2[8] ),
    .B2(\top.julia_calc.z_y2[8] ),
    .A2(\top.julia_calc.z_y2[9] ),
    .A1(\top.julia_calc.z_x2[9] ));
 sg13g2_o21ai_1 _2777_ (.B1(_1930_),
    .Y(_1931_),
    .A1(_1922_),
    .A2(_1925_));
 sg13g2_xnor2_1 _2778_ (.Y(_1932_),
    .A(\top.julia_calc.z_x2[10] ),
    .B(\top.julia_calc.z_y2[10] ));
 sg13g2_nor3_1 _2779_ (.A(_1926_),
    .B(_1928_),
    .C(_1932_),
    .Y(_1933_));
 sg13g2_a221oi_1 _2780_ (.B2(_1933_),
    .C1(_1929_),
    .B1(_1931_),
    .A1(\top.julia_calc.z_x2[11] ),
    .Y(_1934_),
    .A2(\top.julia_calc.z_y2[11] ));
 sg13g2_xnor2_1 _2781_ (.Y(_1935_),
    .A(\top.julia_calc.z_x2[12] ),
    .B(\top.julia_calc.z_y2[12] ));
 sg13g2_xnor2_1 _2782_ (.Y(_1936_),
    .A(_1934_),
    .B(_1935_));
 sg13g2_a21oi_2 _2783_ (.B1(_1906_),
    .Y(_1937_),
    .A2(_1936_),
    .A1(_1907_));
 sg13g2_nand3_1 _2784_ (.B(\top.julia_calc.dest_x[0] ),
    .C(_1937_),
    .A(net843),
    .Y(_1938_));
 sg13g2_nand4_1 _2785_ (.B(\top.julia_calc.dest_x[1] ),
    .C(\top.julia_calc.dest_x[0] ),
    .A(\top.julia_calc.dest_x[2] ),
    .Y(_1939_),
    .D(_1937_));
 sg13g2_inv_2 _2786_ (.Y(\top.julia_calc.new_pixel_group ),
    .A(net440));
 sg13g2_nand2_1 _2787_ (.Y(_1940_),
    .A(net380),
    .B(_1889_));
 sg13g2_nand2_1 _2788_ (.Y(_1941_),
    .A(net583),
    .B(_1889_));
 sg13g2_nand2_1 _2789_ (.Y(_1942_),
    .A(_1890_),
    .B(_1941_));
 sg13g2_a22oi_1 _2790_ (.Y(\uio_out0[4] ),
    .B1(_1940_),
    .B2(_1942_),
    .A2(_1845_),
    .A1(net575));
 sg13g2_nand2_1 _2791_ (.Y(_1943_),
    .A(net370),
    .B(_1889_));
 sg13g2_a22oi_1 _2792_ (.Y(\uio_out0[5] ),
    .B1(_1942_),
    .B2(_1943_),
    .A2(_1851_),
    .A1(net575));
 sg13g2_or2_1 _2793_ (.X(_1944_),
    .B(_1887_),
    .A(net740));
 sg13g2_mux2_1 _2794_ (.A0(net433),
    .A1(_1944_),
    .S(net447),
    .X(_0001_));
 sg13g2_nor2_1 _2795_ (.A(net427),
    .B(net446),
    .Y(_1945_));
 sg13g2_a21oi_1 _2796_ (.A1(_1885_),
    .A2(net446),
    .Y(_0012_),
    .B1(_1945_));
 sg13g2_mux2_1 _2797_ (.A0(net598),
    .A1(_1882_),
    .S(net447),
    .X(_0013_));
 sg13g2_or2_1 _2798_ (.X(_1946_),
    .B(\top.julia_calc.w_addr[0] ),
    .A(net563));
 sg13g2_o21ai_1 _2799_ (.B1(_1946_),
    .Y(_1947_),
    .A1(_1830_),
    .A2(\top.julia_calc.pixel_sreg[0] ));
 sg13g2_nor2_1 _2800_ (.A(net466),
    .B(_1947_),
    .Y(_1948_));
 sg13g2_a21oi_1 _2801_ (.A1(net556),
    .A2(net466),
    .Y(_1949_),
    .B1(_1948_));
 sg13g2_nor2_1 _2802_ (.A(net407),
    .B(net446),
    .Y(_1950_));
 sg13g2_a21oi_1 _2803_ (.A1(net446),
    .A2(_1949_),
    .Y(_0014_),
    .B1(_1950_));
 sg13g2_mux2_1 _2804_ (.A0(\top.julia_calc.w_addr[1] ),
    .A1(\top.julia_calc.pixel_sreg[1] ),
    .S(net564),
    .X(_1951_));
 sg13g2_nor2_1 _2805_ (.A(\top.rs.x[6] ),
    .B(net462),
    .Y(_1952_));
 sg13g2_a21oi_1 _2806_ (.A1(_1882_),
    .A2(_1951_),
    .Y(_1953_),
    .B1(_1952_));
 sg13g2_nor2_1 _2807_ (.A(net403),
    .B(net446),
    .Y(_1954_));
 sg13g2_a21oi_1 _2808_ (.A1(net446),
    .A2(_1953_),
    .Y(_0015_),
    .B1(_1954_));
 sg13g2_a21oi_1 _2809_ (.A1(_1898_),
    .A2(_1902_),
    .Y(_1955_),
    .B1(net462));
 sg13g2_nor2b_1 _2810_ (.A(net563),
    .B_N(\top.julia_calc.w_addr[2] ),
    .Y(_1956_));
 sg13g2_a21oi_1 _2811_ (.A1(net563),
    .A2(net886),
    .Y(_1957_),
    .B1(_1956_));
 sg13g2_a21oi_1 _2812_ (.A1(net462),
    .A2(_1957_),
    .Y(_1958_),
    .B1(_1955_));
 sg13g2_mux2_1 _2813_ (.A0(net620),
    .A1(_1958_),
    .S(net446),
    .X(_0016_));
 sg13g2_nor2_1 _2814_ (.A(net640),
    .B(net445),
    .Y(_1959_));
 sg13g2_nor2_1 _2815_ (.A(\top.rs.x[5] ),
    .B(net558),
    .Y(_1960_));
 sg13g2_inv_1 _2816_ (.Y(_1961_),
    .A(_1960_));
 sg13g2_nor2_1 _2817_ (.A(_1902_),
    .B(net542),
    .Y(_1962_));
 sg13g2_xor2_1 _2818_ (.B(_1962_),
    .A(\top.rs.x[8] ),
    .X(_1963_));
 sg13g2_or2_1 _2819_ (.X(_1964_),
    .B(\top.julia_calc.w_addr[3] ),
    .A(net563));
 sg13g2_o21ai_1 _2820_ (.B1(_1964_),
    .Y(_1965_),
    .A1(_1830_),
    .A2(\top.julia_calc.pixel_sreg[3] ));
 sg13g2_nor2_1 _2821_ (.A(net466),
    .B(_1965_),
    .Y(_1966_));
 sg13g2_a21oi_1 _2822_ (.A1(net466),
    .A2(_1963_),
    .Y(_1967_),
    .B1(_1966_));
 sg13g2_a21oi_1 _2823_ (.A1(net446),
    .A2(_1967_),
    .Y(_0017_),
    .B1(_1959_));
 sg13g2_or2_1 _2824_ (.X(_1968_),
    .B(\top.julia_calc.w_addr[4] ),
    .A(net563));
 sg13g2_o21ai_1 _2825_ (.B1(_1968_),
    .Y(_1969_),
    .A1(_1830_),
    .A2(\top.julia_calc.pixel_sreg[4] ));
 sg13g2_nor3_1 _2826_ (.A(_0022_),
    .B(_1902_),
    .C(net542),
    .Y(_1970_));
 sg13g2_xnor2_1 _2827_ (.Y(_1971_),
    .A(_1842_),
    .B(_1970_));
 sg13g2_nor2_1 _2828_ (.A(net462),
    .B(_1971_),
    .Y(_1972_));
 sg13g2_a21oi_1 _2829_ (.A1(net462),
    .A2(_1969_),
    .Y(_1973_),
    .B1(_1972_));
 sg13g2_mux2_1 _2830_ (.A0(net365),
    .A1(_1973_),
    .S(net445),
    .X(_0018_));
 sg13g2_mux2_1 _2831_ (.A0(\top.julia_calc.w_addr[5] ),
    .A1(\top.julia_calc.pixel_sreg[5] ),
    .S(net563),
    .X(_1974_));
 sg13g2_nor2_1 _2832_ (.A(net466),
    .B(_1974_),
    .Y(_1975_));
 sg13g2_nand3_1 _2833_ (.B(\top.rs.x[9] ),
    .C(_1962_),
    .A(\top.rs.x[8] ),
    .Y(_1976_));
 sg13g2_xnor2_1 _2834_ (.Y(_1977_),
    .A(_1841_),
    .B(_1976_));
 sg13g2_a21oi_1 _2835_ (.A1(net466),
    .A2(_1977_),
    .Y(_1978_),
    .B1(_1975_));
 sg13g2_mux2_1 _2836_ (.A0(net418),
    .A1(_1978_),
    .S(net445),
    .X(_0019_));
 sg13g2_nor2b_1 _2837_ (.A(net562),
    .B_N(\top.julia_calc.w_addr[6] ),
    .Y(_1979_));
 sg13g2_a21oi_1 _2838_ (.A1(net562),
    .A2(\top.julia_calc.pixel_sreg[6] ),
    .Y(_1980_),
    .B1(_1979_));
 sg13g2_nor2_1 _2839_ (.A(net465),
    .B(_1980_),
    .Y(_1981_));
 sg13g2_a21oi_1 _2840_ (.A1(\top.next_read_addr[6] ),
    .A2(net466),
    .Y(_1982_),
    .B1(_1981_));
 sg13g2_nor2_1 _2841_ (.A(net621),
    .B(net445),
    .Y(_1983_));
 sg13g2_a21oi_1 _2842_ (.A1(net445),
    .A2(_1982_),
    .Y(_0002_),
    .B1(_1983_));
 sg13g2_nor2b_1 _2843_ (.A(net562),
    .B_N(net675),
    .Y(_1984_));
 sg13g2_a21oi_1 _2844_ (.A1(net565),
    .A2(net686),
    .Y(_1985_),
    .B1(_1984_));
 sg13g2_nor2_1 _2845_ (.A(net465),
    .B(_1985_),
    .Y(_1986_));
 sg13g2_a21oi_1 _2846_ (.A1(\top.next_read_addr[7] ),
    .A2(net465),
    .Y(_1987_),
    .B1(_1986_));
 sg13g2_nor2_1 _2847_ (.A(net773),
    .B(net442),
    .Y(_1988_));
 sg13g2_a21oi_1 _2848_ (.A1(net444),
    .A2(_1987_),
    .Y(_0003_),
    .B1(_1988_));
 sg13g2_nor2b_1 _2849_ (.A(net562),
    .B_N(\top.julia_calc.w_addr[8] ),
    .Y(_1989_));
 sg13g2_a21oi_1 _2850_ (.A1(net565),
    .A2(\top.julia_calc.pixel_sreg[8] ),
    .Y(_1990_),
    .B1(_1989_));
 sg13g2_nor2_1 _2851_ (.A(net463),
    .B(_1990_),
    .Y(_1991_));
 sg13g2_a21oi_1 _2852_ (.A1(\top.next_read_addr[8] ),
    .A2(net465),
    .Y(_1992_),
    .B1(_1991_));
 sg13g2_nor2_1 _2853_ (.A(net425),
    .B(net443),
    .Y(_1993_));
 sg13g2_a21oi_1 _2854_ (.A1(net444),
    .A2(_1992_),
    .Y(_0004_),
    .B1(_1993_));
 sg13g2_nor2b_1 _2855_ (.A(net562),
    .B_N(\top.julia_calc.w_addr[9] ),
    .Y(_1994_));
 sg13g2_a21oi_1 _2856_ (.A1(net562),
    .A2(\top.julia_calc.pixel_sreg[9] ),
    .Y(_1995_),
    .B1(_1994_));
 sg13g2_nor2_1 _2857_ (.A(net463),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_a21oi_1 _2858_ (.A1(\top.next_read_addr[9] ),
    .A2(net464),
    .Y(_1997_),
    .B1(_1996_));
 sg13g2_nor2_1 _2859_ (.A(net395),
    .B(net442),
    .Y(_1998_));
 sg13g2_a21oi_1 _2860_ (.A1(net442),
    .A2(_1997_),
    .Y(_0005_),
    .B1(_1998_));
 sg13g2_nor2b_1 _2861_ (.A(net561),
    .B_N(\top.julia_calc.w_addr[10] ),
    .Y(_1999_));
 sg13g2_a21oi_1 _2862_ (.A1(net562),
    .A2(\top.julia_calc.pixel_sreg[10] ),
    .Y(_2000_),
    .B1(_1999_));
 sg13g2_nor2_1 _2863_ (.A(net463),
    .B(_2000_),
    .Y(_2001_));
 sg13g2_a21oi_1 _2864_ (.A1(\top.next_read_addr[10] ),
    .A2(net464),
    .Y(_2002_),
    .B1(_2001_));
 sg13g2_nor2_1 _2865_ (.A(net361),
    .B(net442),
    .Y(_2003_));
 sg13g2_a21oi_1 _2866_ (.A1(net442),
    .A2(_2002_),
    .Y(_0006_),
    .B1(_2003_));
 sg13g2_nor2b_1 _2867_ (.A(net561),
    .B_N(\top.julia_calc.w_addr[11] ),
    .Y(_2004_));
 sg13g2_a21oi_1 _2868_ (.A1(net561),
    .A2(\top.julia_calc.pixel_sreg[11] ),
    .Y(_2005_),
    .B1(_2004_));
 sg13g2_nor2_1 _2869_ (.A(net463),
    .B(_2005_),
    .Y(_2006_));
 sg13g2_a21oi_1 _2870_ (.A1(\top.next_read_addr[11] ),
    .A2(net464),
    .Y(_2007_),
    .B1(_2006_));
 sg13g2_nor2_1 _2871_ (.A(net423),
    .B(net442),
    .Y(_2008_));
 sg13g2_a21oi_1 _2872_ (.A1(net442),
    .A2(_2007_),
    .Y(_0007_),
    .B1(_2008_));
 sg13g2_nor2b_1 _2873_ (.A(net561),
    .B_N(\top.julia_calc.w_addr[12] ),
    .Y(_2009_));
 sg13g2_a21oi_1 _2874_ (.A1(net561),
    .A2(\top.julia_calc.pixel_sreg[12] ),
    .Y(_2010_),
    .B1(_2009_));
 sg13g2_nor2_1 _2875_ (.A(net463),
    .B(_2010_),
    .Y(_2011_));
 sg13g2_a21oi_1 _2876_ (.A1(\top.next_read_addr[12] ),
    .A2(net463),
    .Y(_2012_),
    .B1(_2011_));
 sg13g2_nor2_1 _2877_ (.A(net606),
    .B(net444),
    .Y(_2013_));
 sg13g2_a21oi_1 _2878_ (.A1(net442),
    .A2(_2012_),
    .Y(_0008_),
    .B1(_2013_));
 sg13g2_nor2b_1 _2879_ (.A(net561),
    .B_N(\top.julia_calc.w_addr[13] ),
    .Y(_2014_));
 sg13g2_a21oi_1 _2880_ (.A1(net561),
    .A2(\top.julia_calc.pixel_sreg[13] ),
    .Y(_2015_),
    .B1(_2014_));
 sg13g2_nor2_1 _2881_ (.A(net463),
    .B(_2015_),
    .Y(_2016_));
 sg13g2_a21oi_1 _2882_ (.A1(\top.next_read_addr[13] ),
    .A2(net463),
    .Y(_2017_),
    .B1(_2016_));
 sg13g2_nor2_1 _2883_ (.A(net414),
    .B(net443),
    .Y(_2018_));
 sg13g2_a21oi_1 _2884_ (.A1(net443),
    .A2(_2017_),
    .Y(_0009_),
    .B1(_2018_));
 sg13g2_o21ai_1 _2885_ (.B1(net795),
    .Y(_2019_),
    .A1(_1889_),
    .A2(_1890_));
 sg13g2_and2_1 _2886_ (.A(net561),
    .B(\top.julia_calc.pixel_sreg[14] ),
    .X(_2020_));
 sg13g2_a221oi_1 _2887_ (.B2(net557),
    .C1(_2020_),
    .B1(_1880_),
    .A1(_1830_),
    .Y(_2021_),
    .A2(net628));
 sg13g2_o21ai_1 _2888_ (.B1(net445),
    .Y(_2022_),
    .A1(net783),
    .A2(net462));
 sg13g2_o21ai_1 _2889_ (.B1(_2019_),
    .Y(_0010_),
    .A1(_2021_),
    .A2(_2022_));
 sg13g2_nand4_1 _2890_ (.B(net781),
    .C(net462),
    .A(net563),
    .Y(_2023_),
    .D(net445));
 sg13g2_nand2_1 _2891_ (.Y(_0011_),
    .A(_2019_),
    .B(_2023_));
 sg13g2_xor2_1 _2892_ (.B(net860),
    .A(net572),
    .X(_2024_));
 sg13g2_nand2_1 _2893_ (.Y(_0064_),
    .A(net578),
    .B(net861));
 sg13g2_o21ai_1 _2894_ (.B1(net852),
    .Y(_2025_),
    .A1(_1835_),
    .A2(\top.julia_calc.write_data_available ));
 sg13g2_nor2_1 _2895_ (.A(\top.julia_calc.phase[1] ),
    .B(_1835_),
    .Y(_2026_));
 sg13g2_nand2b_1 _2896_ (.Y(_2027_),
    .B(net520),
    .A_N(\top.julia_calc.write_data_available ));
 sg13g2_nand3_1 _2897_ (.B(net853),
    .C(_2027_),
    .A(net578),
    .Y(_0065_));
 sg13g2_and2_2 _2898_ (.A(net736),
    .B(\top.julia_calc.new_pixel_group ),
    .X(_2028_));
 sg13g2_nand3_1 _2899_ (.B(\top.julia_calc.dest_x[4] ),
    .C(_2028_),
    .A(\top.julia_calc.dest_x[5] ),
    .Y(_2029_));
 sg13g2_nor4_2 _2900_ (.A(\top.julia_calc.dest_x[7] ),
    .B(\top.julia_calc.dest_x[6] ),
    .C(_0055_),
    .Y(_2030_),
    .D(_2029_));
 sg13g2_nand2b_2 _2901_ (.Y(_2031_),
    .B(net578),
    .A_N(_2030_));
 sg13g2_nand2b_1 _2902_ (.Y(_2032_),
    .B(\top.julia_calc.dest_x[0] ),
    .A_N(_1937_));
 sg13g2_nand2_1 _2903_ (.Y(_2033_),
    .A(net338),
    .B(_1937_));
 sg13g2_a21oi_1 _2904_ (.A1(_2032_),
    .A2(_2033_),
    .Y(_0066_),
    .B1(_2031_));
 sg13g2_a21oi_1 _2905_ (.A1(\top.julia_calc.dest_x[0] ),
    .A2(_1937_),
    .Y(_2034_),
    .B1(net843));
 sg13g2_nor2_1 _2906_ (.A(_2031_),
    .B(net844),
    .Y(_2035_));
 sg13g2_and2_1 _2907_ (.A(_1938_),
    .B(_2035_),
    .X(_0067_));
 sg13g2_nor2b_1 _2908_ (.A(net662),
    .B_N(_1938_),
    .Y(_2036_));
 sg13g2_nor3_1 _2909_ (.A(\top.julia_calc.new_pixel_group ),
    .B(_2031_),
    .C(net663),
    .Y(_0068_));
 sg13g2_nor2_1 _2910_ (.A(net736),
    .B(net439),
    .Y(_2037_));
 sg13g2_nor3_1 _2911_ (.A(net573),
    .B(_2028_),
    .C(_2037_),
    .Y(_0069_));
 sg13g2_o21ai_1 _2912_ (.B1(net578),
    .Y(_2038_),
    .A1(net814),
    .A2(_2028_));
 sg13g2_a21oi_1 _2913_ (.A1(net814),
    .A2(_2028_),
    .Y(_0070_),
    .B1(_2038_));
 sg13g2_a21oi_1 _2914_ (.A1(net814),
    .A2(_2028_),
    .Y(_2039_),
    .B1(net840));
 sg13g2_nand2_1 _2915_ (.Y(_2040_),
    .A(net578),
    .B(_2029_));
 sg13g2_nor2_1 _2916_ (.A(_2039_),
    .B(_2040_),
    .Y(_0071_));
 sg13g2_and2_1 _2917_ (.A(\top.julia_calc.dest_x[6] ),
    .B(\top.julia_calc.dest_x[5] ),
    .X(_2041_));
 sg13g2_nand4_1 _2918_ (.B(\top.julia_calc.dest_x[5] ),
    .C(\top.julia_calc.dest_x[4] ),
    .A(\top.julia_calc.dest_x[6] ),
    .Y(_2042_),
    .D(_2028_));
 sg13g2_xor2_1 _2919_ (.B(_2029_),
    .A(net865),
    .X(_2043_));
 sg13g2_nor2_1 _2920_ (.A(_2031_),
    .B(net866),
    .Y(_0072_));
 sg13g2_nand4_1 _2921_ (.B(\top.julia_calc.dest_x[4] ),
    .C(_2028_),
    .A(\top.julia_calc.dest_x[7] ),
    .Y(_2044_),
    .D(_2041_));
 sg13g2_xor2_1 _2922_ (.B(_2042_),
    .A(net855),
    .X(_2045_));
 sg13g2_nor2_1 _2923_ (.A(_2031_),
    .B(net856),
    .Y(_0073_));
 sg13g2_xor2_1 _2924_ (.B(_2044_),
    .A(net765),
    .X(_2046_));
 sg13g2_nor2_1 _2925_ (.A(_2031_),
    .B(net766),
    .Y(_0074_));
 sg13g2_nor2_1 _2926_ (.A(net573),
    .B(_1937_),
    .Y(_2047_));
 sg13g2_o21ai_1 _2927_ (.B1(_2047_),
    .Y(_0075_),
    .A1(net523),
    .A2(net544));
 sg13g2_and2_2 _2928_ (.A(\top.julia_calc.phase[1] ),
    .B(net572),
    .X(_2048_));
 sg13g2_nand2_2 _2929_ (.Y(_2049_),
    .A(\top.julia_calc.phase[1] ),
    .B(net572));
 sg13g2_nand2_1 _2930_ (.Y(_2050_),
    .A(net595),
    .B(_2049_));
 sg13g2_and2_1 _2931_ (.A(_0059_),
    .B(_2048_),
    .X(_2051_));
 sg13g2_nand2b_1 _2932_ (.Y(_2052_),
    .B(\top.julia_calc.z_x2[10] ),
    .A_N(\top.julia_calc.z_y2[10] ));
 sg13g2_nand2_1 _2933_ (.Y(_2053_),
    .A(\top.c_x[10] ),
    .B(_1932_));
 sg13g2_xnor2_1 _2934_ (.Y(_2054_),
    .A(\top.c_x[11] ),
    .B(_1928_));
 sg13g2_a21o_1 _2935_ (.A2(_2053_),
    .A1(_2052_),
    .B1(_2054_),
    .X(_2055_));
 sg13g2_nand3_1 _2936_ (.B(_2053_),
    .C(_2054_),
    .A(_2052_),
    .Y(_2056_));
 sg13g2_nand2_1 _2937_ (.Y(_2057_),
    .A(_2055_),
    .B(_2056_));
 sg13g2_xor2_1 _2938_ (.B(_1932_),
    .A(\top.c_x[10] ),
    .X(_2058_));
 sg13g2_xnor2_1 _2939_ (.Y(_2059_),
    .A(\top.julia_calc.z_x2[9] ),
    .B(\top.julia_calc.z_y2[9] ));
 sg13g2_nor2b_1 _2940_ (.A(\top.julia_calc.z_y2[9] ),
    .B_N(\top.julia_calc.z_x2[9] ),
    .Y(_2060_));
 sg13g2_a21oi_1 _2941_ (.A1(\top.c_x[9] ),
    .A2(_2059_),
    .Y(_2061_),
    .B1(_2060_));
 sg13g2_nand2b_1 _2942_ (.Y(_2062_),
    .B(_2058_),
    .A_N(_2061_));
 sg13g2_xor2_1 _2943_ (.B(_2059_),
    .A(\top.c_x[9] ),
    .X(_2063_));
 sg13g2_nor2b_1 _2944_ (.A(\top.julia_calc.z_y2[8] ),
    .B_N(\top.julia_calc.z_x2[8] ),
    .Y(_2064_));
 sg13g2_xnor2_1 _2945_ (.Y(_2065_),
    .A(\top.julia_calc.z_x2[8] ),
    .B(\top.julia_calc.z_y2[8] ));
 sg13g2_a21oi_1 _2946_ (.A1(\top.c_x[8] ),
    .A2(_2065_),
    .Y(_2066_),
    .B1(_2064_));
 sg13g2_nor2b_1 _2947_ (.A(_2066_),
    .B_N(_2063_),
    .Y(_2067_));
 sg13g2_nor2b_1 _2948_ (.A(\top.julia_calc.z_y2[7] ),
    .B_N(\top.julia_calc.z_x2[7] ),
    .Y(_2068_));
 sg13g2_a21oi_1 _2949_ (.A1(\top.c_x[7] ),
    .A2(_1923_),
    .Y(_2069_),
    .B1(_2068_));
 sg13g2_xor2_1 _2950_ (.B(_2065_),
    .A(\top.c_x[8] ),
    .X(_2070_));
 sg13g2_nand2b_1 _2951_ (.Y(_2071_),
    .B(_2070_),
    .A_N(_2069_));
 sg13g2_nor2b_1 _2952_ (.A(\top.julia_calc.z_y2[6] ),
    .B_N(\top.julia_calc.z_x2[6] ),
    .Y(_2072_));
 sg13g2_xnor2_1 _2953_ (.Y(_2073_),
    .A(\top.julia_calc.z_x2[6] ),
    .B(\top.julia_calc.z_y2[6] ));
 sg13g2_a21oi_1 _2954_ (.A1(\top.c_x[6] ),
    .A2(_2073_),
    .Y(_2074_),
    .B1(_2072_));
 sg13g2_xor2_1 _2955_ (.B(_1923_),
    .A(\top.c_x[7] ),
    .X(_2075_));
 sg13g2_nand2b_1 _2956_ (.Y(_2076_),
    .B(_2075_),
    .A_N(_2074_));
 sg13g2_inv_1 _2957_ (.Y(_2077_),
    .A(_2076_));
 sg13g2_xor2_1 _2958_ (.B(_2073_),
    .A(\top.c_x[6] ),
    .X(_2078_));
 sg13g2_nor2b_1 _2959_ (.A(\top.julia_calc.z_y2[5] ),
    .B_N(\top.julia_calc.z_x2[5] ),
    .Y(_2079_));
 sg13g2_xnor2_1 _2960_ (.Y(_2080_),
    .A(\top.julia_calc.z_x2[5] ),
    .B(\top.julia_calc.z_y2[5] ));
 sg13g2_a21oi_1 _2961_ (.A1(\top.c_x[5] ),
    .A2(_2080_),
    .Y(_2081_),
    .B1(_2079_));
 sg13g2_nand2b_1 _2962_ (.Y(_2082_),
    .B(_2078_),
    .A_N(_2081_));
 sg13g2_nor2b_1 _2963_ (.A(\top.julia_calc.z_y2[4] ),
    .B_N(\top.julia_calc.z_x2[4] ),
    .Y(_2083_));
 sg13g2_xnor2_1 _2964_ (.Y(_2084_),
    .A(\top.julia_calc.z_x2[4] ),
    .B(\top.julia_calc.z_y2[4] ));
 sg13g2_a21oi_1 _2965_ (.A1(\top.c_x[4] ),
    .A2(_2084_),
    .Y(_2085_),
    .B1(_2083_));
 sg13g2_xor2_1 _2966_ (.B(_2080_),
    .A(\top.c_x[5] ),
    .X(_2086_));
 sg13g2_nand2b_1 _2967_ (.Y(_2087_),
    .B(_2086_),
    .A_N(_2085_));
 sg13g2_inv_1 _2968_ (.Y(_2088_),
    .A(_2087_));
 sg13g2_xor2_1 _2969_ (.B(_2084_),
    .A(\top.c_x[4] ),
    .X(_2089_));
 sg13g2_nor2b_1 _2970_ (.A(\top.julia_calc.z_y2[3] ),
    .B_N(\top.julia_calc.z_x2[3] ),
    .Y(_2090_));
 sg13g2_a21oi_1 _2971_ (.A1(\top.c_x[3] ),
    .A2(_1915_),
    .Y(_2091_),
    .B1(_2090_));
 sg13g2_nand2b_1 _2972_ (.Y(_2092_),
    .B(_2089_),
    .A_N(_2091_));
 sg13g2_xnor2_1 _2973_ (.Y(_2093_),
    .A(\top.julia_calc.z_x2[2] ),
    .B(\top.julia_calc.z_y2[2] ));
 sg13g2_nor2b_1 _2974_ (.A(\top.julia_calc.z_y2[2] ),
    .B_N(\top.julia_calc.z_x2[2] ),
    .Y(_2094_));
 sg13g2_a21oi_1 _2975_ (.A1(\top.c_x[2] ),
    .A2(_2093_),
    .Y(_2095_),
    .B1(_2094_));
 sg13g2_xor2_1 _2976_ (.B(_1915_),
    .A(\top.c_x[3] ),
    .X(_2096_));
 sg13g2_nand2b_1 _2977_ (.Y(_2097_),
    .B(_2096_),
    .A_N(_2095_));
 sg13g2_xor2_1 _2978_ (.B(_2093_),
    .A(\top.c_x[2] ),
    .X(_2098_));
 sg13g2_inv_1 _2979_ (.Y(_2099_),
    .A(_2098_));
 sg13g2_nor2b_1 _2980_ (.A(\top.julia_calc.z_y2[1] ),
    .B_N(\top.julia_calc.z_x2[1] ),
    .Y(_2100_));
 sg13g2_a21oi_1 _2981_ (.A1(\top.c_x[1] ),
    .A2(_1912_),
    .Y(_2101_),
    .B1(_2100_));
 sg13g2_xor2_1 _2982_ (.B(_1912_),
    .A(\top.c_x[1] ),
    .X(_2102_));
 sg13g2_nand2b_1 _2983_ (.Y(_2103_),
    .B(\top.julia_calc.z_y2[0] ),
    .A_N(\top.c_x[0] ));
 sg13g2_nand2_1 _2984_ (.Y(_2104_),
    .A(_2102_),
    .B(_2103_));
 sg13g2_xor2_1 _2985_ (.B(\top.c_x[0] ),
    .A(\top.julia_calc.z_y2[0] ),
    .X(_2105_));
 sg13g2_nand2_1 _2986_ (.Y(_2106_),
    .A(\top.julia_calc.z_x2[0] ),
    .B(_2105_));
 sg13g2_xor2_1 _2987_ (.B(_2103_),
    .A(_2102_),
    .X(_2107_));
 sg13g2_nand2b_1 _2988_ (.Y(_2108_),
    .B(_2107_),
    .A_N(_2106_));
 sg13g2_xor2_1 _2989_ (.B(_2101_),
    .A(_2098_),
    .X(_2109_));
 sg13g2_a21o_1 _2990_ (.A2(_2108_),
    .A1(_2104_),
    .B1(_2109_),
    .X(_2110_));
 sg13g2_o21ai_1 _2991_ (.B1(_2110_),
    .Y(_2111_),
    .A1(_2099_),
    .A2(_2101_));
 sg13g2_xnor2_1 _2992_ (.Y(_2112_),
    .A(_2095_),
    .B(_2096_));
 sg13g2_nand2_1 _2993_ (.Y(_2113_),
    .A(_2111_),
    .B(_2112_));
 sg13g2_xor2_1 _2994_ (.B(_2091_),
    .A(_2089_),
    .X(_2114_));
 sg13g2_a21o_1 _2995_ (.A2(_2113_),
    .A1(_2097_),
    .B1(_2114_),
    .X(_2115_));
 sg13g2_xnor2_1 _2996_ (.Y(_2116_),
    .A(_2085_),
    .B(_2086_));
 sg13g2_inv_1 _2997_ (.Y(_2117_),
    .A(_2116_));
 sg13g2_a21oi_1 _2998_ (.A1(_2092_),
    .A2(_2115_),
    .Y(_2118_),
    .B1(_2117_));
 sg13g2_a21o_1 _2999_ (.A2(_2115_),
    .A1(_2092_),
    .B1(_2117_),
    .X(_2119_));
 sg13g2_nand2_1 _3000_ (.Y(_2120_),
    .A(_2087_),
    .B(_2119_));
 sg13g2_xnor2_1 _3001_ (.Y(_2121_),
    .A(_2078_),
    .B(_2081_));
 sg13g2_o21ai_1 _3002_ (.B1(_2121_),
    .Y(_2122_),
    .A1(_2088_),
    .A2(_2118_));
 sg13g2_xnor2_1 _3003_ (.Y(_2123_),
    .A(_2074_),
    .B(_2075_));
 sg13g2_inv_1 _3004_ (.Y(_2124_),
    .A(_2123_));
 sg13g2_a21oi_1 _3005_ (.A1(_2082_),
    .A2(_2122_),
    .Y(_2125_),
    .B1(_2124_));
 sg13g2_nor2_1 _3006_ (.A(_2077_),
    .B(_2125_),
    .Y(_2126_));
 sg13g2_xnor2_1 _3007_ (.Y(_2127_),
    .A(_2069_),
    .B(_2070_));
 sg13g2_o21ai_1 _3008_ (.B1(_2127_),
    .Y(_2128_),
    .A1(_2077_),
    .A2(_2125_));
 sg13g2_xor2_1 _3009_ (.B(_2066_),
    .A(_2063_),
    .X(_2129_));
 sg13g2_a21oi_1 _3010_ (.A1(_2071_),
    .A2(_2128_),
    .Y(_2130_),
    .B1(_2129_));
 sg13g2_xnor2_1 _3011_ (.Y(_2131_),
    .A(_2058_),
    .B(_2061_));
 sg13g2_o21ai_1 _3012_ (.B1(_2131_),
    .Y(_2132_),
    .A1(_2067_),
    .A2(_2130_));
 sg13g2_and2_1 _3013_ (.A(_2062_),
    .B(_2132_),
    .X(_2133_));
 sg13g2_o21ai_1 _3014_ (.B1(_2055_),
    .Y(_2134_),
    .A1(_2057_),
    .A2(_2133_));
 sg13g2_xnor2_1 _3015_ (.Y(_2135_),
    .A(_1935_),
    .B(_2134_));
 sg13g2_xnor2_1 _3016_ (.Y(_2136_),
    .A(_2057_),
    .B(_2133_));
 sg13g2_a21oi_1 _3017_ (.A1(\top.julia_calc.z_x2[11] ),
    .A2(_1837_),
    .Y(_2137_),
    .B1(\top.c_x[11] ));
 sg13g2_o21ai_1 _3018_ (.B1(\top.c_x[11] ),
    .Y(_2138_),
    .A1(\top.julia_calc.z_x2[11] ),
    .A2(_1837_));
 sg13g2_nor2b_1 _3019_ (.A(_2137_),
    .B_N(_2138_),
    .Y(_2139_));
 sg13g2_xnor2_1 _3020_ (.Y(_2140_),
    .A(_2136_),
    .B(_2139_));
 sg13g2_nor2b_1 _3021_ (.A(\top.c_y[11] ),
    .B_N(\top.julia_calc.z_xy[10] ),
    .Y(_2141_));
 sg13g2_nand2b_1 _3022_ (.Y(_2142_),
    .B(\top.c_y[11] ),
    .A_N(\top.julia_calc.z_xy[10] ));
 sg13g2_nor2_1 _3023_ (.A(\top.julia_calc.z_xy[9] ),
    .B(\top.c_y[10] ),
    .Y(_2143_));
 sg13g2_nand2_1 _3024_ (.Y(_2144_),
    .A(\top.julia_calc.z_xy[9] ),
    .B(\top.c_y[10] ));
 sg13g2_nand2_1 _3025_ (.Y(_2145_),
    .A(\top.julia_calc.z_xy[7] ),
    .B(\top.c_y[8] ));
 sg13g2_and2_1 _3026_ (.A(\top.julia_calc.z_xy[6] ),
    .B(\top.c_y[7] ),
    .X(_2146_));
 sg13g2_nand2_1 _3027_ (.Y(_2147_),
    .A(\top.julia_calc.z_xy[5] ),
    .B(\top.c_y[6] ));
 sg13g2_and2_1 _3028_ (.A(\top.julia_calc.z_xy[4] ),
    .B(\top.c_y[5] ),
    .X(_2148_));
 sg13g2_nand2_1 _3029_ (.Y(_2149_),
    .A(\top.julia_calc.z_xy[3] ),
    .B(\top.c_y[4] ));
 sg13g2_nand2_1 _3030_ (.Y(_2150_),
    .A(\top.julia_calc.z_xy[2] ),
    .B(\top.c_y[3] ));
 sg13g2_nand2_1 _3031_ (.Y(_2151_),
    .A(\top.julia_calc.z_xy[1] ),
    .B(\top.c_y[2] ));
 sg13g2_or2_1 _3032_ (.X(_2152_),
    .B(\top.c_y[2] ),
    .A(\top.julia_calc.z_xy[1] ));
 sg13g2_nand4_1 _3033_ (.B(\top.c_y[1] ),
    .C(_2151_),
    .A(\top.julia_calc.z_xy[0] ),
    .Y(_2153_),
    .D(_2152_));
 sg13g2_xnor2_1 _3034_ (.Y(_2154_),
    .A(\top.julia_calc.z_xy[2] ),
    .B(\top.c_y[3] ));
 sg13g2_a21o_1 _3035_ (.A2(_2153_),
    .A1(_2151_),
    .B1(_2154_),
    .X(_2155_));
 sg13g2_xnor2_1 _3036_ (.Y(_2156_),
    .A(\top.julia_calc.z_xy[3] ),
    .B(\top.c_y[4] ));
 sg13g2_a21o_1 _3037_ (.A2(_2155_),
    .A1(_2150_),
    .B1(_2156_),
    .X(_2157_));
 sg13g2_xnor2_1 _3038_ (.Y(_2158_),
    .A(\top.julia_calc.z_xy[4] ),
    .B(\top.c_y[5] ));
 sg13g2_a21oi_1 _3039_ (.A1(_2149_),
    .A2(_2157_),
    .Y(_2159_),
    .B1(_2158_));
 sg13g2_xor2_1 _3040_ (.B(\top.c_y[6] ),
    .A(\top.julia_calc.z_xy[5] ),
    .X(_2160_));
 sg13g2_o21ai_1 _3041_ (.B1(_2160_),
    .Y(_2161_),
    .A1(_2148_),
    .A2(_2159_));
 sg13g2_xnor2_1 _3042_ (.Y(_2162_),
    .A(\top.julia_calc.z_xy[6] ),
    .B(\top.c_y[7] ));
 sg13g2_a21oi_1 _3043_ (.A1(_2147_),
    .A2(_2161_),
    .Y(_2163_),
    .B1(_2162_));
 sg13g2_xor2_1 _3044_ (.B(\top.c_y[8] ),
    .A(\top.julia_calc.z_xy[7] ),
    .X(_2164_));
 sg13g2_o21ai_1 _3045_ (.B1(_2164_),
    .Y(_2165_),
    .A1(_2146_),
    .A2(_2163_));
 sg13g2_xnor2_1 _3046_ (.Y(_2166_),
    .A(\top.julia_calc.z_xy[8] ),
    .B(\top.c_y[9] ));
 sg13g2_a21o_1 _3047_ (.A2(_2165_),
    .A1(_2145_),
    .B1(_2166_),
    .X(_2167_));
 sg13g2_inv_1 _3048_ (.Y(_2168_),
    .A(_2167_));
 sg13g2_a21oi_1 _3049_ (.A1(\top.julia_calc.z_xy[8] ),
    .A2(\top.c_y[9] ),
    .Y(_2169_),
    .B1(_2168_));
 sg13g2_o21ai_1 _3050_ (.B1(_2144_),
    .Y(_2170_),
    .A1(_2143_),
    .A2(_2169_));
 sg13g2_o21ai_1 _3051_ (.B1(_2142_),
    .Y(_2171_),
    .A1(_2141_),
    .A2(_2170_));
 sg13g2_xnor2_1 _3052_ (.Y(_2172_),
    .A(\top.julia_calc.z_xy[11] ),
    .B(_2171_));
 sg13g2_xnor2_1 _3053_ (.Y(_2173_),
    .A(_2135_),
    .B(_2140_));
 sg13g2_o21ai_1 _3054_ (.B1(_2051_),
    .Y(_2174_),
    .A1(_2172_),
    .A2(_2173_));
 sg13g2_a21oi_1 _3055_ (.A1(_2050_),
    .A2(_2174_),
    .Y(_0076_),
    .B1(net573));
 sg13g2_nand2_1 _3056_ (.Y(_0314_),
    .A(_1878_),
    .B(net542));
 sg13g2_inv_1 _3057_ (.Y(_0315_),
    .A(_0314_));
 sg13g2_nor2b_2 _3058_ (.A(\top.early_x[3] ),
    .B_N(\top.early_x[2] ),
    .Y(_0316_));
 sg13g2_nand2b_1 _3059_ (.Y(_0317_),
    .B(\top.early_x[2] ),
    .A_N(net559));
 sg13g2_nand2b_2 _3060_ (.Y(_0318_),
    .B(net558),
    .A_N(net556));
 sg13g2_nor2_1 _3061_ (.A(_0317_),
    .B(_0318_),
    .Y(_0319_));
 sg13g2_and2_1 _3062_ (.A(net556),
    .B(net558),
    .X(_0320_));
 sg13g2_nand2_2 _3063_ (.Y(_0321_),
    .A(net556),
    .B(net558));
 sg13g2_nand2_2 _3064_ (.Y(_0322_),
    .A(net559),
    .B(net560));
 sg13g2_nor2_2 _3065_ (.A(_0321_),
    .B(_0322_),
    .Y(_0323_));
 sg13g2_a22oi_1 _3066_ (.Y(_0324_),
    .B1(_0323_),
    .B2(net586),
    .A2(_0319_),
    .A1(\top.pixel_buffer[5][0] ));
 sg13g2_nor2_1 _3067_ (.A(_0317_),
    .B(_0321_),
    .Y(_0325_));
 sg13g2_nand2b_2 _3068_ (.Y(_0326_),
    .B(net556),
    .A_N(net557));
 sg13g2_nor3_2 _3069_ (.A(net559),
    .B(\top.early_x[2] ),
    .C(_0326_),
    .Y(_0327_));
 sg13g2_a22oi_1 _3070_ (.Y(_0328_),
    .B1(_0327_),
    .B2(\top.pixel_buffer[8][0] ),
    .A2(_0325_),
    .A1(\top.pixel_buffer[13][0] ));
 sg13g2_nand2_1 _3071_ (.Y(_0329_),
    .A(_0324_),
    .B(_0328_));
 sg13g2_nand3_1 _3072_ (.B(_1878_),
    .C(_0320_),
    .A(\top.pixel_buffer[12][0] ),
    .Y(_0330_));
 sg13g2_nand2b_1 _3073_ (.Y(_0331_),
    .B(net559),
    .A_N(net560));
 sg13g2_nor2_1 _3074_ (.A(_0318_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_nor2_1 _3075_ (.A(_0322_),
    .B(_0326_),
    .Y(_0333_));
 sg13g2_a22oi_1 _3076_ (.Y(_0334_),
    .B1(_0333_),
    .B2(\top.pixel_buffer[11][0] ),
    .A2(_0332_),
    .A1(\top.pixel_buffer[6][0] ));
 sg13g2_nand3_1 _3077_ (.B(_0330_),
    .C(_0334_),
    .A(_0314_),
    .Y(_0335_));
 sg13g2_nor2_1 _3078_ (.A(_0321_),
    .B(_0331_),
    .Y(_0336_));
 sg13g2_nor2_1 _3079_ (.A(_1961_),
    .B(_0331_),
    .Y(_0337_));
 sg13g2_a22oi_1 _3080_ (.Y(_0338_),
    .B1(_0337_),
    .B2(\top.pixel_buffer[2][0] ),
    .A2(_0336_),
    .A1(\top.pixel_buffer[14][0] ));
 sg13g2_nor2_1 _3081_ (.A(_0326_),
    .B(_0331_),
    .Y(_0339_));
 sg13g2_nand2_1 _3082_ (.Y(_0340_),
    .A(\top.pixel_buffer[10][0] ),
    .B(_0339_));
 sg13g2_nand3_1 _3083_ (.B(net542),
    .C(_0316_),
    .A(\top.pixel_buffer[1][0] ),
    .Y(_0341_));
 sg13g2_nor2_1 _3084_ (.A(_0317_),
    .B(_0326_),
    .Y(_0342_));
 sg13g2_nand2_1 _3085_ (.Y(_0343_),
    .A(\top.pixel_buffer[9][0] ),
    .B(_0342_));
 sg13g2_or2_2 _3086_ (.X(_0344_),
    .B(_0322_),
    .A(_0318_));
 sg13g2_o21ai_1 _3087_ (.B1(_0343_),
    .Y(_0345_),
    .A1(_1834_),
    .A2(_0344_));
 sg13g2_nor3_2 _3088_ (.A(net559),
    .B(net560),
    .C(_0318_),
    .Y(_0346_));
 sg13g2_nor2_1 _3089_ (.A(_1961_),
    .B(_0322_),
    .Y(_0347_));
 sg13g2_a221oi_1 _3090_ (.B2(\top.pixel_buffer[3][0] ),
    .C1(_0345_),
    .B1(_0347_),
    .A1(\top.pixel_buffer[4][0] ),
    .Y(_0348_),
    .A2(_0346_));
 sg13g2_nand4_1 _3091_ (.B(_0340_),
    .C(_0341_),
    .A(_0338_),
    .Y(_0349_),
    .D(_0348_));
 sg13g2_nor3_1 _3092_ (.A(_0329_),
    .B(_0335_),
    .C(_0349_),
    .Y(_0350_));
 sg13g2_a21oi_1 _3093_ (.A1(net731),
    .A2(_0315_),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_a22oi_1 _3094_ (.Y(_0352_),
    .B1(_0342_),
    .B2(\top.pixel_buffer[9][1] ),
    .A2(_0332_),
    .A1(\top.pixel_buffer[6][1] ));
 sg13g2_nand3_1 _3095_ (.B(_1878_),
    .C(_0320_),
    .A(\top.pixel_buffer[12][1] ),
    .Y(_0353_));
 sg13g2_nand3_1 _3096_ (.B(net542),
    .C(_0316_),
    .A(\top.pixel_buffer[1][1] ),
    .Y(_0354_));
 sg13g2_nand4_1 _3097_ (.B(net560),
    .C(\top.pixel_buffer[3][1] ),
    .A(net559),
    .Y(_0355_),
    .D(net542));
 sg13g2_o21ai_1 _3098_ (.B1(_0355_),
    .Y(_0356_),
    .A1(_1832_),
    .A2(_0344_));
 sg13g2_a221oi_1 _3099_ (.B2(\top.pixel_buffer[14][1] ),
    .C1(_0356_),
    .B1(_0336_),
    .A1(_1878_),
    .Y(_0357_),
    .A2(net542));
 sg13g2_nand4_1 _3100_ (.B(_0353_),
    .C(_0354_),
    .A(_0352_),
    .Y(_0358_),
    .D(_0357_));
 sg13g2_a22oi_1 _3101_ (.Y(_0359_),
    .B1(_0325_),
    .B2(\top.pixel_buffer[13][1] ),
    .A2(_0319_),
    .A1(\top.pixel_buffer[5][1] ));
 sg13g2_a22oi_1 _3102_ (.Y(_0360_),
    .B1(_0346_),
    .B2(\top.pixel_buffer[4][1] ),
    .A2(_0337_),
    .A1(\top.pixel_buffer[2][1] ));
 sg13g2_a22oi_1 _3103_ (.Y(_0361_),
    .B1(_0333_),
    .B2(\top.pixel_buffer[11][1] ),
    .A2(_0323_),
    .A1(\top.pixel_buffer[15][1] ));
 sg13g2_a22oi_1 _3104_ (.Y(_0362_),
    .B1(_0339_),
    .B2(\top.pixel_buffer[10][1] ),
    .A2(_0327_),
    .A1(\top.pixel_buffer[8][1] ));
 sg13g2_nand4_1 _3105_ (.B(_0360_),
    .C(_0361_),
    .A(_0359_),
    .Y(_0363_),
    .D(_0362_));
 sg13g2_nor2_1 _3106_ (.A(\top.rs.x[8] ),
    .B(\top.rs.x[9] ),
    .Y(_0364_));
 sg13g2_nand2_1 _3107_ (.Y(_0365_),
    .A(\top.rs.x[10] ),
    .B(_0058_));
 sg13g2_o21ai_1 _3108_ (.B1(_1893_),
    .Y(_0366_),
    .A1(_0364_),
    .A2(_0365_));
 sg13g2_nor2_2 _3109_ (.A(net744),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_o21ai_1 _3110_ (.B1(_0367_),
    .Y(_0368_),
    .A1(_0358_),
    .A2(_0363_));
 sg13g2_a21oi_2 _3111_ (.B1(_0368_),
    .Y(_0080_),
    .A2(_0315_),
    .A1(_1833_));
 sg13g2_and2_1 _3112_ (.A(_0351_),
    .B(_0080_),
    .X(_0077_));
 sg13g2_and2_1 _3113_ (.A(_0351_),
    .B(_0367_),
    .X(_0294_));
 sg13g2_or2_1 _3114_ (.X(_0078_),
    .B(_0294_),
    .A(_0080_));
 sg13g2_nor2b_1 _3115_ (.A(_0351_),
    .B_N(_0080_),
    .Y(_0079_));
 sg13g2_nand2_1 _3116_ (.Y(_0369_),
    .A(net577),
    .B(_1944_));
 sg13g2_a21oi_1 _3117_ (.A1(_1830_),
    .A2(_1884_),
    .Y(_0081_),
    .B1(_0369_));
 sg13g2_xor2_1 _3118_ (.B(\top.debouncer_inst.last_data[3] ),
    .A(net4),
    .X(_0370_));
 sg13g2_xor2_1 _3119_ (.B(\top.debouncer_inst.last_data[4] ),
    .A(net5),
    .X(_0371_));
 sg13g2_xor2_1 _3120_ (.B(\top.debouncer_inst.last_data[5] ),
    .A(net6),
    .X(_0372_));
 sg13g2_nor3_1 _3121_ (.A(_0370_),
    .B(_0371_),
    .C(_0372_),
    .Y(_0373_));
 sg13g2_nand2b_1 _3122_ (.Y(_0374_),
    .B(\top.debouncer_inst.last_data[2] ),
    .A_N(net3));
 sg13g2_xnor2_1 _3123_ (.Y(_0375_),
    .A(net2),
    .B(\top.debouncer_inst.last_data[1] ));
 sg13g2_o21ai_1 _3124_ (.B1(net581),
    .Y(_0376_),
    .A1(net1),
    .A2(_1846_));
 sg13g2_a221oi_1 _3125_ (.B2(_1847_),
    .C1(_0376_),
    .B1(net3),
    .A1(net1),
    .Y(_0377_),
    .A2(_1846_));
 sg13g2_nand4_1 _3126_ (.B(_0374_),
    .C(_0375_),
    .A(_0373_),
    .Y(_0378_),
    .D(_0377_));
 sg13g2_nor2b_1 _3127_ (.A(\top.buttons_stable ),
    .B_N(net386),
    .Y(_0379_));
 sg13g2_nor2b_1 _3128_ (.A(net386),
    .B_N(\top.buttons_stable ),
    .Y(_0380_));
 sg13g2_nor3_1 _3129_ (.A(net456),
    .B(_0379_),
    .C(net387),
    .Y(_0082_));
 sg13g2_and2_1 _3130_ (.A(net584),
    .B(_0379_),
    .X(_0381_));
 sg13g2_nor2_1 _3131_ (.A(net584),
    .B(_0379_),
    .Y(_0382_));
 sg13g2_nor3_1 _3132_ (.A(net455),
    .B(_0381_),
    .C(_0382_),
    .Y(_0083_));
 sg13g2_xnor2_1 _3133_ (.Y(_0383_),
    .A(net680),
    .B(_0381_));
 sg13g2_nor2_1 _3134_ (.A(net456),
    .B(_0383_),
    .Y(_0084_));
 sg13g2_and3_1 _3135_ (.X(_0384_),
    .A(net680),
    .B(net383),
    .C(_0381_));
 sg13g2_a21oi_1 _3136_ (.A1(\top.debouncer_inst.timer[2] ),
    .A2(_0381_),
    .Y(_0385_),
    .B1(net383));
 sg13g2_nor3_1 _3137_ (.A(net456),
    .B(_0384_),
    .C(net384),
    .Y(_0085_));
 sg13g2_a21oi_1 _3138_ (.A1(net802),
    .A2(_0384_),
    .Y(_0386_),
    .B1(net454));
 sg13g2_o21ai_1 _3139_ (.B1(_0386_),
    .Y(_0387_),
    .A1(net802),
    .A2(_0384_));
 sg13g2_inv_1 _3140_ (.Y(_0086_),
    .A(_0387_));
 sg13g2_a21oi_1 _3141_ (.A1(\top.debouncer_inst.timer[4] ),
    .A2(_0384_),
    .Y(_0388_),
    .B1(net400));
 sg13g2_and3_1 _3142_ (.X(_0389_),
    .A(\top.debouncer_inst.timer[4] ),
    .B(net400),
    .C(_0384_));
 sg13g2_nor3_1 _3143_ (.A(net454),
    .B(net401),
    .C(_0389_),
    .Y(_0087_));
 sg13g2_nor2_1 _3144_ (.A(net612),
    .B(_0389_),
    .Y(_0390_));
 sg13g2_and2_1 _3145_ (.A(net612),
    .B(_0389_),
    .X(_0391_));
 sg13g2_nor3_1 _3146_ (.A(net454),
    .B(net613),
    .C(_0391_),
    .Y(_0088_));
 sg13g2_xnor2_1 _3147_ (.Y(_0392_),
    .A(net760),
    .B(_0391_));
 sg13g2_nor2_1 _3148_ (.A(net454),
    .B(_0392_),
    .Y(_0089_));
 sg13g2_a21oi_1 _3149_ (.A1(\top.debouncer_inst.timer[7] ),
    .A2(_0391_),
    .Y(_0393_),
    .B1(net371));
 sg13g2_and3_1 _3150_ (.X(_0394_),
    .A(\top.debouncer_inst.timer[7] ),
    .B(net371),
    .C(_0391_));
 sg13g2_nor3_1 _3151_ (.A(net454),
    .B(net372),
    .C(_0394_),
    .Y(_0090_));
 sg13g2_xnor2_1 _3152_ (.Y(_0395_),
    .A(net715),
    .B(_0394_));
 sg13g2_nor2_1 _3153_ (.A(net454),
    .B(net716),
    .Y(_0091_));
 sg13g2_a21oi_1 _3154_ (.A1(\top.debouncer_inst.timer[9] ),
    .A2(_0394_),
    .Y(_0396_),
    .B1(net409));
 sg13g2_and3_1 _3155_ (.X(_0397_),
    .A(\top.debouncer_inst.timer[9] ),
    .B(net409),
    .C(_0394_));
 sg13g2_nor3_1 _3156_ (.A(net454),
    .B(net410),
    .C(_0397_),
    .Y(_0092_));
 sg13g2_nor2_1 _3157_ (.A(net648),
    .B(_0397_),
    .Y(_0398_));
 sg13g2_and2_1 _3158_ (.A(net648),
    .B(_0397_),
    .X(_0399_));
 sg13g2_nor3_1 _3159_ (.A(net454),
    .B(net649),
    .C(_0399_),
    .Y(_0093_));
 sg13g2_nor2_1 _3160_ (.A(net652),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_and2_1 _3161_ (.A(net652),
    .B(_0399_),
    .X(_0401_));
 sg13g2_nor3_1 _3162_ (.A(net455),
    .B(_0400_),
    .C(_0401_),
    .Y(_0094_));
 sg13g2_xnor2_1 _3163_ (.Y(_0402_),
    .A(net710),
    .B(_0401_));
 sg13g2_nor2_1 _3164_ (.A(net455),
    .B(_0402_),
    .Y(_0095_));
 sg13g2_a21oi_1 _3165_ (.A1(\top.debouncer_inst.timer[13] ),
    .A2(_0401_),
    .Y(_0403_),
    .B1(net367));
 sg13g2_and3_2 _3166_ (.X(_0404_),
    .A(net710),
    .B(net367),
    .C(_0401_));
 sg13g2_nor3_1 _3167_ (.A(net455),
    .B(net368),
    .C(_0404_),
    .Y(_0096_));
 sg13g2_a21oi_1 _3168_ (.A1(net738),
    .A2(_0404_),
    .Y(_0405_),
    .B1(net455));
 sg13g2_o21ai_1 _3169_ (.B1(_0405_),
    .Y(_0406_),
    .A1(net738),
    .A2(_0404_));
 sg13g2_inv_1 _3170_ (.Y(_0097_),
    .A(_0406_));
 sg13g2_a21oi_1 _3171_ (.A1(\top.debouncer_inst.timer[15] ),
    .A2(_0404_),
    .Y(_0407_),
    .B1(net397));
 sg13g2_and3_1 _3172_ (.X(_0408_),
    .A(\top.debouncer_inst.timer[15] ),
    .B(net397),
    .C(_0404_));
 sg13g2_nor3_1 _3173_ (.A(net455),
    .B(net398),
    .C(_0408_),
    .Y(_0098_));
 sg13g2_nor2_1 _3174_ (.A(net646),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_and2_1 _3175_ (.A(net646),
    .B(_0408_),
    .X(_0410_));
 sg13g2_nor3_1 _3176_ (.A(net456),
    .B(net647),
    .C(_0410_),
    .Y(_0099_));
 sg13g2_a21oi_1 _3177_ (.A1(net689),
    .A2(_0410_),
    .Y(_0411_),
    .B1(net455));
 sg13g2_o21ai_1 _3178_ (.B1(_0411_),
    .Y(_0412_),
    .A1(net689),
    .A2(_0410_));
 sg13g2_inv_1 _3179_ (.Y(_0100_),
    .A(_0412_));
 sg13g2_a21oi_1 _3180_ (.A1(net689),
    .A2(_0410_),
    .Y(_0413_),
    .B1(\top.buttons_stable ));
 sg13g2_nor2_1 _3181_ (.A(net455),
    .B(net690),
    .Y(_0101_));
 sg13g2_o21ai_1 _3182_ (.B1(net631),
    .Y(_0414_),
    .A1(net563),
    .A2(_1884_));
 sg13g2_a21oi_1 _3183_ (.A1(net441),
    .A2(_0414_),
    .Y(_0102_),
    .B1(net573));
 sg13g2_a21oi_1 _3184_ (.A1(\top.julia_calc.write_data_available ),
    .A2(_1944_),
    .Y(_0415_),
    .B1(net347));
 sg13g2_nor2_1 _3185_ (.A(net573),
    .B(net348),
    .Y(_0103_));
 sg13g2_nand2_1 _3186_ (.Y(_0416_),
    .A(net577),
    .B(_2048_));
 sg13g2_nor2_1 _3187_ (.A(net566),
    .B(_2049_),
    .Y(_0417_));
 sg13g2_nor2_2 _3188_ (.A(net567),
    .B(net514),
    .Y(_0418_));
 sg13g2_xor2_1 _3189_ (.B(_2105_),
    .A(\top.julia_calc.z_x2[0] ),
    .X(_0419_));
 sg13g2_a22oi_1 _3190_ (.Y(_0420_),
    .B1(_0418_),
    .B2(_0419_),
    .A2(net513),
    .A1(net378));
 sg13g2_inv_1 _3191_ (.Y(_0104_),
    .A(net379));
 sg13g2_xnor2_1 _3192_ (.Y(_0421_),
    .A(_2106_),
    .B(_2107_));
 sg13g2_a22oi_1 _3193_ (.Y(_0422_),
    .B1(_0418_),
    .B2(_0421_),
    .A2(net513),
    .A1(net359));
 sg13g2_inv_1 _3194_ (.Y(_0105_),
    .A(net360));
 sg13g2_nand3_1 _3195_ (.B(_2108_),
    .C(_2109_),
    .A(_2104_),
    .Y(_0423_));
 sg13g2_and2_1 _3196_ (.A(_2110_),
    .B(_0418_),
    .X(_0424_));
 sg13g2_a22oi_1 _3197_ (.Y(_0425_),
    .B1(_0423_),
    .B2(_0424_),
    .A2(net514),
    .A1(net356));
 sg13g2_inv_1 _3198_ (.Y(_0106_),
    .A(_0425_));
 sg13g2_a22oi_1 _3199_ (.Y(_0426_),
    .B1(_0418_),
    .B2(\top.c_y[0] ),
    .A2(net513),
    .A1(net374));
 sg13g2_inv_1 _3200_ (.Y(_0107_),
    .A(net375));
 sg13g2_xor2_1 _3201_ (.B(\top.c_y[1] ),
    .A(\top.julia_calc.z_xy[0] ),
    .X(_0427_));
 sg13g2_a22oi_1 _3202_ (.Y(_0428_),
    .B1(_0418_),
    .B2(_0427_),
    .A2(net513),
    .A1(net357));
 sg13g2_inv_1 _3203_ (.Y(_0108_),
    .A(net358));
 sg13g2_nand2_1 _3204_ (.Y(_0429_),
    .A(net363),
    .B(net513));
 sg13g2_a22oi_1 _3205_ (.Y(_0430_),
    .B1(_2151_),
    .B2(_2152_),
    .A2(\top.c_y[1] ),
    .A1(\top.julia_calc.z_xy[0] ));
 sg13g2_nand2_1 _3206_ (.Y(_0431_),
    .A(_2153_),
    .B(_0418_));
 sg13g2_o21ai_1 _3207_ (.B1(_0429_),
    .Y(_0109_),
    .A1(_0430_),
    .A2(_0431_));
 sg13g2_nor3_2 _3208_ (.A(net523),
    .B(\top.julia_calc.write_data_available ),
    .C(_2049_),
    .Y(_0432_));
 sg13g2_mux2_1 _3209_ (.A0(net625),
    .A1(\top.julia_calc.pixel_sreg[2] ),
    .S(net507),
    .X(_0110_));
 sg13g2_mux2_1 _3210_ (.A0(net693),
    .A1(\top.julia_calc.pixel_sreg[3] ),
    .S(net507),
    .X(_0111_));
 sg13g2_mux2_1 _3211_ (.A0(net713),
    .A1(\top.julia_calc.pixel_sreg[4] ),
    .S(net507),
    .X(_0112_));
 sg13g2_mux2_1 _3212_ (.A0(net711),
    .A1(\top.julia_calc.pixel_sreg[5] ),
    .S(_0432_),
    .X(_0113_));
 sg13g2_mux2_1 _3213_ (.A0(\top.julia_calc.pixel_sreg[4] ),
    .A1(net655),
    .S(net507),
    .X(_0114_));
 sg13g2_mux2_1 _3214_ (.A0(net730),
    .A1(net686),
    .S(net507),
    .X(_0115_));
 sg13g2_mux2_1 _3215_ (.A0(net655),
    .A1(net688),
    .S(net507),
    .X(_0116_));
 sg13g2_mux2_1 _3216_ (.A0(net686),
    .A1(\top.julia_calc.pixel_sreg[9] ),
    .S(net507),
    .X(_0117_));
 sg13g2_mux2_1 _3217_ (.A0(\top.julia_calc.pixel_sreg[8] ),
    .A1(net650),
    .S(net506),
    .X(_0118_));
 sg13g2_mux2_1 _3218_ (.A0(net748),
    .A1(net653),
    .S(net506),
    .X(_0119_));
 sg13g2_mux2_1 _3219_ (.A0(net650),
    .A1(net644),
    .S(net506),
    .X(_0120_));
 sg13g2_mux2_1 _3220_ (.A0(net653),
    .A1(\top.julia_calc.pixel_sreg[13] ),
    .S(net506),
    .X(_0121_));
 sg13g2_mux2_1 _3221_ (.A0(net644),
    .A1(\top.julia_calc.pixel_sreg[14] ),
    .S(net506),
    .X(_0122_));
 sg13g2_mux2_1 _3222_ (.A0(net702),
    .A1(\top.julia_calc.pixel_sreg[15] ),
    .S(net506),
    .X(_0123_));
 sg13g2_mux2_1 _3223_ (.A0(net657),
    .A1(\top.julia_calc.iter[0] ),
    .S(net506),
    .X(_0124_));
 sg13g2_mux2_1 _3224_ (.A0(net781),
    .A1(net707),
    .S(net506),
    .X(_0125_));
 sg13g2_nor2_2 _3225_ (.A(\top.julia_calc.phase[1] ),
    .B(net572),
    .Y(_0433_));
 sg13g2_xnor2_1 _3226_ (.Y(_0434_),
    .A(\top.julia_calc.phase[1] ),
    .B(net572));
 sg13g2_mux2_1 _3227_ (.A0(_0049_),
    .A1(_0048_),
    .S(net536),
    .X(_0435_));
 sg13g2_nor2_1 _3228_ (.A(net571),
    .B(_0048_),
    .Y(_0436_));
 sg13g2_nand2b_1 _3229_ (.Y(_0437_),
    .B(net571),
    .A_N(_0049_));
 sg13g2_nor2b_2 _3230_ (.A(_0436_),
    .B_N(_0437_),
    .Y(_0438_));
 sg13g2_nand2b_2 _3231_ (.Y(_0439_),
    .B(_0437_),
    .A_N(_0436_));
 sg13g2_nor2_1 _3232_ (.A(net505),
    .B(net502),
    .Y(_0440_));
 sg13g2_mux2_2 _3233_ (.A0(_0042_),
    .A1(_0043_),
    .S(net571),
    .X(_0441_));
 sg13g2_inv_2 _3234_ (.Y(_0442_),
    .A(net533));
 sg13g2_mux2_1 _3235_ (.A0(_0051_),
    .A1(_0050_),
    .S(net537),
    .X(_0443_));
 sg13g2_mux2_2 _3236_ (.A0(_1874_),
    .A1(_1875_),
    .S(net536),
    .X(_0444_));
 sg13g2_mux2_2 _3237_ (.A0(_0047_),
    .A1(_0046_),
    .S(net537),
    .X(_0445_));
 sg13g2_mux2_2 _3238_ (.A0(_1871_),
    .A1(_1872_),
    .S(net535),
    .X(_0446_));
 sg13g2_nor2_1 _3239_ (.A(net569),
    .B(_0032_),
    .Y(_0447_));
 sg13g2_nand2b_1 _3240_ (.Y(_0448_),
    .B(net569),
    .A_N(_0033_));
 sg13g2_nor2b_2 _3241_ (.A(_0447_),
    .B_N(_0448_),
    .Y(_0449_));
 sg13g2_nand2b_2 _3242_ (.Y(_0450_),
    .B(_0448_),
    .A_N(_0447_));
 sg13g2_nor2_1 _3243_ (.A(net534),
    .B(_0445_),
    .Y(_0451_));
 sg13g2_nor2_1 _3244_ (.A(net501),
    .B(net498),
    .Y(_0452_));
 sg13g2_and2_1 _3245_ (.A(_0451_),
    .B(_0452_),
    .X(_0453_));
 sg13g2_or2_1 _3246_ (.X(_0454_),
    .B(_0452_),
    .A(_0451_));
 sg13g2_xor2_1 _3247_ (.B(_0452_),
    .A(_0451_),
    .X(_0455_));
 sg13g2_xnor2_1 _3248_ (.Y(_0456_),
    .A(_0440_),
    .B(_0455_));
 sg13g2_nor2_1 _3249_ (.A(net569),
    .B(_0038_),
    .Y(_0457_));
 sg13g2_nand2b_1 _3250_ (.Y(_0458_),
    .B(net569),
    .A_N(_0039_));
 sg13g2_nor2b_1 _3251_ (.A(_0457_),
    .B_N(_0458_),
    .Y(_0459_));
 sg13g2_nand2b_2 _3252_ (.Y(_0460_),
    .B(_0458_),
    .A_N(_0457_));
 sg13g2_nor4_2 _3253_ (.A(net534),
    .B(net501),
    .C(_0445_),
    .Y(_0461_),
    .D(net497));
 sg13g2_nand2b_1 _3254_ (.Y(_0462_),
    .B(_0450_),
    .A_N(net504));
 sg13g2_a22oi_1 _3255_ (.Y(_0463_),
    .B1(_0446_),
    .B2(_0460_),
    .A2(_0444_),
    .A1(_0442_));
 sg13g2_or3_1 _3256_ (.A(_0461_),
    .B(_0462_),
    .C(_0463_),
    .X(_0464_));
 sg13g2_nor2b_1 _3257_ (.A(_0461_),
    .B_N(_0464_),
    .Y(_0465_));
 sg13g2_or2_1 _3258_ (.X(_0466_),
    .B(_0465_),
    .A(_0456_));
 sg13g2_mux2_1 _3259_ (.A0(_0043_),
    .A1(_0042_),
    .S(net536),
    .X(_0467_));
 sg13g2_mux2_2 _3260_ (.A0(_1867_),
    .A1(_1868_),
    .S(net536),
    .X(_0468_));
 sg13g2_mux2_1 _3261_ (.A0(_0030_),
    .A1(_0031_),
    .S(net570),
    .X(_0469_));
 sg13g2_nor2_1 _3262_ (.A(net494),
    .B(net532),
    .Y(_0470_));
 sg13g2_mux2_1 _3263_ (.A0(_0046_),
    .A1(_0047_),
    .S(net570),
    .X(_0471_));
 sg13g2_inv_2 _3264_ (.Y(_0472_),
    .A(net530));
 sg13g2_mux2_1 _3265_ (.A0(_0039_),
    .A1(_0038_),
    .S(net537),
    .X(_0473_));
 sg13g2_mux2_2 _3266_ (.A0(_1861_),
    .A1(_1862_),
    .S(net536),
    .X(_0474_));
 sg13g2_nor2_1 _3267_ (.A(net530),
    .B(net493),
    .Y(_0475_));
 sg13g2_nor2_1 _3268_ (.A(net494),
    .B(net530),
    .Y(_0476_));
 sg13g2_nor2_1 _3269_ (.A(net532),
    .B(net493),
    .Y(_0477_));
 sg13g2_nor2_1 _3270_ (.A(net570),
    .B(_0044_),
    .Y(_0478_));
 sg13g2_nand2b_1 _3271_ (.Y(_0479_),
    .B(net570),
    .A_N(_0045_));
 sg13g2_nor2b_1 _3272_ (.A(_0478_),
    .B_N(_0479_),
    .Y(_0480_));
 sg13g2_nand2b_2 _3273_ (.Y(_0481_),
    .B(_0479_),
    .A_N(_0478_));
 sg13g2_mux2_1 _3274_ (.A0(_0035_),
    .A1(_0034_),
    .S(net536),
    .X(_0482_));
 sg13g2_nor2_1 _3275_ (.A(net491),
    .B(net490),
    .Y(_0483_));
 sg13g2_xor2_1 _3276_ (.B(_0477_),
    .A(_0476_),
    .X(_0484_));
 sg13g2_a22oi_1 _3277_ (.Y(_0485_),
    .B1(_0483_),
    .B2(_0484_),
    .A2(_0475_),
    .A1(_0470_));
 sg13g2_mux2_1 _3278_ (.A0(_0040_),
    .A1(_0041_),
    .S(net570),
    .X(_0486_));
 sg13g2_inv_2 _3279_ (.Y(_0487_),
    .A(net527));
 sg13g2_nor2_1 _3280_ (.A(net489),
    .B(net528),
    .Y(_0488_));
 sg13g2_nor2_1 _3281_ (.A(net493),
    .B(net491),
    .Y(_0489_));
 sg13g2_xnor2_1 _3282_ (.Y(_0490_),
    .A(_0470_),
    .B(_0489_));
 sg13g2_nor3_1 _3283_ (.A(net490),
    .B(net528),
    .C(_0490_),
    .Y(_0491_));
 sg13g2_xor2_1 _3284_ (.B(_0490_),
    .A(_0488_),
    .X(_0492_));
 sg13g2_or2_1 _3285_ (.X(_0493_),
    .B(_0492_),
    .A(_0485_));
 sg13g2_xor2_1 _3286_ (.B(_0492_),
    .A(_0485_),
    .X(_0494_));
 sg13g2_inv_1 _3287_ (.Y(_0495_),
    .A(_0494_));
 sg13g2_nor2_1 _3288_ (.A(net569),
    .B(_0050_),
    .Y(_0496_));
 sg13g2_nand2b_1 _3289_ (.Y(_0497_),
    .B(net569),
    .A_N(_0051_));
 sg13g2_nor2b_2 _3290_ (.A(_0496_),
    .B_N(_0497_),
    .Y(_0498_));
 sg13g2_nand2b_2 _3291_ (.Y(_0499_),
    .B(_0497_),
    .A_N(_0496_));
 sg13g2_nor4_2 _3292_ (.A(net494),
    .B(net530),
    .C(net492),
    .Y(_0500_),
    .D(_0498_));
 sg13g2_or2_1 _3293_ (.X(_0501_),
    .B(net489),
    .A(net531));
 sg13g2_a22oi_1 _3294_ (.Y(_0502_),
    .B1(_0499_),
    .B2(_0468_),
    .A2(_0474_),
    .A1(_0472_));
 sg13g2_or3_1 _3295_ (.A(_0500_),
    .B(_0501_),
    .C(_0502_),
    .X(_0503_));
 sg13g2_nor2b_1 _3296_ (.A(_0500_),
    .B_N(_0503_),
    .Y(_0504_));
 sg13g2_xnor2_1 _3297_ (.Y(_0505_),
    .A(_0483_),
    .B(_0484_));
 sg13g2_or2_1 _3298_ (.X(_0506_),
    .B(_0505_),
    .A(_0504_));
 sg13g2_xnor2_1 _3299_ (.Y(_0507_),
    .A(_0466_),
    .B(_0494_));
 sg13g2_nand2b_1 _3300_ (.Y(_0508_),
    .B(_0507_),
    .A_N(_0506_));
 sg13g2_o21ai_1 _3301_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0466_),
    .A2(_0495_));
 sg13g2_mux2_1 _3302_ (.A0(_0031_),
    .A1(_0030_),
    .S(net537),
    .X(_0510_));
 sg13g2_nor2_1 _3303_ (.A(net569),
    .B(_0034_),
    .Y(_0511_));
 sg13g2_nand2b_1 _3304_ (.Y(_0512_),
    .B(net569),
    .A_N(_0035_));
 sg13g2_nor2b_2 _3305_ (.A(_0511_),
    .B_N(_0512_),
    .Y(_0513_));
 sg13g2_nand2b_2 _3306_ (.Y(_0514_),
    .B(_0512_),
    .A_N(_0511_));
 sg13g2_nor2_1 _3307_ (.A(net487),
    .B(net485),
    .Y(_0515_));
 sg13g2_mux2_1 _3308_ (.A0(_0045_),
    .A1(_0044_),
    .S(net535),
    .X(_0516_));
 sg13g2_mux2_2 _3309_ (.A0(_1869_),
    .A1(_1870_),
    .S(net535),
    .X(_0517_));
 sg13g2_nor2_1 _3310_ (.A(net497),
    .B(net484),
    .Y(_0518_));
 sg13g2_nand2_1 _3311_ (.Y(_0519_),
    .A(_0514_),
    .B(_0517_));
 sg13g2_nor4_2 _3312_ (.A(net497),
    .B(net487),
    .C(net485),
    .Y(_0520_),
    .D(net484));
 sg13g2_or2_1 _3313_ (.X(_0521_),
    .B(net487),
    .A(net496));
 sg13g2_a21oi_1 _3314_ (.A1(_0519_),
    .A2(_0521_),
    .Y(_0522_),
    .B1(_0520_));
 sg13g2_mux2_1 _3315_ (.A0(_0033_),
    .A1(_0032_),
    .S(net536),
    .X(_0523_));
 sg13g2_mux2_1 _3316_ (.A0(_1857_),
    .A1(_1858_),
    .S(net536),
    .X(_0524_));
 sg13g2_nor2_1 _3317_ (.A(net488),
    .B(net482),
    .Y(_0525_));
 sg13g2_and2_1 _3318_ (.A(_0522_),
    .B(_0525_),
    .X(_0526_));
 sg13g2_xnor2_1 _3319_ (.Y(_0527_),
    .A(_0522_),
    .B(_0525_));
 sg13g2_nand2_2 _3320_ (.Y(_0528_),
    .A(_0514_),
    .B(_0524_));
 sg13g2_nor2_2 _3321_ (.A(net502),
    .B(net487),
    .Y(_0529_));
 sg13g2_nor2b_1 _3322_ (.A(_0528_),
    .B_N(_0529_),
    .Y(_0530_));
 sg13g2_nor2b_1 _3323_ (.A(_0527_),
    .B_N(_0530_),
    .Y(_0531_));
 sg13g2_xor2_1 _3324_ (.B(_0465_),
    .A(_0456_),
    .X(_0532_));
 sg13g2_xnor2_1 _3325_ (.Y(_0533_),
    .A(_0527_),
    .B(_0530_));
 sg13g2_a21oi_1 _3326_ (.A1(_0532_),
    .A2(_0533_),
    .Y(_0534_),
    .B1(_0531_));
 sg13g2_or2_1 _3327_ (.X(_0535_),
    .B(net487),
    .A(net534));
 sg13g2_mux2_2 _3328_ (.A0(_0041_),
    .A1(_0040_),
    .S(net535),
    .X(_0536_));
 sg13g2_mux2_2 _3329_ (.A0(_1865_),
    .A1(_1866_),
    .S(net535),
    .X(_0537_));
 sg13g2_nor4_2 _3330_ (.A(net497),
    .B(_0513_),
    .C(net484),
    .Y(_0538_),
    .D(_0536_));
 sg13g2_a22oi_1 _3331_ (.Y(_0539_),
    .B1(_0537_),
    .B2(_0514_),
    .A2(_0517_),
    .A1(_0460_));
 sg13g2_or3_1 _3332_ (.A(_0535_),
    .B(_0538_),
    .C(_0539_),
    .X(_0540_));
 sg13g2_o21ai_1 _3333_ (.B1(_0535_),
    .Y(_0541_),
    .A1(_0538_),
    .A2(_0539_));
 sg13g2_nor2_1 _3334_ (.A(net530),
    .B(net482),
    .Y(_0542_));
 sg13g2_nand3_1 _3335_ (.B(_0541_),
    .C(_0542_),
    .A(_0540_),
    .Y(_0543_));
 sg13g2_a21o_1 _3336_ (.A2(_0541_),
    .A1(_0540_),
    .B1(_0542_),
    .X(_0544_));
 sg13g2_and2_1 _3337_ (.A(_0543_),
    .B(_0544_),
    .X(_0545_));
 sg13g2_nand3_1 _3338_ (.B(_0543_),
    .C(_0544_),
    .A(_0526_),
    .Y(_0546_));
 sg13g2_a21o_1 _3339_ (.A2(_0544_),
    .A1(_0543_),
    .B1(_0526_),
    .X(_0547_));
 sg13g2_a21oi_1 _3340_ (.A1(_0440_),
    .A2(_0454_),
    .Y(_0548_),
    .B1(_0453_));
 sg13g2_nand2b_1 _3341_ (.Y(_0549_),
    .B(_0499_),
    .A_N(net505));
 sg13g2_nor4_2 _3342_ (.A(net503),
    .B(net501),
    .C(net499),
    .Y(_0550_),
    .D(net498));
 sg13g2_a22oi_1 _3343_ (.Y(_0551_),
    .B1(_0446_),
    .B2(_0450_),
    .A2(_0444_),
    .A1(_0439_));
 sg13g2_or3_1 _3344_ (.A(_0549_),
    .B(_0550_),
    .C(_0551_),
    .X(_0552_));
 sg13g2_o21ai_1 _3345_ (.B1(_0549_),
    .Y(_0553_),
    .A1(_0550_),
    .A2(_0551_));
 sg13g2_and3_1 _3346_ (.X(_0554_),
    .A(_0520_),
    .B(_0552_),
    .C(_0553_));
 sg13g2_a21oi_1 _3347_ (.A1(_0552_),
    .A2(_0553_),
    .Y(_0555_),
    .B1(_0520_));
 sg13g2_or3_1 _3348_ (.A(_0548_),
    .B(_0554_),
    .C(_0555_),
    .X(_0556_));
 sg13g2_o21ai_1 _3349_ (.B1(_0548_),
    .Y(_0557_),
    .A1(_0554_),
    .A2(_0555_));
 sg13g2_and4_1 _3350_ (.A(_0546_),
    .B(_0547_),
    .C(_0556_),
    .D(_0557_),
    .X(_0558_));
 sg13g2_a22oi_1 _3351_ (.Y(_0559_),
    .B1(_0556_),
    .B2(_0557_),
    .A2(_0547_),
    .A1(_0546_));
 sg13g2_or3_1 _3352_ (.A(_0534_),
    .B(_0558_),
    .C(_0559_),
    .X(_0560_));
 sg13g2_o21ai_1 _3353_ (.B1(_0534_),
    .Y(_0561_),
    .A1(_0558_),
    .A2(_0559_));
 sg13g2_xnor2_1 _3354_ (.Y(_0562_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_nand3_1 _3355_ (.B(_0561_),
    .C(_0562_),
    .A(_0560_),
    .Y(_0563_));
 sg13g2_and2_1 _3356_ (.A(_0560_),
    .B(_0563_),
    .X(_0564_));
 sg13g2_nand2b_1 _3357_ (.Y(_0565_),
    .B(_0556_),
    .A_N(_0554_));
 sg13g2_a21oi_1 _3358_ (.A1(_0470_),
    .A2(_0489_),
    .Y(_0566_),
    .B1(_0491_));
 sg13g2_mux2_1 _3359_ (.A0(_0036_),
    .A1(_0037_),
    .S(net570),
    .X(_0567_));
 sg13g2_inv_1 _3360_ (.Y(_0568_),
    .A(net525));
 sg13g2_nor2_1 _3361_ (.A(net490),
    .B(net526),
    .Y(_0569_));
 sg13g2_nor2_1 _3362_ (.A(net495),
    .B(net527),
    .Y(_0570_));
 sg13g2_nand2_2 _3363_ (.Y(_0571_),
    .A(_0474_),
    .B(_0487_));
 sg13g2_and2_1 _3364_ (.A(_0489_),
    .B(_0570_),
    .X(_0572_));
 sg13g2_o21ai_1 _3365_ (.B1(_0571_),
    .Y(_0573_),
    .A1(net495),
    .A2(net491));
 sg13g2_nand2b_1 _3366_ (.Y(_0574_),
    .B(_0573_),
    .A_N(_0572_));
 sg13g2_xor2_1 _3367_ (.B(_0574_),
    .A(_0569_),
    .X(_0575_));
 sg13g2_or2_1 _3368_ (.X(_0576_),
    .B(_0575_),
    .A(_0566_));
 sg13g2_xor2_1 _3369_ (.B(_0575_),
    .A(_0566_),
    .X(_0577_));
 sg13g2_nand2_1 _3370_ (.Y(_0578_),
    .A(_0565_),
    .B(_0577_));
 sg13g2_xnor2_1 _3371_ (.Y(_0579_),
    .A(_0565_),
    .B(_0577_));
 sg13g2_xor2_1 _3372_ (.B(_0579_),
    .A(_0493_),
    .X(_0580_));
 sg13g2_a21oi_2 _3373_ (.B1(_0558_),
    .Y(_0581_),
    .A2(_0545_),
    .A1(_0526_));
 sg13g2_nor2b_1 _3374_ (.A(_0550_),
    .B_N(_0552_),
    .Y(_0582_));
 sg13g2_nor2b_1 _3375_ (.A(_0538_),
    .B_N(_0540_),
    .Y(_0583_));
 sg13g2_nor2_1 _3376_ (.A(net505),
    .B(net529),
    .Y(_0584_));
 sg13g2_nor2_1 _3377_ (.A(net501),
    .B(_0498_),
    .Y(_0585_));
 sg13g2_nor4_1 _3378_ (.A(net503),
    .B(net501),
    .C(net499),
    .D(_0498_),
    .Y(_0586_));
 sg13g2_a22oi_1 _3379_ (.Y(_0587_),
    .B1(_0499_),
    .B2(_0444_),
    .A2(_0446_),
    .A1(_0439_));
 sg13g2_nor2_1 _3380_ (.A(_0586_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_xnor2_1 _3381_ (.Y(_0589_),
    .A(_0584_),
    .B(_0588_));
 sg13g2_or2_1 _3382_ (.X(_0590_),
    .B(_0589_),
    .A(_0583_));
 sg13g2_xnor2_1 _3383_ (.Y(_0591_),
    .A(_0583_),
    .B(_0589_));
 sg13g2_xor2_1 _3384_ (.B(_0591_),
    .A(_0582_),
    .X(_0592_));
 sg13g2_nor2_1 _3385_ (.A(_0449_),
    .B(net486),
    .Y(_0593_));
 sg13g2_nor2_2 _3386_ (.A(net534),
    .B(net477),
    .Y(_0594_));
 sg13g2_nor2_1 _3387_ (.A(net534),
    .B(net484),
    .Y(_0595_));
 sg13g2_a22oi_1 _3388_ (.Y(_0596_),
    .B1(_0537_),
    .B2(_0460_),
    .A2(_0517_),
    .A1(_0442_));
 sg13g2_a21oi_1 _3389_ (.A1(_0518_),
    .A2(_0594_),
    .Y(_0597_),
    .B1(_0596_));
 sg13g2_xnor2_1 _3390_ (.Y(_0598_),
    .A(_0593_),
    .B(_0597_));
 sg13g2_mux2_1 _3391_ (.A0(_0037_),
    .A1(_0036_),
    .S(net535),
    .X(_0599_));
 sg13g2_inv_1 _3392_ (.Y(_0600_),
    .A(net475));
 sg13g2_or2_1 _3393_ (.X(_0601_),
    .B(net476),
    .A(net531));
 sg13g2_nor2_1 _3394_ (.A(net531),
    .B(net482),
    .Y(_0602_));
 sg13g2_nor2_2 _3395_ (.A(_0528_),
    .B(_0601_),
    .Y(_0603_));
 sg13g2_a21oi_1 _3396_ (.A1(_0514_),
    .A2(_0600_),
    .Y(_0604_),
    .B1(_0602_));
 sg13g2_nor2_2 _3397_ (.A(_0603_),
    .B(_0604_),
    .Y(_0605_));
 sg13g2_nand2b_1 _3398_ (.Y(_0606_),
    .B(_0605_),
    .A_N(_0598_));
 sg13g2_xnor2_1 _3399_ (.Y(_0607_),
    .A(_0598_),
    .B(_0605_));
 sg13g2_nor2b_1 _3400_ (.A(_0543_),
    .B_N(_0607_),
    .Y(_0608_));
 sg13g2_xnor2_1 _3401_ (.Y(_0609_),
    .A(_0543_),
    .B(_0607_));
 sg13g2_xnor2_1 _3402_ (.Y(_0610_),
    .A(_0592_),
    .B(_0609_));
 sg13g2_nor2_1 _3403_ (.A(_0581_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_xor2_1 _3404_ (.B(_0610_),
    .A(_0581_),
    .X(_0612_));
 sg13g2_xnor2_1 _3405_ (.Y(_0613_),
    .A(_0580_),
    .B(_0612_));
 sg13g2_nor2_1 _3406_ (.A(_0564_),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_xor2_1 _3407_ (.B(_0613_),
    .A(_0564_),
    .X(_0615_));
 sg13g2_xor2_1 _3408_ (.B(_0615_),
    .A(_0509_),
    .X(_0616_));
 sg13g2_a21oi_1 _3409_ (.A1(_0439_),
    .A2(net480),
    .Y(_0617_),
    .B1(_0515_));
 sg13g2_or2_1 _3410_ (.X(_0618_),
    .B(_0617_),
    .A(_0530_));
 sg13g2_o21ai_1 _3411_ (.B1(_0462_),
    .Y(_0619_),
    .A1(_0461_),
    .A2(_0463_));
 sg13g2_nand2_1 _3412_ (.Y(_0620_),
    .A(_0444_),
    .B(_0514_));
 sg13g2_nor4_2 _3413_ (.A(net500),
    .B(_0445_),
    .C(net497),
    .Y(_0621_),
    .D(net485));
 sg13g2_nand4_1 _3414_ (.B(_0446_),
    .C(_0460_),
    .A(_0444_),
    .Y(_0622_),
    .D(_0514_));
 sg13g2_nand2b_1 _3415_ (.Y(_0623_),
    .B(_0442_),
    .A_N(net504));
 sg13g2_a22oi_1 _3416_ (.Y(_0624_),
    .B1(_0514_),
    .B2(_0446_),
    .A2(_0460_),
    .A1(_0444_));
 sg13g2_or3_1 _3417_ (.A(_0621_),
    .B(_0623_),
    .C(_0624_),
    .X(_0625_));
 sg13g2_o21ai_1 _3418_ (.B1(_0622_),
    .Y(_0626_),
    .A1(_0623_),
    .A2(_0624_));
 sg13g2_and3_1 _3419_ (.X(_0627_),
    .A(_0464_),
    .B(_0619_),
    .C(_0626_));
 sg13g2_a21oi_1 _3420_ (.A1(_0464_),
    .A2(_0619_),
    .Y(_0628_),
    .B1(_0626_));
 sg13g2_or3_2 _3421_ (.A(_0618_),
    .B(_0627_),
    .C(_0628_),
    .X(_0629_));
 sg13g2_xnor2_1 _3422_ (.Y(_0630_),
    .A(_0532_),
    .B(_0533_));
 sg13g2_nor2_1 _3423_ (.A(_0629_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_nand2_1 _3424_ (.Y(_0632_),
    .A(_0629_),
    .B(_0630_));
 sg13g2_xnor2_1 _3425_ (.Y(_0633_),
    .A(_0629_),
    .B(_0630_));
 sg13g2_nor4_1 _3426_ (.A(net502),
    .B(net494),
    .C(net492),
    .D(net488),
    .Y(_0634_));
 sg13g2_nand4_1 _3427_ (.B(_0468_),
    .C(_0474_),
    .A(_0439_),
    .Y(_0635_),
    .D(_0499_));
 sg13g2_or2_1 _3428_ (.X(_0636_),
    .B(net489),
    .A(net529));
 sg13g2_a22oi_1 _3429_ (.Y(_0637_),
    .B1(_0474_),
    .B2(_0499_),
    .A2(_0468_),
    .A1(_0439_));
 sg13g2_nor3_1 _3430_ (.A(_0634_),
    .B(_0636_),
    .C(_0637_),
    .Y(_0638_));
 sg13g2_o21ai_1 _3431_ (.B1(_0635_),
    .Y(_0639_),
    .A1(_0636_),
    .A2(_0637_));
 sg13g2_o21ai_1 _3432_ (.B1(_0501_),
    .Y(_0640_),
    .A1(_0500_),
    .A2(_0502_));
 sg13g2_nand3_1 _3433_ (.B(_0639_),
    .C(_0640_),
    .A(_0503_),
    .Y(_0641_));
 sg13g2_xor2_1 _3434_ (.B(_0505_),
    .A(_0504_),
    .X(_0642_));
 sg13g2_xor2_1 _3435_ (.B(_0642_),
    .A(_0627_),
    .X(_0643_));
 sg13g2_nor2b_1 _3436_ (.A(_0641_),
    .B_N(_0643_),
    .Y(_0644_));
 sg13g2_xnor2_1 _3437_ (.Y(_0645_),
    .A(_0641_),
    .B(_0643_));
 sg13g2_a21o_1 _3438_ (.A2(_0645_),
    .A1(_0632_),
    .B1(_0631_),
    .X(_0646_));
 sg13g2_a21o_1 _3439_ (.A2(_0561_),
    .A1(_0560_),
    .B1(_0562_),
    .X(_0647_));
 sg13g2_nand3_1 _3440_ (.B(_0646_),
    .C(_0647_),
    .A(_0563_),
    .Y(_0648_));
 sg13g2_a21oi_1 _3441_ (.A1(_0627_),
    .A2(_0642_),
    .Y(_0649_),
    .B1(_0644_));
 sg13g2_inv_1 _3442_ (.Y(_0650_),
    .A(_0649_));
 sg13g2_a21oi_1 _3443_ (.A1(_0563_),
    .A2(_0647_),
    .Y(_0651_),
    .B1(_0646_));
 sg13g2_a21o_1 _3444_ (.A2(_0647_),
    .A1(_0563_),
    .B1(_0646_),
    .X(_0652_));
 sg13g2_and3_1 _3445_ (.X(_0653_),
    .A(_0648_),
    .B(_0650_),
    .C(_0652_));
 sg13g2_o21ai_1 _3446_ (.B1(_0648_),
    .Y(_0654_),
    .A1(_0649_),
    .A2(_0651_));
 sg13g2_nand2_1 _3447_ (.Y(_0655_),
    .A(_0616_),
    .B(_0654_));
 sg13g2_xor2_1 _3448_ (.B(_0654_),
    .A(_0616_),
    .X(_0656_));
 sg13g2_xnor2_1 _3449_ (.Y(_0657_),
    .A(_0616_),
    .B(_0654_));
 sg13g2_nor2_1 _3450_ (.A(net504),
    .B(net485),
    .Y(_0658_));
 sg13g2_nor3_2 _3451_ (.A(net504),
    .B(net496),
    .C(_0620_),
    .Y(_0659_));
 sg13g2_o21ai_1 _3452_ (.B1(_0623_),
    .Y(_0660_),
    .A1(_0621_),
    .A2(_0624_));
 sg13g2_and3_1 _3453_ (.X(_0661_),
    .A(_0625_),
    .B(_0659_),
    .C(_0660_));
 sg13g2_nand3_1 _3454_ (.B(_0659_),
    .C(_0660_),
    .A(_0625_),
    .Y(_0662_));
 sg13g2_a21o_1 _3455_ (.A2(_0660_),
    .A1(_0625_),
    .B1(_0659_),
    .X(_0663_));
 sg13g2_and4_2 _3456_ (.A(_0450_),
    .B(net480),
    .C(_0662_),
    .D(_0663_),
    .X(_0664_));
 sg13g2_o21ai_1 _3457_ (.B1(_0618_),
    .Y(_0665_),
    .A1(_0627_),
    .A2(_0628_));
 sg13g2_nand3_1 _3458_ (.B(_0664_),
    .C(_0665_),
    .A(_0629_),
    .Y(_0666_));
 sg13g2_a21o_1 _3459_ (.A2(_0665_),
    .A1(_0629_),
    .B1(_0664_),
    .X(_0667_));
 sg13g2_o21ai_1 _3460_ (.B1(_0636_),
    .Y(_0668_),
    .A1(_0634_),
    .A2(_0637_));
 sg13g2_nor2b_1 _3461_ (.A(_0638_),
    .B_N(_0668_),
    .Y(_0669_));
 sg13g2_nor2_1 _3462_ (.A(net498),
    .B(net492),
    .Y(_0670_));
 sg13g2_nor4_2 _3463_ (.A(net502),
    .B(net498),
    .C(net494),
    .Y(_0671_),
    .D(net492));
 sg13g2_nand2b_1 _3464_ (.Y(_0672_),
    .B(_0499_),
    .A_N(net489));
 sg13g2_a22oi_1 _3465_ (.Y(_0673_),
    .B1(_0474_),
    .B2(_0439_),
    .A2(_0468_),
    .A1(_0450_));
 sg13g2_nor3_1 _3466_ (.A(_0671_),
    .B(_0672_),
    .C(_0673_),
    .Y(_0674_));
 sg13g2_nor2_1 _3467_ (.A(_0671_),
    .B(_0674_),
    .Y(_0675_));
 sg13g2_nand2b_1 _3468_ (.Y(_0676_),
    .B(_0669_),
    .A_N(_0675_));
 sg13g2_a21o_1 _3469_ (.A2(_0640_),
    .A1(_0503_),
    .B1(_0639_),
    .X(_0677_));
 sg13g2_and3_1 _3470_ (.X(_0678_),
    .A(_0641_),
    .B(_0661_),
    .C(_0677_));
 sg13g2_a21oi_1 _3471_ (.A1(_0641_),
    .A2(_0677_),
    .Y(_0679_),
    .B1(_0661_));
 sg13g2_or3_1 _3472_ (.A(_0676_),
    .B(_0678_),
    .C(_0679_),
    .X(_0680_));
 sg13g2_o21ai_1 _3473_ (.B1(_0676_),
    .Y(_0681_),
    .A1(_0678_),
    .A2(_0679_));
 sg13g2_and4_1 _3474_ (.A(_0666_),
    .B(_0667_),
    .C(_0680_),
    .D(_0681_),
    .X(_0682_));
 sg13g2_nand4_1 _3475_ (.B(_0667_),
    .C(_0680_),
    .A(_0666_),
    .Y(_0683_),
    .D(_0681_));
 sg13g2_nand2_1 _3476_ (.Y(_0684_),
    .A(_0666_),
    .B(_0683_));
 sg13g2_xnor2_1 _3477_ (.Y(_0685_),
    .A(_0633_),
    .B(_0645_));
 sg13g2_and2_1 _3478_ (.A(_0684_),
    .B(_0685_),
    .X(_0686_));
 sg13g2_nor2b_1 _3479_ (.A(_0678_),
    .B_N(_0680_),
    .Y(_0687_));
 sg13g2_inv_1 _3480_ (.Y(_0688_),
    .A(_0687_));
 sg13g2_xor2_1 _3481_ (.B(_0685_),
    .A(_0684_),
    .X(_0689_));
 sg13g2_a21oi_1 _3482_ (.A1(_0688_),
    .A2(_0689_),
    .Y(_0690_),
    .B1(_0686_));
 sg13g2_a21oi_1 _3483_ (.A1(_0648_),
    .A2(_0652_),
    .Y(_0691_),
    .B1(_0650_));
 sg13g2_o21ai_1 _3484_ (.B1(_0690_),
    .Y(_0692_),
    .A1(_0653_),
    .A2(_0691_));
 sg13g2_nor2_1 _3485_ (.A(net533),
    .B(net492),
    .Y(_0693_));
 sg13g2_nor2_2 _3486_ (.A(net533),
    .B(net494),
    .Y(_0694_));
 sg13g2_and2_1 _3487_ (.A(_0670_),
    .B(_0694_),
    .X(_0695_));
 sg13g2_nor2_1 _3488_ (.A(net502),
    .B(net489),
    .Y(_0696_));
 sg13g2_or2_1 _3489_ (.X(_0697_),
    .B(_0694_),
    .A(_0670_));
 sg13g2_xnor2_1 _3490_ (.Y(_0698_),
    .A(_0670_),
    .B(_0694_));
 sg13g2_a21oi_1 _3491_ (.A1(_0696_),
    .A2(_0697_),
    .Y(_0699_),
    .B1(_0695_));
 sg13g2_o21ai_1 _3492_ (.B1(_0672_),
    .Y(_0700_),
    .A1(_0671_),
    .A2(_0673_));
 sg13g2_nor2b_1 _3493_ (.A(_0674_),
    .B_N(_0700_),
    .Y(_0701_));
 sg13g2_nand2b_1 _3494_ (.Y(_0702_),
    .B(_0701_),
    .A_N(_0699_));
 sg13g2_xnor2_1 _3495_ (.Y(_0703_),
    .A(_0669_),
    .B(_0675_));
 sg13g2_nor2b_1 _3496_ (.A(_0702_),
    .B_N(_0703_),
    .Y(_0704_));
 sg13g2_xnor2_1 _3497_ (.Y(_0705_),
    .A(_0702_),
    .B(_0703_));
 sg13g2_nor2_1 _3498_ (.A(net533),
    .B(net482),
    .Y(_0706_));
 sg13g2_nand2b_1 _3499_ (.Y(_0707_),
    .B(_0460_),
    .A_N(net504));
 sg13g2_a21oi_1 _3500_ (.A1(_0620_),
    .A2(_0707_),
    .Y(_0708_),
    .B1(_0659_));
 sg13g2_nand2_1 _3501_ (.Y(_0709_),
    .A(_0706_),
    .B(_0708_));
 sg13g2_a22oi_1 _3502_ (.Y(_0710_),
    .B1(_0662_),
    .B2(_0663_),
    .A2(net480),
    .A1(_0450_));
 sg13g2_nor3_1 _3503_ (.A(_0664_),
    .B(_0709_),
    .C(_0710_),
    .Y(_0711_));
 sg13g2_or3_1 _3504_ (.A(_0664_),
    .B(_0709_),
    .C(_0710_),
    .X(_0712_));
 sg13g2_o21ai_1 _3505_ (.B1(_0709_),
    .Y(_0713_),
    .A1(_0664_),
    .A2(_0710_));
 sg13g2_nand3_1 _3506_ (.B(_0712_),
    .C(_0713_),
    .A(_0705_),
    .Y(_0714_));
 sg13g2_a21o_1 _3507_ (.A2(_0713_),
    .A1(_0712_),
    .B1(_0705_),
    .X(_0715_));
 sg13g2_xnor2_1 _3508_ (.Y(_0716_),
    .A(_0706_),
    .B(_0708_));
 sg13g2_nor2_1 _3509_ (.A(_0528_),
    .B(_0707_),
    .Y(_0717_));
 sg13g2_nor2b_1 _3510_ (.A(_0716_),
    .B_N(_0717_),
    .Y(_0718_));
 sg13g2_xnor2_1 _3511_ (.Y(_0719_),
    .A(_0696_),
    .B(_0698_));
 sg13g2_nor2_1 _3512_ (.A(net496),
    .B(net492),
    .Y(_0720_));
 sg13g2_nor2_1 _3513_ (.A(net496),
    .B(net494),
    .Y(_0721_));
 sg13g2_nor2_1 _3514_ (.A(net498),
    .B(net489),
    .Y(_0722_));
 sg13g2_xor2_1 _3515_ (.B(_0721_),
    .A(_0693_),
    .X(_0723_));
 sg13g2_a22oi_1 _3516_ (.Y(_0724_),
    .B1(_0722_),
    .B2(_0723_),
    .A2(_0720_),
    .A1(_0694_));
 sg13g2_nand2b_1 _3517_ (.Y(_0725_),
    .B(_0719_),
    .A_N(_0724_));
 sg13g2_xnor2_1 _3518_ (.Y(_0726_),
    .A(_0699_),
    .B(_0701_));
 sg13g2_nand2b_1 _3519_ (.Y(_0727_),
    .B(_0726_),
    .A_N(_0725_));
 sg13g2_xnor2_1 _3520_ (.Y(_0728_),
    .A(_0725_),
    .B(_0726_));
 sg13g2_xnor2_1 _3521_ (.Y(_0729_),
    .A(_0716_),
    .B(_0717_));
 sg13g2_a21o_1 _3522_ (.A2(_0729_),
    .A1(_0728_),
    .B1(_0718_),
    .X(_0730_));
 sg13g2_and3_1 _3523_ (.X(_0731_),
    .A(_0714_),
    .B(_0715_),
    .C(_0730_));
 sg13g2_nand3_1 _3524_ (.B(_0715_),
    .C(_0730_),
    .A(_0714_),
    .Y(_0732_));
 sg13g2_a21oi_1 _3525_ (.A1(_0714_),
    .A2(_0715_),
    .Y(_0733_),
    .B1(_0730_));
 sg13g2_or3_1 _3526_ (.A(_0727_),
    .B(_0731_),
    .C(_0733_),
    .X(_0734_));
 sg13g2_o21ai_1 _3527_ (.B1(_0732_),
    .Y(_0735_),
    .A1(_0727_),
    .A2(_0733_));
 sg13g2_a21oi_1 _3528_ (.A1(_0705_),
    .A2(_0713_),
    .Y(_0736_),
    .B1(_0711_));
 sg13g2_a22oi_1 _3529_ (.Y(_0737_),
    .B1(_0680_),
    .B2(_0681_),
    .A2(_0667_),
    .A1(_0666_));
 sg13g2_or3_1 _3530_ (.A(_0682_),
    .B(_0736_),
    .C(_0737_),
    .X(_0738_));
 sg13g2_o21ai_1 _3531_ (.B1(_0736_),
    .Y(_0739_),
    .A1(_0682_),
    .A2(_0737_));
 sg13g2_nand3_1 _3532_ (.B(_0738_),
    .C(_0739_),
    .A(_0704_),
    .Y(_0740_));
 sg13g2_a21o_1 _3533_ (.A2(_0739_),
    .A1(_0738_),
    .B1(_0704_),
    .X(_0741_));
 sg13g2_nand3_1 _3534_ (.B(_0740_),
    .C(_0741_),
    .A(_0735_),
    .Y(_0742_));
 sg13g2_o21ai_1 _3535_ (.B1(_0727_),
    .Y(_0743_),
    .A1(_0731_),
    .A2(_0733_));
 sg13g2_a21oi_1 _3536_ (.A1(_0460_),
    .A2(net480),
    .Y(_0744_),
    .B1(_0658_));
 sg13g2_nor2_1 _3537_ (.A(_0717_),
    .B(_0744_),
    .Y(_0745_));
 sg13g2_xnor2_1 _3538_ (.Y(_0746_),
    .A(_0719_),
    .B(_0724_));
 sg13g2_nand2_1 _3539_ (.Y(_0747_),
    .A(_0745_),
    .B(_0746_));
 sg13g2_xor2_1 _3540_ (.B(_0729_),
    .A(_0728_),
    .X(_0748_));
 sg13g2_xnor2_1 _3541_ (.Y(_0749_),
    .A(_0722_),
    .B(_0723_));
 sg13g2_nor2_1 _3542_ (.A(net533),
    .B(net489),
    .Y(_0750_));
 sg13g2_nand2_1 _3543_ (.Y(_0751_),
    .A(_0720_),
    .B(_0750_));
 sg13g2_o21ai_1 _3544_ (.B1(_0751_),
    .Y(_0752_),
    .A1(net494),
    .A2(net485));
 sg13g2_o21ai_1 _3545_ (.B1(_0752_),
    .Y(_0753_),
    .A1(_0720_),
    .A2(_0750_));
 sg13g2_or2_1 _3546_ (.X(_0754_),
    .B(_0753_),
    .A(_0749_));
 sg13g2_nor4_1 _3547_ (.A(net496),
    .B(net492),
    .C(net489),
    .D(net485),
    .Y(_0755_));
 sg13g2_nand2b_1 _3548_ (.Y(_0756_),
    .B(_0755_),
    .A_N(_0723_));
 sg13g2_nand3_1 _3549_ (.B(_0754_),
    .C(_0756_),
    .A(_0528_),
    .Y(_0757_));
 sg13g2_nand2b_1 _3550_ (.Y(_0758_),
    .B(net480),
    .A_N(_0756_));
 sg13g2_nand3_1 _3551_ (.B(_0753_),
    .C(_0758_),
    .A(_0749_),
    .Y(_0759_));
 sg13g2_nand3_1 _3552_ (.B(_0757_),
    .C(_0759_),
    .A(_0748_),
    .Y(_0760_));
 sg13g2_nand2_1 _3553_ (.Y(_0761_),
    .A(_0747_),
    .B(_0760_));
 sg13g2_o21ai_1 _3554_ (.B1(_0748_),
    .Y(_0762_),
    .A1(_0745_),
    .A2(_0746_));
 sg13g2_o21ai_1 _3555_ (.B1(_0762_),
    .Y(_0763_),
    .A1(_0754_),
    .A2(_0758_));
 sg13g2_nand4_1 _3556_ (.B(_0743_),
    .C(_0761_),
    .A(_0734_),
    .Y(_0764_),
    .D(_0763_));
 sg13g2_a21oi_1 _3557_ (.A1(_0740_),
    .A2(_0741_),
    .Y(_0765_),
    .B1(_0735_));
 sg13g2_and2_1 _3558_ (.A(_0738_),
    .B(_0740_),
    .X(_0766_));
 sg13g2_xnor2_1 _3559_ (.Y(_0767_),
    .A(_0688_),
    .B(_0689_));
 sg13g2_a221oi_1 _3560_ (.B2(_0767_),
    .C1(_0765_),
    .B1(_0766_),
    .A1(_0742_),
    .Y(_0768_),
    .A2(_0764_));
 sg13g2_or3_1 _3561_ (.A(_0653_),
    .B(_0690_),
    .C(_0691_),
    .X(_0769_));
 sg13g2_nor2_1 _3562_ (.A(_0766_),
    .B(_0767_),
    .Y(_0770_));
 sg13g2_o21ai_1 _3563_ (.B1(_0692_),
    .Y(_0771_),
    .A1(_0768_),
    .A2(_0770_));
 sg13g2_nand2_1 _3564_ (.Y(_0772_),
    .A(_0769_),
    .B(_0771_));
 sg13g2_nand2_1 _3565_ (.Y(_0773_),
    .A(_0656_),
    .B(_0772_));
 sg13g2_xnor2_1 _3566_ (.Y(_0774_),
    .A(_0656_),
    .B(_0772_));
 sg13g2_nor2_1 _3567_ (.A(net786),
    .B(net540),
    .Y(_0775_));
 sg13g2_a21oi_1 _3568_ (.A1(net540),
    .A2(_0774_),
    .Y(_0126_),
    .B1(_0775_));
 sg13g2_nor2_1 _3569_ (.A(net770),
    .B(net540),
    .Y(_0776_));
 sg13g2_nand2_1 _3570_ (.Y(_0777_),
    .A(_0655_),
    .B(_0773_));
 sg13g2_a21oi_1 _3571_ (.A1(_0509_),
    .A2(_0615_),
    .Y(_0778_),
    .B1(_0614_));
 sg13g2_a21o_1 _3572_ (.A2(_0615_),
    .A1(_0509_),
    .B1(_0614_),
    .X(_0779_));
 sg13g2_o21ai_1 _3573_ (.B1(_0578_),
    .Y(_0780_),
    .A1(_0493_),
    .A2(_0579_));
 sg13g2_a21oi_2 _3574_ (.B1(_0611_),
    .Y(_0781_),
    .A2(_0612_),
    .A1(_0580_));
 sg13g2_o21ai_1 _3575_ (.B1(_0590_),
    .Y(_0782_),
    .A1(_0582_),
    .A2(_0591_));
 sg13g2_a21oi_1 _3576_ (.A1(_0569_),
    .A2(_0573_),
    .Y(_0783_),
    .B1(_0572_));
 sg13g2_nor2_1 _3577_ (.A(net570),
    .B(_0052_),
    .Y(_0784_));
 sg13g2_nand2b_1 _3578_ (.Y(_0785_),
    .B(net570),
    .A_N(_0053_));
 sg13g2_nor2b_1 _3579_ (.A(_0784_),
    .B_N(_0785_),
    .Y(_0786_));
 sg13g2_nand2b_2 _3580_ (.Y(_0787_),
    .B(_0785_),
    .A_N(_0784_));
 sg13g2_nor2_2 _3581_ (.A(net490),
    .B(net474),
    .Y(_0788_));
 sg13g2_nor2_1 _3582_ (.A(net495),
    .B(net526),
    .Y(_0789_));
 sg13g2_nor2_1 _3583_ (.A(net493),
    .B(net526),
    .Y(_0790_));
 sg13g2_xnor2_1 _3584_ (.Y(_0791_),
    .A(_0570_),
    .B(_0790_));
 sg13g2_nor3_1 _3585_ (.A(net490),
    .B(net474),
    .C(_0791_),
    .Y(_0792_));
 sg13g2_xor2_1 _3586_ (.B(_0791_),
    .A(_0788_),
    .X(_0793_));
 sg13g2_xor2_1 _3587_ (.B(_0793_),
    .A(_0783_),
    .X(_0794_));
 sg13g2_mux2_1 _3588_ (.A0(_0053_),
    .A1(_0052_),
    .S(net535),
    .X(_0795_));
 sg13g2_mux2_1 _3589_ (.A0(_1876_),
    .A1(_1877_),
    .S(net535),
    .X(_0796_));
 sg13g2_nand2_1 _3590_ (.Y(_0797_),
    .A(_0794_),
    .B(_0796_));
 sg13g2_xnor2_1 _3591_ (.Y(_0798_),
    .A(_0794_),
    .B(net470));
 sg13g2_nand2_1 _3592_ (.Y(_0799_),
    .A(_0782_),
    .B(_0798_));
 sg13g2_xnor2_1 _3593_ (.Y(_0800_),
    .A(_0782_),
    .B(_0798_));
 sg13g2_xor2_1 _3594_ (.B(_0800_),
    .A(_0576_),
    .X(_0801_));
 sg13g2_a21oi_2 _3595_ (.B1(_0608_),
    .Y(_0802_),
    .A2(_0609_),
    .A1(_0592_));
 sg13g2_a21oi_1 _3596_ (.A1(_0584_),
    .A2(_0588_),
    .Y(_0803_),
    .B1(_0586_));
 sg13g2_a22oi_1 _3597_ (.Y(_0804_),
    .B1(_0597_),
    .B2(_0593_),
    .A2(_0594_),
    .A1(_0518_));
 sg13g2_nor2_1 _3598_ (.A(net505),
    .B(net532),
    .Y(_0805_));
 sg13g2_nor2_2 _3599_ (.A(net499),
    .B(net530),
    .Y(_0806_));
 sg13g2_nor2_1 _3600_ (.A(net500),
    .B(net529),
    .Y(_0807_));
 sg13g2_a22oi_1 _3601_ (.Y(_0808_),
    .B1(_0499_),
    .B2(_0446_),
    .A2(_0472_),
    .A1(_0444_));
 sg13g2_a21oi_1 _3602_ (.A1(_0585_),
    .A2(_0806_),
    .Y(_0809_),
    .B1(_0808_));
 sg13g2_xnor2_1 _3603_ (.Y(_0810_),
    .A(_0805_),
    .B(_0809_));
 sg13g2_or2_1 _3604_ (.X(_0811_),
    .B(_0810_),
    .A(_0804_));
 sg13g2_and2_1 _3605_ (.A(_0804_),
    .B(_0810_),
    .X(_0812_));
 sg13g2_xor2_1 _3606_ (.B(_0810_),
    .A(_0804_),
    .X(_0813_));
 sg13g2_xnor2_1 _3607_ (.Y(_0814_),
    .A(_0803_),
    .B(_0813_));
 sg13g2_nor2_1 _3608_ (.A(_0449_),
    .B(_0536_),
    .Y(_0815_));
 sg13g2_nor2_2 _3609_ (.A(_0449_),
    .B(net483),
    .Y(_0816_));
 sg13g2_xor2_1 _3610_ (.B(_0816_),
    .A(_0594_),
    .X(_0817_));
 sg13g2_xnor2_1 _3611_ (.Y(_0818_),
    .A(_0594_),
    .B(_0816_));
 sg13g2_xnor2_1 _3612_ (.Y(_0819_),
    .A(_0529_),
    .B(_0818_));
 sg13g2_xnor2_1 _3613_ (.Y(_0820_),
    .A(_0529_),
    .B(_0817_));
 sg13g2_or2_1 _3614_ (.X(_0821_),
    .B(net476),
    .A(net496));
 sg13g2_nor4_1 _3615_ (.A(net491),
    .B(_0514_),
    .C(net481),
    .D(net470),
    .Y(_0822_));
 sg13g2_nand4_1 _3616_ (.B(net485),
    .C(net478),
    .A(_0481_),
    .Y(_0823_),
    .D(net468));
 sg13g2_a22oi_1 _3617_ (.Y(_0824_),
    .B1(net468),
    .B2(net485),
    .A2(net478),
    .A1(_0481_));
 sg13g2_or3_1 _3618_ (.A(_0821_),
    .B(_0822_),
    .C(_0824_),
    .X(_0825_));
 sg13g2_o21ai_1 _3619_ (.B1(_0821_),
    .Y(_0826_),
    .A1(_0822_),
    .A2(_0824_));
 sg13g2_nand3_1 _3620_ (.B(_0825_),
    .C(_0826_),
    .A(_0603_),
    .Y(_0827_));
 sg13g2_a21oi_1 _3621_ (.A1(_0825_),
    .A2(_0826_),
    .Y(_0828_),
    .B1(_0603_));
 sg13g2_a21o_1 _3622_ (.A2(_0826_),
    .A1(_0825_),
    .B1(_0603_),
    .X(_0829_));
 sg13g2_and3_1 _3623_ (.X(_0830_),
    .A(_0819_),
    .B(_0827_),
    .C(_0829_));
 sg13g2_a21oi_2 _3624_ (.B1(_0819_),
    .Y(_0831_),
    .A2(_0829_),
    .A1(_0827_));
 sg13g2_nor3_1 _3625_ (.A(_0606_),
    .B(_0830_),
    .C(_0831_),
    .Y(_0832_));
 sg13g2_or3_1 _3626_ (.A(_0606_),
    .B(_0830_),
    .C(_0831_),
    .X(_0833_));
 sg13g2_o21ai_1 _3627_ (.B1(_0606_),
    .Y(_0834_),
    .A1(_0830_),
    .A2(_0831_));
 sg13g2_and3_1 _3628_ (.X(_0835_),
    .A(_0814_),
    .B(_0833_),
    .C(_0834_));
 sg13g2_a21oi_2 _3629_ (.B1(_0814_),
    .Y(_0836_),
    .A2(_0834_),
    .A1(_0833_));
 sg13g2_nor3_1 _3630_ (.A(_0802_),
    .B(_0835_),
    .C(_0836_),
    .Y(_0837_));
 sg13g2_or3_1 _3631_ (.A(_0802_),
    .B(_0835_),
    .C(_0836_),
    .X(_0838_));
 sg13g2_o21ai_1 _3632_ (.B1(_0802_),
    .Y(_0839_),
    .A1(_0835_),
    .A2(_0836_));
 sg13g2_and3_1 _3633_ (.X(_0840_),
    .A(_0801_),
    .B(_0838_),
    .C(_0839_));
 sg13g2_a21oi_1 _3634_ (.A1(_0838_),
    .A2(_0839_),
    .Y(_0841_),
    .B1(_0801_));
 sg13g2_nor3_1 _3635_ (.A(_0781_),
    .B(_0840_),
    .C(_0841_),
    .Y(_0842_));
 sg13g2_or3_1 _3636_ (.A(_0781_),
    .B(_0840_),
    .C(_0841_),
    .X(_0843_));
 sg13g2_o21ai_1 _3637_ (.B1(_0781_),
    .Y(_0844_),
    .A1(_0840_),
    .A2(_0841_));
 sg13g2_nand3_1 _3638_ (.B(_0843_),
    .C(_0844_),
    .A(_0780_),
    .Y(_0845_));
 sg13g2_a21o_1 _3639_ (.A2(_0844_),
    .A1(_0843_),
    .B1(_0780_),
    .X(_0846_));
 sg13g2_a21oi_1 _3640_ (.A1(_0845_),
    .A2(_0846_),
    .Y(_0847_),
    .B1(_0779_));
 sg13g2_nand3_1 _3641_ (.B(_0845_),
    .C(_0846_),
    .A(_0779_),
    .Y(_0848_));
 sg13g2_a21o_1 _3642_ (.A2(_0846_),
    .A1(_0845_),
    .B1(_0778_),
    .X(_0849_));
 sg13g2_nand3_1 _3643_ (.B(_0845_),
    .C(_0846_),
    .A(_0778_),
    .Y(_0850_));
 sg13g2_nand2_1 _3644_ (.Y(_0851_),
    .A(_0849_),
    .B(_0850_));
 sg13g2_xnor2_1 _3645_ (.Y(_0852_),
    .A(_0777_),
    .B(_0851_));
 sg13g2_a21oi_1 _3646_ (.A1(net540),
    .A2(_0852_),
    .Y(_0127_),
    .B1(_0776_));
 sg13g2_a21oi_1 _3647_ (.A1(_0780_),
    .A2(_0844_),
    .Y(_0853_),
    .B1(_0842_));
 sg13g2_o21ai_1 _3648_ (.B1(_0799_),
    .Y(_0854_),
    .A1(_0576_),
    .A2(_0800_));
 sg13g2_a21oi_2 _3649_ (.B1(_0837_),
    .Y(_0855_),
    .A2(_0839_),
    .A1(_0801_));
 sg13g2_o21ai_1 _3650_ (.B1(_0797_),
    .Y(_0856_),
    .A1(_0783_),
    .A2(_0793_));
 sg13g2_o21ai_1 _3651_ (.B1(_0811_),
    .Y(_0857_),
    .A1(_0803_),
    .A2(_0812_));
 sg13g2_a21oi_1 _3652_ (.A1(_0570_),
    .A2(_0790_),
    .Y(_0858_),
    .B1(_0792_));
 sg13g2_nor2_1 _3653_ (.A(net493),
    .B(net474),
    .Y(_0859_));
 sg13g2_nand2_1 _3654_ (.Y(_0860_),
    .A(_0468_),
    .B(_0859_));
 sg13g2_xnor2_1 _3655_ (.Y(_0861_),
    .A(_0789_),
    .B(_0859_));
 sg13g2_nor3_1 _3656_ (.A(net490),
    .B(net474),
    .C(_0861_),
    .Y(_0862_));
 sg13g2_xnor2_1 _3657_ (.Y(_0863_),
    .A(_0788_),
    .B(_0861_));
 sg13g2_nand2b_1 _3658_ (.Y(_0864_),
    .B(_0863_),
    .A_N(_0858_));
 sg13g2_xnor2_1 _3659_ (.Y(_0865_),
    .A(_0858_),
    .B(_0863_));
 sg13g2_xnor2_1 _3660_ (.Y(_0866_),
    .A(_0857_),
    .B(_0865_));
 sg13g2_nor2b_1 _3661_ (.A(_0866_),
    .B_N(_0856_),
    .Y(_0867_));
 sg13g2_xnor2_1 _3662_ (.Y(_0868_),
    .A(_0856_),
    .B(_0866_));
 sg13g2_a21oi_2 _3663_ (.B1(_0832_),
    .Y(_0869_),
    .A2(_0834_),
    .A1(_0814_));
 sg13g2_a22oi_1 _3664_ (.Y(_0870_),
    .B1(_0809_),
    .B2(_0805_),
    .A2(_0806_),
    .A1(_0585_));
 sg13g2_a22oi_1 _3665_ (.Y(_0871_),
    .B1(_0817_),
    .B2(_0529_),
    .A2(_0815_),
    .A1(_0595_));
 sg13g2_nor2_1 _3666_ (.A(net505),
    .B(net491),
    .Y(_0872_));
 sg13g2_nor2_1 _3667_ (.A(net499),
    .B(net531),
    .Y(_0873_));
 sg13g2_nor2_1 _3668_ (.A(net500),
    .B(net531),
    .Y(_0874_));
 sg13g2_xor2_1 _3669_ (.B(_0874_),
    .A(_0806_),
    .X(_0875_));
 sg13g2_xnor2_1 _3670_ (.Y(_0876_),
    .A(_0872_),
    .B(_0875_));
 sg13g2_or2_1 _3671_ (.X(_0877_),
    .B(_0876_),
    .A(_0871_));
 sg13g2_and2_1 _3672_ (.A(_0871_),
    .B(_0876_),
    .X(_0878_));
 sg13g2_xor2_1 _3673_ (.B(_0876_),
    .A(_0871_),
    .X(_0879_));
 sg13g2_xnor2_1 _3674_ (.Y(_0880_),
    .A(_0870_),
    .B(_0879_));
 sg13g2_xor2_1 _3675_ (.B(_0879_),
    .A(_0870_),
    .X(_0881_));
 sg13g2_o21ai_1 _3676_ (.B1(_0827_),
    .Y(_0882_),
    .A1(_0820_),
    .A2(_0828_));
 sg13g2_nor2_1 _3677_ (.A(net488),
    .B(net487),
    .Y(_0883_));
 sg13g2_nor2_1 _3678_ (.A(net503),
    .B(net477),
    .Y(_0884_));
 sg13g2_nor2_1 _3679_ (.A(net503),
    .B(net483),
    .Y(_0885_));
 sg13g2_xor2_1 _3680_ (.B(_0885_),
    .A(_0815_),
    .X(_0886_));
 sg13g2_xor2_1 _3681_ (.B(_0886_),
    .A(_0883_),
    .X(_0887_));
 sg13g2_o21ai_1 _3682_ (.B1(_0823_),
    .Y(_0888_),
    .A1(_0821_),
    .A2(_0824_));
 sg13g2_or2_1 _3683_ (.X(_0889_),
    .B(net476),
    .A(net533));
 sg13g2_nor4_1 _3684_ (.A(_0460_),
    .B(net527),
    .C(net481),
    .D(net469),
    .Y(_0890_));
 sg13g2_nand4_1 _3685_ (.B(_0487_),
    .C(net479),
    .A(net496),
    .Y(_0891_),
    .D(net468));
 sg13g2_a22oi_1 _3686_ (.Y(_0892_),
    .B1(net468),
    .B2(net496),
    .A2(_0524_),
    .A1(_0487_));
 sg13g2_or3_1 _3687_ (.A(_0889_),
    .B(_0890_),
    .C(_0892_),
    .X(_0893_));
 sg13g2_o21ai_1 _3688_ (.B1(_0889_),
    .Y(_0894_),
    .A1(_0890_),
    .A2(_0892_));
 sg13g2_and3_1 _3689_ (.X(_0895_),
    .A(_0888_),
    .B(_0893_),
    .C(_0894_));
 sg13g2_nand3_1 _3690_ (.B(_0893_),
    .C(_0894_),
    .A(_0888_),
    .Y(_0896_));
 sg13g2_a21o_1 _3691_ (.A2(_0894_),
    .A1(_0893_),
    .B1(_0888_),
    .X(_0897_));
 sg13g2_nand3_1 _3692_ (.B(_0896_),
    .C(_0897_),
    .A(_0887_),
    .Y(_0898_));
 sg13g2_a21o_1 _3693_ (.A2(_0897_),
    .A1(_0896_),
    .B1(_0887_),
    .X(_0899_));
 sg13g2_nand3_1 _3694_ (.B(_0898_),
    .C(_0899_),
    .A(_0882_),
    .Y(_0900_));
 sg13g2_a21oi_1 _3695_ (.A1(_0898_),
    .A2(_0899_),
    .Y(_0901_),
    .B1(_0882_));
 sg13g2_a21o_1 _3696_ (.A2(_0899_),
    .A1(_0898_),
    .B1(_0882_),
    .X(_0902_));
 sg13g2_and3_1 _3697_ (.X(_0903_),
    .A(_0880_),
    .B(_0900_),
    .C(_0902_));
 sg13g2_a21oi_2 _3698_ (.B1(_0880_),
    .Y(_0904_),
    .A2(_0902_),
    .A1(_0900_));
 sg13g2_nor3_1 _3699_ (.A(_0869_),
    .B(_0903_),
    .C(_0904_),
    .Y(_0905_));
 sg13g2_or3_1 _3700_ (.A(_0869_),
    .B(_0903_),
    .C(_0904_),
    .X(_0906_));
 sg13g2_o21ai_1 _3701_ (.B1(_0869_),
    .Y(_0907_),
    .A1(_0903_),
    .A2(_0904_));
 sg13g2_and3_1 _3702_ (.X(_0908_),
    .A(_0868_),
    .B(_0906_),
    .C(_0907_));
 sg13g2_a21oi_1 _3703_ (.A1(_0906_),
    .A2(_0907_),
    .Y(_0909_),
    .B1(_0868_));
 sg13g2_nor3_1 _3704_ (.A(_0855_),
    .B(_0908_),
    .C(_0909_),
    .Y(_0910_));
 sg13g2_or3_1 _3705_ (.A(_0855_),
    .B(_0908_),
    .C(_0909_),
    .X(_0911_));
 sg13g2_o21ai_1 _3706_ (.B1(_0855_),
    .Y(_0912_),
    .A1(_0908_),
    .A2(_0909_));
 sg13g2_and3_1 _3707_ (.X(_0913_),
    .A(_0854_),
    .B(_0911_),
    .C(_0912_));
 sg13g2_nand3_1 _3708_ (.B(_0911_),
    .C(_0912_),
    .A(_0854_),
    .Y(_0914_));
 sg13g2_a21oi_1 _3709_ (.A1(_0911_),
    .A2(_0912_),
    .Y(_0915_),
    .B1(_0854_));
 sg13g2_a21o_1 _3710_ (.A2(_0912_),
    .A1(_0911_),
    .B1(_0854_),
    .X(_0916_));
 sg13g2_nor3_2 _3711_ (.A(_0853_),
    .B(_0913_),
    .C(_0915_),
    .Y(_0917_));
 sg13g2_a221oi_1 _3712_ (.B2(_0916_),
    .C1(_0842_),
    .B1(_0914_),
    .A1(_0780_),
    .Y(_0918_),
    .A2(_0844_));
 sg13g2_or2_1 _3713_ (.X(_0919_),
    .B(_0918_),
    .A(_0917_));
 sg13g2_inv_1 _3714_ (.Y(_0920_),
    .A(_0919_));
 sg13g2_a221oi_1 _3715_ (.B2(_0850_),
    .C1(_0657_),
    .B1(_0849_),
    .A1(_0769_),
    .Y(_0921_),
    .A2(_0771_));
 sg13g2_a21oi_1 _3716_ (.A1(_0655_),
    .A2(_0848_),
    .Y(_0922_),
    .B1(_0847_));
 sg13g2_or2_1 _3717_ (.X(_0923_),
    .B(_0922_),
    .A(_0921_));
 sg13g2_xnor2_1 _3718_ (.Y(_0924_),
    .A(_0920_),
    .B(_0923_));
 sg13g2_nor2_1 _3719_ (.A(net799),
    .B(net540),
    .Y(_0925_));
 sg13g2_a21oi_1 _3720_ (.A1(net540),
    .A2(_0924_),
    .Y(_0128_),
    .B1(_0925_));
 sg13g2_nor2_1 _3721_ (.A(net741),
    .B(net540),
    .Y(_0926_));
 sg13g2_a21oi_1 _3722_ (.A1(_0854_),
    .A2(_0912_),
    .Y(_0927_),
    .B1(_0910_));
 sg13g2_a21o_1 _3723_ (.A2(_0865_),
    .A1(_0857_),
    .B1(_0867_),
    .X(_0928_));
 sg13g2_inv_1 _3724_ (.Y(_0929_),
    .A(_0928_));
 sg13g2_a21o_1 _3725_ (.A2(_0907_),
    .A1(_0868_),
    .B1(_0905_),
    .X(_0930_));
 sg13g2_o21ai_1 _3726_ (.B1(_0877_),
    .Y(_0931_),
    .A1(_0870_),
    .A2(_0878_));
 sg13g2_nor2_1 _3727_ (.A(net490),
    .B(_0860_),
    .Y(_0932_));
 sg13g2_a21oi_2 _3728_ (.B1(net474),
    .Y(_0933_),
    .A2(net492),
    .A1(net495));
 sg13g2_nand2_1 _3729_ (.Y(_0934_),
    .A(_0860_),
    .B(_0933_));
 sg13g2_a21oi_1 _3730_ (.A1(_0789_),
    .A2(_0859_),
    .Y(_0935_),
    .B1(_0862_));
 sg13g2_xor2_1 _3731_ (.B(_0934_),
    .A(_0788_),
    .X(_0936_));
 sg13g2_a21oi_1 _3732_ (.A1(_0935_),
    .A2(_0936_),
    .Y(_0937_),
    .B1(_0932_));
 sg13g2_nand2_1 _3733_ (.Y(_0938_),
    .A(_0931_),
    .B(_0937_));
 sg13g2_xnor2_1 _3734_ (.Y(_0939_),
    .A(_0931_),
    .B(_0937_));
 sg13g2_xnor2_1 _3735_ (.Y(_0940_),
    .A(_0864_),
    .B(_0939_));
 sg13g2_o21ai_1 _3736_ (.B1(_0900_),
    .Y(_0941_),
    .A1(_0881_),
    .A2(_0901_));
 sg13g2_a22oi_1 _3737_ (.Y(_0942_),
    .B1(_0875_),
    .B2(_0872_),
    .A2(_0873_),
    .A1(_0807_));
 sg13g2_a22oi_1 _3738_ (.Y(_0943_),
    .B1(_0886_),
    .B2(_0883_),
    .A2(_0884_),
    .A1(_0816_));
 sg13g2_nor2_1 _3739_ (.A(net504),
    .B(net527),
    .Y(_0944_));
 sg13g2_nor2_1 _3740_ (.A(net499),
    .B(_0480_),
    .Y(_0945_));
 sg13g2_nor2_1 _3741_ (.A(net500),
    .B(_0480_),
    .Y(_0946_));
 sg13g2_xor2_1 _3742_ (.B(_0946_),
    .A(_0873_),
    .X(_0947_));
 sg13g2_xnor2_1 _3743_ (.Y(_0948_),
    .A(_0944_),
    .B(_0947_));
 sg13g2_xor2_1 _3744_ (.B(_0948_),
    .A(_0943_),
    .X(_0949_));
 sg13g2_nand2b_1 _3745_ (.Y(_0950_),
    .B(_0949_),
    .A_N(_0942_));
 sg13g2_xor2_1 _3746_ (.B(_0949_),
    .A(_0942_),
    .X(_0951_));
 sg13g2_a21o_1 _3747_ (.A2(_0897_),
    .A1(_0887_),
    .B1(_0895_),
    .X(_0952_));
 sg13g2_nor2_1 _3748_ (.A(net529),
    .B(net487),
    .Y(_0953_));
 sg13g2_nor2_1 _3749_ (.A(net488),
    .B(net477),
    .Y(_0954_));
 sg13g2_nor2_1 _3750_ (.A(net488),
    .B(net483),
    .Y(_0955_));
 sg13g2_xor2_1 _3751_ (.B(_0955_),
    .A(_0884_),
    .X(_0956_));
 sg13g2_xnor2_1 _3752_ (.Y(_0957_),
    .A(_0953_),
    .B(_0956_));
 sg13g2_o21ai_1 _3753_ (.B1(_0891_),
    .Y(_0958_),
    .A1(_0889_),
    .A2(_0892_));
 sg13g2_or2_1 _3754_ (.X(_0959_),
    .B(net476),
    .A(net498));
 sg13g2_nor4_1 _3755_ (.A(_0442_),
    .B(net482),
    .C(net525),
    .D(net470),
    .Y(_0960_));
 sg13g2_nand4_1 _3756_ (.B(net479),
    .C(_0568_),
    .A(net533),
    .Y(_0961_),
    .D(net467));
 sg13g2_a22oi_1 _3757_ (.Y(_0962_),
    .B1(net467),
    .B2(net533),
    .A2(_0568_),
    .A1(net479));
 sg13g2_or3_1 _3758_ (.A(_0959_),
    .B(_0960_),
    .C(_0962_),
    .X(_0963_));
 sg13g2_o21ai_1 _3759_ (.B1(_0959_),
    .Y(_0964_),
    .A1(_0960_),
    .A2(_0962_));
 sg13g2_and3_1 _3760_ (.X(_0965_),
    .A(_0958_),
    .B(_0963_),
    .C(_0964_));
 sg13g2_nand3_1 _3761_ (.B(_0963_),
    .C(_0964_),
    .A(_0958_),
    .Y(_0966_));
 sg13g2_a21oi_2 _3762_ (.B1(_0958_),
    .Y(_0967_),
    .A2(_0964_),
    .A1(_0963_));
 sg13g2_or3_1 _3763_ (.A(_0957_),
    .B(_0965_),
    .C(_0967_),
    .X(_0968_));
 sg13g2_o21ai_1 _3764_ (.B1(_0957_),
    .Y(_0969_),
    .A1(_0965_),
    .A2(_0967_));
 sg13g2_and3_1 _3765_ (.X(_0970_),
    .A(_0952_),
    .B(_0968_),
    .C(_0969_));
 sg13g2_nand3_1 _3766_ (.B(_0968_),
    .C(_0969_),
    .A(_0952_),
    .Y(_0971_));
 sg13g2_a21oi_1 _3767_ (.A1(_0968_),
    .A2(_0969_),
    .Y(_0972_),
    .B1(_0952_));
 sg13g2_or3_2 _3768_ (.A(_0951_),
    .B(_0970_),
    .C(_0972_),
    .X(_0973_));
 sg13g2_o21ai_1 _3769_ (.B1(_0951_),
    .Y(_0974_),
    .A1(_0970_),
    .A2(_0972_));
 sg13g2_and3_1 _3770_ (.X(_0975_),
    .A(_0941_),
    .B(_0973_),
    .C(_0974_));
 sg13g2_nand3_1 _3771_ (.B(_0973_),
    .C(_0974_),
    .A(_0941_),
    .Y(_0976_));
 sg13g2_a21oi_1 _3772_ (.A1(_0973_),
    .A2(_0974_),
    .Y(_0977_),
    .B1(_0941_));
 sg13g2_or3_1 _3773_ (.A(_0940_),
    .B(_0975_),
    .C(_0977_),
    .X(_0978_));
 sg13g2_o21ai_1 _3774_ (.B1(_0940_),
    .Y(_0979_),
    .A1(_0975_),
    .A2(_0977_));
 sg13g2_and3_1 _3775_ (.X(_0980_),
    .A(_0930_),
    .B(_0978_),
    .C(_0979_));
 sg13g2_nand3_1 _3776_ (.B(_0978_),
    .C(_0979_),
    .A(_0930_),
    .Y(_0981_));
 sg13g2_a21oi_1 _3777_ (.A1(_0978_),
    .A2(_0979_),
    .Y(_0982_),
    .B1(_0930_));
 sg13g2_a21o_1 _3778_ (.A2(_0979_),
    .A1(_0978_),
    .B1(_0930_),
    .X(_0983_));
 sg13g2_nor3_1 _3779_ (.A(_0929_),
    .B(_0980_),
    .C(_0982_),
    .Y(_0984_));
 sg13g2_a21oi_1 _3780_ (.A1(_0981_),
    .A2(_0983_),
    .Y(_0985_),
    .B1(_0928_));
 sg13g2_a21oi_1 _3781_ (.A1(_0981_),
    .A2(_0983_),
    .Y(_0986_),
    .B1(_0929_));
 sg13g2_nor3_1 _3782_ (.A(_0928_),
    .B(_0980_),
    .C(_0982_),
    .Y(_0987_));
 sg13g2_nor4_1 _3783_ (.A(_0910_),
    .B(_0913_),
    .C(_0986_),
    .D(_0987_),
    .Y(_0988_));
 sg13g2_o21ai_1 _3784_ (.B1(_0927_),
    .Y(_0989_),
    .A1(_0984_),
    .A2(_0985_));
 sg13g2_nor3_1 _3785_ (.A(_0927_),
    .B(_0984_),
    .C(_0985_),
    .Y(_0990_));
 sg13g2_or2_1 _3786_ (.X(_0991_),
    .B(_0990_),
    .A(_0988_));
 sg13g2_a21oi_1 _3787_ (.A1(_0920_),
    .A2(_0923_),
    .Y(_0992_),
    .B1(_0917_));
 sg13g2_xnor2_1 _3788_ (.Y(_0993_),
    .A(_0991_),
    .B(_0992_));
 sg13g2_a21oi_1 _3789_ (.A1(net540),
    .A2(_0993_),
    .Y(_0129_),
    .B1(_0926_));
 sg13g2_o21ai_1 _3790_ (.B1(_0981_),
    .Y(_0994_),
    .A1(_0929_),
    .A2(_0982_));
 sg13g2_o21ai_1 _3791_ (.B1(_0938_),
    .Y(_0995_),
    .A1(_0864_),
    .A2(_0939_));
 sg13g2_inv_1 _3792_ (.Y(_0996_),
    .A(_0995_));
 sg13g2_o21ai_1 _3793_ (.B1(_0976_),
    .Y(_0997_),
    .A1(_0940_),
    .A2(_0977_));
 sg13g2_o21ai_1 _3794_ (.B1(_0950_),
    .Y(_0998_),
    .A1(_0943_),
    .A2(_0948_));
 sg13g2_nor2_2 _3795_ (.A(_0788_),
    .B(_0933_),
    .Y(_0999_));
 sg13g2_or2_1 _3796_ (.X(_1000_),
    .B(_0933_),
    .A(_0788_));
 sg13g2_nand2_1 _3797_ (.Y(_1001_),
    .A(_0998_),
    .B(net453));
 sg13g2_xnor2_1 _3798_ (.Y(_1002_),
    .A(_0998_),
    .B(net453));
 sg13g2_o21ai_1 _3799_ (.B1(_0971_),
    .Y(_1003_),
    .A1(_0951_),
    .A2(_0972_));
 sg13g2_a22oi_1 _3800_ (.Y(_1004_),
    .B1(_0947_),
    .B2(_0944_),
    .A2(_0945_),
    .A1(_0874_));
 sg13g2_a22oi_1 _3801_ (.Y(_1005_),
    .B1(_0956_),
    .B2(_0953_),
    .A2(_0954_),
    .A1(_0885_));
 sg13g2_nor2_1 _3802_ (.A(net504),
    .B(net525),
    .Y(_1006_));
 sg13g2_nor2_1 _3803_ (.A(net499),
    .B(net528),
    .Y(_1007_));
 sg13g2_nor2_1 _3804_ (.A(net500),
    .B(net528),
    .Y(_1008_));
 sg13g2_xor2_1 _3805_ (.B(_1008_),
    .A(_0945_),
    .X(_1009_));
 sg13g2_xnor2_1 _3806_ (.Y(_1010_),
    .A(_1006_),
    .B(_1009_));
 sg13g2_xor2_1 _3807_ (.B(_1010_),
    .A(_1005_),
    .X(_1011_));
 sg13g2_nand2b_1 _3808_ (.Y(_1012_),
    .B(_1011_),
    .A_N(_1004_));
 sg13g2_xnor2_1 _3809_ (.Y(_1013_),
    .A(_1004_),
    .B(_1011_));
 sg13g2_o21ai_1 _3810_ (.B1(_0966_),
    .Y(_1014_),
    .A1(_0957_),
    .A2(_0967_));
 sg13g2_nor2_1 _3811_ (.A(net532),
    .B(net486),
    .Y(_1015_));
 sg13g2_nor2_1 _3812_ (.A(net529),
    .B(net477),
    .Y(_1016_));
 sg13g2_nor2_1 _3813_ (.A(net529),
    .B(net483),
    .Y(_1017_));
 sg13g2_xor2_1 _3814_ (.B(_1017_),
    .A(_0954_),
    .X(_1018_));
 sg13g2_xnor2_1 _3815_ (.Y(_1019_),
    .A(_1015_),
    .B(_1018_));
 sg13g2_o21ai_1 _3816_ (.B1(_0961_),
    .Y(_1020_),
    .A1(_0959_),
    .A2(_0962_));
 sg13g2_or2_1 _3817_ (.X(_1021_),
    .B(net476),
    .A(net502));
 sg13g2_nor2_2 _3818_ (.A(net481),
    .B(net472),
    .Y(_1022_));
 sg13g2_nor4_1 _3819_ (.A(_0450_),
    .B(net481),
    .C(net473),
    .D(net470),
    .Y(_1023_));
 sg13g2_nand4_1 _3820_ (.B(net479),
    .C(_0787_),
    .A(net498),
    .Y(_1024_),
    .D(net467));
 sg13g2_a22oi_1 _3821_ (.Y(_1025_),
    .B1(net467),
    .B2(net498),
    .A2(_0787_),
    .A1(net478));
 sg13g2_or3_1 _3822_ (.A(_1021_),
    .B(_1023_),
    .C(_1025_),
    .X(_1026_));
 sg13g2_o21ai_1 _3823_ (.B1(_1021_),
    .Y(_1027_),
    .A1(_1023_),
    .A2(_1025_));
 sg13g2_and3_1 _3824_ (.X(_1028_),
    .A(_1020_),
    .B(_1026_),
    .C(_1027_));
 sg13g2_nand3_1 _3825_ (.B(_1026_),
    .C(_1027_),
    .A(_1020_),
    .Y(_1029_));
 sg13g2_a21oi_1 _3826_ (.A1(_1026_),
    .A2(_1027_),
    .Y(_1030_),
    .B1(_1020_));
 sg13g2_or3_2 _3827_ (.A(_1019_),
    .B(_1028_),
    .C(_1030_),
    .X(_1031_));
 sg13g2_o21ai_1 _3828_ (.B1(_1019_),
    .Y(_1032_),
    .A1(_1028_),
    .A2(_1030_));
 sg13g2_and3_1 _3829_ (.X(_1033_),
    .A(_1014_),
    .B(_1031_),
    .C(_1032_));
 sg13g2_nand3_1 _3830_ (.B(_1031_),
    .C(_1032_),
    .A(_1014_),
    .Y(_1034_));
 sg13g2_a21o_1 _3831_ (.A2(_1032_),
    .A1(_1031_),
    .B1(_1014_),
    .X(_1035_));
 sg13g2_nand3_1 _3832_ (.B(_1034_),
    .C(_1035_),
    .A(_1013_),
    .Y(_1036_));
 sg13g2_a21o_1 _3833_ (.A2(_1035_),
    .A1(_1034_),
    .B1(_1013_),
    .X(_1037_));
 sg13g2_and3_1 _3834_ (.X(_1038_),
    .A(_1003_),
    .B(_1036_),
    .C(_1037_));
 sg13g2_nand3_1 _3835_ (.B(_1036_),
    .C(_1037_),
    .A(_1003_),
    .Y(_1039_));
 sg13g2_a21oi_1 _3836_ (.A1(_1036_),
    .A2(_1037_),
    .Y(_1040_),
    .B1(_1003_));
 sg13g2_or3_1 _3837_ (.A(_1002_),
    .B(_1038_),
    .C(_1040_),
    .X(_1041_));
 sg13g2_o21ai_1 _3838_ (.B1(_1002_),
    .Y(_1042_),
    .A1(_1038_),
    .A2(_1040_));
 sg13g2_nand3_1 _3839_ (.B(_1041_),
    .C(_1042_),
    .A(_0997_),
    .Y(_1043_));
 sg13g2_a21oi_1 _3840_ (.A1(_1041_),
    .A2(_1042_),
    .Y(_1044_),
    .B1(_0997_));
 sg13g2_a21o_1 _3841_ (.A2(_1042_),
    .A1(_1041_),
    .B1(_0997_),
    .X(_1045_));
 sg13g2_nand3_1 _3842_ (.B(_1043_),
    .C(_1045_),
    .A(_0995_),
    .Y(_1046_));
 sg13g2_a21o_1 _3843_ (.A2(_1045_),
    .A1(_1043_),
    .B1(_0995_),
    .X(_1047_));
 sg13g2_nand3_1 _3844_ (.B(_1046_),
    .C(_1047_),
    .A(_0994_),
    .Y(_1048_));
 sg13g2_a21o_1 _3845_ (.A2(_1047_),
    .A1(_1046_),
    .B1(_0994_),
    .X(_1049_));
 sg13g2_and2_1 _3846_ (.A(_1048_),
    .B(_1049_),
    .X(_1050_));
 sg13g2_nor4_1 _3847_ (.A(_0917_),
    .B(_0918_),
    .C(_0988_),
    .D(_0990_),
    .Y(_1051_));
 sg13g2_and2_1 _3848_ (.A(_0923_),
    .B(_1051_),
    .X(_1052_));
 sg13g2_o21ai_1 _3849_ (.B1(_1051_),
    .Y(_1053_),
    .A1(_0921_),
    .A2(_0922_));
 sg13g2_a21o_1 _3850_ (.A2(_0989_),
    .A1(_0917_),
    .B1(_0990_),
    .X(_1054_));
 sg13g2_nor2_1 _3851_ (.A(_1052_),
    .B(_1054_),
    .Y(_1055_));
 sg13g2_o21ai_1 _3852_ (.B1(_1050_),
    .Y(_1056_),
    .A1(_1052_),
    .A2(_1054_));
 sg13g2_xor2_1 _3853_ (.B(_1055_),
    .A(_1050_),
    .X(_1057_));
 sg13g2_nor2_1 _3854_ (.A(net807),
    .B(net541),
    .Y(_1058_));
 sg13g2_a21oi_1 _3855_ (.A1(net541),
    .A2(_1057_),
    .Y(_0130_),
    .B1(_1058_));
 sg13g2_nor2_1 _3856_ (.A(net788),
    .B(net541),
    .Y(_1059_));
 sg13g2_o21ai_1 _3857_ (.B1(_1043_),
    .Y(_1060_),
    .A1(_0996_),
    .A2(_1044_));
 sg13g2_o21ai_1 _3858_ (.B1(_1039_),
    .Y(_1061_),
    .A1(_1002_),
    .A2(_1040_));
 sg13g2_o21ai_1 _3859_ (.B1(_1012_),
    .Y(_1062_),
    .A1(_1005_),
    .A2(_1010_));
 sg13g2_nand2_1 _3860_ (.Y(_1063_),
    .A(net453),
    .B(_1062_));
 sg13g2_xnor2_1 _3861_ (.Y(_1064_),
    .A(net452),
    .B(_1062_));
 sg13g2_a21o_1 _3862_ (.A2(_1035_),
    .A1(_1013_),
    .B1(_1033_),
    .X(_1065_));
 sg13g2_a22oi_1 _3863_ (.Y(_1066_),
    .B1(_1009_),
    .B2(_1006_),
    .A2(_1007_),
    .A1(_0946_));
 sg13g2_a22oi_1 _3864_ (.Y(_1067_),
    .B1(_1018_),
    .B2(_1015_),
    .A2(_1016_),
    .A1(_0955_));
 sg13g2_nor2_2 _3865_ (.A(net504),
    .B(net472),
    .Y(_1068_));
 sg13g2_nor2_1 _3866_ (.A(net499),
    .B(net525),
    .Y(_1069_));
 sg13g2_nor2_1 _3867_ (.A(net500),
    .B(net526),
    .Y(_1070_));
 sg13g2_xor2_1 _3868_ (.B(_1070_),
    .A(_1007_),
    .X(_1071_));
 sg13g2_xnor2_1 _3869_ (.Y(_1072_),
    .A(_1068_),
    .B(_1071_));
 sg13g2_xor2_1 _3870_ (.B(_1072_),
    .A(_1067_),
    .X(_1073_));
 sg13g2_nand2b_1 _3871_ (.Y(_1074_),
    .B(_1073_),
    .A_N(_1066_));
 sg13g2_xor2_1 _3872_ (.B(_1073_),
    .A(_1066_),
    .X(_1075_));
 sg13g2_o21ai_1 _3873_ (.B1(_1029_),
    .Y(_1076_),
    .A1(_1019_),
    .A2(_1030_));
 sg13g2_nor2_1 _3874_ (.A(net491),
    .B(net486),
    .Y(_1077_));
 sg13g2_nor2_1 _3875_ (.A(net531),
    .B(net477),
    .Y(_1078_));
 sg13g2_nor2_1 _3876_ (.A(net531),
    .B(net483),
    .Y(_1079_));
 sg13g2_xor2_1 _3877_ (.B(_1079_),
    .A(_1016_),
    .X(_1080_));
 sg13g2_xnor2_1 _3878_ (.Y(_1081_),
    .A(_1077_),
    .B(_1080_));
 sg13g2_o21ai_1 _3879_ (.B1(_1024_),
    .Y(_1082_),
    .A1(_1021_),
    .A2(_1025_));
 sg13g2_or2_1 _3880_ (.X(_1083_),
    .B(net475),
    .A(net488));
 sg13g2_nor4_1 _3881_ (.A(_0439_),
    .B(net481),
    .C(net473),
    .D(net469),
    .Y(_1084_));
 sg13g2_nand4_1 _3882_ (.B(net478),
    .C(_0787_),
    .A(net502),
    .Y(_1085_),
    .D(net468));
 sg13g2_a22oi_1 _3883_ (.Y(_1086_),
    .B1(net468),
    .B2(net502),
    .A2(_0787_),
    .A1(net478));
 sg13g2_or3_1 _3884_ (.A(_1083_),
    .B(_1084_),
    .C(_1086_),
    .X(_1087_));
 sg13g2_o21ai_1 _3885_ (.B1(_1083_),
    .Y(_1088_),
    .A1(_1084_),
    .A2(_1086_));
 sg13g2_and3_1 _3886_ (.X(_1089_),
    .A(_1082_),
    .B(_1087_),
    .C(_1088_));
 sg13g2_nand3_1 _3887_ (.B(_1087_),
    .C(_1088_),
    .A(_1082_),
    .Y(_1090_));
 sg13g2_a21oi_1 _3888_ (.A1(_1087_),
    .A2(_1088_),
    .Y(_1091_),
    .B1(_1082_));
 sg13g2_or3_1 _3889_ (.A(_1081_),
    .B(_1089_),
    .C(_1091_),
    .X(_1092_));
 sg13g2_o21ai_1 _3890_ (.B1(_1081_),
    .Y(_1093_),
    .A1(_1089_),
    .A2(_1091_));
 sg13g2_and3_1 _3891_ (.X(_1094_),
    .A(_1076_),
    .B(_1092_),
    .C(_1093_));
 sg13g2_nand3_1 _3892_ (.B(_1092_),
    .C(_1093_),
    .A(_1076_),
    .Y(_1095_));
 sg13g2_a21oi_1 _3893_ (.A1(_1092_),
    .A2(_1093_),
    .Y(_1096_),
    .B1(_1076_));
 sg13g2_or3_1 _3894_ (.A(_1075_),
    .B(_1094_),
    .C(_1096_),
    .X(_1097_));
 sg13g2_o21ai_1 _3895_ (.B1(_1075_),
    .Y(_1098_),
    .A1(_1094_),
    .A2(_1096_));
 sg13g2_and3_1 _3896_ (.X(_1099_),
    .A(_1065_),
    .B(_1097_),
    .C(_1098_));
 sg13g2_nand3_1 _3897_ (.B(_1097_),
    .C(_1098_),
    .A(_1065_),
    .Y(_1100_));
 sg13g2_a21oi_1 _3898_ (.A1(_1097_),
    .A2(_1098_),
    .Y(_1101_),
    .B1(_1065_));
 sg13g2_or3_1 _3899_ (.A(_1064_),
    .B(_1099_),
    .C(_1101_),
    .X(_1102_));
 sg13g2_o21ai_1 _3900_ (.B1(_1064_),
    .Y(_1103_),
    .A1(_1099_),
    .A2(_1101_));
 sg13g2_and3_1 _3901_ (.X(_1104_),
    .A(_1061_),
    .B(_1102_),
    .C(_1103_));
 sg13g2_nand3_1 _3902_ (.B(_1102_),
    .C(_1103_),
    .A(_1061_),
    .Y(_1105_));
 sg13g2_a21oi_1 _3903_ (.A1(_1102_),
    .A2(_1103_),
    .Y(_1106_),
    .B1(_1061_));
 sg13g2_or3_1 _3904_ (.A(_1001_),
    .B(_1104_),
    .C(_1106_),
    .X(_1107_));
 sg13g2_o21ai_1 _3905_ (.B1(_1001_),
    .Y(_1108_),
    .A1(_1104_),
    .A2(_1106_));
 sg13g2_a21oi_1 _3906_ (.A1(_1107_),
    .A2(_1108_),
    .Y(_1109_),
    .B1(_1060_));
 sg13g2_nand3_1 _3907_ (.B(_1107_),
    .C(_1108_),
    .A(_1060_),
    .Y(_1110_));
 sg13g2_nor2b_1 _3908_ (.A(_1109_),
    .B_N(_1110_),
    .Y(_1111_));
 sg13g2_nand2_1 _3909_ (.Y(_1112_),
    .A(_1048_),
    .B(_1056_));
 sg13g2_xnor2_1 _3910_ (.Y(_1113_),
    .A(_1111_),
    .B(_1112_));
 sg13g2_a21oi_1 _3911_ (.A1(net541),
    .A2(_1113_),
    .Y(_0131_),
    .B1(_1059_));
 sg13g2_o21ai_1 _3912_ (.B1(_1100_),
    .Y(_1114_),
    .A1(_1064_),
    .A2(_1101_));
 sg13g2_o21ai_1 _3913_ (.B1(_1074_),
    .Y(_1115_),
    .A1(_1067_),
    .A2(_1072_));
 sg13g2_nand2_1 _3914_ (.Y(_1116_),
    .A(net452),
    .B(_1115_));
 sg13g2_inv_1 _3915_ (.Y(_1117_),
    .A(_1116_));
 sg13g2_xnor2_1 _3916_ (.Y(_1118_),
    .A(net453),
    .B(_1115_));
 sg13g2_o21ai_1 _3917_ (.B1(_1095_),
    .Y(_1119_),
    .A1(_1075_),
    .A2(_1096_));
 sg13g2_a22oi_1 _3918_ (.Y(_1120_),
    .B1(_1071_),
    .B2(_1068_),
    .A2(_1069_),
    .A1(_1008_));
 sg13g2_a22oi_1 _3919_ (.Y(_1121_),
    .B1(_1080_),
    .B2(_1077_),
    .A2(_1078_),
    .A1(_1017_));
 sg13g2_nor2_1 _3920_ (.A(net500),
    .B(net472),
    .Y(_1122_));
 sg13g2_nor2_1 _3921_ (.A(net499),
    .B(net472),
    .Y(_1123_));
 sg13g2_xor2_1 _3922_ (.B(_1122_),
    .A(_1069_),
    .X(_1124_));
 sg13g2_xnor2_1 _3923_ (.Y(_1125_),
    .A(_1068_),
    .B(_1124_));
 sg13g2_xor2_1 _3924_ (.B(_1125_),
    .A(_1121_),
    .X(_1126_));
 sg13g2_nand2b_1 _3925_ (.Y(_1127_),
    .B(_1126_),
    .A_N(_1120_));
 sg13g2_xnor2_1 _3926_ (.Y(_1128_),
    .A(_1120_),
    .B(_1126_));
 sg13g2_xor2_1 _3927_ (.B(_1126_),
    .A(_1120_),
    .X(_1129_));
 sg13g2_o21ai_1 _3928_ (.B1(_1090_),
    .Y(_1130_),
    .A1(_1081_),
    .A2(_1091_));
 sg13g2_nor2_1 _3929_ (.A(net527),
    .B(net486),
    .Y(_1131_));
 sg13g2_nor2_2 _3930_ (.A(net491),
    .B(net477),
    .Y(_1132_));
 sg13g2_nand2_1 _3931_ (.Y(_1133_),
    .A(_0481_),
    .B(_0517_));
 sg13g2_xnor2_1 _3932_ (.Y(_1134_),
    .A(_1078_),
    .B(_1133_));
 sg13g2_xnor2_1 _3933_ (.Y(_1135_),
    .A(_1131_),
    .B(_1134_));
 sg13g2_o21ai_1 _3934_ (.B1(_1085_),
    .Y(_1136_),
    .A1(_1083_),
    .A2(_1086_));
 sg13g2_or2_1 _3935_ (.X(_1137_),
    .B(net475),
    .A(net529));
 sg13g2_nor4_1 _3936_ (.A(_0499_),
    .B(net481),
    .C(net473),
    .D(net469),
    .Y(_1138_));
 sg13g2_nand4_1 _3937_ (.B(net478),
    .C(_0787_),
    .A(net488),
    .Y(_1139_),
    .D(net467));
 sg13g2_a22oi_1 _3938_ (.Y(_1140_),
    .B1(net467),
    .B2(net488),
    .A2(_0787_),
    .A1(net478));
 sg13g2_or3_1 _3939_ (.A(_1137_),
    .B(_1138_),
    .C(_1140_),
    .X(_1141_));
 sg13g2_o21ai_1 _3940_ (.B1(_1137_),
    .Y(_1142_),
    .A1(_1138_),
    .A2(_1140_));
 sg13g2_and3_1 _3941_ (.X(_1143_),
    .A(_1136_),
    .B(_1141_),
    .C(_1142_));
 sg13g2_nand3_1 _3942_ (.B(_1141_),
    .C(_1142_),
    .A(_1136_),
    .Y(_1144_));
 sg13g2_a21oi_1 _3943_ (.A1(_1141_),
    .A2(_1142_),
    .Y(_1145_),
    .B1(_1136_));
 sg13g2_or3_1 _3944_ (.A(_1135_),
    .B(_1143_),
    .C(_1145_),
    .X(_1146_));
 sg13g2_o21ai_1 _3945_ (.B1(_1135_),
    .Y(_1147_),
    .A1(_1143_),
    .A2(_1145_));
 sg13g2_nand3_1 _3946_ (.B(_1146_),
    .C(_1147_),
    .A(_1130_),
    .Y(_1148_));
 sg13g2_a21oi_1 _3947_ (.A1(_1146_),
    .A2(_1147_),
    .Y(_1149_),
    .B1(_1130_));
 sg13g2_a21o_1 _3948_ (.A2(_1147_),
    .A1(_1146_),
    .B1(_1130_),
    .X(_1150_));
 sg13g2_nand3_1 _3949_ (.B(_1148_),
    .C(_1150_),
    .A(_1128_),
    .Y(_1151_));
 sg13g2_a21o_1 _3950_ (.A2(_1150_),
    .A1(_1148_),
    .B1(_1128_),
    .X(_1152_));
 sg13g2_and3_1 _3951_ (.X(_1153_),
    .A(_1119_),
    .B(_1151_),
    .C(_1152_));
 sg13g2_nand3_1 _3952_ (.B(_1151_),
    .C(_1152_),
    .A(_1119_),
    .Y(_1154_));
 sg13g2_a21oi_1 _3953_ (.A1(_1151_),
    .A2(_1152_),
    .Y(_1155_),
    .B1(_1119_));
 sg13g2_or3_1 _3954_ (.A(_1118_),
    .B(_1153_),
    .C(_1155_),
    .X(_1156_));
 sg13g2_o21ai_1 _3955_ (.B1(_1118_),
    .Y(_1157_),
    .A1(_1153_),
    .A2(_1155_));
 sg13g2_and3_1 _3956_ (.X(_1158_),
    .A(_1114_),
    .B(_1156_),
    .C(_1157_));
 sg13g2_nand3_1 _3957_ (.B(_1156_),
    .C(_1157_),
    .A(_1114_),
    .Y(_1159_));
 sg13g2_a21oi_1 _3958_ (.A1(_1156_),
    .A2(_1157_),
    .Y(_1160_),
    .B1(_1114_));
 sg13g2_or3_1 _3959_ (.A(_1063_),
    .B(_1158_),
    .C(_1160_),
    .X(_1161_));
 sg13g2_o21ai_1 _3960_ (.B1(_1063_),
    .Y(_1162_),
    .A1(_1158_),
    .A2(_1160_));
 sg13g2_o21ai_1 _3961_ (.B1(_1105_),
    .Y(_1163_),
    .A1(_1001_),
    .A2(_1106_));
 sg13g2_a21oi_1 _3962_ (.A1(_1161_),
    .A2(_1162_),
    .Y(_1164_),
    .B1(_1163_));
 sg13g2_nand3_1 _3963_ (.B(_1162_),
    .C(_1163_),
    .A(_1161_),
    .Y(_1165_));
 sg13g2_nor2b_2 _3964_ (.A(_1164_),
    .B_N(_1165_),
    .Y(_1166_));
 sg13g2_nand2_1 _3965_ (.Y(_1167_),
    .A(_1050_),
    .B(_1111_));
 sg13g2_a21o_1 _3966_ (.A2(_1110_),
    .A1(_1048_),
    .B1(_1109_),
    .X(_1168_));
 sg13g2_nor2b_1 _3967_ (.A(_1054_),
    .B_N(_1168_),
    .Y(_1169_));
 sg13g2_a22oi_1 _3968_ (.Y(_1170_),
    .B1(_1169_),
    .B2(_1053_),
    .A2(_1168_),
    .A1(_1167_));
 sg13g2_nand2_1 _3969_ (.Y(_1171_),
    .A(_1166_),
    .B(_1170_));
 sg13g2_xnor2_1 _3970_ (.Y(_1172_),
    .A(_1166_),
    .B(_1170_));
 sg13g2_nor2_1 _3971_ (.A(net798),
    .B(net541),
    .Y(_1173_));
 sg13g2_a21oi_1 _3972_ (.A1(net539),
    .A2(_1172_),
    .Y(_0132_),
    .B1(_1173_));
 sg13g2_nor2_1 _3973_ (.A(net739),
    .B(net539),
    .Y(_1174_));
 sg13g2_o21ai_1 _3974_ (.B1(_1154_),
    .Y(_1175_),
    .A1(_1118_),
    .A2(_1155_));
 sg13g2_o21ai_1 _3975_ (.B1(_1127_),
    .Y(_1176_),
    .A1(_1121_),
    .A2(_1125_));
 sg13g2_nand2_1 _3976_ (.Y(_1177_),
    .A(net453),
    .B(_1176_));
 sg13g2_xnor2_1 _3977_ (.Y(_1178_),
    .A(net453),
    .B(_1176_));
 sg13g2_o21ai_1 _3978_ (.B1(_1148_),
    .Y(_1179_),
    .A1(_1129_),
    .A2(_1149_));
 sg13g2_a22oi_1 _3979_ (.Y(_1180_),
    .B1(_1124_),
    .B2(_1068_),
    .A2(_1123_),
    .A1(_1070_));
 sg13g2_a22oi_1 _3980_ (.Y(_1181_),
    .B1(_1134_),
    .B2(_1131_),
    .A2(_1132_),
    .A1(_1079_));
 sg13g2_mux2_1 _3981_ (.A0(_1122_),
    .A1(net500),
    .S(_1123_),
    .X(_1182_));
 sg13g2_xnor2_1 _3982_ (.Y(_1183_),
    .A(_1068_),
    .B(_1182_));
 sg13g2_nor2_1 _3983_ (.A(_1181_),
    .B(_1183_),
    .Y(_1184_));
 sg13g2_xor2_1 _3984_ (.B(net450),
    .A(_1181_),
    .X(_1185_));
 sg13g2_nor2b_1 _3985_ (.A(_1180_),
    .B_N(_1185_),
    .Y(_1186_));
 sg13g2_xnor2_1 _3986_ (.Y(_1187_),
    .A(_1180_),
    .B(_1185_));
 sg13g2_o21ai_1 _3987_ (.B1(_1144_),
    .Y(_1188_),
    .A1(_1135_),
    .A2(_1145_));
 sg13g2_nor2_1 _3988_ (.A(net486),
    .B(net525),
    .Y(_1189_));
 sg13g2_nor2_1 _3989_ (.A(net527),
    .B(net477),
    .Y(_1190_));
 sg13g2_nor2_1 _3990_ (.A(net527),
    .B(net483),
    .Y(_1191_));
 sg13g2_xnor2_1 _3991_ (.Y(_1192_),
    .A(_1132_),
    .B(_1191_));
 sg13g2_nor3_1 _3992_ (.A(net486),
    .B(net525),
    .C(_1192_),
    .Y(_1193_));
 sg13g2_xor2_1 _3993_ (.B(_1192_),
    .A(_1189_),
    .X(_1194_));
 sg13g2_o21ai_1 _3994_ (.B1(_1139_),
    .Y(_1195_),
    .A1(_1137_),
    .A2(_1140_));
 sg13g2_nor4_2 _3995_ (.A(_0472_),
    .B(net481),
    .C(net473),
    .Y(_1196_),
    .D(net469));
 sg13g2_a22oi_1 _3996_ (.Y(_1197_),
    .B1(net467),
    .B2(net529),
    .A2(_0787_),
    .A1(net478));
 sg13g2_or3_1 _3997_ (.A(_0601_),
    .B(_1196_),
    .C(_1197_),
    .X(_1198_));
 sg13g2_o21ai_1 _3998_ (.B1(_0601_),
    .Y(_1199_),
    .A1(_1196_),
    .A2(_1197_));
 sg13g2_and3_1 _3999_ (.X(_1200_),
    .A(_1195_),
    .B(_1198_),
    .C(_1199_));
 sg13g2_a21oi_1 _4000_ (.A1(_1198_),
    .A2(_1199_),
    .Y(_1201_),
    .B1(_1195_));
 sg13g2_or3_1 _4001_ (.A(_1194_),
    .B(_1200_),
    .C(_1201_),
    .X(_1202_));
 sg13g2_o21ai_1 _4002_ (.B1(_1194_),
    .Y(_1203_),
    .A1(_1200_),
    .A2(_1201_));
 sg13g2_nand3_1 _4003_ (.B(_1202_),
    .C(_1203_),
    .A(_1188_),
    .Y(_1204_));
 sg13g2_a21o_1 _4004_ (.A2(_1203_),
    .A1(_1202_),
    .B1(_1188_),
    .X(_1205_));
 sg13g2_nand3_1 _4005_ (.B(_1204_),
    .C(_1205_),
    .A(_1187_),
    .Y(_1206_));
 sg13g2_a21o_1 _4006_ (.A2(_1205_),
    .A1(_1204_),
    .B1(_1187_),
    .X(_1207_));
 sg13g2_and3_1 _4007_ (.X(_1208_),
    .A(_1179_),
    .B(_1206_),
    .C(_1207_));
 sg13g2_a21oi_1 _4008_ (.A1(_1206_),
    .A2(_1207_),
    .Y(_1209_),
    .B1(_1179_));
 sg13g2_or3_1 _4009_ (.A(_1178_),
    .B(_1208_),
    .C(_1209_),
    .X(_1210_));
 sg13g2_o21ai_1 _4010_ (.B1(_1178_),
    .Y(_1211_),
    .A1(_1208_),
    .A2(_1209_));
 sg13g2_nand3_1 _4011_ (.B(_1210_),
    .C(_1211_),
    .A(_1175_),
    .Y(_1212_));
 sg13g2_a21o_1 _4012_ (.A2(_1211_),
    .A1(_1210_),
    .B1(_1175_),
    .X(_1213_));
 sg13g2_nand3_1 _4013_ (.B(_1212_),
    .C(_1213_),
    .A(_1117_),
    .Y(_1214_));
 sg13g2_a21o_1 _4014_ (.A2(_1213_),
    .A1(_1212_),
    .B1(_1117_),
    .X(_1215_));
 sg13g2_o21ai_1 _4015_ (.B1(_1159_),
    .Y(_1216_),
    .A1(_1063_),
    .A2(_1160_));
 sg13g2_a21oi_1 _4016_ (.A1(_1214_),
    .A2(_1215_),
    .Y(_1217_),
    .B1(_1216_));
 sg13g2_nand3_1 _4017_ (.B(_1215_),
    .C(_1216_),
    .A(_1214_),
    .Y(_1218_));
 sg13g2_nor2b_1 _4018_ (.A(_1217_),
    .B_N(_1218_),
    .Y(_1219_));
 sg13g2_nand2_1 _4019_ (.Y(_1220_),
    .A(_1165_),
    .B(_1171_));
 sg13g2_xnor2_1 _4020_ (.Y(_1221_),
    .A(_1219_),
    .B(_1220_));
 sg13g2_a21oi_1 _4021_ (.A1(net539),
    .A2(_1221_),
    .Y(_0133_),
    .B1(_1174_));
 sg13g2_nand2b_1 _4022_ (.Y(_1222_),
    .B(_1210_),
    .A_N(_1208_));
 sg13g2_o21ai_1 _4023_ (.B1(net452),
    .Y(_1223_),
    .A1(_1184_),
    .A2(_1186_));
 sg13g2_or3_1 _4024_ (.A(net452),
    .B(_1184_),
    .C(_1186_),
    .X(_1224_));
 sg13g2_nand2_1 _4025_ (.Y(_1225_),
    .A(_1223_),
    .B(_1224_));
 sg13g2_nand2_1 _4026_ (.Y(_1226_),
    .A(_1204_),
    .B(_1206_));
 sg13g2_a22oi_1 _4027_ (.Y(_1227_),
    .B1(_1182_),
    .B2(_1068_),
    .A2(_1122_),
    .A1(_0446_));
 sg13g2_a21oi_1 _4028_ (.A1(_1132_),
    .A2(_1191_),
    .Y(_1228_),
    .B1(_1193_));
 sg13g2_nor2_1 _4029_ (.A(net450),
    .B(_1228_),
    .Y(_1229_));
 sg13g2_xnor2_1 _4030_ (.Y(_1230_),
    .A(_1183_),
    .B(_1228_));
 sg13g2_nor2_1 _4031_ (.A(_1227_),
    .B(_1230_),
    .Y(_1231_));
 sg13g2_xnor2_1 _4032_ (.Y(_1232_),
    .A(net449),
    .B(_1230_));
 sg13g2_nand2b_1 _4033_ (.Y(_1233_),
    .B(_1202_),
    .A_N(_1200_));
 sg13g2_nor2b_1 _4034_ (.A(_1196_),
    .B_N(_1198_),
    .Y(_1234_));
 sg13g2_nor2_1 _4035_ (.A(net491),
    .B(net475),
    .Y(_1235_));
 sg13g2_nand2_1 _4036_ (.Y(_1236_),
    .A(net531),
    .B(net467));
 sg13g2_nor3_1 _4037_ (.A(net481),
    .B(net471),
    .C(_1236_),
    .Y(_1237_));
 sg13g2_xnor2_1 _4038_ (.Y(_1238_),
    .A(_1022_),
    .B(_1236_));
 sg13g2_xnor2_1 _4039_ (.Y(_1239_),
    .A(_1235_),
    .B(_1238_));
 sg13g2_or2_1 _4040_ (.X(_1240_),
    .B(_1239_),
    .A(_1234_));
 sg13g2_and2_1 _4041_ (.A(_1234_),
    .B(_1239_),
    .X(_1241_));
 sg13g2_xor2_1 _4042_ (.B(_1239_),
    .A(_1234_),
    .X(_1242_));
 sg13g2_nor2_2 _4043_ (.A(net486),
    .B(net471),
    .Y(_1243_));
 sg13g2_nor2_2 _4044_ (.A(net483),
    .B(net525),
    .Y(_1244_));
 sg13g2_nand2_1 _4045_ (.Y(_1245_),
    .A(_1190_),
    .B(_1244_));
 sg13g2_xor2_1 _4046_ (.B(_1244_),
    .A(_1190_),
    .X(_1246_));
 sg13g2_nand2_1 _4047_ (.Y(_1247_),
    .A(_1243_),
    .B(_1246_));
 sg13g2_xnor2_1 _4048_ (.Y(_1248_),
    .A(_1243_),
    .B(_1246_));
 sg13g2_xnor2_1 _4049_ (.Y(_1249_),
    .A(_1242_),
    .B(_1248_));
 sg13g2_nand2_1 _4050_ (.Y(_1250_),
    .A(_1233_),
    .B(_1249_));
 sg13g2_xnor2_1 _4051_ (.Y(_1251_),
    .A(_1233_),
    .B(_1249_));
 sg13g2_xor2_1 _4052_ (.B(_1251_),
    .A(_1232_),
    .X(_1252_));
 sg13g2_nand2_1 _4053_ (.Y(_1253_),
    .A(_1226_),
    .B(_1252_));
 sg13g2_xnor2_1 _4054_ (.Y(_1254_),
    .A(_1226_),
    .B(_1252_));
 sg13g2_xor2_1 _4055_ (.B(_1254_),
    .A(_1225_),
    .X(_1255_));
 sg13g2_nand2_1 _4056_ (.Y(_1256_),
    .A(_1222_),
    .B(_1255_));
 sg13g2_xnor2_1 _4057_ (.Y(_1257_),
    .A(_1222_),
    .B(_1255_));
 sg13g2_xor2_1 _4058_ (.B(_1257_),
    .A(_1177_),
    .X(_1258_));
 sg13g2_nand2_1 _4059_ (.Y(_1259_),
    .A(_1212_),
    .B(_1214_));
 sg13g2_nand2_1 _4060_ (.Y(_1260_),
    .A(_1258_),
    .B(_1259_));
 sg13g2_xor2_1 _4061_ (.B(_1259_),
    .A(_1258_),
    .X(_1261_));
 sg13g2_inv_1 _4062_ (.Y(_1262_),
    .A(_1261_));
 sg13g2_and2_1 _4063_ (.A(_1166_),
    .B(_1219_),
    .X(_1263_));
 sg13g2_a21oi_1 _4064_ (.A1(_1165_),
    .A2(_1218_),
    .Y(_1264_),
    .B1(_1217_));
 sg13g2_a21oi_1 _4065_ (.A1(_1170_),
    .A2(_1263_),
    .Y(_1265_),
    .B1(_1264_));
 sg13g2_xnor2_1 _4066_ (.Y(_1266_),
    .A(_1262_),
    .B(_1265_));
 sg13g2_nor2_1 _4067_ (.A(net794),
    .B(net539),
    .Y(_1267_));
 sg13g2_a21oi_1 _4068_ (.A1(net538),
    .A2(_1266_),
    .Y(_0134_),
    .B1(_1267_));
 sg13g2_nor2_1 _4069_ (.A(net803),
    .B(net538),
    .Y(_1268_));
 sg13g2_o21ai_1 _4070_ (.B1(_1256_),
    .Y(_1269_),
    .A1(_1177_),
    .A2(_1257_));
 sg13g2_o21ai_1 _4071_ (.B1(_1253_),
    .Y(_1270_),
    .A1(_1225_),
    .A2(_1254_));
 sg13g2_o21ai_1 _4072_ (.B1(net452),
    .Y(_1271_),
    .A1(_1229_),
    .A2(_1231_));
 sg13g2_or3_1 _4073_ (.A(net452),
    .B(_1229_),
    .C(_1231_),
    .X(_1272_));
 sg13g2_nand2_1 _4074_ (.Y(_1273_),
    .A(_1271_),
    .B(_1272_));
 sg13g2_o21ai_1 _4075_ (.B1(_1250_),
    .Y(_1274_),
    .A1(_1232_),
    .A2(_1251_));
 sg13g2_o21ai_1 _4076_ (.B1(_1240_),
    .Y(_1275_),
    .A1(_1241_),
    .A2(_1248_));
 sg13g2_a21oi_2 _4077_ (.B1(_1237_),
    .Y(_1276_),
    .A2(_1238_),
    .A1(_1235_));
 sg13g2_nor2_1 _4078_ (.A(_0481_),
    .B(net469),
    .Y(_1277_));
 sg13g2_xnor2_1 _4079_ (.Y(_1278_),
    .A(_1022_),
    .B(_1277_));
 sg13g2_nor2_1 _4080_ (.A(net527),
    .B(net475),
    .Y(_1279_));
 sg13g2_nor2b_1 _4081_ (.A(_1278_),
    .B_N(_1279_),
    .Y(_1280_));
 sg13g2_xnor2_1 _4082_ (.Y(_1281_),
    .A(_1278_),
    .B(_1279_));
 sg13g2_nand2b_1 _4083_ (.Y(_1282_),
    .B(_1281_),
    .A_N(_1276_));
 sg13g2_nor2b_1 _4084_ (.A(_1281_),
    .B_N(_1276_),
    .Y(_1283_));
 sg13g2_xnor2_1 _4085_ (.Y(_1284_),
    .A(_1276_),
    .B(_1281_));
 sg13g2_nor2_1 _4086_ (.A(net483),
    .B(net471),
    .Y(_1285_));
 sg13g2_a21oi_1 _4087_ (.A1(_0537_),
    .A2(_0568_),
    .Y(_1286_),
    .B1(_1285_));
 sg13g2_nor2_2 _4088_ (.A(net477),
    .B(net471),
    .Y(_1287_));
 sg13g2_a21oi_1 _4089_ (.A1(_1244_),
    .A2(_1287_),
    .Y(_1288_),
    .B1(_1286_));
 sg13g2_xnor2_1 _4090_ (.Y(_1289_),
    .A(_1243_),
    .B(_1288_));
 sg13g2_xnor2_1 _4091_ (.Y(_1290_),
    .A(_1284_),
    .B(_1289_));
 sg13g2_nand2_1 _4092_ (.Y(_1291_),
    .A(_1275_),
    .B(_1290_));
 sg13g2_xnor2_1 _4093_ (.Y(_1292_),
    .A(_1275_),
    .B(_1290_));
 sg13g2_a21oi_1 _4094_ (.A1(_1245_),
    .A2(_1247_),
    .Y(_1293_),
    .B1(net450));
 sg13g2_nand3_1 _4095_ (.B(_1245_),
    .C(_1247_),
    .A(net450),
    .Y(_1294_));
 sg13g2_nand2b_1 _4096_ (.Y(_1295_),
    .B(_1294_),
    .A_N(_1293_));
 sg13g2_nor2_1 _4097_ (.A(net449),
    .B(_1295_),
    .Y(_1296_));
 sg13g2_xor2_1 _4098_ (.B(_1295_),
    .A(net449),
    .X(_1297_));
 sg13g2_inv_1 _4099_ (.Y(_1298_),
    .A(_1297_));
 sg13g2_xnor2_1 _4100_ (.Y(_1299_),
    .A(_1292_),
    .B(_1297_));
 sg13g2_nand2_1 _4101_ (.Y(_1300_),
    .A(_1274_),
    .B(_1299_));
 sg13g2_xnor2_1 _4102_ (.Y(_1301_),
    .A(_1274_),
    .B(_1299_));
 sg13g2_xor2_1 _4103_ (.B(_1301_),
    .A(_1273_),
    .X(_1302_));
 sg13g2_xnor2_1 _4104_ (.Y(_1303_),
    .A(_1270_),
    .B(_1302_));
 sg13g2_nor2_1 _4105_ (.A(_1223_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_xor2_1 _4106_ (.B(_1303_),
    .A(_1223_),
    .X(_1305_));
 sg13g2_nor2_1 _4107_ (.A(_1269_),
    .B(_1305_),
    .Y(_1306_));
 sg13g2_xor2_1 _4108_ (.B(_1305_),
    .A(_1269_),
    .X(_1307_));
 sg13g2_o21ai_1 _4109_ (.B1(_1260_),
    .Y(_1308_),
    .A1(_1262_),
    .A2(_1265_));
 sg13g2_xnor2_1 _4110_ (.Y(_1309_),
    .A(_1307_),
    .B(_1308_));
 sg13g2_a21oi_1 _4111_ (.A1(net538),
    .A2(_1309_),
    .Y(_0135_),
    .B1(_1268_));
 sg13g2_nor2_1 _4112_ (.A(net767),
    .B(net539),
    .Y(_1310_));
 sg13g2_o21ai_1 _4113_ (.B1(_1300_),
    .Y(_1311_),
    .A1(_1273_),
    .A2(_1301_));
 sg13g2_o21ai_1 _4114_ (.B1(net452),
    .Y(_1312_),
    .A1(_1293_),
    .A2(_1296_));
 sg13g2_or3_1 _4115_ (.A(net452),
    .B(_1293_),
    .C(_1296_),
    .X(_1313_));
 sg13g2_nand2_1 _4116_ (.Y(_1314_),
    .A(_1312_),
    .B(_1313_));
 sg13g2_o21ai_1 _4117_ (.B1(_1291_),
    .Y(_1315_),
    .A1(_1292_),
    .A2(_1298_));
 sg13g2_o21ai_1 _4118_ (.B1(_1282_),
    .Y(_1316_),
    .A1(_1283_),
    .A2(_1289_));
 sg13g2_a21oi_1 _4119_ (.A1(_1022_),
    .A2(_1277_),
    .Y(_1317_),
    .B1(_1280_));
 sg13g2_nor2_1 _4120_ (.A(_0487_),
    .B(net469),
    .Y(_1318_));
 sg13g2_xnor2_1 _4121_ (.Y(_1319_),
    .A(_1022_),
    .B(_1318_));
 sg13g2_nor2_1 _4122_ (.A(net525),
    .B(net475),
    .Y(_1320_));
 sg13g2_nor2b_1 _4123_ (.A(_1319_),
    .B_N(_1320_),
    .Y(_1321_));
 sg13g2_xnor2_1 _4124_ (.Y(_1322_),
    .A(_1319_),
    .B(_1320_));
 sg13g2_nor2b_1 _4125_ (.A(_1317_),
    .B_N(_1322_),
    .Y(_1323_));
 sg13g2_xnor2_1 _4126_ (.Y(_1324_),
    .A(_1317_),
    .B(_1322_));
 sg13g2_nand2_1 _4127_ (.Y(_1325_),
    .A(_0517_),
    .B(_1287_));
 sg13g2_o21ai_1 _4128_ (.B1(_1325_),
    .Y(_1326_),
    .A1(_1285_),
    .A2(_1287_));
 sg13g2_or3_1 _4129_ (.A(net486),
    .B(net471),
    .C(_1326_),
    .X(_1327_));
 sg13g2_xor2_1 _4130_ (.B(_1326_),
    .A(_1243_),
    .X(_1328_));
 sg13g2_inv_1 _4131_ (.Y(_1329_),
    .A(_1328_));
 sg13g2_xnor2_1 _4132_ (.Y(_1330_),
    .A(_1324_),
    .B(_1328_));
 sg13g2_nand2_1 _4133_ (.Y(_1331_),
    .A(_1316_),
    .B(_1330_));
 sg13g2_xnor2_1 _4134_ (.Y(_1332_),
    .A(_1316_),
    .B(_1330_));
 sg13g2_a22oi_1 _4135_ (.Y(_1333_),
    .B1(_1288_),
    .B2(_1243_),
    .A2(_1287_),
    .A1(_1244_));
 sg13g2_nor2_1 _4136_ (.A(net450),
    .B(_1333_),
    .Y(_1334_));
 sg13g2_xnor2_1 _4137_ (.Y(_1335_),
    .A(net450),
    .B(_1333_));
 sg13g2_nor2_1 _4138_ (.A(net449),
    .B(_1335_),
    .Y(_1336_));
 sg13g2_xor2_1 _4139_ (.B(_1335_),
    .A(net449),
    .X(_1337_));
 sg13g2_inv_1 _4140_ (.Y(_1338_),
    .A(_1337_));
 sg13g2_xnor2_1 _4141_ (.Y(_1339_),
    .A(_1332_),
    .B(_1337_));
 sg13g2_nand2_1 _4142_ (.Y(_1340_),
    .A(_1315_),
    .B(_1339_));
 sg13g2_xnor2_1 _4143_ (.Y(_1341_),
    .A(_1315_),
    .B(_1339_));
 sg13g2_xor2_1 _4144_ (.B(_1341_),
    .A(_1314_),
    .X(_1342_));
 sg13g2_and2_1 _4145_ (.A(_1311_),
    .B(_1342_),
    .X(_1343_));
 sg13g2_xnor2_1 _4146_ (.Y(_1344_),
    .A(_1311_),
    .B(_1342_));
 sg13g2_nor2_1 _4147_ (.A(_1271_),
    .B(_1344_),
    .Y(_1345_));
 sg13g2_xor2_1 _4148_ (.B(_1344_),
    .A(_1271_),
    .X(_1346_));
 sg13g2_a21oi_1 _4149_ (.A1(_1270_),
    .A2(_1302_),
    .Y(_1347_),
    .B1(_1304_));
 sg13g2_nand2b_1 _4150_ (.Y(_1348_),
    .B(_1346_),
    .A_N(_1347_));
 sg13g2_inv_1 _4151_ (.Y(_1349_),
    .A(_1348_));
 sg13g2_xnor2_1 _4152_ (.Y(_1350_),
    .A(_1346_),
    .B(_1347_));
 sg13g2_and3_1 _4153_ (.X(_1351_),
    .A(_1261_),
    .B(_1263_),
    .C(_1307_));
 sg13g2_nand3_1 _4154_ (.B(_1264_),
    .C(_1307_),
    .A(_1261_),
    .Y(_1352_));
 sg13g2_a22oi_1 _4155_ (.Y(_1353_),
    .B1(_1269_),
    .B2(_1305_),
    .A2(_1259_),
    .A1(_1258_));
 sg13g2_o21ai_1 _4156_ (.B1(_1352_),
    .Y(_1354_),
    .A1(_1306_),
    .A2(_1353_));
 sg13g2_a21o_1 _4157_ (.A2(_1351_),
    .A1(_1170_),
    .B1(_1354_),
    .X(_1355_));
 sg13g2_xnor2_1 _4158_ (.Y(_1356_),
    .A(_1350_),
    .B(_1355_));
 sg13g2_a21oi_1 _4159_ (.A1(net538),
    .A2(_1356_),
    .Y(_0136_),
    .B1(_1310_));
 sg13g2_nor2_1 _4160_ (.A(net804),
    .B(net538),
    .Y(_1357_));
 sg13g2_o21ai_1 _4161_ (.B1(_1340_),
    .Y(_1358_),
    .A1(_1314_),
    .A2(_1341_));
 sg13g2_nor2_1 _4162_ (.A(_1334_),
    .B(_1336_),
    .Y(_1359_));
 sg13g2_nor2_1 _4163_ (.A(_0999_),
    .B(_1359_),
    .Y(_1360_));
 sg13g2_xnor2_1 _4164_ (.Y(_1361_),
    .A(_0999_),
    .B(_1359_));
 sg13g2_o21ai_1 _4165_ (.B1(_1331_),
    .Y(_1362_),
    .A1(_1332_),
    .A2(_1338_));
 sg13g2_a21o_1 _4166_ (.A2(_1329_),
    .A1(_1324_),
    .B1(_1323_),
    .X(_1363_));
 sg13g2_a21oi_2 _4167_ (.B1(_1321_),
    .Y(_1364_),
    .A2(_1318_),
    .A1(_1022_));
 sg13g2_nor2_1 _4168_ (.A(_0568_),
    .B(net469),
    .Y(_1365_));
 sg13g2_nand2_1 _4169_ (.Y(_1366_),
    .A(_1022_),
    .B(_1365_));
 sg13g2_xnor2_1 _4170_ (.Y(_1367_),
    .A(_1022_),
    .B(_1365_));
 sg13g2_nor2_1 _4171_ (.A(net475),
    .B(net471),
    .Y(_1368_));
 sg13g2_nand2b_1 _4172_ (.Y(_1369_),
    .B(_1368_),
    .A_N(_1367_));
 sg13g2_xnor2_1 _4173_ (.Y(_1370_),
    .A(_1367_),
    .B(_1368_));
 sg13g2_nand2b_1 _4174_ (.Y(_1371_),
    .B(_1370_),
    .A_N(_1364_));
 sg13g2_xnor2_1 _4175_ (.Y(_1372_),
    .A(_1364_),
    .B(_1370_));
 sg13g2_xnor2_1 _4176_ (.Y(_1373_),
    .A(_1328_),
    .B(_1372_));
 sg13g2_xnor2_1 _4177_ (.Y(_1374_),
    .A(_1363_),
    .B(_1373_));
 sg13g2_a21oi_1 _4178_ (.A1(_1325_),
    .A2(_1327_),
    .Y(_1375_),
    .B1(net450));
 sg13g2_nand3_1 _4179_ (.B(_1325_),
    .C(_1327_),
    .A(net450),
    .Y(_1376_));
 sg13g2_nor2b_1 _4180_ (.A(_1375_),
    .B_N(_1376_),
    .Y(_1377_));
 sg13g2_xnor2_1 _4181_ (.Y(_1378_),
    .A(net449),
    .B(_1377_));
 sg13g2_nor2b_1 _4182_ (.A(_1374_),
    .B_N(_1378_),
    .Y(_1379_));
 sg13g2_xnor2_1 _4183_ (.Y(_1380_),
    .A(_1374_),
    .B(_1378_));
 sg13g2_xnor2_1 _4184_ (.Y(_1381_),
    .A(_1362_),
    .B(_1380_));
 sg13g2_nor2_1 _4185_ (.A(_1361_),
    .B(_1381_),
    .Y(_1382_));
 sg13g2_xor2_1 _4186_ (.B(_1381_),
    .A(_1361_),
    .X(_1383_));
 sg13g2_nand2_1 _4187_ (.Y(_1384_),
    .A(_1358_),
    .B(_1383_));
 sg13g2_xnor2_1 _4188_ (.Y(_1385_),
    .A(_1358_),
    .B(_1383_));
 sg13g2_xor2_1 _4189_ (.B(_1385_),
    .A(_1312_),
    .X(_1386_));
 sg13g2_nor3_1 _4190_ (.A(_1343_),
    .B(_1345_),
    .C(_1386_),
    .Y(_1387_));
 sg13g2_o21ai_1 _4191_ (.B1(_1386_),
    .Y(_1388_),
    .A1(_1343_),
    .A2(_1345_));
 sg13g2_nor2b_1 _4192_ (.A(_1387_),
    .B_N(_1388_),
    .Y(_1389_));
 sg13g2_a21oi_1 _4193_ (.A1(_1350_),
    .A2(_1355_),
    .Y(_1390_),
    .B1(_1349_));
 sg13g2_xor2_1 _4194_ (.B(_1390_),
    .A(_1389_),
    .X(_1391_));
 sg13g2_a21oi_1 _4195_ (.A1(net538),
    .A2(_1391_),
    .Y(_0137_),
    .B1(_1357_));
 sg13g2_and2_1 _4196_ (.A(_1350_),
    .B(_1389_),
    .X(_1392_));
 sg13g2_o21ai_1 _4197_ (.B1(_1388_),
    .Y(_1393_),
    .A1(_1348_),
    .A2(_1387_));
 sg13g2_a21oi_1 _4198_ (.A1(_1355_),
    .A2(_1392_),
    .Y(_1394_),
    .B1(_1393_));
 sg13g2_o21ai_1 _4199_ (.B1(_1384_),
    .Y(_1395_),
    .A1(_1312_),
    .A2(_1385_));
 sg13g2_a21oi_1 _4200_ (.A1(_1362_),
    .A2(_1380_),
    .Y(_1396_),
    .B1(_1382_));
 sg13g2_a21oi_1 _4201_ (.A1(_1363_),
    .A2(_1373_),
    .Y(_1397_),
    .B1(_1379_));
 sg13g2_nor2_1 _4202_ (.A(net449),
    .B(_1375_),
    .Y(_1398_));
 sg13g2_a21oi_1 _4203_ (.A1(net449),
    .A2(_1376_),
    .Y(_1399_),
    .B1(_1398_));
 sg13g2_a22oi_1 _4204_ (.Y(_1400_),
    .B1(_1366_),
    .B2(_1369_),
    .A2(_1022_),
    .A1(_0600_));
 sg13g2_nor2_1 _4205_ (.A(net480),
    .B(net471),
    .Y(_1401_));
 sg13g2_a221oi_1 _4206_ (.B2(net475),
    .C1(_1400_),
    .B1(_1401_),
    .A1(net471),
    .Y(_1402_),
    .A2(net469));
 sg13g2_xnor2_1 _4207_ (.Y(_1403_),
    .A(_1399_),
    .B(_1402_));
 sg13g2_nand2_1 _4208_ (.Y(_1404_),
    .A(_1329_),
    .B(_1364_));
 sg13g2_a22oi_1 _4209_ (.Y(_1405_),
    .B1(_1371_),
    .B2(_1404_),
    .A2(_1370_),
    .A1(_1329_));
 sg13g2_xnor2_1 _4210_ (.Y(_1406_),
    .A(_0999_),
    .B(_1405_));
 sg13g2_xnor2_1 _4211_ (.Y(_1407_),
    .A(_1403_),
    .B(_1406_));
 sg13g2_xnor2_1 _4212_ (.Y(_1408_),
    .A(_1397_),
    .B(_1407_));
 sg13g2_xnor2_1 _4213_ (.Y(_1409_),
    .A(_1396_),
    .B(_1408_));
 sg13g2_xnor2_1 _4214_ (.Y(_1410_),
    .A(_1360_),
    .B(_1409_));
 sg13g2_xnor2_1 _4215_ (.Y(_1411_),
    .A(_1395_),
    .B(_1410_));
 sg13g2_xnor2_1 _4216_ (.Y(_1412_),
    .A(_1394_),
    .B(_1411_));
 sg13g2_nor2_1 _4217_ (.A(net664),
    .B(net538),
    .Y(_1413_));
 sg13g2_a21oi_1 _4218_ (.A1(net538),
    .A2(_1412_),
    .Y(_0138_),
    .B1(_1413_));
 sg13g2_nor2_1 _4219_ (.A(net801),
    .B(net518),
    .Y(_1414_));
 sg13g2_a21oi_1 _4220_ (.A1(net518),
    .A2(_0774_),
    .Y(_0139_),
    .B1(_1414_));
 sg13g2_nor2_1 _4221_ (.A(net704),
    .B(net518),
    .Y(_1415_));
 sg13g2_a21oi_1 _4222_ (.A1(net518),
    .A2(_0852_),
    .Y(_0140_),
    .B1(_1415_));
 sg13g2_nor2_1 _4223_ (.A(net787),
    .B(net518),
    .Y(_1416_));
 sg13g2_a21oi_1 _4224_ (.A1(net518),
    .A2(_0924_),
    .Y(_0141_),
    .B1(_1416_));
 sg13g2_nor2_1 _4225_ (.A(net776),
    .B(net519),
    .Y(_1417_));
 sg13g2_a21oi_1 _4226_ (.A1(net519),
    .A2(_0993_),
    .Y(_0142_),
    .B1(_1417_));
 sg13g2_nor2_1 _4227_ (.A(net782),
    .B(net519),
    .Y(_1418_));
 sg13g2_a21oi_1 _4228_ (.A1(net519),
    .A2(_1057_),
    .Y(_0143_),
    .B1(_1418_));
 sg13g2_nor2_1 _4229_ (.A(net777),
    .B(net518),
    .Y(_1419_));
 sg13g2_a21oi_1 _4230_ (.A1(net518),
    .A2(_1113_),
    .Y(_0144_),
    .B1(_1419_));
 sg13g2_nor2_1 _4231_ (.A(net808),
    .B(net519),
    .Y(_1420_));
 sg13g2_a21oi_1 _4232_ (.A1(net517),
    .A2(_1172_),
    .Y(_0145_),
    .B1(_1420_));
 sg13g2_nor2_1 _4233_ (.A(net700),
    .B(net517),
    .Y(_1421_));
 sg13g2_a21oi_1 _4234_ (.A1(net517),
    .A2(_1221_),
    .Y(_0146_),
    .B1(_1421_));
 sg13g2_nor2_1 _4235_ (.A(net758),
    .B(net517),
    .Y(_1422_));
 sg13g2_a21oi_1 _4236_ (.A1(net516),
    .A2(_1266_),
    .Y(_0147_),
    .B1(_1422_));
 sg13g2_nor2_1 _4237_ (.A(net759),
    .B(net516),
    .Y(_1423_));
 sg13g2_a21oi_1 _4238_ (.A1(net516),
    .A2(_1309_),
    .Y(_0148_),
    .B1(_1423_));
 sg13g2_nor2_1 _4239_ (.A(net768),
    .B(net517),
    .Y(_1424_));
 sg13g2_a21oi_1 _4240_ (.A1(net516),
    .A2(_1356_),
    .Y(_0149_),
    .B1(_1424_));
 sg13g2_nor2_1 _4241_ (.A(net751),
    .B(net516),
    .Y(_1425_));
 sg13g2_a21oi_1 _4242_ (.A1(net516),
    .A2(_1391_),
    .Y(_0150_),
    .B1(_1425_));
 sg13g2_nor2_1 _4243_ (.A(net610),
    .B(net516),
    .Y(_1426_));
 sg13g2_a21oi_1 _4244_ (.A1(net516),
    .A2(_1412_),
    .Y(_0151_),
    .B1(_1426_));
 sg13g2_nor2_1 _4245_ (.A(net764),
    .B(net545),
    .Y(_1427_));
 sg13g2_a21oi_1 _4246_ (.A1(net545),
    .A2(_0774_),
    .Y(_0152_),
    .B1(_1427_));
 sg13g2_nor2_1 _4247_ (.A(net661),
    .B(net545),
    .Y(_1428_));
 sg13g2_a21oi_1 _4248_ (.A1(net545),
    .A2(_0852_),
    .Y(_0153_),
    .B1(_1428_));
 sg13g2_nor2_1 _4249_ (.A(net724),
    .B(net545),
    .Y(_1429_));
 sg13g2_a21oi_1 _4250_ (.A1(net545),
    .A2(_0924_),
    .Y(_0154_),
    .B1(_1429_));
 sg13g2_nor2_1 _4251_ (.A(net778),
    .B(net545),
    .Y(_1430_));
 sg13g2_a21oi_1 _4252_ (.A1(net545),
    .A2(_0993_),
    .Y(_0155_),
    .B1(_1430_));
 sg13g2_nor2_1 _4253_ (.A(net753),
    .B(net546),
    .Y(_1431_));
 sg13g2_a21oi_1 _4254_ (.A1(net546),
    .A2(_1057_),
    .Y(_0156_),
    .B1(net754));
 sg13g2_nor2_1 _4255_ (.A(net745),
    .B(net546),
    .Y(_1432_));
 sg13g2_a21oi_1 _4256_ (.A1(net546),
    .A2(_1113_),
    .Y(_0157_),
    .B1(net746));
 sg13g2_nor2_1 _4257_ (.A(net769),
    .B(net544),
    .Y(_1433_));
 sg13g2_a21oi_1 _4258_ (.A1(net544),
    .A2(_1172_),
    .Y(_0158_),
    .B1(_1433_));
 sg13g2_nor2_1 _4259_ (.A(net719),
    .B(net544),
    .Y(_1434_));
 sg13g2_a21oi_1 _4260_ (.A1(net543),
    .A2(_1221_),
    .Y(_0159_),
    .B1(_1434_));
 sg13g2_nor2_1 _4261_ (.A(net735),
    .B(net544),
    .Y(_1435_));
 sg13g2_a21oi_1 _4262_ (.A1(net543),
    .A2(_1266_),
    .Y(_0160_),
    .B1(_1435_));
 sg13g2_nor2_1 _4263_ (.A(net637),
    .B(net543),
    .Y(_1436_));
 sg13g2_a21oi_1 _4264_ (.A1(net543),
    .A2(_1309_),
    .Y(_0161_),
    .B1(_1436_));
 sg13g2_nor2_1 _4265_ (.A(net639),
    .B(net543),
    .Y(_1437_));
 sg13g2_a21oi_1 _4266_ (.A1(net543),
    .A2(_1356_),
    .Y(_0162_),
    .B1(_1437_));
 sg13g2_nor2_1 _4267_ (.A(net615),
    .B(net543),
    .Y(_1438_));
 sg13g2_a21oi_1 _4268_ (.A1(net543),
    .A2(_1391_),
    .Y(_0163_),
    .B1(_1438_));
 sg13g2_o21ai_1 _4269_ (.B1(net577),
    .Y(_1439_),
    .A1(net752),
    .A2(_0417_));
 sg13g2_a21oi_1 _4270_ (.A1(net752),
    .A2(_2048_),
    .Y(_0164_),
    .B1(_1439_));
 sg13g2_o21ai_1 _4271_ (.B1(net577),
    .Y(_1440_),
    .A1(_0059_),
    .A2(_2049_));
 sg13g2_and3_1 _4272_ (.X(_1441_),
    .A(net707),
    .B(\top.julia_calc.iter[0] ),
    .C(_2048_));
 sg13g2_a21oi_1 _4273_ (.A1(\top.julia_calc.iter[0] ),
    .A2(_2048_),
    .Y(_1442_),
    .B1(net707));
 sg13g2_nor3_1 _4274_ (.A(_1440_),
    .B(_1441_),
    .C(net708),
    .Y(_0165_));
 sg13g2_nor2_1 _4275_ (.A(net705),
    .B(_1441_),
    .Y(_1443_));
 sg13g2_and2_1 _4276_ (.A(net705),
    .B(_1441_),
    .X(_1444_));
 sg13g2_nor3_1 _4277_ (.A(_1440_),
    .B(net706),
    .C(_1444_),
    .Y(_0166_));
 sg13g2_xnor2_1 _4278_ (.Y(_1445_),
    .A(net800),
    .B(_1444_));
 sg13g2_nor2_1 _4279_ (.A(_1440_),
    .B(_1445_),
    .Y(_0167_));
 sg13g2_a21oi_1 _4280_ (.A1(\top.julia_calc.iter[3] ),
    .A2(_1444_),
    .Y(_1446_),
    .B1(net668));
 sg13g2_and3_1 _4281_ (.X(_1447_),
    .A(net668),
    .B(\top.julia_calc.iter[3] ),
    .C(_1444_));
 sg13g2_nor3_1 _4282_ (.A(_1440_),
    .B(net669),
    .C(_1447_),
    .Y(_0168_));
 sg13g2_nor2_1 _4283_ (.A(net722),
    .B(_1447_),
    .Y(_1448_));
 sg13g2_and2_1 _4284_ (.A(net722),
    .B(_1447_),
    .X(_1449_));
 sg13g2_nor3_1 _4285_ (.A(_1440_),
    .B(net723),
    .C(_1449_),
    .Y(_0169_));
 sg13g2_nand2_1 _4286_ (.Y(_1450_),
    .A(net737),
    .B(_1449_));
 sg13g2_xnor2_1 _4287_ (.Y(_1451_),
    .A(net737),
    .B(_1449_));
 sg13g2_nor2_1 _4288_ (.A(_1440_),
    .B(_1451_),
    .Y(_0170_));
 sg13g2_xor2_1 _4289_ (.B(_1450_),
    .A(net775),
    .X(_1452_));
 sg13g2_nor2_1 _4290_ (.A(_1440_),
    .B(_1452_),
    .Y(_0171_));
 sg13g2_nand4_1 _4291_ (.B(\top.julia_calc.iter[4] ),
    .C(\top.julia_calc.iter[3] ),
    .A(\top.julia_calc.iter[5] ),
    .Y(_1453_),
    .D(\top.julia_calc.iter[0] ));
 sg13g2_nand4_1 _4292_ (.B(\top.julia_calc.iter[6] ),
    .C(\top.julia_calc.iter[2] ),
    .A(\top.julia_calc.iter[7] ),
    .Y(_1454_),
    .D(\top.julia_calc.iter[1] ));
 sg13g2_nor2_2 _4293_ (.A(_1453_),
    .B(_1454_),
    .Y(_1455_));
 sg13g2_xnor2_1 _4294_ (.Y(_1456_),
    .A(_0056_),
    .B(_1455_));
 sg13g2_a22oi_1 _4295_ (.Y(_1457_),
    .B1(_2051_),
    .B2(_1456_),
    .A2(_2049_),
    .A1(net381));
 sg13g2_nor2_1 _4296_ (.A(net573),
    .B(net382),
    .Y(_0172_));
 sg13g2_nand3_1 _4297_ (.B(net756),
    .C(net857),
    .A(\top.receiver.receiver.counter[0] ),
    .Y(_1458_));
 sg13g2_or2_2 _4298_ (.X(_1459_),
    .B(_1458_),
    .A(\top.receiver.receiver.counter[3] ));
 sg13g2_nor2b_1 _4299_ (.A(\top.receiver.receiver.counter[1] ),
    .B_N(\top.receiver.receiver.counter[0] ),
    .Y(_1460_));
 sg13g2_nand4_1 _4300_ (.B(net884),
    .C(\rx_pins[0] ),
    .A(net642),
    .Y(_1461_),
    .D(_1460_));
 sg13g2_nand3_1 _4301_ (.B(_1459_),
    .C(_1461_),
    .A(net583),
    .Y(_1462_));
 sg13g2_or2_1 _4302_ (.X(_0173_),
    .B(_1462_),
    .A(net340));
 sg13g2_xnor2_1 _4303_ (.Y(_1463_),
    .A(\top.receiver.receiver.counter[0] ),
    .B(net756));
 sg13g2_nor2_1 _4304_ (.A(_1462_),
    .B(net757),
    .Y(_0174_));
 sg13g2_a21o_1 _4305_ (.A2(net756),
    .A1(\top.receiver.receiver.counter[0] ),
    .B1(net857),
    .X(_1464_));
 sg13g2_a21o_1 _4306_ (.A2(net858),
    .A1(_1458_),
    .B1(_1462_),
    .X(_0175_));
 sg13g2_a21o_1 _4307_ (.A2(_1458_),
    .A1(net642),
    .B1(_1462_),
    .X(_0176_));
 sg13g2_and2_2 _4308_ (.A(net871),
    .B(net761),
    .X(_1465_));
 sg13g2_nand2b_2 _4309_ (.Y(_1466_),
    .B(_1465_),
    .A_N(_1902_));
 sg13g2_nor4_2 _4310_ (.A(\top.rs.x[11] ),
    .B(_1901_),
    .C(_0344_),
    .Y(_1467_),
    .D(_1466_));
 sg13g2_nor4_2 _4311_ (.A(\top.rs.x[11] ),
    .B(_1901_),
    .C(_0344_),
    .Y(_1468_),
    .D(_1466_));
 sg13g2_nor2_1 _4312_ (.A(net576),
    .B(_1468_),
    .Y(_1469_));
 sg13g2_nand2b_1 _4313_ (.Y(_1470_),
    .B(net583),
    .A_N(_1468_));
 sg13g2_and2_1 _4314_ (.A(net328),
    .B(net451),
    .X(_0177_));
 sg13g2_nor3_1 _4315_ (.A(net575),
    .B(net762),
    .C(_1465_),
    .Y(_0178_));
 sg13g2_o21ai_1 _4316_ (.B1(net451),
    .Y(_1471_),
    .A1(net560),
    .A2(_1465_));
 sg13g2_a21oi_1 _4317_ (.A1(net560),
    .A2(_1465_),
    .Y(_0179_),
    .B1(_1471_));
 sg13g2_nor2b_1 _4318_ (.A(_0322_),
    .B_N(_1465_),
    .Y(_1472_));
 sg13g2_a21oi_1 _4319_ (.A1(net560),
    .A2(_1465_),
    .Y(_1473_),
    .B1(net559));
 sg13g2_nor3_1 _4320_ (.A(_1470_),
    .B(_1472_),
    .C(net848),
    .Y(_0180_));
 sg13g2_o21ai_1 _4321_ (.B1(_1469_),
    .Y(_1474_),
    .A1(net557),
    .A2(_1472_));
 sg13g2_a21oi_1 _4322_ (.A1(net557),
    .A2(_1472_),
    .Y(_0181_),
    .B1(_1474_));
 sg13g2_and2_1 _4323_ (.A(_0323_),
    .B(_1465_),
    .X(_1475_));
 sg13g2_a21oi_1 _4324_ (.A1(net557),
    .A2(_1472_),
    .Y(_1476_),
    .B1(net556));
 sg13g2_o21ai_1 _4325_ (.B1(net451),
    .Y(_0182_),
    .A1(_1475_),
    .A2(_1476_));
 sg13g2_o21ai_1 _4326_ (.B1(_1469_),
    .Y(_1477_),
    .A1(net805),
    .A2(_1475_));
 sg13g2_a21oi_1 _4327_ (.A1(net805),
    .A2(_1475_),
    .Y(_0183_),
    .B1(_1477_));
 sg13g2_a21oi_1 _4328_ (.A1(net805),
    .A2(_1475_),
    .Y(_1478_),
    .B1(net806));
 sg13g2_nor3_2 _4329_ (.A(_0321_),
    .B(_0322_),
    .C(_1466_),
    .Y(_1479_));
 sg13g2_o21ai_1 _4330_ (.B1(net451),
    .Y(_0184_),
    .A1(_1478_),
    .A2(_1479_));
 sg13g2_xor2_1 _4331_ (.B(_1479_),
    .A(net732),
    .X(_1480_));
 sg13g2_nand2_1 _4332_ (.Y(_0185_),
    .A(net451),
    .B(_1480_));
 sg13g2_nand2_1 _4333_ (.Y(_1481_),
    .A(net874),
    .B(_1479_));
 sg13g2_xnor2_1 _4334_ (.Y(_1482_),
    .A(_1842_),
    .B(_1481_));
 sg13g2_nand2_1 _4335_ (.Y(_0186_),
    .A(net451),
    .B(_1482_));
 sg13g2_o21ai_1 _4336_ (.B1(_1841_),
    .Y(_1483_),
    .A1(_1842_),
    .A2(_1481_));
 sg13g2_nand4_1 _4337_ (.B(\top.rs.x[8] ),
    .C(\top.rs.x[9] ),
    .A(net850),
    .Y(_1484_),
    .D(_1479_));
 sg13g2_a21o_1 _4338_ (.A2(net851),
    .A1(_1483_),
    .B1(_1470_),
    .X(_0187_));
 sg13g2_xor2_1 _4339_ (.B(net851),
    .A(net744),
    .X(_1485_));
 sg13g2_nand2_1 _4340_ (.Y(_0188_),
    .A(net451),
    .B(_1485_));
 sg13g2_nor2_2 _4341_ (.A(net574),
    .B(\top.buttons_stable ),
    .Y(_1486_));
 sg13g2_nand2_1 _4342_ (.Y(_1487_),
    .A(net412),
    .B(_1486_));
 sg13g2_o21ai_1 _4343_ (.B1(_1487_),
    .Y(_0189_),
    .A1(_1846_),
    .A2(_1486_));
 sg13g2_mux2_1 _4344_ (.A0(\top.debouncer_inst.last_data[1] ),
    .A1(net725),
    .S(_1486_),
    .X(_0190_));
 sg13g2_nand2_1 _4345_ (.Y(_1488_),
    .A(net592),
    .B(_1486_));
 sg13g2_o21ai_1 _4346_ (.B1(_1488_),
    .Y(_0191_),
    .A1(_1847_),
    .A2(_1486_));
 sg13g2_mux2_1 _4347_ (.A0(\top.debouncer_inst.last_data[3] ),
    .A1(net695),
    .S(_1486_),
    .X(_0192_));
 sg13g2_mux2_1 _4348_ (.A0(\top.debouncer_inst.last_data[4] ),
    .A1(net742),
    .S(_1486_),
    .X(_0193_));
 sg13g2_mux2_1 _4349_ (.A0(\top.debouncer_inst.last_data[5] ),
    .A1(net727),
    .S(_1486_),
    .X(_0194_));
 sg13g2_nor2b_2 _4350_ (.A(_0024_),
    .B_N(net7),
    .Y(_1489_));
 sg13g2_nand2_1 _4351_ (.Y(_1490_),
    .A(\top.debouncer_inst.last_data[4] ),
    .B(_1489_));
 sg13g2_nand3b_1 _4352_ (.B(\top.buttons_stable ),
    .C(\top.last_stable_buttons[4] ),
    .Y(_1491_),
    .A_N(\top.debouncer_inst.last_data[4] ));
 sg13g2_o21ai_1 _4353_ (.B1(_1491_),
    .Y(_1492_),
    .A1(\top.last_stable_buttons[4] ),
    .A2(_1490_));
 sg13g2_nor2_1 _4354_ (.A(net555),
    .B(net551),
    .Y(_1493_));
 sg13g2_nand3_1 _4355_ (.B(net554),
    .C(_1493_),
    .A(net549),
    .Y(_1494_));
 sg13g2_nand2_1 _4356_ (.Y(_1495_),
    .A(_1492_),
    .B(_1494_));
 sg13g2_nand2_1 _4357_ (.Y(_1496_),
    .A(\top.debouncer_inst.last_data[5] ),
    .B(_1489_));
 sg13g2_nand3b_1 _4358_ (.B(\top.buttons_stable ),
    .C(\top.last_stable_buttons[5] ),
    .Y(_1497_),
    .A_N(\top.debouncer_inst.last_data[5] ));
 sg13g2_o21ai_1 _4359_ (.B1(_1497_),
    .Y(_1498_),
    .A1(\top.last_stable_buttons[5] ),
    .A2(_1496_));
 sg13g2_nand2b_1 _4360_ (.Y(_1499_),
    .B(_1493_),
    .A_N(net549));
 sg13g2_o21ai_1 _4361_ (.B1(_1498_),
    .Y(_1500_),
    .A1(net554),
    .A2(_1499_));
 sg13g2_nor2b_2 _4362_ (.A(_1500_),
    .B_N(_1495_),
    .Y(_1501_));
 sg13g2_xnor2_1 _4363_ (.Y(_1502_),
    .A(_1495_),
    .B(_1500_));
 sg13g2_and2_1 _4364_ (.A(_1852_),
    .B(_1502_),
    .X(_1503_));
 sg13g2_nor2_1 _4365_ (.A(_1852_),
    .B(_1502_),
    .Y(_1504_));
 sg13g2_nor3_1 _4366_ (.A(net574),
    .B(_1503_),
    .C(_1504_),
    .Y(_0195_));
 sg13g2_and2_1 _4367_ (.A(net553),
    .B(_1501_),
    .X(_1505_));
 sg13g2_xnor2_1 _4368_ (.Y(_1506_),
    .A(_1853_),
    .B(_1501_));
 sg13g2_nor2_1 _4369_ (.A(_1504_),
    .B(_1506_),
    .Y(_1507_));
 sg13g2_and2_1 _4370_ (.A(_1504_),
    .B(_1506_),
    .X(_1508_));
 sg13g2_nor3_1 _4371_ (.A(net574),
    .B(_1507_),
    .C(_1508_),
    .Y(_0196_));
 sg13g2_nor2_1 _4372_ (.A(_0026_),
    .B(_1501_),
    .Y(_1509_));
 sg13g2_xnor2_1 _4373_ (.Y(_1510_),
    .A(net881),
    .B(_1501_));
 sg13g2_o21ai_1 _4374_ (.B1(_1510_),
    .Y(_1511_),
    .A1(_1505_),
    .A2(_1508_));
 sg13g2_or3_1 _4375_ (.A(_1505_),
    .B(_1508_),
    .C(_1510_),
    .X(_1512_));
 sg13g2_a21o_1 _4376_ (.A2(_1512_),
    .A1(_1511_),
    .B1(net574),
    .X(_0197_));
 sg13g2_and2_1 _4377_ (.A(net521),
    .B(_1501_),
    .X(_1513_));
 sg13g2_a22oi_1 _4378_ (.Y(_1514_),
    .B1(_1511_),
    .B2(_1513_),
    .A2(_1509_),
    .A1(_1508_));
 sg13g2_o21ai_1 _4379_ (.B1(net579),
    .Y(_1515_),
    .A1(net548),
    .A2(_1514_));
 sg13g2_a21oi_1 _4380_ (.A1(net548),
    .A2(_1514_),
    .Y(_0198_),
    .B1(_1515_));
 sg13g2_nor3_1 _4381_ (.A(net542),
    .B(_0320_),
    .C(_1459_),
    .Y(_1516_));
 sg13g2_mux2_1 _4382_ (.A0(\top.pixel_buffer[8][0] ),
    .A1(net691),
    .S(net460),
    .X(_0199_));
 sg13g2_mux2_1 _4383_ (.A0(\top.pixel_buffer[8][1] ),
    .A1(net677),
    .S(net460),
    .X(_0200_));
 sg13g2_mux2_1 _4384_ (.A0(net729),
    .A1(net322),
    .S(net460),
    .X(_0201_));
 sg13g2_mux2_1 _4385_ (.A0(net679),
    .A1(net323),
    .S(net460),
    .X(_0202_));
 sg13g2_mux2_1 _4386_ (.A0(net681),
    .A1(net329),
    .S(net460),
    .X(_0203_));
 sg13g2_mux2_1 _4387_ (.A0(net588),
    .A1(net333),
    .S(net459),
    .X(_0204_));
 sg13g2_mux2_1 _4388_ (.A0(net587),
    .A1(net332),
    .S(net459),
    .X(_0205_));
 sg13g2_mux2_1 _4389_ (.A0(net604),
    .A1(net326),
    .S(net459),
    .X(_0206_));
 sg13g2_mux2_1 _4390_ (.A0(net430),
    .A1(net331),
    .S(net459),
    .X(_0207_));
 sg13g2_mux2_1 _4391_ (.A0(net585),
    .A1(net337),
    .S(net459),
    .X(_0208_));
 sg13g2_mux2_1 _4392_ (.A0(net594),
    .A1(net324),
    .S(net460),
    .X(_0209_));
 sg13g2_mux2_1 _4393_ (.A0(net611),
    .A1(net334),
    .S(net461),
    .X(_0210_));
 sg13g2_mux2_1 _4394_ (.A0(net627),
    .A1(net325),
    .S(net460),
    .X(_0211_));
 sg13g2_mux2_1 _4395_ (.A0(net614),
    .A1(net327),
    .S(net459),
    .X(_0212_));
 sg13g2_nor2_1 _4396_ (.A(net586),
    .B(net461),
    .Y(_1517_));
 sg13g2_a21oi_1 _4397_ (.A1(_1845_),
    .A2(net460),
    .Y(_0213_),
    .B1(_1517_));
 sg13g2_nor2_1 _4398_ (.A(net633),
    .B(net459),
    .Y(_1518_));
 sg13g2_a21oi_1 _4399_ (.A1(_1851_),
    .A2(net459),
    .Y(_0214_),
    .B1(_1518_));
 sg13g2_a21o_1 _4400_ (.A2(net441),
    .A1(net659),
    .B1(_2028_),
    .X(_0215_));
 sg13g2_mux2_1 _4401_ (.A0(\top.julia_calc.dest_x[4] ),
    .A1(net629),
    .S(net441),
    .X(_0216_));
 sg13g2_mux2_1 _4402_ (.A0(\top.julia_calc.dest_x[5] ),
    .A1(net684),
    .S(net440),
    .X(_0217_));
 sg13g2_mux2_1 _4403_ (.A0(\top.julia_calc.dest_x[6] ),
    .A1(net665),
    .S(net441),
    .X(_0218_));
 sg13g2_mux2_1 _4404_ (.A0(\top.julia_calc.dest_x[7] ),
    .A1(net717),
    .S(net441),
    .X(_0219_));
 sg13g2_mux2_1 _4405_ (.A0(\top.julia_calc.dest_x[8] ),
    .A1(net618),
    .S(net441),
    .X(_0220_));
 sg13g2_mux2_1 _4406_ (.A0(\top.julia_calc.dest_y[0] ),
    .A1(net671),
    .S(net440),
    .X(_0221_));
 sg13g2_mux2_1 _4407_ (.A0(\top.julia_calc.dest_y[1] ),
    .A1(net675),
    .S(net440),
    .X(_0222_));
 sg13g2_nor2_1 _4408_ (.A(net599),
    .B(net439),
    .Y(_1519_));
 sg13g2_a21oi_1 _4409_ (.A1(_1838_),
    .A2(net439),
    .Y(_0223_),
    .B1(_1519_));
 sg13g2_mux2_1 _4410_ (.A0(\top.julia_calc.dest_y[3] ),
    .A1(net682),
    .S(net440),
    .X(_0224_));
 sg13g2_nor2_1 _4411_ (.A(net616),
    .B(net439),
    .Y(_1520_));
 sg13g2_a21oi_1 _4412_ (.A1(_1839_),
    .A2(net439),
    .Y(_0225_),
    .B1(_1520_));
 sg13g2_mux2_1 _4413_ (.A0(\top.julia_calc.dest_y[5] ),
    .A1(net733),
    .S(net440),
    .X(_0226_));
 sg13g2_nor2_1 _4414_ (.A(net635),
    .B(net439),
    .Y(_1521_));
 sg13g2_a21oi_1 _4415_ (.A1(_1840_),
    .A2(net439),
    .Y(_0227_),
    .B1(_1521_));
 sg13g2_mux2_1 _4416_ (.A0(\top.julia_calc.dest_y[7] ),
    .A1(net673),
    .S(net440),
    .X(_0228_));
 sg13g2_mux2_1 _4417_ (.A0(net624),
    .A1(net628),
    .S(net440),
    .X(_0229_));
 sg13g2_a21oi_1 _4418_ (.A1(\top.debouncer_inst.last_data[1] ),
    .A2(net7),
    .Y(_1522_),
    .B1(\top.last_stable_buttons[1] ));
 sg13g2_a21oi_1 _4419_ (.A1(\top.debouncer_inst.last_data[1] ),
    .A2(\top.last_stable_buttons[1] ),
    .Y(_1523_),
    .B1(_0024_));
 sg13g2_nand2b_2 _4420_ (.Y(_1524_),
    .B(_1523_),
    .A_N(_1522_));
 sg13g2_nor2b_1 _4421_ (.A(\top.last_stable_buttons[0] ),
    .B_N(\top.debouncer_inst.last_data[0] ),
    .Y(_1525_));
 sg13g2_nor2b_1 _4422_ (.A(\top.debouncer_inst.last_data[0] ),
    .B_N(\top.last_stable_buttons[0] ),
    .Y(_1526_));
 sg13g2_a22oi_1 _4423_ (.Y(_1527_),
    .B1(_1526_),
    .B2(\top.buttons_stable ),
    .A2(_1525_),
    .A1(_1489_));
 sg13g2_nor2b_2 _4424_ (.A(_1524_),
    .B_N(_1527_),
    .Y(_1528_));
 sg13g2_xnor2_1 _4425_ (.Y(_1529_),
    .A(_1524_),
    .B(_1527_));
 sg13g2_nor2_1 _4426_ (.A(\top.step_size[0] ),
    .B(_1529_),
    .Y(_1530_));
 sg13g2_nor4_2 _4427_ (.A(net555),
    .B(net554),
    .C(net551),
    .Y(_1531_),
    .D(_1529_));
 sg13g2_inv_1 _4428_ (.Y(_1532_),
    .A(_1531_));
 sg13g2_a21oi_1 _4429_ (.A1(net548),
    .A2(_1531_),
    .Y(_1533_),
    .B1(net771));
 sg13g2_and3_1 _4430_ (.X(_1534_),
    .A(net771),
    .B(net548),
    .C(_1531_));
 sg13g2_nor3_1 _4431_ (.A(net575),
    .B(net772),
    .C(_1534_),
    .Y(_0230_));
 sg13g2_nand3b_1 _4432_ (.B(net555),
    .C(_1524_),
    .Y(_1535_),
    .A_N(_1527_));
 sg13g2_nor2b_1 _4433_ (.A(_1528_),
    .B_N(_1535_),
    .Y(_1536_));
 sg13g2_nand3b_1 _4434_ (.B(_1854_),
    .C(_1853_),
    .Y(_1537_),
    .A_N(_1536_));
 sg13g2_nor3_1 _4435_ (.A(_1849_),
    .B(_1855_),
    .C(_1537_),
    .Y(_1538_));
 sg13g2_o21ai_1 _4436_ (.B1(_1849_),
    .Y(_1539_),
    .A1(_1855_),
    .A2(_1537_));
 sg13g2_nor2b_1 _4437_ (.A(_1538_),
    .B_N(_1539_),
    .Y(_1540_));
 sg13g2_xnor2_1 _4438_ (.Y(_1541_),
    .A(_1534_),
    .B(_1540_));
 sg13g2_nand2_1 _4439_ (.Y(_0231_),
    .A(net581),
    .B(_1541_));
 sg13g2_a21oi_2 _4440_ (.B1(_1538_),
    .Y(_1542_),
    .A2(_1539_),
    .A1(_1534_));
 sg13g2_or2_1 _4441_ (.X(_1543_),
    .B(_1528_),
    .A(net554));
 sg13g2_o21ai_1 _4442_ (.B1(_1543_),
    .Y(_1544_),
    .A1(_1853_),
    .A2(_1530_));
 sg13g2_nand3b_1 _4443_ (.B(net521),
    .C(net548),
    .Y(_1545_),
    .A_N(_1544_));
 sg13g2_or2_1 _4444_ (.X(_1546_),
    .B(_1545_),
    .A(_1848_));
 sg13g2_xnor2_1 _4445_ (.Y(_1547_),
    .A(_1848_),
    .B(_1545_));
 sg13g2_o21ai_1 _4446_ (.B1(net579),
    .Y(_1548_),
    .A1(_1542_),
    .A2(_1547_));
 sg13g2_a21oi_1 _4447_ (.A1(_1542_),
    .A2(_1547_),
    .Y(_0232_),
    .B1(_1548_));
 sg13g2_nor2b_2 _4448_ (.A(_1536_),
    .B_N(_1543_),
    .Y(_1549_));
 sg13g2_nand2_1 _4449_ (.Y(_1550_),
    .A(net521),
    .B(_1549_));
 sg13g2_nand3_1 _4450_ (.B(net548),
    .C(_1549_),
    .A(net521),
    .Y(_1551_));
 sg13g2_nor2_1 _4451_ (.A(net862),
    .B(_1551_),
    .Y(_1552_));
 sg13g2_xor2_1 _4452_ (.B(_1551_),
    .A(net862),
    .X(_1553_));
 sg13g2_o21ai_1 _4453_ (.B1(_1546_),
    .Y(_1554_),
    .A1(_1542_),
    .A2(_1547_));
 sg13g2_xnor2_1 _4454_ (.Y(_1555_),
    .A(_1553_),
    .B(_1554_));
 sg13g2_nand2_1 _4455_ (.Y(_0233_),
    .A(net579),
    .B(_1555_));
 sg13g2_a21oi_2 _4456_ (.B1(_1552_),
    .Y(_1556_),
    .A2(_1554_),
    .A1(_1553_));
 sg13g2_o21ai_1 _4457_ (.B1(net548),
    .Y(_1557_),
    .A1(net552),
    .A2(_1528_));
 sg13g2_inv_1 _4458_ (.Y(_1558_),
    .A(_1557_));
 sg13g2_a21oi_1 _4459_ (.A1(_1853_),
    .A2(_1530_),
    .Y(_1559_),
    .B1(_1854_));
 sg13g2_nor2_1 _4460_ (.A(_1557_),
    .B(_1559_),
    .Y(_1560_));
 sg13g2_nand2_1 _4461_ (.Y(_1561_),
    .A(\top.c_y[4] ),
    .B(_1560_));
 sg13g2_xnor2_1 _4462_ (.Y(_1562_),
    .A(\top.c_y[4] ),
    .B(_1560_));
 sg13g2_xnor2_1 _4463_ (.Y(_1563_),
    .A(_1556_),
    .B(_1562_));
 sg13g2_nand2_1 _4464_ (.Y(_0234_),
    .A(net580),
    .B(_1563_));
 sg13g2_o21ai_1 _4465_ (.B1(net552),
    .Y(_1564_),
    .A1(net554),
    .A2(_1536_));
 sg13g2_and2_1 _4466_ (.A(_1558_),
    .B(_1564_),
    .X(_1565_));
 sg13g2_nor2b_1 _4467_ (.A(net867),
    .B_N(_1565_),
    .Y(_1566_));
 sg13g2_xnor2_1 _4468_ (.Y(_1567_),
    .A(net867),
    .B(_1565_));
 sg13g2_o21ai_1 _4469_ (.B1(_1561_),
    .Y(_1568_),
    .A1(_1556_),
    .A2(_1562_));
 sg13g2_xnor2_1 _4470_ (.Y(_1569_),
    .A(_1567_),
    .B(_1568_));
 sg13g2_nand2_1 _4471_ (.Y(_0235_),
    .A(net580),
    .B(_1569_));
 sg13g2_a21oi_1 _4472_ (.A1(_1567_),
    .A2(_1568_),
    .Y(_1570_),
    .B1(_1566_));
 sg13g2_a21oi_1 _4473_ (.A1(net552),
    .A2(_1544_),
    .Y(_1571_),
    .B1(_1557_));
 sg13g2_xnor2_1 _4474_ (.Y(_1572_),
    .A(\top.c_y[6] ),
    .B(_1571_));
 sg13g2_nor2_1 _4475_ (.A(_1570_),
    .B(_1572_),
    .Y(_1573_));
 sg13g2_and2_1 _4476_ (.A(_1570_),
    .B(_1572_),
    .X(_1574_));
 sg13g2_o21ai_1 _4477_ (.B1(net579),
    .Y(_0236_),
    .A1(_1573_),
    .A2(_1574_));
 sg13g2_a21oi_1 _4478_ (.A1(net870),
    .A2(_1571_),
    .Y(_1575_),
    .B1(_1573_));
 sg13g2_nand3_1 _4479_ (.B(_1549_),
    .C(_1558_),
    .A(\top.c_y[7] ),
    .Y(_1576_));
 sg13g2_a21o_1 _4480_ (.A2(_1558_),
    .A1(_1549_),
    .B1(\top.c_y[7] ),
    .X(_1577_));
 sg13g2_nand2_1 _4481_ (.Y(_1578_),
    .A(_1576_),
    .B(_1577_));
 sg13g2_or2_1 _4482_ (.X(_1579_),
    .B(_1578_),
    .A(_1575_));
 sg13g2_nand2_1 _4483_ (.Y(_1580_),
    .A(net579),
    .B(_1579_));
 sg13g2_a21oi_1 _4484_ (.A1(_1575_),
    .A2(_1578_),
    .Y(_0237_),
    .B1(_1580_));
 sg13g2_nor2_1 _4485_ (.A(net550),
    .B(_1528_),
    .Y(_1581_));
 sg13g2_or2_1 _4486_ (.X(_1582_),
    .B(_1528_),
    .A(net550));
 sg13g2_a21oi_1 _4487_ (.A1(net550),
    .A2(_1532_),
    .Y(_1583_),
    .B1(_1581_));
 sg13g2_nand2_1 _4488_ (.Y(_1584_),
    .A(\top.c_y[8] ),
    .B(_1583_));
 sg13g2_xnor2_1 _4489_ (.Y(_1585_),
    .A(\top.c_y[8] ),
    .B(_1583_));
 sg13g2_nand3_1 _4490_ (.B(_1579_),
    .C(_1585_),
    .A(_1576_),
    .Y(_1586_));
 sg13g2_a21o_1 _4491_ (.A2(_1579_),
    .A1(_1576_),
    .B1(_1585_),
    .X(_1587_));
 sg13g2_and3_1 _4492_ (.X(_0238_),
    .A(net579),
    .B(_1586_),
    .C(_1587_));
 sg13g2_and2_1 _4493_ (.A(_1584_),
    .B(_1587_),
    .X(_1588_));
 sg13g2_nand2_1 _4494_ (.Y(_1589_),
    .A(net550),
    .B(_1537_));
 sg13g2_a21oi_1 _4495_ (.A1(_1582_),
    .A2(_1589_),
    .Y(_1590_),
    .B1(\top.c_y[9] ));
 sg13g2_and3_1 _4496_ (.X(_1591_),
    .A(\top.c_y[9] ),
    .B(_1582_),
    .C(_1589_));
 sg13g2_nor2_1 _4497_ (.A(_1590_),
    .B(_1591_),
    .Y(_1592_));
 sg13g2_a21oi_1 _4498_ (.A1(_1588_),
    .A2(_1592_),
    .Y(_1593_),
    .B1(net574));
 sg13g2_o21ai_1 _4499_ (.B1(_1593_),
    .Y(_0239_),
    .A1(_1588_),
    .A2(_1592_));
 sg13g2_o21ai_1 _4500_ (.B1(net550),
    .Y(_1594_),
    .A1(net552),
    .A2(_1544_));
 sg13g2_and2_1 _4501_ (.A(_1582_),
    .B(_1594_),
    .X(_1595_));
 sg13g2_nand2_1 _4502_ (.Y(_1596_),
    .A(\top.c_y[10] ),
    .B(_1595_));
 sg13g2_xor2_1 _4503_ (.B(_1595_),
    .A(\top.c_y[10] ),
    .X(_1597_));
 sg13g2_a21oi_1 _4504_ (.A1(_1584_),
    .A2(_1587_),
    .Y(_1598_),
    .B1(_1590_));
 sg13g2_nor3_1 _4505_ (.A(_1591_),
    .B(_1597_),
    .C(_1598_),
    .Y(_1599_));
 sg13g2_o21ai_1 _4506_ (.B1(_1597_),
    .Y(_1600_),
    .A1(_1591_),
    .A2(_1598_));
 sg13g2_nand2_1 _4507_ (.Y(_1601_),
    .A(net579),
    .B(_1600_));
 sg13g2_nor2_1 _4508_ (.A(_1599_),
    .B(_1601_),
    .Y(_0240_));
 sg13g2_and2_1 _4509_ (.A(_1596_),
    .B(_1600_),
    .X(_1602_));
 sg13g2_a21oi_1 _4510_ (.A1(net550),
    .A2(_1550_),
    .Y(_1603_),
    .B1(_1581_));
 sg13g2_xnor2_1 _4511_ (.Y(_1604_),
    .A(net863),
    .B(_1603_));
 sg13g2_o21ai_1 _4512_ (.B1(net579),
    .Y(_1605_),
    .A1(_1602_),
    .A2(_1604_));
 sg13g2_a21oi_1 _4513_ (.A1(_1602_),
    .A2(_1604_),
    .Y(_0241_),
    .B1(_1605_));
 sg13g2_a21oi_1 _4514_ (.A1(\top.debouncer_inst.last_data[2] ),
    .A2(net7),
    .Y(_1606_),
    .B1(\top.last_stable_buttons[2] ));
 sg13g2_a21oi_1 _4515_ (.A1(\top.debouncer_inst.last_data[2] ),
    .A2(\top.last_stable_buttons[2] ),
    .Y(_1607_),
    .B1(_0024_));
 sg13g2_nor2b_1 _4516_ (.A(_1606_),
    .B_N(_1607_),
    .Y(_1608_));
 sg13g2_nor2b_1 _4517_ (.A(\top.last_stable_buttons[3] ),
    .B_N(\top.debouncer_inst.last_data[3] ),
    .Y(_1609_));
 sg13g2_nor2b_1 _4518_ (.A(\top.debouncer_inst.last_data[3] ),
    .B_N(\top.last_stable_buttons[3] ),
    .Y(_1610_));
 sg13g2_a22oi_1 _4519_ (.Y(_1611_),
    .B1(_1610_),
    .B2(\top.buttons_stable ),
    .A2(_1609_),
    .A1(_1489_));
 sg13g2_and2_1 _4520_ (.A(_1608_),
    .B(_1611_),
    .X(_1612_));
 sg13g2_xor2_1 _4521_ (.B(_1611_),
    .A(_1608_),
    .X(_1613_));
 sg13g2_or3_1 _4522_ (.A(net555),
    .B(net553),
    .C(_1613_),
    .X(_1614_));
 sg13g2_nor4_2 _4523_ (.A(net555),
    .B(net553),
    .C(net551),
    .Y(_1615_),
    .D(_1613_));
 sg13g2_and3_1 _4524_ (.X(_1616_),
    .A(net824),
    .B(net547),
    .C(_1615_));
 sg13g2_a21oi_1 _4525_ (.A1(net547),
    .A2(_1615_),
    .Y(_1617_),
    .B1(net824));
 sg13g2_o21ai_1 _4526_ (.B1(net581),
    .Y(_0242_),
    .A1(_1616_),
    .A2(net825));
 sg13g2_a21oi_1 _4527_ (.A1(_1608_),
    .A2(_1611_),
    .Y(_1618_),
    .B1(net555));
 sg13g2_or2_1 _4528_ (.X(_1619_),
    .B(_1618_),
    .A(_1613_));
 sg13g2_nor4_2 _4529_ (.A(net553),
    .B(net551),
    .C(_1613_),
    .Y(_1620_),
    .D(_1618_));
 sg13g2_and3_1 _4530_ (.X(_1621_),
    .A(\top.c_x[1] ),
    .B(net547),
    .C(_1620_));
 sg13g2_nand3_1 _4531_ (.B(net547),
    .C(_1620_),
    .A(net876),
    .Y(_1622_));
 sg13g2_a21o_1 _4532_ (.A2(_1620_),
    .A1(net547),
    .B1(\top.c_x[1] ),
    .X(_1623_));
 sg13g2_a21oi_1 _4533_ (.A1(_1622_),
    .A2(_1623_),
    .Y(_1624_),
    .B1(_1616_));
 sg13g2_and3_1 _4534_ (.X(_1625_),
    .A(_1616_),
    .B(_1622_),
    .C(_1623_));
 sg13g2_nor3_1 _4535_ (.A(net574),
    .B(_1624_),
    .C(_1625_),
    .Y(_0243_));
 sg13g2_nor2_1 _4536_ (.A(net553),
    .B(_1612_),
    .Y(_1626_));
 sg13g2_or2_1 _4537_ (.X(_1627_),
    .B(_1612_),
    .A(net553));
 sg13g2_o21ai_1 _4538_ (.B1(net553),
    .Y(_1628_),
    .A1(net555),
    .A2(_1613_));
 sg13g2_nand3_1 _4539_ (.B(_1627_),
    .C(_1628_),
    .A(net521),
    .Y(_1629_));
 sg13g2_and4_1 _4540_ (.A(net521),
    .B(net547),
    .C(_1627_),
    .D(_1628_),
    .X(_1630_));
 sg13g2_nand2_1 _4541_ (.Y(_1631_),
    .A(\top.c_x[2] ),
    .B(_1630_));
 sg13g2_xnor2_1 _4542_ (.Y(_1632_),
    .A(net875),
    .B(_1630_));
 sg13g2_a21oi_1 _4543_ (.A1(_1616_),
    .A2(_1623_),
    .Y(_1633_),
    .B1(_1621_));
 sg13g2_o21ai_1 _4544_ (.B1(net581),
    .Y(_1634_),
    .A1(_1632_),
    .A2(_1633_));
 sg13g2_a21oi_1 _4545_ (.A1(_1632_),
    .A2(_1633_),
    .Y(_0244_),
    .B1(_1634_));
 sg13g2_nor2_2 _4546_ (.A(_1619_),
    .B(_1626_),
    .Y(_1635_));
 sg13g2_inv_1 _4547_ (.Y(_1636_),
    .A(_1635_));
 sg13g2_nand3_1 _4548_ (.B(net547),
    .C(_1635_),
    .A(net521),
    .Y(_1637_));
 sg13g2_nor2_1 _4549_ (.A(net869),
    .B(_1637_),
    .Y(_1638_));
 sg13g2_xor2_1 _4550_ (.B(_1637_),
    .A(net869),
    .X(_1639_));
 sg13g2_o21ai_1 _4551_ (.B1(_1631_),
    .Y(_1640_),
    .A1(_1632_),
    .A2(_1633_));
 sg13g2_xnor2_1 _4552_ (.Y(_1641_),
    .A(_1639_),
    .B(_1640_));
 sg13g2_nand2_1 _4553_ (.Y(_0245_),
    .A(net582),
    .B(_1641_));
 sg13g2_o21ai_1 _4554_ (.B1(net547),
    .Y(_1642_),
    .A1(net551),
    .A2(_1612_));
 sg13g2_inv_1 _4555_ (.Y(_1643_),
    .A(_1642_));
 sg13g2_a21oi_1 _4556_ (.A1(net551),
    .A2(_1614_),
    .Y(_1644_),
    .B1(_1642_));
 sg13g2_nand2_1 _4557_ (.Y(_1645_),
    .A(\top.c_x[4] ),
    .B(_1644_));
 sg13g2_xnor2_1 _4558_ (.Y(_1646_),
    .A(\top.c_x[4] ),
    .B(_1644_));
 sg13g2_a21oi_1 _4559_ (.A1(_1639_),
    .A2(_1640_),
    .Y(_1647_),
    .B1(_1638_));
 sg13g2_xnor2_1 _4560_ (.Y(_1648_),
    .A(_1646_),
    .B(_1647_));
 sg13g2_nand2_1 _4561_ (.Y(_0246_),
    .A(net582),
    .B(_1648_));
 sg13g2_o21ai_1 _4562_ (.B1(_1645_),
    .Y(_1649_),
    .A1(_1646_),
    .A2(_1647_));
 sg13g2_o21ai_1 _4563_ (.B1(net551),
    .Y(_1650_),
    .A1(net553),
    .A2(_1619_));
 sg13g2_and2_1 _4564_ (.A(_1643_),
    .B(_1650_),
    .X(_1651_));
 sg13g2_nor2b_1 _4565_ (.A(net883),
    .B_N(_1651_),
    .Y(_1652_));
 sg13g2_xnor2_1 _4566_ (.Y(_1653_),
    .A(net841),
    .B(_1651_));
 sg13g2_o21ai_1 _4567_ (.B1(net582),
    .Y(_1654_),
    .A1(_1649_),
    .A2(_1653_));
 sg13g2_a21oi_1 _4568_ (.A1(_1649_),
    .A2(_1653_),
    .Y(_0247_),
    .B1(_1654_));
 sg13g2_a21o_1 _4569_ (.A2(_1653_),
    .A1(_1649_),
    .B1(_1652_),
    .X(_1655_));
 sg13g2_a21oi_1 _4570_ (.A1(_1627_),
    .A2(_1628_),
    .Y(_1656_),
    .B1(net521));
 sg13g2_nor2_1 _4571_ (.A(_1642_),
    .B(_1656_),
    .Y(_1657_));
 sg13g2_nand2_1 _4572_ (.Y(_1658_),
    .A(\top.c_x[6] ),
    .B(_1657_));
 sg13g2_xnor2_1 _4573_ (.Y(_1659_),
    .A(\top.c_x[6] ),
    .B(_1657_));
 sg13g2_nand2b_1 _4574_ (.Y(_1660_),
    .B(_1659_),
    .A_N(_1655_));
 sg13g2_nand2b_1 _4575_ (.Y(_1661_),
    .B(_1655_),
    .A_N(_1659_));
 sg13g2_and3_1 _4576_ (.X(_0248_),
    .A(net582),
    .B(_1660_),
    .C(_1661_));
 sg13g2_nand2_1 _4577_ (.Y(_1662_),
    .A(_1658_),
    .B(_1661_));
 sg13g2_inv_1 _4578_ (.Y(_1663_),
    .A(_1662_));
 sg13g2_nand3_1 _4579_ (.B(_1635_),
    .C(_1643_),
    .A(\top.c_x[7] ),
    .Y(_1664_));
 sg13g2_a21o_1 _4580_ (.A2(_1643_),
    .A1(_1635_),
    .B1(\top.c_x[7] ),
    .X(_1665_));
 sg13g2_nand2_1 _4581_ (.Y(_1666_),
    .A(_1664_),
    .B(_1665_));
 sg13g2_xor2_1 _4582_ (.B(_1666_),
    .A(_1662_),
    .X(_1667_));
 sg13g2_nand2_1 _4583_ (.Y(_0249_),
    .A(net582),
    .B(_1667_));
 sg13g2_o21ai_1 _4584_ (.B1(_1664_),
    .Y(_1668_),
    .A1(_1663_),
    .A2(_1666_));
 sg13g2_nor2_1 _4585_ (.A(net549),
    .B(_1612_),
    .Y(_1669_));
 sg13g2_or2_1 _4586_ (.X(_1670_),
    .B(_1612_),
    .A(net549));
 sg13g2_nor2b_1 _4587_ (.A(_1615_),
    .B_N(net549),
    .Y(_1671_));
 sg13g2_nor2_1 _4588_ (.A(_1669_),
    .B(_1671_),
    .Y(_1672_));
 sg13g2_nand2_1 _4589_ (.Y(_1673_),
    .A(\top.c_x[8] ),
    .B(_1672_));
 sg13g2_xnor2_1 _4590_ (.Y(_1674_),
    .A(net882),
    .B(_1672_));
 sg13g2_nand2b_1 _4591_ (.Y(_1675_),
    .B(_1674_),
    .A_N(_1668_));
 sg13g2_nand2b_1 _4592_ (.Y(_1676_),
    .B(_1668_),
    .A_N(_1674_));
 sg13g2_and3_1 _4593_ (.X(_0250_),
    .A(net582),
    .B(_1675_),
    .C(_1676_));
 sg13g2_nand2_1 _4594_ (.Y(_1677_),
    .A(_1673_),
    .B(_1676_));
 sg13g2_nand2b_1 _4595_ (.Y(_1678_),
    .B(net549),
    .A_N(_1620_));
 sg13g2_a21oi_1 _4596_ (.A1(_1670_),
    .A2(_1678_),
    .Y(_1679_),
    .B1(net878));
 sg13g2_nand3_1 _4597_ (.B(_1670_),
    .C(_1678_),
    .A(\top.c_x[9] ),
    .Y(_1680_));
 sg13g2_nand2b_1 _4598_ (.Y(_1681_),
    .B(_1680_),
    .A_N(_1679_));
 sg13g2_a21oi_1 _4599_ (.A1(_1677_),
    .A2(_1681_),
    .Y(_1682_),
    .B1(net574));
 sg13g2_o21ai_1 _4600_ (.B1(_1682_),
    .Y(_0251_),
    .A1(_1677_),
    .A2(_1681_));
 sg13g2_a21oi_2 _4601_ (.B1(_1669_),
    .Y(_1683_),
    .A2(_1629_),
    .A1(net549));
 sg13g2_and2_1 _4602_ (.A(\top.c_x[10] ),
    .B(_1683_),
    .X(_1684_));
 sg13g2_xor2_1 _4603_ (.B(_1683_),
    .A(\top.c_x[10] ),
    .X(_1685_));
 sg13g2_nand3_1 _4604_ (.B(_1676_),
    .C(_1680_),
    .A(_1673_),
    .Y(_1686_));
 sg13g2_nor2b_1 _4605_ (.A(_1679_),
    .B_N(_1686_),
    .Y(_1687_));
 sg13g2_xnor2_1 _4606_ (.Y(_1688_),
    .A(_1685_),
    .B(_1687_));
 sg13g2_nand2_1 _4607_ (.Y(_0252_),
    .A(net580),
    .B(_1688_));
 sg13g2_a21o_1 _4608_ (.A2(_1687_),
    .A1(_1685_),
    .B1(_1684_),
    .X(_1689_));
 sg13g2_o21ai_1 _4609_ (.B1(net549),
    .Y(_1690_),
    .A1(net551),
    .A2(_1636_));
 sg13g2_nand2_1 _4610_ (.Y(_1691_),
    .A(_1670_),
    .B(_1690_));
 sg13g2_xor2_1 _4611_ (.B(_1691_),
    .A(net873),
    .X(_1692_));
 sg13g2_a21oi_1 _4612_ (.A1(_1689_),
    .A2(_1692_),
    .Y(_1693_),
    .B1(net574));
 sg13g2_o21ai_1 _4613_ (.B1(_1693_),
    .Y(_0253_),
    .A1(_1689_),
    .A2(_1692_));
 sg13g2_nor3_1 _4614_ (.A(\top.transmitter.transmitter.counter[0] ),
    .B(_1844_),
    .C(net836),
    .Y(_1694_));
 sg13g2_a22oi_1 _4615_ (.Y(_1695_),
    .B1(_1694_),
    .B2(net833),
    .A2(_1941_),
    .A1(_1890_));
 sg13g2_nand2b_1 _4616_ (.Y(_0254_),
    .B(_1695_),
    .A_N(net335));
 sg13g2_xnor2_1 _4617_ (.Y(_1696_),
    .A(\top.transmitter.transmitter.counter[0] ),
    .B(net817));
 sg13g2_nand2_1 _4618_ (.Y(_0255_),
    .A(_1942_),
    .B(net818));
 sg13g2_a21o_1 _4619_ (.A2(net817),
    .A1(\top.transmitter.transmitter.counter[0] ),
    .B1(net836),
    .X(_1697_));
 sg13g2_nand2_1 _4620_ (.Y(_1698_),
    .A(_1888_),
    .B(net837));
 sg13g2_nand2_1 _4621_ (.Y(_0256_),
    .A(_1695_),
    .B(net838));
 sg13g2_xor2_1 _4622_ (.B(_1888_),
    .A(net833),
    .X(_1699_));
 sg13g2_nand2_1 _4623_ (.Y(_0257_),
    .A(_1695_),
    .B(net834));
 sg13g2_or2_1 _4624_ (.X(_0258_),
    .B(net447),
    .A(net429));
 sg13g2_a21oi_2 _4625_ (.B1(_1459_),
    .Y(_1700_),
    .A2(_0321_),
    .A1(_1961_));
 sg13g2_mux2_1 _4626_ (.A0(net393),
    .A1(\top.receiver.data[0] ),
    .S(net458),
    .X(_0259_));
 sg13g2_mux2_1 _4627_ (.A0(net590),
    .A1(\top.receiver.data[1] ),
    .S(net458),
    .X(_0260_));
 sg13g2_mux2_1 _4628_ (.A0(net701),
    .A1(net322),
    .S(net458),
    .X(_0261_));
 sg13g2_mux2_1 _4629_ (.A0(net667),
    .A1(net323),
    .S(net458),
    .X(_0262_));
 sg13g2_mux2_1 _4630_ (.A0(net697),
    .A1(net329),
    .S(net458),
    .X(_0263_));
 sg13g2_mux2_1 _4631_ (.A0(net589),
    .A1(net333),
    .S(net457),
    .X(_0264_));
 sg13g2_mux2_1 _4632_ (.A0(net623),
    .A1(net332),
    .S(net457),
    .X(_0265_));
 sg13g2_mux2_1 _4633_ (.A0(net597),
    .A1(net326),
    .S(net457),
    .X(_0266_));
 sg13g2_mux2_1 _4634_ (.A0(net608),
    .A1(net331),
    .S(net457),
    .X(_0267_));
 sg13g2_mux2_1 _4635_ (.A0(net605),
    .A1(net337),
    .S(net457),
    .X(_0268_));
 sg13g2_mux2_1 _4636_ (.A0(net609),
    .A1(net324),
    .S(_1700_),
    .X(_0269_));
 sg13g2_mux2_1 _4637_ (.A0(net432),
    .A1(net334),
    .S(net458),
    .X(_0270_));
 sg13g2_mux2_1 _4638_ (.A0(net638),
    .A1(net325),
    .S(_1700_),
    .X(_0271_));
 sg13g2_mux2_1 _4639_ (.A0(net603),
    .A1(net327),
    .S(_1700_),
    .X(_0272_));
 sg13g2_nor2_1 _4640_ (.A(net634),
    .B(net458),
    .Y(_1701_));
 sg13g2_a21oi_1 _4641_ (.A1(_1845_),
    .A2(net457),
    .Y(_0273_),
    .B1(_1701_));
 sg13g2_nor2_1 _4642_ (.A(net431),
    .B(net457),
    .Y(_1702_));
 sg13g2_a21oi_1 _4643_ (.A1(_1851_),
    .A2(net457),
    .Y(_0274_),
    .B1(_1702_));
 sg13g2_nand2_1 _4644_ (.Y(_1703_),
    .A(net349),
    .B(net513));
 sg13g2_xor2_1 _4645_ (.B(_2112_),
    .A(_2111_),
    .X(_1704_));
 sg13g2_a21oi_1 _4646_ (.A1(net568),
    .A2(_1831_),
    .Y(_1705_),
    .B1(net512));
 sg13g2_o21ai_1 _4647_ (.B1(_1705_),
    .Y(_1706_),
    .A1(net567),
    .A2(_1704_));
 sg13g2_nand2_1 _4648_ (.Y(_0275_),
    .A(_1703_),
    .B(_1706_));
 sg13g2_nand2_1 _4649_ (.Y(_1707_),
    .A(net343),
    .B(net513));
 sg13g2_nand3_1 _4650_ (.B(_2113_),
    .C(_2114_),
    .A(_2097_),
    .Y(_1708_));
 sg13g2_and2_1 _4651_ (.A(_2115_),
    .B(_1708_),
    .X(_1709_));
 sg13g2_nand2b_1 _4652_ (.Y(_1710_),
    .B(net567),
    .A_N(\top.julia_calc.dest_x[1] ));
 sg13g2_o21ai_1 _4653_ (.B1(_1710_),
    .Y(_1711_),
    .A1(net567),
    .A2(_1709_));
 sg13g2_o21ai_1 _4654_ (.B1(_1707_),
    .Y(_0276_),
    .A1(net514),
    .A2(_1711_));
 sg13g2_nand3_1 _4655_ (.B(_2115_),
    .C(_2117_),
    .A(_2092_),
    .Y(_1712_));
 sg13g2_a21oi_1 _4656_ (.A1(_2119_),
    .A2(_1712_),
    .Y(_1713_),
    .B1(net567));
 sg13g2_nor2_1 _4657_ (.A(net523),
    .B(\top.julia_calc.dest_x[2] ),
    .Y(_1714_));
 sg13g2_nor3_1 _4658_ (.A(net514),
    .B(_1713_),
    .C(_1714_),
    .Y(_1715_));
 sg13g2_a21o_1 _4659_ (.A2(net514),
    .A1(net391),
    .B1(_1715_),
    .X(_0277_));
 sg13g2_nand2_1 _4660_ (.Y(_1716_),
    .A(net354),
    .B(net511));
 sg13g2_xnor2_1 _4661_ (.Y(_1717_),
    .A(_2120_),
    .B(_2121_));
 sg13g2_nand2_1 _4662_ (.Y(_1718_),
    .A(net522),
    .B(_1717_));
 sg13g2_o21ai_1 _4663_ (.B1(_1718_),
    .Y(_1719_),
    .A1(net522),
    .A2(\top.julia_calc.dest_x[3] ));
 sg13g2_o21ai_1 _4664_ (.B1(_1716_),
    .Y(_0278_),
    .A1(net511),
    .A2(_1719_));
 sg13g2_nand2_1 _4665_ (.Y(_1720_),
    .A(net345),
    .B(net511));
 sg13g2_nand3_1 _4666_ (.B(_2122_),
    .C(_2124_),
    .A(_2082_),
    .Y(_1721_));
 sg13g2_nor2b_1 _4667_ (.A(_2125_),
    .B_N(_1721_),
    .Y(_1722_));
 sg13g2_nand2b_1 _4668_ (.Y(_1723_),
    .B(net568),
    .A_N(\top.julia_calc.dest_x[4] ));
 sg13g2_o21ai_1 _4669_ (.B1(_1723_),
    .Y(_1724_),
    .A1(net568),
    .A2(_1722_));
 sg13g2_o21ai_1 _4670_ (.B1(_1720_),
    .Y(_0279_),
    .A1(net511),
    .A2(_1724_));
 sg13g2_nand2_1 _4671_ (.Y(_1725_),
    .A(net341),
    .B(net512));
 sg13g2_xnor2_1 _4672_ (.Y(_1726_),
    .A(_2126_),
    .B(_2127_));
 sg13g2_a21oi_1 _4673_ (.A1(net568),
    .A2(_1850_),
    .Y(_1727_),
    .B1(net511));
 sg13g2_o21ai_1 _4674_ (.B1(_1727_),
    .Y(_1728_),
    .A1(net567),
    .A2(_1726_));
 sg13g2_nand2_1 _4675_ (.Y(_0280_),
    .A(_1725_),
    .B(_1728_));
 sg13g2_nand3_1 _4676_ (.B(_2128_),
    .C(_2129_),
    .A(_2071_),
    .Y(_1729_));
 sg13g2_nor2_1 _4677_ (.A(net567),
    .B(_2130_),
    .Y(_1730_));
 sg13g2_nand2_1 _4678_ (.Y(_1731_),
    .A(_1729_),
    .B(_1730_));
 sg13g2_xnor2_1 _4679_ (.Y(_1732_),
    .A(\top.julia_calc.dest_x[6] ),
    .B(\top.julia_calc.dest_x[5] ));
 sg13g2_a21oi_1 _4680_ (.A1(net568),
    .A2(_1732_),
    .Y(_1733_),
    .B1(net512));
 sg13g2_a22oi_1 _4681_ (.Y(_0281_),
    .B1(_1731_),
    .B2(_1733_),
    .A2(net512),
    .A1(_1863_));
 sg13g2_or3_1 _4682_ (.A(_2067_),
    .B(_2130_),
    .C(_2131_),
    .X(_1734_));
 sg13g2_and2_1 _4683_ (.A(net522),
    .B(_2132_),
    .X(_1735_));
 sg13g2_o21ai_1 _4684_ (.B1(\top.julia_calc.dest_x[7] ),
    .Y(_1736_),
    .A1(\top.julia_calc.dest_x[6] ),
    .A2(\top.julia_calc.dest_x[5] ));
 sg13g2_or3_1 _4685_ (.A(\top.julia_calc.dest_x[7] ),
    .B(\top.julia_calc.dest_x[6] ),
    .C(\top.julia_calc.dest_x[5] ),
    .X(_1737_));
 sg13g2_nand3_1 _4686_ (.B(_1736_),
    .C(_1737_),
    .A(net568),
    .Y(_1738_));
 sg13g2_a21oi_1 _4687_ (.A1(_1734_),
    .A2(_1735_),
    .Y(_1739_),
    .B1(net512));
 sg13g2_a22oi_1 _4688_ (.Y(_0282_),
    .B1(_1738_),
    .B2(_1739_),
    .A2(net512),
    .A1(_1859_));
 sg13g2_or2_1 _4689_ (.X(_1740_),
    .B(_1736_),
    .A(_0055_));
 sg13g2_a21oi_1 _4690_ (.A1(_0055_),
    .A2(_1736_),
    .Y(_1741_),
    .B1(net523));
 sg13g2_a221oi_1 _4691_ (.B2(_1741_),
    .C1(net511),
    .B1(_1740_),
    .A1(net523),
    .Y(_1742_),
    .A2(_2136_));
 sg13g2_a21o_1 _4692_ (.A2(net511),
    .A1(net419),
    .B1(_1742_),
    .X(_0283_));
 sg13g2_nand3_1 _4693_ (.B(_2153_),
    .C(_2154_),
    .A(_2151_),
    .Y(_1743_));
 sg13g2_nand3_1 _4694_ (.B(_2155_),
    .C(_1743_),
    .A(net522),
    .Y(_1744_));
 sg13g2_a21oi_1 _4695_ (.A1(\top.julia_calc.iter_done_reg ),
    .A2(\top.julia_calc.dest_y[0] ),
    .Y(_1745_),
    .B1(net511));
 sg13g2_a22oi_1 _4696_ (.Y(_0284_),
    .B1(_1744_),
    .B2(_1745_),
    .A2(net513),
    .A1(_1856_));
 sg13g2_nand3_1 _4697_ (.B(_2155_),
    .C(_2156_),
    .A(_2150_),
    .Y(_1746_));
 sg13g2_nand3_1 _4698_ (.B(_2157_),
    .C(_1746_),
    .A(net522),
    .Y(_1747_));
 sg13g2_a21oi_1 _4699_ (.A1(net566),
    .A2(\top.julia_calc.dest_y[1] ),
    .Y(_1748_),
    .B1(net510));
 sg13g2_a22oi_1 _4700_ (.Y(_0285_),
    .B1(_1747_),
    .B2(_1748_),
    .A2(net510),
    .A1(_1873_));
 sg13g2_and2_1 _4701_ (.A(net785),
    .B(net510),
    .X(_1749_));
 sg13g2_and3_1 _4702_ (.X(_1750_),
    .A(_2149_),
    .B(_2157_),
    .C(_2158_));
 sg13g2_o21ai_1 _4703_ (.B1(net522),
    .Y(_1751_),
    .A1(_2159_),
    .A2(_1750_));
 sg13g2_a21oi_1 _4704_ (.A1(net566),
    .A2(_1838_),
    .Y(_1752_),
    .B1(net510));
 sg13g2_a21o_1 _4705_ (.A2(_1752_),
    .A1(_1751_),
    .B1(_1749_),
    .X(_0286_));
 sg13g2_or3_1 _4706_ (.A(_2148_),
    .B(_2159_),
    .C(_2160_),
    .X(_1753_));
 sg13g2_a21o_1 _4707_ (.A2(_1753_),
    .A1(_2161_),
    .B1(net567),
    .X(_1754_));
 sg13g2_o21ai_1 _4708_ (.B1(_1754_),
    .Y(_1755_),
    .A1(net524),
    .A2(\top.julia_calc.dest_y[3] ));
 sg13g2_nand2_1 _4709_ (.Y(_1756_),
    .A(net351),
    .B(net509));
 sg13g2_o21ai_1 _4710_ (.B1(_1756_),
    .Y(_0287_),
    .A1(net509),
    .A2(_1755_));
 sg13g2_nand2_1 _4711_ (.Y(_1757_),
    .A(net376),
    .B(net508));
 sg13g2_and3_1 _4712_ (.X(_1758_),
    .A(_2147_),
    .B(_2161_),
    .C(_2162_));
 sg13g2_o21ai_1 _4713_ (.B1(net522),
    .Y(_1759_),
    .A1(_2163_),
    .A2(_1758_));
 sg13g2_nand2b_1 _4714_ (.Y(_1760_),
    .B(net566),
    .A_N(_0020_));
 sg13g2_nand4_1 _4715_ (.B(_2048_),
    .C(_1759_),
    .A(net577),
    .Y(_1761_),
    .D(_1760_));
 sg13g2_nand2_1 _4716_ (.Y(_0288_),
    .A(_1757_),
    .B(_1761_));
 sg13g2_nand2_1 _4717_ (.Y(_1762_),
    .A(net353),
    .B(net508));
 sg13g2_or3_1 _4718_ (.A(_2146_),
    .B(_2163_),
    .C(_2164_),
    .X(_1763_));
 sg13g2_and2_1 _4719_ (.A(_2165_),
    .B(_1763_),
    .X(_1764_));
 sg13g2_or2_1 _4720_ (.X(_1765_),
    .B(\top.julia_calc.dest_y[5] ),
    .A(\top.julia_calc.dest_y[4] ));
 sg13g2_nand2_1 _4721_ (.Y(_1766_),
    .A(\top.julia_calc.dest_y[4] ),
    .B(\top.julia_calc.dest_y[5] ));
 sg13g2_a21o_1 _4722_ (.A2(_1766_),
    .A1(_1765_),
    .B1(net524),
    .X(_1767_));
 sg13g2_o21ai_1 _4723_ (.B1(_1767_),
    .Y(_1768_),
    .A1(net566),
    .A2(_1764_));
 sg13g2_o21ai_1 _4724_ (.B1(_1762_),
    .Y(_0289_),
    .A1(net508),
    .A2(_1768_));
 sg13g2_nand3_1 _4725_ (.B(_2165_),
    .C(_2166_),
    .A(_2145_),
    .Y(_1769_));
 sg13g2_nand3_1 _4726_ (.B(_2167_),
    .C(_1769_),
    .A(net522),
    .Y(_1770_));
 sg13g2_nand3_1 _4727_ (.B(\top.julia_calc.dest_y[5] ),
    .C(\top.julia_calc.dest_y[6] ),
    .A(\top.julia_calc.dest_y[4] ),
    .Y(_1771_));
 sg13g2_a21oi_1 _4728_ (.A1(_1840_),
    .A2(_1766_),
    .Y(_1772_),
    .B1(net524));
 sg13g2_a21oi_1 _4729_ (.A1(_1771_),
    .A2(_1772_),
    .Y(_1773_),
    .B1(net508));
 sg13g2_a22oi_1 _4730_ (.Y(_0290_),
    .B1(_1770_),
    .B2(_1773_),
    .A2(net508),
    .A1(_1864_));
 sg13g2_nor2b_1 _4731_ (.A(_2143_),
    .B_N(_2144_),
    .Y(_1774_));
 sg13g2_xnor2_1 _4732_ (.Y(_1775_),
    .A(_2169_),
    .B(_1774_));
 sg13g2_nand2b_1 _4733_ (.Y(_1776_),
    .B(_1771_),
    .A_N(\top.julia_calc.dest_y[7] ));
 sg13g2_nand4_1 _4734_ (.B(\top.julia_calc.dest_y[5] ),
    .C(\top.julia_calc.dest_y[7] ),
    .A(\top.julia_calc.dest_y[4] ),
    .Y(_1777_),
    .D(\top.julia_calc.dest_y[6] ));
 sg13g2_nand3_1 _4735_ (.B(_1776_),
    .C(_1777_),
    .A(net566),
    .Y(_1778_));
 sg13g2_a21oi_1 _4736_ (.A1(net524),
    .A2(_1775_),
    .Y(_1779_),
    .B1(net509));
 sg13g2_a22oi_1 _4737_ (.Y(_0291_),
    .B1(_1778_),
    .B2(_1779_),
    .A2(net508),
    .A1(_1860_));
 sg13g2_nor2b_1 _4738_ (.A(_2141_),
    .B_N(_2142_),
    .Y(_1780_));
 sg13g2_o21ai_1 _4739_ (.B1(net523),
    .Y(_1781_),
    .A1(_2170_),
    .A2(_1780_));
 sg13g2_a21oi_2 _4740_ (.B1(_1781_),
    .Y(_1782_),
    .A2(_1780_),
    .A1(_2170_));
 sg13g2_o21ai_1 _4741_ (.B1(net566),
    .Y(_1783_),
    .A1(_0057_),
    .A2(_1777_));
 sg13g2_a21oi_1 _4742_ (.A1(_0057_),
    .A2(_1777_),
    .Y(_1784_),
    .B1(_1783_));
 sg13g2_nor3_1 _4743_ (.A(net508),
    .B(_1782_),
    .C(_1784_),
    .Y(_1785_));
 sg13g2_a21o_1 _4744_ (.A2(net508),
    .A1(net416),
    .B1(_1785_),
    .X(_0292_));
 sg13g2_nor2_1 _4745_ (.A(net779),
    .B(_2030_),
    .Y(_1786_));
 sg13g2_and2_1 _4746_ (.A(net779),
    .B(_2030_),
    .X(_1787_));
 sg13g2_nor3_1 _4747_ (.A(net573),
    .B(net780),
    .C(_1787_),
    .Y(_0295_));
 sg13g2_and2_1 _4748_ (.A(net796),
    .B(_1787_),
    .X(_1788_));
 sg13g2_o21ai_1 _4749_ (.B1(net577),
    .Y(_1789_),
    .A1(net796),
    .A2(_1787_));
 sg13g2_nor2_1 _4750_ (.A(_1788_),
    .B(net797),
    .Y(_0296_));
 sg13g2_nor3_1 _4751_ (.A(_1839_),
    .B(\top.julia_calc.dest_y[5] ),
    .C(_0057_),
    .Y(_1790_));
 sg13g2_nand3_1 _4752_ (.B(\top.julia_calc.dest_y[6] ),
    .C(_1790_),
    .A(\top.julia_calc.dest_y[7] ),
    .Y(_1791_));
 sg13g2_and2_1 _4753_ (.A(net698),
    .B(_1788_),
    .X(_1792_));
 sg13g2_nand2_1 _4754_ (.Y(_1793_),
    .A(net868),
    .B(_1792_));
 sg13g2_nand3_1 _4755_ (.B(net698),
    .C(_1788_),
    .A(net868),
    .Y(_1794_));
 sg13g2_o21ai_1 _4756_ (.B1(net577),
    .Y(_1795_),
    .A1(_1791_),
    .A2(_1794_));
 sg13g2_nor2_1 _4757_ (.A(net698),
    .B(_1788_),
    .Y(_1796_));
 sg13g2_nor3_1 _4758_ (.A(net573),
    .B(_1792_),
    .C(net699),
    .Y(_0297_));
 sg13g2_or2_1 _4759_ (.X(_1797_),
    .B(_1792_),
    .A(net868));
 sg13g2_and3_1 _4760_ (.X(_0298_),
    .A(net577),
    .B(_1793_),
    .C(_1797_));
 sg13g2_xnor2_1 _4761_ (.Y(_1798_),
    .A(_1839_),
    .B(_1794_));
 sg13g2_nor2_1 _4762_ (.A(_1795_),
    .B(_1798_),
    .Y(_0299_));
 sg13g2_nor2_1 _4763_ (.A(net789),
    .B(_1794_),
    .Y(_1799_));
 sg13g2_xnor2_1 _4764_ (.Y(_1800_),
    .A(\top.julia_calc.dest_y[5] ),
    .B(_1799_));
 sg13g2_nor2_1 _4765_ (.A(_1795_),
    .B(net790),
    .Y(_0300_));
 sg13g2_nor2_1 _4766_ (.A(_1766_),
    .B(_1793_),
    .Y(_1801_));
 sg13g2_xnor2_1 _4767_ (.Y(_1802_),
    .A(net831),
    .B(_1801_));
 sg13g2_nor2_1 _4768_ (.A(_1795_),
    .B(net832),
    .Y(_0301_));
 sg13g2_a21oi_1 _4769_ (.A1(\top.julia_calc.dest_y[6] ),
    .A2(_1801_),
    .Y(_1803_),
    .B1(net749));
 sg13g2_nor2_1 _4770_ (.A(_1777_),
    .B(_1794_),
    .Y(_1804_));
 sg13g2_nor3_1 _4771_ (.A(_1795_),
    .B(net750),
    .C(_1804_),
    .Y(_0302_));
 sg13g2_xnor2_1 _4772_ (.Y(_1805_),
    .A(net624),
    .B(_1804_));
 sg13g2_nor2_1 _4773_ (.A(_1795_),
    .B(_1805_),
    .Y(_0303_));
 sg13g2_nor4_1 _4774_ (.A(\top.next_read_addr[11] ),
    .B(\top.next_read_addr[10] ),
    .C(\top.next_read_addr[7] ),
    .D(\top.next_read_addr[6] ),
    .Y(_1806_));
 sg13g2_nor4_1 _4775_ (.A(\top.next_read_addr[14] ),
    .B(_1843_),
    .C(\top.next_read_addr[13] ),
    .D(\top.next_read_addr[12] ),
    .Y(_1807_));
 sg13g2_nand4_1 _4776_ (.B(\top.next_read_addr[8] ),
    .C(_1806_),
    .A(\top.next_read_addr[9] ),
    .Y(_1808_),
    .D(_1807_));
 sg13g2_a21oi_2 _4777_ (.B1(net451),
    .Y(_1809_),
    .A2(_1808_),
    .A1(net578));
 sg13g2_nor2_1 _4778_ (.A(net815),
    .B(_1468_),
    .Y(_1810_));
 sg13g2_and2_1 _4779_ (.A(net815),
    .B(_1468_),
    .X(_1811_));
 sg13g2_nor3_1 _4780_ (.A(net448),
    .B(net816),
    .C(_1811_),
    .Y(_0304_));
 sg13g2_nor2_1 _4781_ (.A(net826),
    .B(_1811_),
    .Y(_1812_));
 sg13g2_nand2_1 _4782_ (.Y(_1813_),
    .A(net826),
    .B(_1811_));
 sg13g2_inv_1 _4783_ (.Y(_1814_),
    .A(_1813_));
 sg13g2_nor3_1 _4784_ (.A(net448),
    .B(_1812_),
    .C(_1814_),
    .Y(_0305_));
 sg13g2_nor2_1 _4785_ (.A(net821),
    .B(_1814_),
    .Y(_1815_));
 sg13g2_and4_1 _4786_ (.A(\top.next_read_addr[8] ),
    .B(\top.next_read_addr[7] ),
    .C(\top.next_read_addr[6] ),
    .D(_1467_),
    .X(_1816_));
 sg13g2_nor3_1 _4787_ (.A(_1809_),
    .B(net822),
    .C(_1816_),
    .Y(_0306_));
 sg13g2_nor2_1 _4788_ (.A(net819),
    .B(_1816_),
    .Y(_1817_));
 sg13g2_and3_1 _4789_ (.X(_1818_),
    .A(net819),
    .B(net885),
    .C(_1814_));
 sg13g2_nor3_1 _4790_ (.A(net448),
    .B(net820),
    .C(_1818_),
    .Y(_0307_));
 sg13g2_nor2_1 _4791_ (.A(net812),
    .B(_1818_),
    .Y(_1819_));
 sg13g2_and2_1 _4792_ (.A(net812),
    .B(_1818_),
    .X(_1820_));
 sg13g2_nor3_1 _4793_ (.A(net448),
    .B(net813),
    .C(_1820_),
    .Y(_0308_));
 sg13g2_nor2_1 _4794_ (.A(net810),
    .B(_1820_),
    .Y(_1821_));
 sg13g2_and4_1 _4795_ (.A(net810),
    .B(\top.next_read_addr[10] ),
    .C(\top.next_read_addr[9] ),
    .D(_1816_),
    .X(_1822_));
 sg13g2_nor3_1 _4796_ (.A(net448),
    .B(net811),
    .C(_1822_),
    .Y(_0309_));
 sg13g2_xnor2_1 _4797_ (.Y(_1823_),
    .A(net829),
    .B(_1822_));
 sg13g2_nor2_1 _4798_ (.A(net448),
    .B(net830),
    .Y(_0310_));
 sg13g2_a21oi_1 _4799_ (.A1(\top.next_read_addr[12] ),
    .A2(_1822_),
    .Y(_1824_),
    .B1(net720));
 sg13g2_and2_1 _4800_ (.A(_1891_),
    .B(_1820_),
    .X(_1825_));
 sg13g2_nor3_1 _4801_ (.A(net448),
    .B(net721),
    .C(_1825_),
    .Y(_0311_));
 sg13g2_nand2_1 _4802_ (.Y(_1826_),
    .A(net783),
    .B(_1825_));
 sg13g2_xnor2_1 _4803_ (.Y(_1827_),
    .A(net783),
    .B(_1825_));
 sg13g2_nor2_1 _4804_ (.A(net448),
    .B(_1827_),
    .Y(_0312_));
 sg13g2_xnor2_1 _4805_ (.Y(_1828_),
    .A(_1843_),
    .B(_1826_));
 sg13g2_nor2_1 _4806_ (.A(_1809_),
    .B(_1828_),
    .Y(_0313_));
 sg13g2_a21oi_1 _4807_ (.A1(_1833_),
    .A2(_0315_),
    .Y(_0293_),
    .B1(_0368_));
 sg13g2_inv_1 _4808_ (.Y(_1829_),
    .A(net566));
 sg13g2_inv_2 _4809_ (.Y(_1830_),
    .A(net564));
 sg13g2_inv_1 _4810_ (.Y(_1831_),
    .A(\top.julia_calc.dest_x[0] ));
 sg13g2_inv_1 _4811_ (.Y(_1832_),
    .A(\top.pixel_buffer[7][1] ));
 sg13g2_inv_1 _4812_ (.Y(_1833_),
    .A(net590));
 sg13g2_inv_1 _4813_ (.Y(_1834_),
    .A(\top.pixel_buffer[7][0] ));
 sg13g2_inv_1 _4814_ (.Y(_1835_),
    .A(net572));
 sg13g2_inv_1 _4815_ (.Y(_1836_),
    .A(net583));
 sg13g2_inv_1 _4816_ (.Y(_1837_),
    .A(\top.julia_calc.z_y2[11] ));
 sg13g2_inv_1 _4817_ (.Y(_1838_),
    .A(net698));
 sg13g2_inv_1 _4818_ (.Y(_1839_),
    .A(net877));
 sg13g2_inv_1 _4819_ (.Y(_1840_),
    .A(\top.julia_calc.dest_y[6] ));
 sg13g2_inv_1 _4820_ (.Y(_1841_),
    .A(net850));
 sg13g2_inv_1 _4821_ (.Y(_1842_),
    .A(net880));
 sg13g2_inv_1 _4822_ (.Y(_1843_),
    .A(net809));
 sg13g2_inv_1 _4823_ (.Y(_1844_),
    .A(net817));
 sg13g2_inv_1 _4824_ (.Y(_1845_),
    .A(net330));
 sg13g2_inv_1 _4825_ (.Y(_1846_),
    .A(\top.debouncer_inst.last_data[0] ));
 sg13g2_inv_1 _4826_ (.Y(_1847_),
    .A(\top.debouncer_inst.last_data[2] ));
 sg13g2_inv_1 _4827_ (.Y(_1848_),
    .A(\top.c_y[2] ));
 sg13g2_inv_1 _4828_ (.Y(_1849_),
    .A(\top.c_y[1] ));
 sg13g2_inv_1 _4829_ (.Y(_1850_),
    .A(_0021_));
 sg13g2_inv_1 _4830_ (.Y(_1851_),
    .A(net321));
 sg13g2_inv_1 _4831_ (.Y(_1852_),
    .A(net555));
 sg13g2_inv_1 _4832_ (.Y(_1853_),
    .A(net554));
 sg13g2_inv_1 _4833_ (.Y(_1854_),
    .A(net552));
 sg13g2_inv_1 _4834_ (.Y(_1855_),
    .A(net548));
 sg13g2_inv_1 _4835_ (.Y(_1856_),
    .A(net389));
 sg13g2_inv_1 _4836_ (.Y(_1857_),
    .A(_0033_));
 sg13g2_inv_1 _4837_ (.Y(_1858_),
    .A(_0032_));
 sg13g2_inv_1 _4838_ (.Y(_1859_),
    .A(net435));
 sg13g2_inv_1 _4839_ (.Y(_1860_),
    .A(net437));
 sg13g2_inv_1 _4840_ (.Y(_1861_),
    .A(_0039_));
 sg13g2_inv_1 _4841_ (.Y(_1862_),
    .A(_0038_));
 sg13g2_inv_1 _4842_ (.Y(_1863_),
    .A(net601));
 sg13g2_inv_1 _4843_ (.Y(_1864_),
    .A(net421));
 sg13g2_inv_1 _4844_ (.Y(_1865_),
    .A(_0041_));
 sg13g2_inv_1 _4845_ (.Y(_1866_),
    .A(_0040_));
 sg13g2_inv_1 _4846_ (.Y(_1867_),
    .A(_0043_));
 sg13g2_inv_1 _4847_ (.Y(_1868_),
    .A(_0042_));
 sg13g2_inv_1 _4848_ (.Y(_1869_),
    .A(_0045_));
 sg13g2_inv_1 _4849_ (.Y(_1870_),
    .A(_0044_));
 sg13g2_inv_1 _4850_ (.Y(_1871_),
    .A(_0047_));
 sg13g2_inv_1 _4851_ (.Y(_1872_),
    .A(_0046_));
 sg13g2_inv_1 _4852_ (.Y(_1873_),
    .A(net405));
 sg13g2_inv_1 _4853_ (.Y(_1874_),
    .A(_0051_));
 sg13g2_inv_1 _4854_ (.Y(_1875_),
    .A(_0050_));
 sg13g2_inv_1 _4855_ (.Y(_1876_),
    .A(_0053_));
 sg13g2_inv_1 _4856_ (.Y(_1877_),
    .A(_0052_));
 sg13g2_nor2_2 _4857_ (.A(net559),
    .B(net560),
    .Y(_1878_));
 sg13g2_nor2_1 _4858_ (.A(\top.early_x[0] ),
    .B(net761),
    .Y(_1879_));
 sg13g2_and2_2 _4859_ (.A(_1878_),
    .B(_1879_),
    .X(_1880_));
 sg13g2_dfrbp_1 _4860_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net33),
    .D(_0064_),
    .Q_N(_2381_),
    .Q(\top.julia_calc.phase[0] ));
 sg13g2_dfrbp_1 _4861_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net119),
    .D(net854),
    .Q_N(_2380_),
    .Q(\top.julia_calc.phase[1] ));
 sg13g2_dfrbp_1 _4862_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net118),
    .D(net339),
    .Q_N(_0063_),
    .Q(\top.julia_calc.dest_x[0] ));
 sg13g2_dfrbp_1 _4863_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net116),
    .D(net845),
    .Q_N(_2379_),
    .Q(\top.julia_calc.dest_x[1] ));
 sg13g2_dfrbp_1 _4864_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net114),
    .D(_0068_),
    .Q_N(_2378_),
    .Q(\top.julia_calc.dest_x[2] ));
 sg13g2_dfrbp_1 _4865_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net112),
    .D(_0069_),
    .Q_N(_2377_),
    .Q(\top.julia_calc.dest_x[3] ));
 sg13g2_dfrbp_1 _4866_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net110),
    .D(_0070_),
    .Q_N(_2376_),
    .Q(\top.julia_calc.dest_x[4] ));
 sg13g2_dfrbp_1 _4867_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net108),
    .D(_0071_),
    .Q_N(_0021_),
    .Q(\top.julia_calc.dest_x[5] ));
 sg13g2_dfrbp_1 _4868_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net106),
    .D(_0072_),
    .Q_N(_2375_),
    .Q(\top.julia_calc.dest_x[6] ));
 sg13g2_dfrbp_1 _4869_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net104),
    .D(_0073_),
    .Q_N(_2374_),
    .Q(\top.julia_calc.dest_x[7] ));
 sg13g2_dfrbp_1 _4870_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net40),
    .D(_0074_),
    .Q_N(_0055_),
    .Q(\top.julia_calc.dest_x[8] ));
 sg13g2_dfrbp_1 _4871_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net102),
    .D(net439),
    .Q_N(_2373_),
    .Q(\top.julia_calc.new_pixel_group1 ));
 sg13g2_dfrbp_1 _4872_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net100),
    .D(_0075_),
    .Q_N(_0059_),
    .Q(\top.julia_calc.iter_done_reg ));
 sg13g2_dfrbp_1 _4873_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net98),
    .D(net596),
    .Q_N(_2372_),
    .Q(\top.julia_calc.far_outside_reg ));
 sg13g2_dfrbp_1 _4874_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net96),
    .D(_0077_),
    .Q_N(_2371_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _4875_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net95),
    .D(_0078_),
    .Q_N(_2370_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _4876_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net94),
    .D(_0079_),
    .Q_N(_2369_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _4877_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net41),
    .D(_0080_),
    .Q_N(_2382_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _4878_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net156),
    .D(\uio_out0[4] ),
    .Q_N(_2383_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _4879_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net93),
    .D(\uio_out0[5] ),
    .Q_N(_2368_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _4880_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net92),
    .D(_0081_),
    .Q_N(_0000_),
    .Q(\top.julia_calc.write_mode_data ));
 sg13g2_dfrbp_1 _4881_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net90),
    .D(net388),
    .Q_N(_2367_),
    .Q(\top.debouncer_inst.timer[0] ));
 sg13g2_dfrbp_1 _4882_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net89),
    .D(_0083_),
    .Q_N(_2366_),
    .Q(\top.debouncer_inst.timer[1] ));
 sg13g2_dfrbp_1 _4883_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net88),
    .D(_0084_),
    .Q_N(_2365_),
    .Q(\top.debouncer_inst.timer[2] ));
 sg13g2_dfrbp_1 _4884_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net87),
    .D(net385),
    .Q_N(_2364_),
    .Q(\top.debouncer_inst.timer[3] ));
 sg13g2_dfrbp_1 _4885_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net86),
    .D(_0086_),
    .Q_N(_2363_),
    .Q(\top.debouncer_inst.timer[4] ));
 sg13g2_dfrbp_1 _4886_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net85),
    .D(net402),
    .Q_N(_2362_),
    .Q(\top.debouncer_inst.timer[5] ));
 sg13g2_dfrbp_1 _4887_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net84),
    .D(_0088_),
    .Q_N(_2361_),
    .Q(\top.debouncer_inst.timer[6] ));
 sg13g2_dfrbp_1 _4888_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net83),
    .D(_0089_),
    .Q_N(_2360_),
    .Q(\top.debouncer_inst.timer[7] ));
 sg13g2_dfrbp_1 _4889_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net82),
    .D(net373),
    .Q_N(_2359_),
    .Q(\top.debouncer_inst.timer[8] ));
 sg13g2_dfrbp_1 _4890_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net81),
    .D(_0091_),
    .Q_N(_2358_),
    .Q(\top.debouncer_inst.timer[9] ));
 sg13g2_dfrbp_1 _4891_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net80),
    .D(net411),
    .Q_N(_2357_),
    .Q(\top.debouncer_inst.timer[10] ));
 sg13g2_dfrbp_1 _4892_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net79),
    .D(_0093_),
    .Q_N(_2356_),
    .Q(\top.debouncer_inst.timer[11] ));
 sg13g2_dfrbp_1 _4893_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net78),
    .D(_0094_),
    .Q_N(_2355_),
    .Q(\top.debouncer_inst.timer[12] ));
 sg13g2_dfrbp_1 _4894_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net77),
    .D(_0095_),
    .Q_N(_2354_),
    .Q(\top.debouncer_inst.timer[13] ));
 sg13g2_dfrbp_1 _4895_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net76),
    .D(net369),
    .Q_N(_2353_),
    .Q(\top.debouncer_inst.timer[14] ));
 sg13g2_dfrbp_1 _4896_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net75),
    .D(_0097_),
    .Q_N(_2352_),
    .Q(\top.debouncer_inst.timer[15] ));
 sg13g2_dfrbp_1 _4897_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net74),
    .D(net399),
    .Q_N(_2351_),
    .Q(\top.debouncer_inst.timer[16] ));
 sg13g2_dfrbp_1 _4898_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net73),
    .D(_0099_),
    .Q_N(_2350_),
    .Q(\top.debouncer_inst.timer[17] ));
 sg13g2_dfrbp_1 _4899_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net72),
    .D(_0100_),
    .Q_N(_2349_),
    .Q(\top.debouncer_inst.timer[18] ));
 sg13g2_dfrbp_1 _4900_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net71),
    .D(_0101_),
    .Q_N(_0024_),
    .Q(\top.buttons_stable ));
 sg13g2_dfrbp_1 _4901_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net70),
    .D(net632),
    .Q_N(_2348_),
    .Q(\top.julia_calc.write_addr_available ));
 sg13g2_dfrbp_1 _4902_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net69),
    .D(_0103_),
    .Q_N(_2347_),
    .Q(\top.julia_calc.write_data_available ));
 sg13g2_dfrbp_1 _4903_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net68),
    .D(_0104_),
    .Q_N(_0034_),
    .Q(\top.julia_calc.z_x[0] ));
 sg13g2_dfrbp_1 _4904_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net66),
    .D(_0105_),
    .Q_N(_0038_),
    .Q(\top.julia_calc.z_x[1] ));
 sg13g2_dfrbp_1 _4905_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net64),
    .D(_0106_),
    .Q_N(_0042_),
    .Q(\top.julia_calc.z_x[2] ));
 sg13g2_dfrbp_1 _4906_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net62),
    .D(_0107_),
    .Q_N(_0035_),
    .Q(\top.julia_calc.z_y[0] ));
 sg13g2_dfrbp_1 _4907_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net60),
    .D(_0108_),
    .Q_N(_0039_),
    .Q(\top.julia_calc.z_y[1] ));
 sg13g2_dfrbp_1 _4908_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net58),
    .D(net364),
    .Q_N(_0043_),
    .Q(\top.julia_calc.z_y[2] ));
 sg13g2_dfrbp_1 _4909_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net56),
    .D(net626),
    .Q_N(_2346_),
    .Q(\top.julia_calc.pixel_sreg[0] ));
 sg13g2_dfrbp_1 _4910_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net55),
    .D(net694),
    .Q_N(_2345_),
    .Q(\top.julia_calc.pixel_sreg[1] ));
 sg13g2_dfrbp_1 _4911_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net54),
    .D(net714),
    .Q_N(_2344_),
    .Q(\top.julia_calc.pixel_sreg[2] ));
 sg13g2_dfrbp_1 _4912_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net53),
    .D(net712),
    .Q_N(_2343_),
    .Q(\top.julia_calc.pixel_sreg[3] ));
 sg13g2_dfrbp_1 _4913_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net52),
    .D(net656),
    .Q_N(_2342_),
    .Q(\top.julia_calc.pixel_sreg[4] ));
 sg13g2_dfrbp_1 _4914_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net51),
    .D(_0115_),
    .Q_N(_2341_),
    .Q(\top.julia_calc.pixel_sreg[5] ));
 sg13g2_dfrbp_1 _4915_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net50),
    .D(_0116_),
    .Q_N(_2340_),
    .Q(\top.julia_calc.pixel_sreg[6] ));
 sg13g2_dfrbp_1 _4916_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net49),
    .D(net687),
    .Q_N(_2339_),
    .Q(\top.julia_calc.pixel_sreg[7] ));
 sg13g2_dfrbp_1 _4917_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net48),
    .D(net651),
    .Q_N(_2338_),
    .Q(\top.julia_calc.pixel_sreg[8] ));
 sg13g2_dfrbp_1 _4918_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net47),
    .D(_0119_),
    .Q_N(_2337_),
    .Q(\top.julia_calc.pixel_sreg[9] ));
 sg13g2_dfrbp_1 _4919_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net46),
    .D(_0120_),
    .Q_N(_2336_),
    .Q(\top.julia_calc.pixel_sreg[10] ));
 sg13g2_dfrbp_1 _4920_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net45),
    .D(net654),
    .Q_N(_2335_),
    .Q(\top.julia_calc.pixel_sreg[11] ));
 sg13g2_dfrbp_1 _4921_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net44),
    .D(net645),
    .Q_N(_2334_),
    .Q(\top.julia_calc.pixel_sreg[12] ));
 sg13g2_dfrbp_1 _4922_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net43),
    .D(net703),
    .Q_N(_2333_),
    .Q(\top.julia_calc.pixel_sreg[13] ));
 sg13g2_dfrbp_1 _4923_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net42),
    .D(net658),
    .Q_N(_2332_),
    .Q(\top.julia_calc.pixel_sreg[14] ));
 sg13g2_dfrbp_1 _4924_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net39),
    .D(_0125_),
    .Q_N(_2331_),
    .Q(\top.julia_calc.pixel_sreg[15] ));
 sg13g2_dfrbp_1 _4925_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net38),
    .D(_0126_),
    .Q_N(_2330_),
    .Q(\top.julia_calc.z_x2[0] ));
 sg13g2_dfrbp_1 _4926_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net37),
    .D(_0127_),
    .Q_N(_2329_),
    .Q(\top.julia_calc.z_x2[1] ));
 sg13g2_dfrbp_1 _4927_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net36),
    .D(_0128_),
    .Q_N(_2328_),
    .Q(\top.julia_calc.z_x2[2] ));
 sg13g2_dfrbp_1 _4928_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net35),
    .D(_0129_),
    .Q_N(_2327_),
    .Q(\top.julia_calc.z_x2[3] ));
 sg13g2_dfrbp_1 _4929_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net34),
    .D(_0130_),
    .Q_N(_2326_),
    .Q(\top.julia_calc.z_x2[4] ));
 sg13g2_dfrbp_1 _4930_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net32),
    .D(_0131_),
    .Q_N(_2325_),
    .Q(\top.julia_calc.z_x2[5] ));
 sg13g2_dfrbp_1 _4931_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net31),
    .D(_0132_),
    .Q_N(_2324_),
    .Q(\top.julia_calc.z_x2[6] ));
 sg13g2_dfrbp_1 _4932_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net30),
    .D(_0133_),
    .Q_N(_2323_),
    .Q(\top.julia_calc.z_x2[7] ));
 sg13g2_dfrbp_1 _4933_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net29),
    .D(_0134_),
    .Q_N(_2322_),
    .Q(\top.julia_calc.z_x2[8] ));
 sg13g2_dfrbp_1 _4934_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net28),
    .D(_0135_),
    .Q_N(_2321_),
    .Q(\top.julia_calc.z_x2[9] ));
 sg13g2_dfrbp_1 _4935_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net27),
    .D(_0136_),
    .Q_N(_2320_),
    .Q(\top.julia_calc.z_x2[10] ));
 sg13g2_dfrbp_1 _4936_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net26),
    .D(_0137_),
    .Q_N(_2319_),
    .Q(\top.julia_calc.z_x2[11] ));
 sg13g2_dfrbp_1 _4937_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net25),
    .D(_0138_),
    .Q_N(_2318_),
    .Q(\top.julia_calc.z_x2[12] ));
 sg13g2_dfrbp_1 _4938_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net24),
    .D(_0139_),
    .Q_N(_2317_),
    .Q(\top.julia_calc.z_y2[0] ));
 sg13g2_dfrbp_1 _4939_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net23),
    .D(_0140_),
    .Q_N(_2316_),
    .Q(\top.julia_calc.z_y2[1] ));
 sg13g2_dfrbp_1 _4940_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net22),
    .D(_0141_),
    .Q_N(_2315_),
    .Q(\top.julia_calc.z_y2[2] ));
 sg13g2_dfrbp_1 _4941_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net318),
    .D(_0142_),
    .Q_N(_2314_),
    .Q(\top.julia_calc.z_y2[3] ));
 sg13g2_dfrbp_1 _4942_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net317),
    .D(_0143_),
    .Q_N(_2313_),
    .Q(\top.julia_calc.z_y2[4] ));
 sg13g2_dfrbp_1 _4943_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net316),
    .D(_0144_),
    .Q_N(_2312_),
    .Q(\top.julia_calc.z_y2[5] ));
 sg13g2_dfrbp_1 _4944_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net315),
    .D(_0145_),
    .Q_N(_2311_),
    .Q(\top.julia_calc.z_y2[6] ));
 sg13g2_dfrbp_1 _4945_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net314),
    .D(_0146_),
    .Q_N(_2310_),
    .Q(\top.julia_calc.z_y2[7] ));
 sg13g2_dfrbp_1 _4946_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net313),
    .D(_0147_),
    .Q_N(_2309_),
    .Q(\top.julia_calc.z_y2[8] ));
 sg13g2_dfrbp_1 _4947_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net312),
    .D(_0148_),
    .Q_N(_2308_),
    .Q(\top.julia_calc.z_y2[9] ));
 sg13g2_dfrbp_1 _4948_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net311),
    .D(_0149_),
    .Q_N(_2307_),
    .Q(\top.julia_calc.z_y2[10] ));
 sg13g2_dfrbp_1 _4949_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net310),
    .D(_0150_),
    .Q_N(_2306_),
    .Q(\top.julia_calc.z_y2[11] ));
 sg13g2_dfrbp_1 _4950_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net309),
    .D(_0151_),
    .Q_N(_2305_),
    .Q(\top.julia_calc.z_y2[12] ));
 sg13g2_dfrbp_1 _4951_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net294),
    .D(_0152_),
    .Q_N(_2304_),
    .Q(\top.julia_calc.z_xy[0] ));
 sg13g2_dfrbp_1 _4952_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net293),
    .D(_0153_),
    .Q_N(_2303_),
    .Q(\top.julia_calc.z_xy[1] ));
 sg13g2_dfrbp_1 _4953_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net292),
    .D(_0154_),
    .Q_N(_2302_),
    .Q(\top.julia_calc.z_xy[2] ));
 sg13g2_dfrbp_1 _4954_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net291),
    .D(_0155_),
    .Q_N(_2301_),
    .Q(\top.julia_calc.z_xy[3] ));
 sg13g2_dfrbp_1 _4955_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net290),
    .D(net755),
    .Q_N(_2300_),
    .Q(\top.julia_calc.z_xy[4] ));
 sg13g2_dfrbp_1 _4956_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net289),
    .D(net747),
    .Q_N(_2299_),
    .Q(\top.julia_calc.z_xy[5] ));
 sg13g2_dfrbp_1 _4957_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net288),
    .D(_0158_),
    .Q_N(_2298_),
    .Q(\top.julia_calc.z_xy[6] ));
 sg13g2_dfrbp_1 _4958_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net287),
    .D(_0159_),
    .Q_N(_2297_),
    .Q(\top.julia_calc.z_xy[7] ));
 sg13g2_dfrbp_1 _4959_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net286),
    .D(_0160_),
    .Q_N(_2296_),
    .Q(\top.julia_calc.z_xy[8] ));
 sg13g2_dfrbp_1 _4960_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net285),
    .D(_0161_),
    .Q_N(_2295_),
    .Q(\top.julia_calc.z_xy[9] ));
 sg13g2_dfrbp_1 _4961_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net284),
    .D(_0162_),
    .Q_N(_2294_),
    .Q(\top.julia_calc.z_xy[10] ));
 sg13g2_dfrbp_1 _4962_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net283),
    .D(_0163_),
    .Q_N(_2293_),
    .Q(\top.julia_calc.z_xy[11] ));
 sg13g2_dfrbp_1 _4963_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net282),
    .D(_0164_),
    .Q_N(_2292_),
    .Q(\top.julia_calc.iter[0] ));
 sg13g2_dfrbp_1 _4964_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net280),
    .D(net709),
    .Q_N(_2291_),
    .Q(\top.julia_calc.iter[1] ));
 sg13g2_dfrbp_1 _4965_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net278),
    .D(_0166_),
    .Q_N(_2290_),
    .Q(\top.julia_calc.iter[2] ));
 sg13g2_dfrbp_1 _4966_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net276),
    .D(_0167_),
    .Q_N(_2289_),
    .Q(\top.julia_calc.iter[3] ));
 sg13g2_dfrbp_1 _4967_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net274),
    .D(net670),
    .Q_N(_2288_),
    .Q(\top.julia_calc.iter[4] ));
 sg13g2_dfrbp_1 _4968_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net272),
    .D(_0169_),
    .Q_N(_2287_),
    .Q(\top.julia_calc.iter[5] ));
 sg13g2_dfrbp_1 _4969_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net270),
    .D(_0170_),
    .Q_N(_2286_),
    .Q(\top.julia_calc.iter[6] ));
 sg13g2_dfrbp_1 _4970_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net268),
    .D(_0171_),
    .Q_N(_2285_),
    .Q(\top.julia_calc.iter[7] ));
 sg13g2_dfrbp_1 _4971_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net266),
    .D(_0172_),
    .Q_N(_0056_),
    .Q(\top.julia_calc.iter[8] ));
 sg13g2_dfrbp_1 _4972_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net264),
    .D(_0173_),
    .Q_N(_0062_),
    .Q(\top.receiver.receiver.counter[0] ));
 sg13g2_dfrbp_1 _4973_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net263),
    .D(_0174_),
    .Q_N(_2284_),
    .Q(\top.receiver.receiver.counter[1] ));
 sg13g2_dfrbp_1 _4974_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net262),
    .D(net859),
    .Q_N(_2283_),
    .Q(\top.receiver.receiver.counter[2] ));
 sg13g2_dfrbp_1 _4975_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net261),
    .D(net643),
    .Q_N(_2282_),
    .Q(\top.receiver.receiver.counter[3] ));
 sg13g2_dfrbp_1 _4976_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net260),
    .D(_0177_),
    .Q_N(_0061_),
    .Q(\top.early_x[0] ));
 sg13g2_dfrbp_1 _4977_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net259),
    .D(net763),
    .Q_N(_2281_),
    .Q(\top.early_x[1] ));
 sg13g2_dfrbp_1 _4978_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net258),
    .D(net872),
    .Q_N(_2280_),
    .Q(\top.early_x[2] ));
 sg13g2_dfrbp_1 _4979_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net257),
    .D(_0180_),
    .Q_N(_2279_),
    .Q(\top.early_x[3] ));
 sg13g2_dfrbp_1 _4980_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net256),
    .D(_0181_),
    .Q_N(_2278_),
    .Q(\top.rs.x[4] ));
 sg13g2_dfrbp_1 _4981_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net255),
    .D(_0182_),
    .Q_N(_2277_),
    .Q(\top.rs.x[5] ));
 sg13g2_dfrbp_1 _4982_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net254),
    .D(_0183_),
    .Q_N(_2276_),
    .Q(\top.rs.x[6] ));
 sg13g2_dfrbp_1 _4983_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net253),
    .D(_0184_),
    .Q_N(_2275_),
    .Q(\top.rs.x[7] ));
 sg13g2_dfrbp_1 _4984_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net252),
    .D(_0185_),
    .Q_N(_0022_),
    .Q(\top.rs.x[8] ));
 sg13g2_dfrbp_1 _4985_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net251),
    .D(_0186_),
    .Q_N(_2274_),
    .Q(\top.rs.x[9] ));
 sg13g2_dfrbp_1 _4986_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net250),
    .D(_0187_),
    .Q_N(_2273_),
    .Q(\top.rs.x[10] ));
 sg13g2_dfrbp_1 _4987_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net229),
    .D(_0188_),
    .Q_N(_0058_),
    .Q(\top.rs.x[11] ));
 sg13g2_dfrbp_1 _4988_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net226),
    .D(net413),
    .Q_N(_2272_),
    .Q(\top.last_stable_buttons[0] ));
 sg13g2_dfrbp_1 _4989_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net225),
    .D(net726),
    .Q_N(_2271_),
    .Q(\top.last_stable_buttons[1] ));
 sg13g2_dfrbp_1 _4990_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net224),
    .D(net593),
    .Q_N(_2270_),
    .Q(\top.last_stable_buttons[2] ));
 sg13g2_dfrbp_1 _4991_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net223),
    .D(net696),
    .Q_N(_2269_),
    .Q(\top.last_stable_buttons[3] ));
 sg13g2_dfrbp_1 _4992_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net220),
    .D(net743),
    .Q_N(_2268_),
    .Q(\top.last_stable_buttons[4] ));
 sg13g2_dfrbp_1 _4993_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net157),
    .D(net728),
    .Q_N(_2384_),
    .Q(\top.last_stable_buttons[5] ));
 sg13g2_dfrbp_1 _4994_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net158),
    .D(net1),
    .Q_N(_2385_),
    .Q(\top.debouncer_inst.last_data[0] ));
 sg13g2_dfrbp_1 _4995_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net159),
    .D(net2),
    .Q_N(_2386_),
    .Q(\top.debouncer_inst.last_data[1] ));
 sg13g2_dfrbp_1 _4996_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net160),
    .D(net3),
    .Q_N(_2387_),
    .Q(\top.debouncer_inst.last_data[2] ));
 sg13g2_dfrbp_1 _4997_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net161),
    .D(net4),
    .Q_N(_2388_),
    .Q(\top.debouncer_inst.last_data[3] ));
 sg13g2_dfrbp_1 _4998_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net221),
    .D(net5),
    .Q_N(_2389_),
    .Q(\top.debouncer_inst.last_data[4] ));
 sg13g2_dfrbp_1 _4999_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net219),
    .D(net6),
    .Q_N(_2267_),
    .Q(\top.debouncer_inst.last_data[5] ));
 sg13g2_dfrbp_1 _5000_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net218),
    .D(_0195_),
    .Q_N(_2266_),
    .Q(\top.step_size[0] ));
 sg13g2_dfrbp_1 _5001_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net217),
    .D(_0196_),
    .Q_N(_2265_),
    .Q(\top.step_size[1] ));
 sg13g2_dfrbp_1 _5002_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net216),
    .D(_0197_),
    .Q_N(_0026_),
    .Q(\top.step_size[2] ));
 sg13g2_dfrbp_1 _5003_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net215),
    .D(net828),
    .Q_N(_0023_),
    .Q(\top.step_size[3] ));
 sg13g2_dfrbp_1 _5004_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net214),
    .D(net692),
    .Q_N(_2264_),
    .Q(\top.pixel_buffer[8][0] ));
 sg13g2_dfrbp_1 _5005_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net213),
    .D(net678),
    .Q_N(_2263_),
    .Q(\top.pixel_buffer[8][1] ));
 sg13g2_dfrbp_1 _5006_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net212),
    .D(_0201_),
    .Q_N(_2262_),
    .Q(\top.pixel_buffer[9][0] ));
 sg13g2_dfrbp_1 _5007_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net211),
    .D(_0202_),
    .Q_N(_2261_),
    .Q(\top.pixel_buffer[9][1] ));
 sg13g2_dfrbp_1 _5008_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net210),
    .D(_0203_),
    .Q_N(_2260_),
    .Q(\top.pixel_buffer[10][0] ));
 sg13g2_dfrbp_1 _5009_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net209),
    .D(_0204_),
    .Q_N(_2259_),
    .Q(\top.pixel_buffer[10][1] ));
 sg13g2_dfrbp_1 _5010_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net208),
    .D(_0205_),
    .Q_N(_2258_),
    .Q(\top.pixel_buffer[11][0] ));
 sg13g2_dfrbp_1 _5011_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net207),
    .D(_0206_),
    .Q_N(_2257_),
    .Q(\top.pixel_buffer[11][1] ));
 sg13g2_dfrbp_1 _5012_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net206),
    .D(_0207_),
    .Q_N(_2256_),
    .Q(\top.pixel_buffer[12][0] ));
 sg13g2_dfrbp_1 _5013_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net205),
    .D(_0208_),
    .Q_N(_2255_),
    .Q(\top.pixel_buffer[12][1] ));
 sg13g2_dfrbp_1 _5014_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net204),
    .D(_0209_),
    .Q_N(_2254_),
    .Q(\top.pixel_buffer[13][0] ));
 sg13g2_dfrbp_1 _5015_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net203),
    .D(_0210_),
    .Q_N(_2253_),
    .Q(\top.pixel_buffer[13][1] ));
 sg13g2_dfrbp_1 _5016_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net202),
    .D(_0211_),
    .Q_N(_2252_),
    .Q(\top.pixel_buffer[14][0] ));
 sg13g2_dfrbp_1 _5017_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net201),
    .D(_0212_),
    .Q_N(_2251_),
    .Q(\top.pixel_buffer[14][1] ));
 sg13g2_dfrbp_1 _5018_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net200),
    .D(_0213_),
    .Q_N(_2250_),
    .Q(\top.pixel_buffer[15][0] ));
 sg13g2_dfrbp_1 _5019_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net199),
    .D(_0214_),
    .Q_N(_2249_),
    .Q(\top.pixel_buffer[15][1] ));
 sg13g2_dfrbp_1 _5020_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net198),
    .D(net660),
    .Q_N(_2248_),
    .Q(\top.julia_calc.w_addr[0] ));
 sg13g2_dfrbp_1 _5021_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net197),
    .D(net630),
    .Q_N(_2247_),
    .Q(\top.julia_calc.w_addr[1] ));
 sg13g2_dfrbp_1 _5022_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net196),
    .D(net685),
    .Q_N(_2246_),
    .Q(\top.julia_calc.w_addr[2] ));
 sg13g2_dfrbp_1 _5023_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net195),
    .D(net666),
    .Q_N(_2245_),
    .Q(\top.julia_calc.w_addr[3] ));
 sg13g2_dfrbp_1 _5024_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net194),
    .D(net718),
    .Q_N(_2244_),
    .Q(\top.julia_calc.w_addr[4] ));
 sg13g2_dfrbp_1 _5025_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net193),
    .D(net619),
    .Q_N(_2243_),
    .Q(\top.julia_calc.w_addr[5] ));
 sg13g2_dfrbp_1 _5026_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net192),
    .D(net672),
    .Q_N(_2242_),
    .Q(\top.julia_calc.w_addr[6] ));
 sg13g2_dfrbp_1 _5027_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net191),
    .D(net676),
    .Q_N(_2241_),
    .Q(\top.julia_calc.w_addr[7] ));
 sg13g2_dfrbp_1 _5028_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net190),
    .D(net600),
    .Q_N(_2240_),
    .Q(\top.julia_calc.w_addr[8] ));
 sg13g2_dfrbp_1 _5029_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net189),
    .D(net683),
    .Q_N(_2239_),
    .Q(\top.julia_calc.w_addr[9] ));
 sg13g2_dfrbp_1 _5030_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net188),
    .D(net617),
    .Q_N(_2238_),
    .Q(\top.julia_calc.w_addr[10] ));
 sg13g2_dfrbp_1 _5031_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net187),
    .D(net734),
    .Q_N(_2237_),
    .Q(\top.julia_calc.w_addr[11] ));
 sg13g2_dfrbp_1 _5032_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net186),
    .D(net636),
    .Q_N(_2236_),
    .Q(\top.julia_calc.w_addr[12] ));
 sg13g2_dfrbp_1 _5033_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net185),
    .D(net674),
    .Q_N(_2235_),
    .Q(\top.julia_calc.w_addr[13] ));
 sg13g2_dfrbp_1 _5034_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net184),
    .D(_0229_),
    .Q_N(_2234_),
    .Q(\top.julia_calc.w_addr[14] ));
 sg13g2_dfrbp_1 _5035_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net183),
    .D(_0230_),
    .Q_N(_2233_),
    .Q(\top.c_y[0] ));
 sg13g2_dfrbp_1 _5036_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net182),
    .D(_0231_),
    .Q_N(_2232_),
    .Q(\top.c_y[1] ));
 sg13g2_dfrbp_1 _5037_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net181),
    .D(_0232_),
    .Q_N(_2231_),
    .Q(\top.c_y[2] ));
 sg13g2_dfrbp_1 _5038_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net180),
    .D(_0233_),
    .Q_N(_0028_),
    .Q(\top.c_y[3] ));
 sg13g2_dfrbp_1 _5039_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net179),
    .D(_0234_),
    .Q_N(_2230_),
    .Q(\top.c_y[4] ));
 sg13g2_dfrbp_1 _5040_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net178),
    .D(_0235_),
    .Q_N(_0029_),
    .Q(\top.c_y[5] ));
 sg13g2_dfrbp_1 _5041_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net177),
    .D(_0236_),
    .Q_N(_2229_),
    .Q(\top.c_y[6] ));
 sg13g2_dfrbp_1 _5042_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net176),
    .D(_0237_),
    .Q_N(_2228_),
    .Q(\top.c_y[7] ));
 sg13g2_dfrbp_1 _5043_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net175),
    .D(_0238_),
    .Q_N(_2227_),
    .Q(\top.c_y[8] ));
 sg13g2_dfrbp_1 _5044_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net174),
    .D(_0239_),
    .Q_N(_2226_),
    .Q(\top.c_y[9] ));
 sg13g2_dfrbp_1 _5045_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net173),
    .D(_0240_),
    .Q_N(_2225_),
    .Q(\top.c_y[10] ));
 sg13g2_dfrbp_1 _5046_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net172),
    .D(net864),
    .Q_N(_2224_),
    .Q(\top.c_y[11] ));
 sg13g2_dfrbp_1 _5047_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net171),
    .D(_0242_),
    .Q_N(_2223_),
    .Q(\top.c_x[0] ));
 sg13g2_dfrbp_1 _5048_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net170),
    .D(_0243_),
    .Q_N(_2222_),
    .Q(\top.c_x[1] ));
 sg13g2_dfrbp_1 _5049_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net169),
    .D(_0244_),
    .Q_N(_2221_),
    .Q(\top.c_x[2] ));
 sg13g2_dfrbp_1 _5050_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net168),
    .D(_0245_),
    .Q_N(_0025_),
    .Q(\top.c_x[3] ));
 sg13g2_dfrbp_1 _5051_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net167),
    .D(_0246_),
    .Q_N(_2220_),
    .Q(\top.c_x[4] ));
 sg13g2_dfrbp_1 _5052_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net166),
    .D(net842),
    .Q_N(_0027_),
    .Q(\top.c_x[5] ));
 sg13g2_dfrbp_1 _5053_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net165),
    .D(_0248_),
    .Q_N(_2219_),
    .Q(\top.c_x[6] ));
 sg13g2_dfrbp_1 _5054_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net164),
    .D(_0249_),
    .Q_N(_2218_),
    .Q(\top.c_x[7] ));
 sg13g2_dfrbp_1 _5055_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net163),
    .D(_0250_),
    .Q_N(_2217_),
    .Q(\top.c_x[8] ));
 sg13g2_dfrbp_1 _5056_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net162),
    .D(net879),
    .Q_N(_2216_),
    .Q(\top.c_x[9] ));
 sg13g2_dfrbp_1 _5057_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net155),
    .D(_0252_),
    .Q_N(_2215_),
    .Q(\top.c_x[10] ));
 sg13g2_dfrbp_1 _5058_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net222),
    .D(_0253_),
    .Q_N(_2390_),
    .Q(\top.c_x[11] ));
 sg13g2_dfrbp_1 _5059_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net227),
    .D(net8),
    .Q_N(_2391_),
    .Q(\rx_pins[0] ));
 sg13g2_dfrbp_1 _5060_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net154),
    .D(net9),
    .Q_N(_2214_),
    .Q(\rx_pins[1] ));
 sg13g2_dfrbp_1 _5061_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net153),
    .D(net336),
    .Q_N(_0060_),
    .Q(\top.transmitter.transmitter.counter[0] ));
 sg13g2_dfrbp_1 _5062_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net152),
    .D(_0255_),
    .Q_N(_2213_),
    .Q(\top.transmitter.transmitter.counter[1] ));
 sg13g2_dfrbp_1 _5063_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net151),
    .D(net839),
    .Q_N(_2212_),
    .Q(\top.transmitter.transmitter.counter[2] ));
 sg13g2_dfrbp_1 _5064_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net228),
    .D(net835),
    .Q_N(_2392_),
    .Q(\top.transmitter.transmitter.counter[3] ));
 sg13g2_dfrbp_1 _5065_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net230),
    .D(net784),
    .Q_N(_2393_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _5066_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net150),
    .D(net793),
    .Q_N(_2211_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _5067_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net231),
    .D(_0258_),
    .Q_N(_2394_),
    .Q(\top.transmitter.transmitter.tx_sreg[1] ));
 sg13g2_dfrbp_1 _5068_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net232),
    .D(net434),
    .Q_N(_2395_),
    .Q(\top.transmitter.transmitter.tx_sreg[0] ));
 sg13g2_dfrbp_1 _5069_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net233),
    .D(net428),
    .Q_N(_2396_),
    .Q(\top.transmitter.transmitter.tx_sreg[2] ));
 sg13g2_dfrbp_1 _5070_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net234),
    .D(_0013_),
    .Q_N(_2397_),
    .Q(\top.transmitter.transmitter.tx_sreg[3] ));
 sg13g2_dfrbp_1 _5071_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net235),
    .D(net408),
    .Q_N(_2398_),
    .Q(\top.transmitter.transmitter.tx_sreg[4] ));
 sg13g2_dfrbp_1 _5072_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net236),
    .D(net404),
    .Q_N(_2399_),
    .Q(\top.transmitter.transmitter.tx_sreg[5] ));
 sg13g2_dfrbp_1 _5073_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net237),
    .D(_0016_),
    .Q_N(_2400_),
    .Q(\top.transmitter.transmitter.tx_sreg[6] ));
 sg13g2_dfrbp_1 _5074_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net238),
    .D(net641),
    .Q_N(_2401_),
    .Q(\top.transmitter.transmitter.tx_sreg[7] ));
 sg13g2_dfrbp_1 _5075_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net239),
    .D(net366),
    .Q_N(_2402_),
    .Q(\top.transmitter.transmitter.tx_sreg[8] ));
 sg13g2_dfrbp_1 _5076_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net240),
    .D(_0019_),
    .Q_N(_2403_),
    .Q(\top.transmitter.transmitter.tx_sreg[9] ));
 sg13g2_dfrbp_1 _5077_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net241),
    .D(net622),
    .Q_N(_2404_),
    .Q(\top.transmitter.transmitter.tx_sreg[10] ));
 sg13g2_dfrbp_1 _5078_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net242),
    .D(net774),
    .Q_N(_2405_),
    .Q(\top.transmitter.transmitter.tx_sreg[11] ));
 sg13g2_dfrbp_1 _5079_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net243),
    .D(net426),
    .Q_N(_2406_),
    .Q(\top.transmitter.transmitter.tx_sreg[12] ));
 sg13g2_dfrbp_1 _5080_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net244),
    .D(net396),
    .Q_N(_2407_),
    .Q(\top.transmitter.transmitter.tx_sreg[13] ));
 sg13g2_dfrbp_1 _5081_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net245),
    .D(net362),
    .Q_N(_2408_),
    .Q(\top.transmitter.transmitter.tx_sreg[14] ));
 sg13g2_dfrbp_1 _5082_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net246),
    .D(net424),
    .Q_N(_2409_),
    .Q(\top.transmitter.transmitter.tx_sreg[15] ));
 sg13g2_dfrbp_1 _5083_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net247),
    .D(net607),
    .Q_N(_2410_),
    .Q(\top.transmitter.transmitter.tx_sreg[16] ));
 sg13g2_dfrbp_1 _5084_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net248),
    .D(net415),
    .Q_N(_2411_),
    .Q(\top.transmitter.transmitter.tx_sreg[17] ));
 sg13g2_dfrbp_1 _5085_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net249),
    .D(_0010_),
    .Q_N(_2412_),
    .Q(\top.transmitter.transmitter.tx_sreg[18] ));
 sg13g2_dfrbp_1 _5086_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net295),
    .D(_0011_),
    .Q_N(_2413_),
    .Q(\top.transmitter.transmitter.tx_sreg[19] ));
 sg13g2_dfrbp_1 _5087_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net149),
    .D(net447),
    .Q_N(_2210_),
    .Q(\top.transmitter.transmitter.tx_sreg[20] ));
 sg13g2_dfrbp_1 _5088_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net148),
    .D(net394),
    .Q_N(_0054_),
    .Q(\top.pixel_buffer[0][0] ));
 sg13g2_dfrbp_1 _5089_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net147),
    .D(net591),
    .Q_N(_2209_),
    .Q(\top.pixel_buffer[0][1] ));
 sg13g2_dfrbp_1 _5090_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net146),
    .D(_0261_),
    .Q_N(_2208_),
    .Q(\top.pixel_buffer[1][0] ));
 sg13g2_dfrbp_1 _5091_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net145),
    .D(_0262_),
    .Q_N(_2207_),
    .Q(\top.pixel_buffer[1][1] ));
 sg13g2_dfrbp_1 _5092_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net144),
    .D(_0263_),
    .Q_N(_2206_),
    .Q(\top.pixel_buffer[2][0] ));
 sg13g2_dfrbp_1 _5093_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net143),
    .D(_0264_),
    .Q_N(_2205_),
    .Q(\top.pixel_buffer[2][1] ));
 sg13g2_dfrbp_1 _5094_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net142),
    .D(_0265_),
    .Q_N(_2204_),
    .Q(\top.pixel_buffer[3][0] ));
 sg13g2_dfrbp_1 _5095_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net141),
    .D(_0266_),
    .Q_N(_2203_),
    .Q(\top.pixel_buffer[3][1] ));
 sg13g2_dfrbp_1 _5096_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net140),
    .D(_0267_),
    .Q_N(_2202_),
    .Q(\top.pixel_buffer[4][0] ));
 sg13g2_dfrbp_1 _5097_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net139),
    .D(_0268_),
    .Q_N(_2201_),
    .Q(\top.pixel_buffer[4][1] ));
 sg13g2_dfrbp_1 _5098_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net138),
    .D(_0269_),
    .Q_N(_2200_),
    .Q(\top.pixel_buffer[5][0] ));
 sg13g2_dfrbp_1 _5099_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net137),
    .D(_0270_),
    .Q_N(_2199_),
    .Q(\top.pixel_buffer[5][1] ));
 sg13g2_dfrbp_1 _5100_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net136),
    .D(_0271_),
    .Q_N(_2198_),
    .Q(\top.pixel_buffer[6][0] ));
 sg13g2_dfrbp_1 _5101_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net135),
    .D(_0272_),
    .Q_N(_2197_),
    .Q(\top.pixel_buffer[6][1] ));
 sg13g2_dfrbp_1 _5102_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net134),
    .D(_0273_),
    .Q_N(_2196_),
    .Q(\top.pixel_buffer[7][0] ));
 sg13g2_dfrbp_1 _5103_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net133),
    .D(_0274_),
    .Q_N(_2195_),
    .Q(\top.pixel_buffer[7][1] ));
 sg13g2_dfrbp_1 _5104_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net132),
    .D(net350),
    .Q_N(_0032_),
    .Q(\top.julia_calc.z_x[3] ));
 sg13g2_dfrbp_1 _5105_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net131),
    .D(net344),
    .Q_N(_0048_),
    .Q(\top.julia_calc.z_x[4] ));
 sg13g2_dfrbp_1 _5106_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net130),
    .D(net392),
    .Q_N(_0050_),
    .Q(\top.julia_calc.z_x[5] ));
 sg13g2_dfrbp_1 _5107_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net129),
    .D(net355),
    .Q_N(_0046_),
    .Q(\top.julia_calc.z_x[6] ));
 sg13g2_dfrbp_1 _5108_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net128),
    .D(net346),
    .Q_N(_0030_),
    .Q(\top.julia_calc.z_x[7] ));
 sg13g2_dfrbp_1 _5109_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net127),
    .D(net342),
    .Q_N(_0044_),
    .Q(\top.julia_calc.z_x[8] ));
 sg13g2_dfrbp_1 _5110_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net126),
    .D(net602),
    .Q_N(_0040_),
    .Q(\top.julia_calc.z_x[9] ));
 sg13g2_dfrbp_1 _5111_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net125),
    .D(net436),
    .Q_N(_0036_),
    .Q(\top.julia_calc.z_x[10] ));
 sg13g2_dfrbp_1 _5112_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net124),
    .D(net420),
    .Q_N(_0052_),
    .Q(\top.julia_calc.z_x[11] ));
 sg13g2_dfrbp_1 _5113_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net123),
    .D(net390),
    .Q_N(_0033_),
    .Q(\top.julia_calc.z_y[3] ));
 sg13g2_dfrbp_1 _5114_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net122),
    .D(net406),
    .Q_N(_0049_),
    .Q(\top.julia_calc.z_y[4] ));
 sg13g2_dfrbp_1 _5115_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net121),
    .D(_0286_),
    .Q_N(_0051_),
    .Q(\top.julia_calc.z_y[5] ));
 sg13g2_dfrbp_1 _5116_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net120),
    .D(net352),
    .Q_N(_0047_),
    .Q(\top.julia_calc.z_y[6] ));
 sg13g2_dfrbp_1 _5117_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net117),
    .D(net377),
    .Q_N(_0031_),
    .Q(\top.julia_calc.z_y[7] ));
 sg13g2_dfrbp_1 _5118_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net115),
    .D(_0289_),
    .Q_N(_0045_),
    .Q(\top.julia_calc.z_y[8] ));
 sg13g2_dfrbp_1 _5119_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net113),
    .D(net422),
    .Q_N(_0041_),
    .Q(\top.julia_calc.z_y[9] ));
 sg13g2_dfrbp_1 _5120_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net111),
    .D(net438),
    .Q_N(_0037_),
    .Q(\top.julia_calc.z_y[10] ));
 sg13g2_dfrbp_1 _5121_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net109),
    .D(net417),
    .Q_N(_0053_),
    .Q(\top.julia_calc.z_y[11] ));
 sg13g2_dfrbp_1 _5122_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net107),
    .D(_0293_),
    .Q_N(_2194_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _5123_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net105),
    .D(_0294_),
    .Q_N(_2193_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _5124_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net103),
    .D(_0295_),
    .Q_N(_2192_),
    .Q(\top.julia_calc.dest_y[0] ));
 sg13g2_dfrbp_1 _5125_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net101),
    .D(_0296_),
    .Q_N(_2191_),
    .Q(\top.julia_calc.dest_y[1] ));
 sg13g2_dfrbp_1 _5126_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net99),
    .D(_0297_),
    .Q_N(_2190_),
    .Q(\top.julia_calc.dest_y[2] ));
 sg13g2_dfrbp_1 _5127_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net97),
    .D(_0298_),
    .Q_N(_2189_),
    .Q(\top.julia_calc.dest_y[3] ));
 sg13g2_dfrbp_1 _5128_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net91),
    .D(_0299_),
    .Q_N(_0020_),
    .Q(\top.julia_calc.dest_y[4] ));
 sg13g2_dfrbp_1 _5129_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net67),
    .D(_0300_),
    .Q_N(_2188_),
    .Q(\top.julia_calc.dest_y[5] ));
 sg13g2_dfrbp_1 _5130_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net65),
    .D(_0301_),
    .Q_N(_2187_),
    .Q(\top.julia_calc.dest_y[6] ));
 sg13g2_dfrbp_1 _5131_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net63),
    .D(_0302_),
    .Q_N(_2186_),
    .Q(\top.julia_calc.dest_y[7] ));
 sg13g2_dfrbp_1 _5132_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net296),
    .D(_0303_),
    .Q_N(_0057_),
    .Q(\top.julia_calc.dest_y[8] ));
 sg13g2_dfrbp_1 _5133_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net297),
    .D(net322),
    .Q_N(_2414_),
    .Q(\top.receiver.data[0] ));
 sg13g2_dfrbp_1 _5134_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net298),
    .D(net323),
    .Q_N(_2415_),
    .Q(\top.receiver.data[1] ));
 sg13g2_dfrbp_1 _5135_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net299),
    .D(net329),
    .Q_N(_2416_),
    .Q(\top.receiver.data[2] ));
 sg13g2_dfrbp_1 _5136_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net300),
    .D(net333),
    .Q_N(_2417_),
    .Q(\top.receiver.data[3] ));
 sg13g2_dfrbp_1 _5137_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net301),
    .D(net332),
    .Q_N(_2418_),
    .Q(\top.receiver.data[4] ));
 sg13g2_dfrbp_1 _5138_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net302),
    .D(net326),
    .Q_N(_2419_),
    .Q(\top.receiver.data[5] ));
 sg13g2_dfrbp_1 _5139_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net303),
    .D(net331),
    .Q_N(_2420_),
    .Q(\top.receiver.data[6] ));
 sg13g2_dfrbp_1 _5140_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net304),
    .D(net337),
    .Q_N(_2421_),
    .Q(\top.receiver.data[7] ));
 sg13g2_dfrbp_1 _5141_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net305),
    .D(net324),
    .Q_N(_2422_),
    .Q(\top.receiver.data[8] ));
 sg13g2_dfrbp_1 _5142_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net306),
    .D(net334),
    .Q_N(_2423_),
    .Q(\top.receiver.data[9] ));
 sg13g2_dfrbp_1 _5143_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net307),
    .D(net325),
    .Q_N(_2424_),
    .Q(\top.receiver.data[10] ));
 sg13g2_dfrbp_1 _5144_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net308),
    .D(net327),
    .Q_N(_2425_),
    .Q(\top.receiver.data[11] ));
 sg13g2_dfrbp_1 _5145_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net265),
    .D(net330),
    .Q_N(_2426_),
    .Q(\top.receiver.data[12] ));
 sg13g2_dfrbp_1 _5146_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net61),
    .D(net321),
    .Q_N(_2185_),
    .Q(\top.receiver.data[13] ));
 sg13g2_dfrbp_1 _5147_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net59),
    .D(_0304_),
    .Q_N(_2184_),
    .Q(\top.next_read_addr[6] ));
 sg13g2_dfrbp_1 _5148_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net57),
    .D(_0305_),
    .Q_N(_2183_),
    .Q(\top.next_read_addr[7] ));
 sg13g2_dfrbp_1 _5149_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net281),
    .D(net823),
    .Q_N(_2182_),
    .Q(\top.next_read_addr[8] ));
 sg13g2_dfrbp_1 _5150_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net279),
    .D(_0307_),
    .Q_N(_2181_),
    .Q(\top.next_read_addr[9] ));
 sg13g2_dfrbp_1 _5151_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net277),
    .D(_0308_),
    .Q_N(_2180_),
    .Q(\top.next_read_addr[10] ));
 sg13g2_dfrbp_1 _5152_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net275),
    .D(_0309_),
    .Q_N(_2179_),
    .Q(\top.next_read_addr[11] ));
 sg13g2_dfrbp_1 _5153_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net273),
    .D(_0310_),
    .Q_N(_2178_),
    .Q(\top.next_read_addr[12] ));
 sg13g2_dfrbp_1 _5154_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net271),
    .D(_0311_),
    .Q_N(_2177_),
    .Q(\top.next_read_addr[13] ));
 sg13g2_dfrbp_1 _5155_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net269),
    .D(_0312_),
    .Q_N(_2176_),
    .Q(\top.next_read_addr[14] ));
 sg13g2_dfrbp_1 _5156_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net267),
    .D(_0313_),
    .Q_N(_2175_),
    .Q(\top.rs.y[9] ));
 sg13g2_tiehi _4939__23 (.L_HI(net23));
 sg13g2_tiehi _4938__24 (.L_HI(net24));
 sg13g2_tiehi _4937__25 (.L_HI(net25));
 sg13g2_tiehi _4936__26 (.L_HI(net26));
 sg13g2_tiehi _4935__27 (.L_HI(net27));
 sg13g2_tiehi _4934__28 (.L_HI(net28));
 sg13g2_tiehi _4933__29 (.L_HI(net29));
 sg13g2_tiehi _4932__30 (.L_HI(net30));
 sg13g2_tiehi _4931__31 (.L_HI(net31));
 sg13g2_tiehi _4930__32 (.L_HI(net32));
 sg13g2_tiehi _4860__33 (.L_HI(net33));
 sg13g2_tiehi _4929__34 (.L_HI(net34));
 sg13g2_tiehi _4928__35 (.L_HI(net35));
 sg13g2_tiehi _4927__36 (.L_HI(net36));
 sg13g2_tiehi _4926__37 (.L_HI(net37));
 sg13g2_tiehi _4925__38 (.L_HI(net38));
 sg13g2_tiehi _4924__39 (.L_HI(net39));
 sg13g2_tiehi _4870__40 (.L_HI(net40));
 sg13g2_tiehi _4877__41 (.L_HI(net41));
 sg13g2_tiehi _4923__42 (.L_HI(net42));
 sg13g2_tiehi _4922__43 (.L_HI(net43));
 sg13g2_tiehi _4921__44 (.L_HI(net44));
 sg13g2_tiehi _4920__45 (.L_HI(net45));
 sg13g2_tiehi _4919__46 (.L_HI(net46));
 sg13g2_tiehi _4918__47 (.L_HI(net47));
 sg13g2_tiehi _4917__48 (.L_HI(net48));
 sg13g2_tiehi _4916__49 (.L_HI(net49));
 sg13g2_tiehi _4915__50 (.L_HI(net50));
 sg13g2_tiehi _4914__51 (.L_HI(net51));
 sg13g2_tiehi _4913__52 (.L_HI(net52));
 sg13g2_tiehi _4912__53 (.L_HI(net53));
 sg13g2_tiehi _4911__54 (.L_HI(net54));
 sg13g2_tiehi _4910__55 (.L_HI(net55));
 sg13g2_tiehi _4909__56 (.L_HI(net56));
 sg13g2_tiehi _5148__57 (.L_HI(net57));
 sg13g2_tiehi _4908__58 (.L_HI(net58));
 sg13g2_tiehi _5147__59 (.L_HI(net59));
 sg13g2_tiehi _4907__60 (.L_HI(net60));
 sg13g2_tiehi _5146__61 (.L_HI(net61));
 sg13g2_tiehi _4906__62 (.L_HI(net62));
 sg13g2_tiehi _5131__63 (.L_HI(net63));
 sg13g2_tiehi _4905__64 (.L_HI(net64));
 sg13g2_tiehi _5130__65 (.L_HI(net65));
 sg13g2_tiehi _4904__66 (.L_HI(net66));
 sg13g2_tiehi _5129__67 (.L_HI(net67));
 sg13g2_tiehi _4903__68 (.L_HI(net68));
 sg13g2_tiehi _4902__69 (.L_HI(net69));
 sg13g2_tiehi _4901__70 (.L_HI(net70));
 sg13g2_tiehi _4900__71 (.L_HI(net71));
 sg13g2_tiehi _4899__72 (.L_HI(net72));
 sg13g2_tiehi _4898__73 (.L_HI(net73));
 sg13g2_tiehi _4897__74 (.L_HI(net74));
 sg13g2_tiehi _4896__75 (.L_HI(net75));
 sg13g2_tiehi _4895__76 (.L_HI(net76));
 sg13g2_tiehi _4894__77 (.L_HI(net77));
 sg13g2_tiehi _4893__78 (.L_HI(net78));
 sg13g2_tiehi _4892__79 (.L_HI(net79));
 sg13g2_tiehi _4891__80 (.L_HI(net80));
 sg13g2_tiehi _4890__81 (.L_HI(net81));
 sg13g2_tiehi _4889__82 (.L_HI(net82));
 sg13g2_tiehi _4888__83 (.L_HI(net83));
 sg13g2_tiehi _4887__84 (.L_HI(net84));
 sg13g2_tiehi _4886__85 (.L_HI(net85));
 sg13g2_tiehi _4885__86 (.L_HI(net86));
 sg13g2_tiehi _4884__87 (.L_HI(net87));
 sg13g2_tiehi _4883__88 (.L_HI(net88));
 sg13g2_tiehi _4882__89 (.L_HI(net89));
 sg13g2_tiehi _4881__90 (.L_HI(net90));
 sg13g2_tiehi _5128__91 (.L_HI(net91));
 sg13g2_tiehi _4880__92 (.L_HI(net92));
 sg13g2_tiehi _4879__93 (.L_HI(net93));
 sg13g2_tiehi _4876__94 (.L_HI(net94));
 sg13g2_tiehi _4875__95 (.L_HI(net95));
 sg13g2_tiehi _4874__96 (.L_HI(net96));
 sg13g2_tiehi _5127__97 (.L_HI(net97));
 sg13g2_tiehi _4873__98 (.L_HI(net98));
 sg13g2_tiehi _5126__99 (.L_HI(net99));
 sg13g2_tiehi _4872__100 (.L_HI(net100));
 sg13g2_tiehi _5125__101 (.L_HI(net101));
 sg13g2_tiehi _4871__102 (.L_HI(net102));
 sg13g2_tiehi _5124__103 (.L_HI(net103));
 sg13g2_tiehi _4869__104 (.L_HI(net104));
 sg13g2_tiehi _5123__105 (.L_HI(net105));
 sg13g2_tiehi _4868__106 (.L_HI(net106));
 sg13g2_tiehi _5122__107 (.L_HI(net107));
 sg13g2_tiehi _4867__108 (.L_HI(net108));
 sg13g2_tiehi _5121__109 (.L_HI(net109));
 sg13g2_tiehi _4866__110 (.L_HI(net110));
 sg13g2_tiehi _5120__111 (.L_HI(net111));
 sg13g2_tiehi _4865__112 (.L_HI(net112));
 sg13g2_tiehi _5119__113 (.L_HI(net113));
 sg13g2_tiehi _4864__114 (.L_HI(net114));
 sg13g2_tiehi _5118__115 (.L_HI(net115));
 sg13g2_tiehi _4863__116 (.L_HI(net116));
 sg13g2_tiehi _5117__117 (.L_HI(net117));
 sg13g2_tiehi _4862__118 (.L_HI(net118));
 sg13g2_tiehi _4861__119 (.L_HI(net119));
 sg13g2_tiehi _5116__120 (.L_HI(net120));
 sg13g2_tiehi _5115__121 (.L_HI(net121));
 sg13g2_tiehi _5114__122 (.L_HI(net122));
 sg13g2_tiehi _5113__123 (.L_HI(net123));
 sg13g2_tiehi _5112__124 (.L_HI(net124));
 sg13g2_tiehi _5111__125 (.L_HI(net125));
 sg13g2_tiehi _5110__126 (.L_HI(net126));
 sg13g2_tiehi _5109__127 (.L_HI(net127));
 sg13g2_tiehi _5108__128 (.L_HI(net128));
 sg13g2_tiehi _5107__129 (.L_HI(net129));
 sg13g2_tiehi _5106__130 (.L_HI(net130));
 sg13g2_tiehi _5105__131 (.L_HI(net131));
 sg13g2_tiehi _5104__132 (.L_HI(net132));
 sg13g2_tiehi _5103__133 (.L_HI(net133));
 sg13g2_tiehi _5102__134 (.L_HI(net134));
 sg13g2_tiehi _5101__135 (.L_HI(net135));
 sg13g2_tiehi _5100__136 (.L_HI(net136));
 sg13g2_tiehi _5099__137 (.L_HI(net137));
 sg13g2_tiehi _5098__138 (.L_HI(net138));
 sg13g2_tiehi _5097__139 (.L_HI(net139));
 sg13g2_tiehi _5096__140 (.L_HI(net140));
 sg13g2_tiehi _5095__141 (.L_HI(net141));
 sg13g2_tiehi _5094__142 (.L_HI(net142));
 sg13g2_tiehi _5093__143 (.L_HI(net143));
 sg13g2_tiehi _5092__144 (.L_HI(net144));
 sg13g2_tiehi _5091__145 (.L_HI(net145));
 sg13g2_tiehi _5090__146 (.L_HI(net146));
 sg13g2_tiehi _5089__147 (.L_HI(net147));
 sg13g2_tiehi _5088__148 (.L_HI(net148));
 sg13g2_tiehi _5087__149 (.L_HI(net149));
 sg13g2_tiehi _5066__150 (.L_HI(net150));
 sg13g2_tiehi _5063__151 (.L_HI(net151));
 sg13g2_tiehi _5062__152 (.L_HI(net152));
 sg13g2_tiehi _5061__153 (.L_HI(net153));
 sg13g2_tiehi _5060__154 (.L_HI(net154));
 sg13g2_tiehi _5057__155 (.L_HI(net155));
 sg13g2_tiehi _4878__156 (.L_HI(net156));
 sg13g2_tiehi _4993__157 (.L_HI(net157));
 sg13g2_tiehi _4994__158 (.L_HI(net158));
 sg13g2_tiehi _4995__159 (.L_HI(net159));
 sg13g2_tiehi _4996__160 (.L_HI(net160));
 sg13g2_tiehi _4997__161 (.L_HI(net161));
 sg13g2_tiehi _5056__162 (.L_HI(net162));
 sg13g2_tiehi _5055__163 (.L_HI(net163));
 sg13g2_tiehi _5054__164 (.L_HI(net164));
 sg13g2_tiehi _5053__165 (.L_HI(net165));
 sg13g2_tiehi _5052__166 (.L_HI(net166));
 sg13g2_tiehi _5051__167 (.L_HI(net167));
 sg13g2_tiehi _5050__168 (.L_HI(net168));
 sg13g2_tiehi _5049__169 (.L_HI(net169));
 sg13g2_tiehi _5048__170 (.L_HI(net170));
 sg13g2_tiehi _5047__171 (.L_HI(net171));
 sg13g2_tiehi _5046__172 (.L_HI(net172));
 sg13g2_tiehi _5045__173 (.L_HI(net173));
 sg13g2_tiehi _5044__174 (.L_HI(net174));
 sg13g2_tiehi _5043__175 (.L_HI(net175));
 sg13g2_tiehi _5042__176 (.L_HI(net176));
 sg13g2_tiehi _5041__177 (.L_HI(net177));
 sg13g2_tiehi _5040__178 (.L_HI(net178));
 sg13g2_tiehi _5039__179 (.L_HI(net179));
 sg13g2_tiehi _5038__180 (.L_HI(net180));
 sg13g2_tiehi _5037__181 (.L_HI(net181));
 sg13g2_tiehi _5036__182 (.L_HI(net182));
 sg13g2_tiehi _5035__183 (.L_HI(net183));
 sg13g2_tiehi _5034__184 (.L_HI(net184));
 sg13g2_tiehi _5033__185 (.L_HI(net185));
 sg13g2_tiehi _5032__186 (.L_HI(net186));
 sg13g2_tiehi _5031__187 (.L_HI(net187));
 sg13g2_tiehi _5030__188 (.L_HI(net188));
 sg13g2_tiehi _5029__189 (.L_HI(net189));
 sg13g2_tiehi _5028__190 (.L_HI(net190));
 sg13g2_tiehi _5027__191 (.L_HI(net191));
 sg13g2_tiehi _5026__192 (.L_HI(net192));
 sg13g2_tiehi _5025__193 (.L_HI(net193));
 sg13g2_tiehi _5024__194 (.L_HI(net194));
 sg13g2_tiehi _5023__195 (.L_HI(net195));
 sg13g2_tiehi _5022__196 (.L_HI(net196));
 sg13g2_tiehi _5021__197 (.L_HI(net197));
 sg13g2_tiehi _5020__198 (.L_HI(net198));
 sg13g2_tiehi _5019__199 (.L_HI(net199));
 sg13g2_tiehi _5018__200 (.L_HI(net200));
 sg13g2_tiehi _5017__201 (.L_HI(net201));
 sg13g2_tiehi _5016__202 (.L_HI(net202));
 sg13g2_tiehi _5015__203 (.L_HI(net203));
 sg13g2_tiehi _5014__204 (.L_HI(net204));
 sg13g2_tiehi _5013__205 (.L_HI(net205));
 sg13g2_tiehi _5012__206 (.L_HI(net206));
 sg13g2_tiehi _5011__207 (.L_HI(net207));
 sg13g2_tiehi _5010__208 (.L_HI(net208));
 sg13g2_tiehi _5009__209 (.L_HI(net209));
 sg13g2_tiehi _5008__210 (.L_HI(net210));
 sg13g2_tiehi _5007__211 (.L_HI(net211));
 sg13g2_tiehi _5006__212 (.L_HI(net212));
 sg13g2_tiehi _5005__213 (.L_HI(net213));
 sg13g2_tiehi _5004__214 (.L_HI(net214));
 sg13g2_tiehi _5003__215 (.L_HI(net215));
 sg13g2_tiehi _5002__216 (.L_HI(net216));
 sg13g2_tiehi _5001__217 (.L_HI(net217));
 sg13g2_tiehi _5000__218 (.L_HI(net218));
 sg13g2_tiehi _4999__219 (.L_HI(net219));
 sg13g2_tiehi _4992__220 (.L_HI(net220));
 sg13g2_tiehi _4998__221 (.L_HI(net221));
 sg13g2_tiehi _5058__222 (.L_HI(net222));
 sg13g2_tiehi _4991__223 (.L_HI(net223));
 sg13g2_tiehi _4990__224 (.L_HI(net224));
 sg13g2_tiehi _4989__225 (.L_HI(net225));
 sg13g2_tiehi _4988__226 (.L_HI(net226));
 sg13g2_tiehi _5059__227 (.L_HI(net227));
 sg13g2_tiehi _5064__228 (.L_HI(net228));
 sg13g2_tiehi _4987__229 (.L_HI(net229));
 sg13g2_tiehi _5065__230 (.L_HI(net230));
 sg13g2_tiehi _5067__231 (.L_HI(net231));
 sg13g2_tiehi _5068__232 (.L_HI(net232));
 sg13g2_tiehi _5069__233 (.L_HI(net233));
 sg13g2_tiehi _5070__234 (.L_HI(net234));
 sg13g2_tiehi _5071__235 (.L_HI(net235));
 sg13g2_tiehi _5072__236 (.L_HI(net236));
 sg13g2_tiehi _5073__237 (.L_HI(net237));
 sg13g2_tiehi _5074__238 (.L_HI(net238));
 sg13g2_tiehi _5075__239 (.L_HI(net239));
 sg13g2_tiehi _5076__240 (.L_HI(net240));
 sg13g2_tiehi _5077__241 (.L_HI(net241));
 sg13g2_tiehi _5078__242 (.L_HI(net242));
 sg13g2_tiehi _5079__243 (.L_HI(net243));
 sg13g2_tiehi _5080__244 (.L_HI(net244));
 sg13g2_tiehi _5081__245 (.L_HI(net245));
 sg13g2_tiehi _5082__246 (.L_HI(net246));
 sg13g2_tiehi _5083__247 (.L_HI(net247));
 sg13g2_tiehi _5084__248 (.L_HI(net248));
 sg13g2_tiehi _5085__249 (.L_HI(net249));
 sg13g2_tiehi _4986__250 (.L_HI(net250));
 sg13g2_tiehi _4985__251 (.L_HI(net251));
 sg13g2_tiehi _4984__252 (.L_HI(net252));
 sg13g2_tiehi _4983__253 (.L_HI(net253));
 sg13g2_tiehi _4982__254 (.L_HI(net254));
 sg13g2_tiehi _4981__255 (.L_HI(net255));
 sg13g2_tiehi _4980__256 (.L_HI(net256));
 sg13g2_tiehi _4979__257 (.L_HI(net257));
 sg13g2_tiehi _4978__258 (.L_HI(net258));
 sg13g2_tiehi _4977__259 (.L_HI(net259));
 sg13g2_tiehi _4976__260 (.L_HI(net260));
 sg13g2_tiehi _4975__261 (.L_HI(net261));
 sg13g2_tiehi _4974__262 (.L_HI(net262));
 sg13g2_tiehi _4973__263 (.L_HI(net263));
 sg13g2_tiehi _4972__264 (.L_HI(net264));
 sg13g2_tiehi _5145__265 (.L_HI(net265));
 sg13g2_tiehi _4971__266 (.L_HI(net266));
 sg13g2_tiehi _5156__267 (.L_HI(net267));
 sg13g2_tiehi _4970__268 (.L_HI(net268));
 sg13g2_tiehi _5155__269 (.L_HI(net269));
 sg13g2_tiehi _4969__270 (.L_HI(net270));
 sg13g2_tiehi _5154__271 (.L_HI(net271));
 sg13g2_tiehi _4968__272 (.L_HI(net272));
 sg13g2_tiehi _5153__273 (.L_HI(net273));
 sg13g2_tiehi _4967__274 (.L_HI(net274));
 sg13g2_tiehi _5152__275 (.L_HI(net275));
 sg13g2_tiehi _4966__276 (.L_HI(net276));
 sg13g2_tiehi _5151__277 (.L_HI(net277));
 sg13g2_tiehi _4965__278 (.L_HI(net278));
 sg13g2_tiehi _5150__279 (.L_HI(net279));
 sg13g2_tiehi _4964__280 (.L_HI(net280));
 sg13g2_tiehi _5149__281 (.L_HI(net281));
 sg13g2_tiehi _4963__282 (.L_HI(net282));
 sg13g2_tiehi _4962__283 (.L_HI(net283));
 sg13g2_tiehi _4961__284 (.L_HI(net284));
 sg13g2_tiehi _4960__285 (.L_HI(net285));
 sg13g2_tiehi _4959__286 (.L_HI(net286));
 sg13g2_tiehi _4958__287 (.L_HI(net287));
 sg13g2_tiehi _4957__288 (.L_HI(net288));
 sg13g2_tiehi _4956__289 (.L_HI(net289));
 sg13g2_tiehi _4955__290 (.L_HI(net290));
 sg13g2_tiehi _4954__291 (.L_HI(net291));
 sg13g2_tiehi _4953__292 (.L_HI(net292));
 sg13g2_tiehi _4952__293 (.L_HI(net293));
 sg13g2_tiehi _4951__294 (.L_HI(net294));
 sg13g2_tiehi _5086__295 (.L_HI(net295));
 sg13g2_tiehi _5132__296 (.L_HI(net296));
 sg13g2_tiehi _5133__297 (.L_HI(net297));
 sg13g2_tiehi _5134__298 (.L_HI(net298));
 sg13g2_tiehi _5135__299 (.L_HI(net299));
 sg13g2_tiehi _5136__300 (.L_HI(net300));
 sg13g2_tiehi _5137__301 (.L_HI(net301));
 sg13g2_tiehi _5138__302 (.L_HI(net302));
 sg13g2_tiehi _5139__303 (.L_HI(net303));
 sg13g2_tiehi _5140__304 (.L_HI(net304));
 sg13g2_tiehi _5141__305 (.L_HI(net305));
 sg13g2_tiehi _5142__306 (.L_HI(net306));
 sg13g2_tiehi _5143__307 (.L_HI(net307));
 sg13g2_tiehi _5144__308 (.L_HI(net308));
 sg13g2_tiehi _4950__309 (.L_HI(net309));
 sg13g2_tiehi _4949__310 (.L_HI(net310));
 sg13g2_tiehi _4948__311 (.L_HI(net311));
 sg13g2_tiehi _4947__312 (.L_HI(net312));
 sg13g2_tiehi _4946__313 (.L_HI(net313));
 sg13g2_tiehi _4945__314 (.L_HI(net314));
 sg13g2_tiehi _4944__315 (.L_HI(net315));
 sg13g2_tiehi _4943__316 (.L_HI(net316));
 sg13g2_tiehi _4942__317 (.L_HI(net317));
 sg13g2_tiehi _4941__318 (.L_HI(net318));
 sg13g2_tiehi tt_um_toivoh_pio_ram_emu_example_319 (.L_HI(net319));
 sg13g2_tiehi tt_um_toivoh_pio_ram_emu_example_320 (.L_HI(net320));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_11 (.L_LO(net11));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_12 (.L_LO(net12));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_13 (.L_LO(net13));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_14 (.L_LO(net14));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_15 (.L_LO(net15));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_16 (.L_LO(net16));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_17 (.L_LO(net17));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_18 (.L_LO(net18));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_19 (.L_LO(net19));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_20 (.L_LO(net20));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_21 (.L_LO(net21));
 sg13g2_tiehi _4940__22 (.L_HI(net22));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(\top.julia_calc.new_pixel_group ));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(_1939_));
 sg13g2_buf_2 fanout441 (.A(_1939_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_1 fanout443 (.A(net444),
    .X(net443));
 sg13g2_buf_1 fanout444 (.A(net445),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(\top.transmitter.message_accepted ),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(\top.transmitter.message_accepted ),
    .X(net446));
 sg13g2_buf_1 fanout447 (.A(\top.transmitter.message_accepted ),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_1809_),
    .X(net448));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(_1227_));
 sg13g2_buf_2 fanout450 (.A(_1183_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_1469_),
    .X(net451));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(_1000_));
 sg13g2_buf_2 fanout453 (.A(_1000_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(net456),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(net456),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_0378_),
    .X(net456));
 sg13g2_buf_4 fanout457 (.X(net457),
    .A(net458));
 sg13g2_buf_4 fanout458 (.X(net458),
    .A(_1700_));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(net461));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(net461));
 sg13g2_buf_1 fanout461 (.A(_1516_),
    .X(net461));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(_1882_));
 sg13g2_buf_2 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_1 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_1 fanout465 (.A(net466),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_1881_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(net468),
    .X(net467));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(_0796_));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_4 fanout470 (.X(net470),
    .A(_0795_));
 sg13g2_buf_2 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(net473),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_4 fanout474 (.X(net474),
    .A(_0786_));
 sg13g2_buf_2 fanout475 (.A(_0599_),
    .X(net475));
 sg13g2_buf_1 fanout476 (.A(_0599_),
    .X(net476));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(_0536_));
 sg13g2_buf_2 fanout478 (.A(net480),
    .X(net478));
 sg13g2_buf_1 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_0524_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_0523_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_0523_),
    .X(net482));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(_0516_));
 sg13g2_buf_1 fanout484 (.A(_0516_),
    .X(net484));
 sg13g2_buf_4 fanout485 (.X(net485),
    .A(_0513_));
 sg13g2_buf_4 fanout486 (.X(net486),
    .A(_0510_));
 sg13g2_buf_2 fanout487 (.A(_0510_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_0498_),
    .X(net488));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(_0482_));
 sg13g2_buf_2 fanout490 (.A(_0482_),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(_0480_));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(_0473_));
 sg13g2_buf_1 fanout493 (.A(_0473_),
    .X(net493));
 sg13g2_buf_4 fanout494 (.X(net494),
    .A(_0467_));
 sg13g2_buf_1 fanout495 (.A(_0467_),
    .X(net495));
 sg13g2_buf_4 fanout496 (.X(net496),
    .A(_0459_));
 sg13g2_buf_2 fanout497 (.A(_0459_),
    .X(net497));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(_0449_));
 sg13g2_buf_2 fanout499 (.A(_0445_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_0443_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_0443_),
    .X(net501));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(_0438_));
 sg13g2_buf_2 fanout503 (.A(_0438_),
    .X(net503));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(_0435_));
 sg13g2_buf_1 fanout505 (.A(_0435_),
    .X(net505));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(net507));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(_0432_));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_1 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_1 fanout510 (.A(_0416_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net515),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(net515),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net515),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(net515),
    .X(net514));
 sg13g2_buf_1 fanout515 (.A(_0416_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(net520),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(net520),
    .X(net518));
 sg13g2_buf_1 fanout519 (.A(net520),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_2026_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_1854_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(net523),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(net524),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_1829_),
    .X(net524));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(_0567_));
 sg13g2_buf_2 fanout526 (.A(_0567_),
    .X(net526));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(_0486_));
 sg13g2_buf_2 fanout528 (.A(_0486_),
    .X(net528));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(_0471_));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(_0471_));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(_0469_));
 sg13g2_buf_2 fanout532 (.A(_0469_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_0441_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_0441_),
    .X(net534));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(net537));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net537));
 sg13g2_buf_2 fanout537 (.A(_0434_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(net539),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_0433_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_0433_),
    .X(net540));
 sg13g2_buf_1 fanout541 (.A(_0433_),
    .X(net541));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_1960_));
 sg13g2_buf_2 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_1905_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_1905_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_0023_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net827),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(\top.step_size[3] ),
    .X(net549));
 sg13g2_buf_1 fanout550 (.A(\top.step_size[3] ),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(\top.step_size[2] ),
    .X(net551));
 sg13g2_buf_1 fanout552 (.A(\top.step_size[2] ),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(\top.step_size[1] ),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(\top.step_size[1] ),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(\top.step_size[0] ),
    .X(net555));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(net849));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(net846));
 sg13g2_buf_2 fanout558 (.A(\top.rs.x[4] ),
    .X(net558));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(net847));
 sg13g2_buf_2 fanout560 (.A(\top.early_x[2] ),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net565),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net565),
    .X(net563));
 sg13g2_buf_1 fanout564 (.A(net565),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(\top.julia_calc.write_mode_data ),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(\top.julia_calc.iter_done_reg ),
    .X(net566));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(net568));
 sg13g2_buf_2 fanout568 (.A(\top.julia_calc.iter_done_reg ),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(net571),
    .X(net569));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(net572));
 sg13g2_buf_1 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(\top.julia_calc.phase[0] ));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(net576));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(net575));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net576));
 sg13g2_buf_1 fanout576 (.A(_1836_),
    .X(net576));
 sg13g2_buf_4 fanout577 (.X(net577),
    .A(rst_n));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(rst_n));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[6]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[7]),
    .X(net9));
 sg13g2_tielo tt_um_toivoh_pio_ram_emu_example_10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_20_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_21_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\rx_pins[1] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold2 (.A(\top.receiver.data[2] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold3 (.A(\top.receiver.data[3] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold4 (.A(\top.receiver.data[10] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold5 (.A(\top.receiver.data[12] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold6 (.A(\top.receiver.data[7] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold7 (.A(\top.receiver.data[13] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0061_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold9 (.A(\top.receiver.data[4] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold10 (.A(\rx_pins[0] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold11 (.A(\top.receiver.data[8] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold12 (.A(\top.receiver.data[6] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold13 (.A(\top.receiver.data[5] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold14 (.A(\top.receiver.data[11] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0060_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0254_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold17 (.A(\top.receiver.data[9] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0063_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0066_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0062_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold21 (.A(\top.julia_calc.z_x[8] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0280_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold23 (.A(\top.julia_calc.z_x[4] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0276_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold25 (.A(\top.julia_calc.z_x[7] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0279_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold27 (.A(\top.julia_calc.new_pixel_group1 ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0415_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold29 (.A(\top.julia_calc.z_x[3] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0275_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold31 (.A(\top.julia_calc.z_y[6] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0287_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold33 (.A(\top.julia_calc.z_y[8] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold34 (.A(\top.julia_calc.z_x[6] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0278_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold36 (.A(\top.julia_calc.z_x[2] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold37 (.A(\top.julia_calc.z_y[1] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0428_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold39 (.A(\top.julia_calc.z_x[1] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0422_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold41 (.A(\top.transmitter.transmitter.tx_sreg[16] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0006_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold43 (.A(\top.julia_calc.z_y[2] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0109_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold45 (.A(\top.transmitter.transmitter.tx_sreg[10] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0018_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold47 (.A(\top.debouncer_inst.timer[14] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0403_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0096_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold50 (.A(\top.transmitter.transmitter.tx_sreg[1] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold51 (.A(\top.debouncer_inst.timer[8] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0393_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0090_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold54 (.A(\top.julia_calc.z_y[0] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0426_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold56 (.A(\top.julia_calc.z_y[7] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0288_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold58 (.A(\top.julia_calc.z_x[0] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0420_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold60 (.A(\top.transmitter.transmitter.tx_sreg[0] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold61 (.A(\top.julia_calc.iter[8] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold62 (.A(_1457_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold63 (.A(\top.debouncer_inst.timer[3] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0385_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0085_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold66 (.A(\top.debouncer_inst.timer[0] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0380_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0082_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold69 (.A(\top.julia_calc.z_y[3] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0284_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold71 (.A(\top.julia_calc.z_x[5] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0277_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold73 (.A(\top.pixel_buffer[0][0] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0259_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold75 (.A(\top.transmitter.transmitter.tx_sreg[15] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0005_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold77 (.A(\top.debouncer_inst.timer[16] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0407_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0098_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold80 (.A(\top.debouncer_inst.timer[5] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0388_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0087_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold83 (.A(\top.transmitter.transmitter.tx_sreg[7] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0015_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold85 (.A(\top.julia_calc.z_y[4] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0285_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold87 (.A(\top.transmitter.transmitter.tx_sreg[6] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0014_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold89 (.A(\top.debouncer_inst.timer[10] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0396_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0092_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold92 (.A(\top.last_stable_buttons[0] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0189_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold94 (.A(\top.transmitter.transmitter.tx_sreg[19] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0009_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold96 (.A(\top.julia_calc.z_y[11] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0292_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold98 (.A(\top.transmitter.transmitter.tx_sreg[11] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold99 (.A(\top.julia_calc.z_x[11] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0283_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold101 (.A(\top.julia_calc.z_y[9] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0290_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold103 (.A(\top.transmitter.transmitter.tx_sreg[17] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0007_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold105 (.A(\top.transmitter.transmitter.tx_sreg[14] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0004_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold107 (.A(\top.transmitter.transmitter.tx_sreg[4] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0012_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold109 (.A(\top.transmitter.transmitter.tx_sreg[3] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold110 (.A(\top.pixel_buffer[12][0] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold111 (.A(\top.pixel_buffer[7][1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold112 (.A(\top.pixel_buffer[5][1] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold113 (.A(\top.transmitter.transmitter.tx_sreg[2] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0001_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold115 (.A(\top.julia_calc.z_x[10] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0282_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold117 (.A(\top.julia_calc.z_y[10] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0291_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold119 (.A(\top.debouncer_inst.timer[1] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold120 (.A(\top.pixel_buffer[12][1] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold121 (.A(\top.pixel_buffer[15][0] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold122 (.A(\top.pixel_buffer[11][0] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold123 (.A(\top.pixel_buffer[10][1] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold124 (.A(\top.pixel_buffer[2][1] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold125 (.A(\top.pixel_buffer[0][1] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0260_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold127 (.A(\top.last_stable_buttons[2] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0191_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold129 (.A(\top.pixel_buffer[13][0] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold130 (.A(\top.julia_calc.far_outside_reg ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0076_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold132 (.A(\top.pixel_buffer[3][1] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold133 (.A(\top.transmitter.transmitter.tx_sreg[5] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold134 (.A(\top.julia_calc.w_addr[8] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0223_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold136 (.A(\top.julia_calc.z_x[9] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0281_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold138 (.A(\top.pixel_buffer[6][1] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold139 (.A(\top.pixel_buffer[11][1] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold140 (.A(\top.pixel_buffer[4][1] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold141 (.A(\top.transmitter.transmitter.tx_sreg[18] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0008_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold143 (.A(\top.pixel_buffer[4][0] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold144 (.A(\top.pixel_buffer[5][0] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold145 (.A(\top.julia_calc.z_y2[12] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold146 (.A(\top.pixel_buffer[13][1] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold147 (.A(\top.debouncer_inst.timer[6] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0390_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold149 (.A(\top.pixel_buffer[14][1] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold150 (.A(\top.julia_calc.z_xy[11] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold151 (.A(\top.julia_calc.w_addr[10] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0225_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold153 (.A(\top.julia_calc.w_addr[5] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0220_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold155 (.A(\top.transmitter.transmitter.tx_sreg[8] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold156 (.A(\top.transmitter.transmitter.tx_sreg[12] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0002_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold158 (.A(\top.pixel_buffer[3][0] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold159 (.A(\top.julia_calc.dest_y[8] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold160 (.A(\top.julia_calc.pixel_sreg[0] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0110_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold162 (.A(\top.pixel_buffer[14][0] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold163 (.A(\top.julia_calc.w_addr[14] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold164 (.A(\top.julia_calc.w_addr[1] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0216_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold166 (.A(\top.julia_calc.write_addr_available ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0102_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold168 (.A(\top.pixel_buffer[15][1] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold169 (.A(\top.pixel_buffer[7][0] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold170 (.A(\top.julia_calc.w_addr[12] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0227_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold172 (.A(\top.julia_calc.z_xy[9] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold173 (.A(\top.pixel_buffer[6][0] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold174 (.A(\top.julia_calc.z_xy[10] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold175 (.A(\top.transmitter.transmitter.tx_sreg[9] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0017_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold177 (.A(\top.receiver.receiver.counter[3] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0176_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold179 (.A(\top.julia_calc.pixel_sreg[12] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0122_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold181 (.A(\top.debouncer_inst.timer[17] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0409_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold183 (.A(\top.debouncer_inst.timer[11] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0398_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold185 (.A(\top.julia_calc.pixel_sreg[10] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0118_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold187 (.A(\top.debouncer_inst.timer[12] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold188 (.A(\top.julia_calc.pixel_sreg[11] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0121_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold190 (.A(\top.julia_calc.pixel_sreg[6] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0114_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold192 (.A(\top.julia_calc.pixel_sreg[14] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0124_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold194 (.A(\top.julia_calc.w_addr[0] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0215_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold196 (.A(\top.julia_calc.z_xy[1] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold197 (.A(\top.julia_calc.dest_x[2] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold198 (.A(_2036_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold199 (.A(\top.julia_calc.z_x2[12] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold200 (.A(\top.julia_calc.w_addr[3] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0218_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold202 (.A(\top.pixel_buffer[1][1] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold203 (.A(\top.julia_calc.iter[4] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold204 (.A(_1446_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0168_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold206 (.A(\top.julia_calc.w_addr[6] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0221_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold208 (.A(\top.julia_calc.w_addr[13] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0228_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold210 (.A(\top.julia_calc.w_addr[7] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0222_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold212 (.A(\top.receiver.data[1] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0200_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold214 (.A(\top.pixel_buffer[9][1] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold215 (.A(\top.debouncer_inst.timer[2] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold216 (.A(\top.pixel_buffer[10][0] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold217 (.A(\top.julia_calc.w_addr[9] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0224_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold219 (.A(\top.julia_calc.w_addr[2] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0217_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold221 (.A(\top.julia_calc.pixel_sreg[7] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0117_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold223 (.A(\top.julia_calc.pixel_sreg[8] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold224 (.A(\top.debouncer_inst.timer[18] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0413_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold226 (.A(\top.receiver.data[0] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0199_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold228 (.A(\top.julia_calc.pixel_sreg[1] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0111_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold230 (.A(\top.last_stable_buttons[3] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0192_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold232 (.A(\top.pixel_buffer[2][0] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold233 (.A(\top.julia_calc.dest_y[2] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold234 (.A(_1796_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold235 (.A(\top.julia_calc.z_y2[7] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold236 (.A(\top.pixel_buffer[1][0] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold237 (.A(\top.julia_calc.pixel_sreg[13] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0123_),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold239 (.A(\top.julia_calc.z_y2[1] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold240 (.A(\top.julia_calc.iter[2] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold241 (.A(_1443_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold242 (.A(\top.julia_calc.iter[1] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold243 (.A(_1442_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0165_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold245 (.A(\top.debouncer_inst.timer[13] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold246 (.A(\top.julia_calc.pixel_sreg[3] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0113_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold248 (.A(\top.julia_calc.pixel_sreg[2] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0112_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold250 (.A(\top.debouncer_inst.timer[9] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0395_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold252 (.A(\top.julia_calc.w_addr[4] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0219_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold254 (.A(\top.julia_calc.z_xy[7] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold255 (.A(\top.next_read_addr[13] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold256 (.A(_1824_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold257 (.A(\top.julia_calc.iter[5] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold258 (.A(_1448_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold259 (.A(\top.julia_calc.z_xy[2] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold260 (.A(\top.last_stable_buttons[1] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0190_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold262 (.A(\top.last_stable_buttons[5] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0194_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold264 (.A(\top.pixel_buffer[9][0] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold265 (.A(\top.julia_calc.pixel_sreg[5] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0054_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0022_),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold268 (.A(\top.julia_calc.w_addr[11] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0226_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold270 (.A(\top.julia_calc.z_xy[8] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold271 (.A(\top.julia_calc.dest_x[3] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold272 (.A(\top.julia_calc.iter[6] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold273 (.A(\top.debouncer_inst.timer[15] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold274 (.A(\top.julia_calc.z_x2[7] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0000_),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold276 (.A(\top.julia_calc.z_x2[3] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold277 (.A(\top.last_stable_buttons[4] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0193_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold279 (.A(\top.rs.x[11] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold280 (.A(\top.julia_calc.z_xy[5] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold281 (.A(_1432_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0157_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold283 (.A(\top.julia_calc.pixel_sreg[9] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold284 (.A(\top.julia_calc.dest_y[7] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold285 (.A(_1803_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold286 (.A(\top.julia_calc.z_y2[11] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold287 (.A(\top.julia_calc.iter[0] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold288 (.A(\top.julia_calc.z_xy[4] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold289 (.A(_1431_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0156_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold291 (.A(\top.receiver.receiver.counter[1] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold292 (.A(_1463_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold293 (.A(\top.julia_calc.z_y2[8] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold294 (.A(\top.julia_calc.z_y2[9] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold295 (.A(\top.debouncer_inst.timer[7] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold296 (.A(\top.early_x[1] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold297 (.A(_1879_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0178_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold299 (.A(\top.julia_calc.z_xy[0] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold300 (.A(\top.julia_calc.dest_x[8] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold301 (.A(_2046_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold302 (.A(\top.julia_calc.z_x2[10] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold303 (.A(\top.julia_calc.z_y2[10] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold304 (.A(\top.julia_calc.z_xy[6] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold305 (.A(\top.julia_calc.z_x2[1] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold306 (.A(\top.c_y[0] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold307 (.A(_1533_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold308 (.A(\top.transmitter.transmitter.tx_sreg[13] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0003_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold310 (.A(\top.julia_calc.iter[7] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold311 (.A(\top.julia_calc.z_y2[3] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold312 (.A(\top.julia_calc.z_y2[5] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold313 (.A(\top.julia_calc.z_xy[3] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold314 (.A(\top.julia_calc.dest_y[0] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold315 (.A(_1786_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold316 (.A(\top.julia_calc.pixel_sreg[15] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold317 (.A(\top.julia_calc.z_y2[4] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold318 (.A(\top.next_read_addr[14] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold319 (.A(\uo_out0[3] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold320 (.A(\top.julia_calc.z_y[5] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold321 (.A(\top.julia_calc.z_x2[0] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold322 (.A(\top.julia_calc.z_y2[2] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold323 (.A(\top.julia_calc.z_x2[5] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0020_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold325 (.A(_1800_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0058_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold327 (.A(_1900_),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold328 (.A(\uo_out0[7] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold329 (.A(\top.julia_calc.z_x2[8] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold330 (.A(\top.transmitter.transmitter.tx_sreg[20] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold331 (.A(\top.julia_calc.dest_y[1] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold332 (.A(_1789_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold333 (.A(\top.julia_calc.z_x2[6] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold334 (.A(\top.julia_calc.z_x2[2] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold335 (.A(\top.julia_calc.iter[3] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold336 (.A(\top.julia_calc.z_y2[0] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold337 (.A(\top.debouncer_inst.timer[4] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold338 (.A(\top.julia_calc.z_x2[9] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold339 (.A(\top.julia_calc.z_x2[11] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold340 (.A(\top.rs.x[6] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold341 (.A(\top.rs.x[7] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold342 (.A(\top.julia_calc.z_x2[4] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold343 (.A(\top.julia_calc.z_y2[6] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold344 (.A(\top.rs.y[9] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold345 (.A(\top.next_read_addr[11] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold346 (.A(_1821_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold347 (.A(\top.next_read_addr[10] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold348 (.A(_1819_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold349 (.A(\top.julia_calc.dest_x[4] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold350 (.A(\top.next_read_addr[6] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold351 (.A(_1810_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold352 (.A(\top.transmitter.transmitter.counter[1] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold353 (.A(_1696_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold354 (.A(\top.next_read_addr[9] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold355 (.A(_1817_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold356 (.A(\top.next_read_addr[8] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold357 (.A(_1815_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0306_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold359 (.A(\top.c_x[0] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold360 (.A(_1617_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold361 (.A(\top.next_read_addr[7] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0023_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0198_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold364 (.A(\top.next_read_addr[12] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold365 (.A(_1823_),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold366 (.A(\top.julia_calc.dest_y[6] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold367 (.A(_1802_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold368 (.A(\top.transmitter.transmitter.counter[3] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold369 (.A(_1699_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0257_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold371 (.A(\top.transmitter.transmitter.counter[2] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold372 (.A(_1697_),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold373 (.A(_1698_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0256_),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold375 (.A(\top.julia_calc.dest_x[5] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0027_),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0247_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold378 (.A(\top.julia_calc.dest_x[1] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold379 (.A(_2034_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0067_),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold381 (.A(\top.rs.x[4] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold382 (.A(\top.early_x[3] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold383 (.A(_1473_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold384 (.A(\top.rs.x[5] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold385 (.A(\top.rs.x[10] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold386 (.A(_1484_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold387 (.A(\top.julia_calc.phase[1] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold388 (.A(_2025_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0065_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold390 (.A(\top.julia_calc.dest_x[7] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold391 (.A(_2045_),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold392 (.A(\top.receiver.receiver.counter[2] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold393 (.A(_1464_),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0175_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold395 (.A(\top.julia_calc.write_data_available ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold396 (.A(_2024_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0028_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold398 (.A(\top.c_y[11] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0241_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold400 (.A(\top.julia_calc.dest_x[6] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold401 (.A(_2043_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0029_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold403 (.A(\top.julia_calc.dest_y[3] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0025_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold405 (.A(\top.c_y[6] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold406 (.A(\top.early_x[0] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0179_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold408 (.A(\top.c_x[11] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold409 (.A(\top.rs.x[8] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold410 (.A(\top.c_x[2] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold411 (.A(\top.c_x[1] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold412 (.A(\top.julia_calc.dest_y[4] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold413 (.A(\top.c_x[9] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0251_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold415 (.A(\top.rs.x[9] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0026_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold417 (.A(\top.c_x[8] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0027_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold419 (.A(\top.receiver.receiver.counter[2] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold420 (.A(\top.next_read_addr[8] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold421 (.A(\top.julia_calc.pixel_sreg[2] ),
    .X(net886));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_4 FILLER_0_210 ();
 sg13g2_fill_2 FILLER_0_214 ();
 sg13g2_fill_1 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_4 FILLER_0_245 ();
 sg13g2_fill_1 FILLER_0_249 ();
 sg13g2_fill_2 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_fill_1 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_fill_2 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_235 ();
 sg13g2_fill_1 FILLER_1_242 ();
 sg13g2_decap_4 FILLER_1_288 ();
 sg13g2_fill_2 FILLER_1_292 ();
 sg13g2_decap_8 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_decap_8 FILLER_1_331 ();
 sg13g2_decap_4 FILLER_1_346 ();
 sg13g2_fill_2 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_4 FILLER_2_189 ();
 sg13g2_fill_2 FILLER_2_193 ();
 sg13g2_fill_1 FILLER_2_239 ();
 sg13g2_fill_2 FILLER_2_321 ();
 sg13g2_fill_1 FILLER_2_323 ();
 sg13g2_fill_1 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_fill_2 FILLER_3_211 ();
 sg13g2_fill_1 FILLER_3_233 ();
 sg13g2_fill_1 FILLER_3_239 ();
 sg13g2_fill_1 FILLER_3_255 ();
 sg13g2_fill_2 FILLER_3_264 ();
 sg13g2_fill_1 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_286 ();
 sg13g2_fill_1 FILLER_3_318 ();
 sg13g2_fill_1 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_fill_2 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_257 ();
 sg13g2_decap_8 FILLER_4_264 ();
 sg13g2_fill_2 FILLER_4_271 ();
 sg13g2_fill_2 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_fill_2 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_fill_2 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_209 ();
 sg13g2_decap_8 FILLER_5_216 ();
 sg13g2_decap_4 FILLER_5_223 ();
 sg13g2_fill_1 FILLER_5_227 ();
 sg13g2_fill_2 FILLER_5_244 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_fill_2 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_293 ();
 sg13g2_decap_4 FILLER_5_300 ();
 sg13g2_fill_2 FILLER_5_308 ();
 sg13g2_fill_1 FILLER_5_310 ();
 sg13g2_fill_2 FILLER_5_316 ();
 sg13g2_fill_1 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_4 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_fill_2 FILLER_5_367 ();
 sg13g2_fill_1 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_196 ();
 sg13g2_fill_1 FILLER_6_217 ();
 sg13g2_fill_1 FILLER_6_251 ();
 sg13g2_fill_1 FILLER_6_272 ();
 sg13g2_decap_4 FILLER_6_278 ();
 sg13g2_fill_2 FILLER_6_282 ();
 sg13g2_fill_1 FILLER_6_293 ();
 sg13g2_decap_8 FILLER_6_327 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_decap_4 FILLER_6_341 ();
 sg13g2_fill_2 FILLER_6_345 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_fill_1 FILLER_7_220 ();
 sg13g2_fill_1 FILLER_7_249 ();
 sg13g2_fill_2 FILLER_7_262 ();
 sg13g2_fill_2 FILLER_7_294 ();
 sg13g2_fill_2 FILLER_7_337 ();
 sg13g2_decap_4 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_189 ();
 sg13g2_fill_1 FILLER_8_191 ();
 sg13g2_fill_2 FILLER_8_208 ();
 sg13g2_fill_1 FILLER_8_223 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_4 FILLER_8_263 ();
 sg13g2_fill_2 FILLER_8_267 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_1 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_fill_2 FILLER_9_228 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_decap_8 FILLER_9_244 ();
 sg13g2_decap_8 FILLER_9_251 ();
 sg13g2_fill_1 FILLER_9_258 ();
 sg13g2_fill_2 FILLER_9_264 ();
 sg13g2_fill_1 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_291 ();
 sg13g2_decap_4 FILLER_9_297 ();
 sg13g2_decap_4 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_311 ();
 sg13g2_fill_2 FILLER_9_350 ();
 sg13g2_fill_1 FILLER_9_352 ();
 sg13g2_fill_2 FILLER_9_362 ();
 sg13g2_decap_4 FILLER_9_372 ();
 sg13g2_decap_4 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_4 FILLER_10_56 ();
 sg13g2_fill_2 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_4 FILLER_10_140 ();
 sg13g2_fill_1 FILLER_10_144 ();
 sg13g2_decap_4 FILLER_10_149 ();
 sg13g2_fill_2 FILLER_10_166 ();
 sg13g2_fill_1 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_173 ();
 sg13g2_decap_8 FILLER_10_180 ();
 sg13g2_decap_8 FILLER_10_187 ();
 sg13g2_decap_8 FILLER_10_194 ();
 sg13g2_decap_8 FILLER_10_201 ();
 sg13g2_decap_8 FILLER_10_208 ();
 sg13g2_decap_4 FILLER_10_215 ();
 sg13g2_decap_4 FILLER_10_223 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_decap_4 FILLER_10_288 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_decap_4 FILLER_10_311 ();
 sg13g2_fill_1 FILLER_10_320 ();
 sg13g2_decap_4 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_4 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_fill_2 FILLER_10_379 ();
 sg13g2_fill_1 FILLER_10_381 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_4 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_46 ();
 sg13g2_decap_4 FILLER_11_51 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_95 ();
 sg13g2_decap_4 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_fill_1 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_131 ();
 sg13g2_fill_2 FILLER_11_138 ();
 sg13g2_fill_2 FILLER_11_158 ();
 sg13g2_fill_1 FILLER_11_160 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_176 ();
 sg13g2_decap_4 FILLER_11_185 ();
 sg13g2_fill_2 FILLER_11_189 ();
 sg13g2_fill_2 FILLER_11_204 ();
 sg13g2_fill_1 FILLER_11_206 ();
 sg13g2_fill_2 FILLER_11_214 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_fill_2 FILLER_11_309 ();
 sg13g2_fill_1 FILLER_11_321 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_4 FILLER_11_374 ();
 sg13g2_fill_1 FILLER_11_383 ();
 sg13g2_fill_2 FILLER_11_390 ();
 sg13g2_fill_1 FILLER_11_392 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_4 FILLER_12_28 ();
 sg13g2_fill_2 FILLER_12_32 ();
 sg13g2_fill_2 FILLER_12_60 ();
 sg13g2_fill_1 FILLER_12_62 ();
 sg13g2_fill_2 FILLER_12_93 ();
 sg13g2_fill_2 FILLER_12_125 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_202 ();
 sg13g2_fill_1 FILLER_12_241 ();
 sg13g2_fill_2 FILLER_12_261 ();
 sg13g2_fill_2 FILLER_12_270 ();
 sg13g2_fill_2 FILLER_12_305 ();
 sg13g2_fill_1 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_4 FILLER_12_327 ();
 sg13g2_fill_2 FILLER_12_331 ();
 sg13g2_fill_2 FILLER_12_351 ();
 sg13g2_fill_1 FILLER_12_353 ();
 sg13g2_fill_1 FILLER_12_376 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_21 ();
 sg13g2_fill_1 FILLER_13_62 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_208 ();
 sg13g2_fill_2 FILLER_13_218 ();
 sg13g2_fill_1 FILLER_13_220 ();
 sg13g2_fill_1 FILLER_13_234 ();
 sg13g2_fill_2 FILLER_13_247 ();
 sg13g2_fill_1 FILLER_13_254 ();
 sg13g2_decap_4 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_decap_4 FILLER_13_302 ();
 sg13g2_decap_8 FILLER_13_321 ();
 sg13g2_fill_1 FILLER_13_328 ();
 sg13g2_decap_4 FILLER_13_346 ();
 sg13g2_fill_1 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_18 ();
 sg13g2_fill_2 FILLER_14_51 ();
 sg13g2_fill_2 FILLER_14_79 ();
 sg13g2_fill_2 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_122 ();
 sg13g2_fill_2 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_fill_2 FILLER_14_193 ();
 sg13g2_fill_1 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_decap_4 FILLER_14_242 ();
 sg13g2_fill_1 FILLER_14_246 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_4 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_299 ();
 sg13g2_fill_2 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_fill_2 FILLER_14_350 ();
 sg13g2_fill_1 FILLER_14_352 ();
 sg13g2_fill_2 FILLER_14_370 ();
 sg13g2_decap_4 FILLER_14_377 ();
 sg13g2_fill_1 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_45 ();
 sg13g2_fill_1 FILLER_15_79 ();
 sg13g2_fill_1 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_116 ();
 sg13g2_fill_2 FILLER_15_135 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_decap_8 FILLER_15_272 ();
 sg13g2_decap_8 FILLER_15_279 ();
 sg13g2_decap_4 FILLER_15_286 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_decap_4 FILLER_15_307 ();
 sg13g2_fill_2 FILLER_15_311 ();
 sg13g2_fill_2 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_decap_4 FILLER_15_338 ();
 sg13g2_decap_4 FILLER_15_364 ();
 sg13g2_fill_2 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_4 FILLER_15_387 ();
 sg13g2_fill_2 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_1 FILLER_16_54 ();
 sg13g2_fill_2 FILLER_16_96 ();
 sg13g2_fill_1 FILLER_16_98 ();
 sg13g2_fill_1 FILLER_16_179 ();
 sg13g2_fill_2 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_199 ();
 sg13g2_fill_2 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_286 ();
 sg13g2_decap_4 FILLER_16_304 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_decap_4 FILLER_16_335 ();
 sg13g2_decap_4 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_347 ();
 sg13g2_decap_4 FILLER_16_374 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_2 FILLER_17_65 ();
 sg13g2_fill_2 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_221 ();
 sg13g2_fill_2 FILLER_17_250 ();
 sg13g2_fill_1 FILLER_17_252 ();
 sg13g2_fill_2 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_317 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_fill_2 FILLER_17_332 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_decap_4 FILLER_17_377 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_fill_1 FILLER_18_193 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_decap_8 FILLER_18_213 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_255 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_fill_2 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_decap_4 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_fill_2 FILLER_18_377 ();
 sg13g2_fill_1 FILLER_18_379 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_46 ();
 sg13g2_fill_2 FILLER_19_67 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_fill_2 FILLER_19_79 ();
 sg13g2_fill_1 FILLER_19_118 ();
 sg13g2_fill_2 FILLER_19_138 ();
 sg13g2_fill_2 FILLER_19_166 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_206 ();
 sg13g2_decap_8 FILLER_19_213 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_decap_4 FILLER_19_248 ();
 sg13g2_fill_2 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_fill_1 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_354 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_fill_2 FILLER_19_383 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_30 ();
 sg13g2_fill_1 FILLER_20_32 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_fill_2 FILLER_20_50 ();
 sg13g2_fill_2 FILLER_20_141 ();
 sg13g2_fill_1 FILLER_20_143 ();
 sg13g2_fill_1 FILLER_20_179 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_decap_4 FILLER_20_202 ();
 sg13g2_decap_4 FILLER_20_214 ();
 sg13g2_decap_4 FILLER_20_230 ();
 sg13g2_decap_8 FILLER_20_267 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_1 FILLER_20_294 ();
 sg13g2_fill_1 FILLER_20_323 ();
 sg13g2_fill_2 FILLER_20_361 ();
 sg13g2_decap_4 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_fill_1 FILLER_20_396 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_fill_1 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_55 ();
 sg13g2_fill_2 FILLER_21_74 ();
 sg13g2_fill_1 FILLER_21_76 ();
 sg13g2_fill_2 FILLER_21_97 ();
 sg13g2_fill_1 FILLER_21_155 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_195 ();
 sg13g2_fill_2 FILLER_21_202 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_2 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_357 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_fill_2 FILLER_21_390 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_1 FILLER_22_135 ();
 sg13g2_fill_2 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_191 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_decap_4 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_213 ();
 sg13g2_fill_2 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_237 ();
 sg13g2_fill_1 FILLER_22_244 ();
 sg13g2_decap_8 FILLER_22_267 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_fill_2 FILLER_22_313 ();
 sg13g2_decap_4 FILLER_22_322 ();
 sg13g2_fill_1 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_fill_2 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_54 ();
 sg13g2_fill_2 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_decap_4 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_fill_1 FILLER_23_258 ();
 sg13g2_fill_2 FILLER_23_272 ();
 sg13g2_decap_8 FILLER_23_286 ();
 sg13g2_fill_2 FILLER_23_293 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_fill_2 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_decap_4 FILLER_23_334 ();
 sg13g2_fill_1 FILLER_23_338 ();
 sg13g2_decap_4 FILLER_23_369 ();
 sg13g2_fill_1 FILLER_23_388 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_1 FILLER_24_76 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_1 FILLER_24_89 ();
 sg13g2_fill_2 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_121 ();
 sg13g2_fill_1 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_241 ();
 sg13g2_decap_8 FILLER_24_248 ();
 sg13g2_decap_8 FILLER_24_255 ();
 sg13g2_decap_8 FILLER_24_272 ();
 sg13g2_decap_4 FILLER_24_279 ();
 sg13g2_fill_2 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_decap_4 FILLER_24_298 ();
 sg13g2_decap_4 FILLER_24_319 ();
 sg13g2_fill_1 FILLER_24_323 ();
 sg13g2_decap_4 FILLER_24_341 ();
 sg13g2_fill_2 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_fill_2 FILLER_24_359 ();
 sg13g2_fill_1 FILLER_24_361 ();
 sg13g2_fill_1 FILLER_24_384 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_2 FILLER_25_26 ();
 sg13g2_fill_2 FILLER_25_56 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_fill_2 FILLER_25_114 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_fill_2 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_299 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_decap_4 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_1 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_4 FILLER_25_387 ();
 sg13g2_fill_1 FILLER_25_396 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_2 FILLER_26_67 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_fill_1 FILLER_26_86 ();
 sg13g2_fill_1 FILLER_26_107 ();
 sg13g2_fill_2 FILLER_26_144 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_decap_4 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_334 ();
 sg13g2_fill_1 FILLER_26_336 ();
 sg13g2_fill_2 FILLER_26_372 ();
 sg13g2_fill_1 FILLER_26_374 ();
 sg13g2_decap_4 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_fill_1 FILLER_27_44 ();
 sg13g2_fill_2 FILLER_27_59 ();
 sg13g2_fill_1 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_103 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_180 ();
 sg13g2_fill_2 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_218 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_351 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_fill_2 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_fill_2 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_118 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_decap_4 FILLER_28_181 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_fill_2 FILLER_28_237 ();
 sg13g2_fill_1 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_fill_2 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_fill_2 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_fill_1 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_fill_2 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_fill_2 FILLER_29_86 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_156 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_207 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_244 ();
 sg13g2_decap_8 FILLER_29_251 ();
 sg13g2_decap_4 FILLER_29_258 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_4 FILLER_29_273 ();
 sg13g2_decap_4 FILLER_29_287 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_decap_8 FILLER_29_310 ();
 sg13g2_fill_2 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_325 ();
 sg13g2_decap_4 FILLER_29_335 ();
 sg13g2_decap_4 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_4 FILLER_29_383 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_decap_4 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_decap_4 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_fill_2 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_4 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_decap_4 FILLER_30_387 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_fill_2 FILLER_31_52 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_151 ();
 sg13g2_decap_8 FILLER_31_222 ();
 sg13g2_decap_4 FILLER_31_229 ();
 sg13g2_fill_2 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_4 FILLER_31_343 ();
 sg13g2_fill_2 FILLER_31_359 ();
 sg13g2_fill_2 FILLER_31_393 ();
 sg13g2_fill_1 FILLER_31_395 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_73 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_122 ();
 sg13g2_fill_2 FILLER_32_155 ();
 sg13g2_fill_1 FILLER_32_157 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_293 ();
 sg13g2_decap_4 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_fill_1 FILLER_32_373 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_18 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_fill_1 FILLER_33_146 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_196 ();
 sg13g2_decap_4 FILLER_33_233 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_272 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_311 ();
 sg13g2_fill_2 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_383 ();
 sg13g2_decap_4 FILLER_33_393 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_1 FILLER_34_26 ();
 sg13g2_fill_2 FILLER_34_66 ();
 sg13g2_fill_1 FILLER_34_68 ();
 sg13g2_fill_2 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_fill_1 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_fill_2 FILLER_34_138 ();
 sg13g2_fill_2 FILLER_34_159 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_4 FILLER_34_259 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_271 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_decap_4 FILLER_34_308 ();
 sg13g2_fill_2 FILLER_34_312 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_377 ();
 sg13g2_decap_4 FILLER_34_384 ();
 sg13g2_fill_1 FILLER_34_388 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_1 FILLER_35_19 ();
 sg13g2_fill_1 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_fill_2 FILLER_35_272 ();
 sg13g2_decap_8 FILLER_35_310 ();
 sg13g2_decap_4 FILLER_35_317 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_361 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_2 FILLER_36_65 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_193 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_217 ();
 sg13g2_decap_4 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_331 ();
 sg13g2_fill_1 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_347 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_1 FILLER_37_50 ();
 sg13g2_fill_2 FILLER_37_70 ();
 sg13g2_fill_1 FILLER_37_72 ();
 sg13g2_fill_2 FILLER_37_82 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_fill_2 FILLER_37_143 ();
 sg13g2_fill_1 FILLER_37_150 ();
 sg13g2_fill_2 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_180 ();
 sg13g2_fill_2 FILLER_37_240 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_284 ();
 sg13g2_fill_1 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_4 FILLER_37_365 ();
 sg13g2_fill_2 FILLER_37_369 ();
 sg13g2_decap_4 FILLER_37_376 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_2 FILLER_38_12 ();
 sg13g2_fill_1 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_71 ();
 sg13g2_fill_2 FILLER_38_131 ();
 sg13g2_fill_1 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_180 ();
 sg13g2_fill_2 FILLER_38_199 ();
 sg13g2_fill_2 FILLER_38_209 ();
 sg13g2_decap_8 FILLER_38_225 ();
 sg13g2_decap_4 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_261 ();
 sg13g2_decap_8 FILLER_38_272 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_346 ();
 sg13g2_fill_1 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_4 FILLER_38_382 ();
 sg13g2_fill_2 FILLER_38_386 ();
 sg13g2_fill_2 FILLER_39_87 ();
 sg13g2_fill_1 FILLER_39_94 ();
 sg13g2_fill_1 FILLER_39_182 ();
 sg13g2_fill_1 FILLER_39_226 ();
 sg13g2_decap_8 FILLER_39_233 ();
 sg13g2_fill_2 FILLER_39_240 ();
 sg13g2_fill_1 FILLER_39_242 ();
 sg13g2_decap_8 FILLER_39_263 ();
 sg13g2_fill_1 FILLER_39_270 ();
 sg13g2_fill_2 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_276 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_fill_1 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_335 ();
 sg13g2_decap_8 FILLER_39_342 ();
 sg13g2_decap_8 FILLER_39_349 ();
 sg13g2_decap_8 FILLER_39_380 ();
 sg13g2_decap_8 FILLER_39_387 ();
 sg13g2_decap_8 FILLER_39_394 ();
 sg13g2_decap_8 FILLER_39_401 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_9 ();
 sg13g2_fill_2 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_16 ();
 sg13g2_fill_1 FILLER_40_25 ();
 sg13g2_fill_1 FILLER_40_39 ();
 sg13g2_fill_1 FILLER_40_111 ();
 sg13g2_fill_2 FILLER_40_122 ();
 sg13g2_fill_2 FILLER_40_142 ();
 sg13g2_fill_1 FILLER_40_144 ();
 sg13g2_fill_1 FILLER_40_176 ();
 sg13g2_fill_2 FILLER_40_234 ();
 sg13g2_fill_2 FILLER_40_275 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_1 FILLER_40_325 ();
 sg13g2_decap_8 FILLER_40_341 ();
 sg13g2_decap_4 FILLER_40_348 ();
 sg13g2_fill_1 FILLER_40_352 ();
 sg13g2_decap_4 FILLER_40_361 ();
 sg13g2_fill_1 FILLER_40_365 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_44 ();
 sg13g2_fill_2 FILLER_41_95 ();
 sg13g2_fill_1 FILLER_41_97 ();
 sg13g2_fill_1 FILLER_41_149 ();
 sg13g2_fill_2 FILLER_41_318 ();
 sg13g2_fill_2 FILLER_41_347 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_fill_2 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_398 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_26 ();
 sg13g2_fill_1 FILLER_42_57 ();
 sg13g2_fill_1 FILLER_42_93 ();
 sg13g2_fill_1 FILLER_42_108 ();
 sg13g2_fill_1 FILLER_42_123 ();
 sg13g2_fill_1 FILLER_42_213 ();
 sg13g2_fill_1 FILLER_42_219 ();
 sg13g2_fill_2 FILLER_42_229 ();
 sg13g2_fill_2 FILLER_42_295 ();
 sg13g2_fill_1 FILLER_42_324 ();
 sg13g2_fill_2 FILLER_42_350 ();
 sg13g2_decap_4 FILLER_42_367 ();
 sg13g2_fill_2 FILLER_42_376 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_2 FILLER_43_62 ();
 sg13g2_fill_1 FILLER_43_64 ();
 sg13g2_fill_1 FILLER_43_83 ();
 sg13g2_fill_1 FILLER_43_93 ();
 sg13g2_fill_2 FILLER_43_132 ();
 sg13g2_fill_1 FILLER_43_178 ();
 sg13g2_fill_2 FILLER_43_203 ();
 sg13g2_fill_1 FILLER_43_220 ();
 sg13g2_fill_1 FILLER_43_256 ();
 sg13g2_fill_1 FILLER_43_298 ();
 sg13g2_fill_2 FILLER_43_310 ();
 sg13g2_fill_1 FILLER_43_328 ();
 sg13g2_decap_8 FILLER_43_334 ();
 sg13g2_fill_1 FILLER_43_365 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_4 ();
 sg13g2_fill_1 FILLER_44_49 ();
 sg13g2_fill_2 FILLER_44_76 ();
 sg13g2_fill_2 FILLER_44_127 ();
 sg13g2_fill_1 FILLER_44_129 ();
 sg13g2_fill_1 FILLER_44_139 ();
 sg13g2_fill_1 FILLER_44_208 ();
 sg13g2_fill_1 FILLER_44_260 ();
 sg13g2_fill_2 FILLER_44_271 ();
 sg13g2_fill_2 FILLER_44_287 ();
 sg13g2_fill_1 FILLER_44_298 ();
 sg13g2_fill_2 FILLER_44_307 ();
 sg13g2_fill_1 FILLER_44_309 ();
 sg13g2_decap_8 FILLER_44_327 ();
 sg13g2_decap_8 FILLER_44_334 ();
 sg13g2_decap_8 FILLER_44_341 ();
 sg13g2_fill_1 FILLER_44_348 ();
 sg13g2_fill_2 FILLER_44_369 ();
 sg13g2_fill_1 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_388 ();
 sg13g2_decap_4 FILLER_44_395 ();
 sg13g2_fill_2 FILLER_44_399 ();
 sg13g2_fill_2 FILLER_45_26 ();
 sg13g2_fill_1 FILLER_45_28 ();
 sg13g2_fill_2 FILLER_45_74 ();
 sg13g2_fill_2 FILLER_45_93 ();
 sg13g2_fill_1 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_105 ();
 sg13g2_fill_1 FILLER_45_107 ();
 sg13g2_fill_1 FILLER_45_140 ();
 sg13g2_fill_1 FILLER_45_201 ();
 sg13g2_fill_1 FILLER_45_247 ();
 sg13g2_fill_1 FILLER_45_253 ();
 sg13g2_fill_2 FILLER_45_273 ();
 sg13g2_fill_2 FILLER_45_305 ();
 sg13g2_decap_4 FILLER_45_334 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_decap_8 FILLER_45_349 ();
 sg13g2_decap_8 FILLER_45_356 ();
 sg13g2_decap_4 FILLER_45_363 ();
 sg13g2_fill_1 FILLER_45_367 ();
 sg13g2_decap_8 FILLER_45_386 ();
 sg13g2_fill_2 FILLER_45_397 ();
 sg13g2_fill_2 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_fill_1 FILLER_46_26 ();
 sg13g2_fill_1 FILLER_46_80 ();
 sg13g2_fill_2 FILLER_46_121 ();
 sg13g2_fill_2 FILLER_46_171 ();
 sg13g2_fill_1 FILLER_46_190 ();
 sg13g2_fill_2 FILLER_46_220 ();
 sg13g2_fill_1 FILLER_46_276 ();
 sg13g2_fill_1 FILLER_46_311 ();
 sg13g2_fill_2 FILLER_46_343 ();
 sg13g2_fill_1 FILLER_46_345 ();
 sg13g2_decap_8 FILLER_46_355 ();
 sg13g2_fill_1 FILLER_46_382 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_110 ();
 sg13g2_fill_2 FILLER_47_129 ();
 sg13g2_fill_1 FILLER_47_131 ();
 sg13g2_fill_1 FILLER_47_141 ();
 sg13g2_fill_2 FILLER_47_156 ();
 sg13g2_fill_2 FILLER_47_218 ();
 sg13g2_fill_1 FILLER_47_281 ();
 sg13g2_fill_1 FILLER_47_317 ();
 sg13g2_fill_2 FILLER_47_372 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_4 ();
 sg13g2_fill_1 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_99 ();
 sg13g2_fill_1 FILLER_48_116 ();
 sg13g2_fill_1 FILLER_48_130 ();
 sg13g2_fill_1 FILLER_48_204 ();
 sg13g2_fill_2 FILLER_48_246 ();
 sg13g2_fill_1 FILLER_48_255 ();
 sg13g2_fill_1 FILLER_48_283 ();
 sg13g2_fill_1 FILLER_48_293 ();
 sg13g2_fill_2 FILLER_48_377 ();
 sg13g2_fill_2 FILLER_49_60 ();
 sg13g2_fill_1 FILLER_49_62 ();
 sg13g2_fill_2 FILLER_49_87 ();
 sg13g2_fill_1 FILLER_49_98 ();
 sg13g2_fill_2 FILLER_49_134 ();
 sg13g2_fill_1 FILLER_49_136 ();
 sg13g2_fill_1 FILLER_49_198 ();
 sg13g2_fill_1 FILLER_49_236 ();
 sg13g2_fill_2 FILLER_49_294 ();
 sg13g2_fill_2 FILLER_49_307 ();
 sg13g2_fill_2 FILLER_49_375 ();
 sg13g2_fill_2 FILLER_50_26 ();
 sg13g2_fill_1 FILLER_50_28 ();
 sg13g2_fill_1 FILLER_50_44 ();
 sg13g2_fill_1 FILLER_50_101 ();
 sg13g2_fill_1 FILLER_50_152 ();
 sg13g2_fill_2 FILLER_50_158 ();
 sg13g2_fill_1 FILLER_50_160 ();
 sg13g2_fill_2 FILLER_50_170 ();
 sg13g2_decap_4 FILLER_50_228 ();
 sg13g2_fill_2 FILLER_50_240 ();
 sg13g2_fill_2 FILLER_50_246 ();
 sg13g2_fill_1 FILLER_50_248 ();
 sg13g2_fill_2 FILLER_50_253 ();
 sg13g2_fill_1 FILLER_50_268 ();
 sg13g2_fill_2 FILLER_50_294 ();
 sg13g2_fill_1 FILLER_50_382 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_37 ();
 sg13g2_fill_2 FILLER_51_122 ();
 sg13g2_fill_2 FILLER_51_155 ();
 sg13g2_fill_1 FILLER_51_157 ();
 sg13g2_fill_1 FILLER_51_177 ();
 sg13g2_fill_1 FILLER_51_194 ();
 sg13g2_fill_2 FILLER_51_209 ();
 sg13g2_fill_1 FILLER_51_211 ();
 sg13g2_decap_8 FILLER_51_217 ();
 sg13g2_decap_8 FILLER_51_224 ();
 sg13g2_fill_2 FILLER_51_231 ();
 sg13g2_fill_1 FILLER_51_233 ();
 sg13g2_decap_8 FILLER_51_238 ();
 sg13g2_fill_1 FILLER_51_245 ();
 sg13g2_fill_2 FILLER_51_259 ();
 sg13g2_fill_1 FILLER_51_261 ();
 sg13g2_fill_1 FILLER_51_271 ();
 sg13g2_fill_2 FILLER_51_339 ();
 sg13g2_fill_1 FILLER_51_359 ();
 sg13g2_decap_4 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_47 ();
 sg13g2_fill_1 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_69 ();
 sg13g2_fill_1 FILLER_52_118 ();
 sg13g2_fill_1 FILLER_52_123 ();
 sg13g2_fill_2 FILLER_52_128 ();
 sg13g2_fill_1 FILLER_52_139 ();
 sg13g2_fill_1 FILLER_52_145 ();
 sg13g2_fill_2 FILLER_52_150 ();
 sg13g2_fill_2 FILLER_52_165 ();
 sg13g2_fill_1 FILLER_52_167 ();
 sg13g2_fill_1 FILLER_52_173 ();
 sg13g2_fill_1 FILLER_52_182 ();
 sg13g2_fill_2 FILLER_52_188 ();
 sg13g2_fill_1 FILLER_52_190 ();
 sg13g2_fill_2 FILLER_52_200 ();
 sg13g2_fill_1 FILLER_52_206 ();
 sg13g2_fill_2 FILLER_52_212 ();
 sg13g2_fill_1 FILLER_52_214 ();
 sg13g2_fill_1 FILLER_52_241 ();
 sg13g2_fill_1 FILLER_52_272 ();
 sg13g2_fill_2 FILLER_52_317 ();
 sg13g2_fill_2 FILLER_52_325 ();
 sg13g2_fill_1 FILLER_52_349 ();
 sg13g2_fill_2 FILLER_52_376 ();
 sg13g2_fill_2 FILLER_53_26 ();
 sg13g2_fill_1 FILLER_53_52 ();
 sg13g2_fill_2 FILLER_53_62 ();
 sg13g2_fill_1 FILLER_53_64 ();
 sg13g2_decap_8 FILLER_53_73 ();
 sg13g2_fill_2 FILLER_53_80 ();
 sg13g2_fill_1 FILLER_53_113 ();
 sg13g2_decap_8 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_189 ();
 sg13g2_fill_2 FILLER_53_196 ();
 sg13g2_fill_1 FILLER_53_198 ();
 sg13g2_decap_4 FILLER_53_204 ();
 sg13g2_fill_2 FILLER_53_239 ();
 sg13g2_fill_2 FILLER_53_383 ();
 sg13g2_fill_1 FILLER_53_390 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_9 ();
 sg13g2_fill_2 FILLER_54_27 ();
 sg13g2_fill_2 FILLER_54_34 ();
 sg13g2_fill_1 FILLER_54_44 ();
 sg13g2_fill_1 FILLER_54_56 ();
 sg13g2_fill_1 FILLER_54_60 ();
 sg13g2_fill_2 FILLER_54_87 ();
 sg13g2_fill_2 FILLER_54_158 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_fill_2 FILLER_54_187 ();
 sg13g2_fill_1 FILLER_54_189 ();
 sg13g2_fill_1 FILLER_54_216 ();
 sg13g2_fill_1 FILLER_54_273 ();
 sg13g2_fill_2 FILLER_54_279 ();
 sg13g2_fill_1 FILLER_54_312 ();
 sg13g2_fill_1 FILLER_54_317 ();
 sg13g2_fill_2 FILLER_54_374 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_fill_2 FILLER_55_26 ();
 sg13g2_fill_2 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_87 ();
 sg13g2_fill_2 FILLER_55_93 ();
 sg13g2_fill_2 FILLER_55_104 ();
 sg13g2_fill_1 FILLER_55_106 ();
 sg13g2_fill_2 FILLER_55_137 ();
 sg13g2_fill_2 FILLER_55_174 ();
 sg13g2_fill_1 FILLER_55_176 ();
 sg13g2_fill_2 FILLER_55_186 ();
 sg13g2_fill_1 FILLER_55_244 ();
 sg13g2_fill_2 FILLER_55_250 ();
 sg13g2_fill_1 FILLER_55_262 ();
 sg13g2_fill_1 FILLER_55_272 ();
 sg13g2_fill_1 FILLER_55_316 ();
 sg13g2_fill_2 FILLER_55_353 ();
 sg13g2_fill_1 FILLER_55_355 ();
 sg13g2_fill_2 FILLER_55_378 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_fill_2 FILLER_56_47 ();
 sg13g2_fill_1 FILLER_56_54 ();
 sg13g2_fill_2 FILLER_56_151 ();
 sg13g2_fill_1 FILLER_56_163 ();
 sg13g2_fill_1 FILLER_56_169 ();
 sg13g2_decap_8 FILLER_56_187 ();
 sg13g2_fill_1 FILLER_56_194 ();
 sg13g2_fill_1 FILLER_56_204 ();
 sg13g2_decap_4 FILLER_56_222 ();
 sg13g2_fill_2 FILLER_56_230 ();
 sg13g2_fill_2 FILLER_56_236 ();
 sg13g2_fill_1 FILLER_56_238 ();
 sg13g2_fill_2 FILLER_56_243 ();
 sg13g2_fill_2 FILLER_56_256 ();
 sg13g2_fill_1 FILLER_56_271 ();
 sg13g2_fill_2 FILLER_56_328 ();
 sg13g2_fill_2 FILLER_56_347 ();
 sg13g2_fill_1 FILLER_56_349 ();
 sg13g2_fill_2 FILLER_56_376 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_106 ();
 sg13g2_decap_8 FILLER_57_131 ();
 sg13g2_decap_4 FILLER_57_138 ();
 sg13g2_fill_1 FILLER_57_142 ();
 sg13g2_fill_2 FILLER_57_147 ();
 sg13g2_fill_1 FILLER_57_153 ();
 sg13g2_decap_4 FILLER_57_158 ();
 sg13g2_fill_2 FILLER_57_162 ();
 sg13g2_decap_8 FILLER_57_190 ();
 sg13g2_decap_8 FILLER_57_197 ();
 sg13g2_fill_2 FILLER_57_204 ();
 sg13g2_fill_1 FILLER_57_206 ();
 sg13g2_fill_2 FILLER_57_235 ();
 sg13g2_fill_2 FILLER_57_293 ();
 sg13g2_fill_1 FILLER_57_303 ();
 sg13g2_fill_2 FILLER_57_308 ();
 sg13g2_fill_1 FILLER_57_338 ();
 sg13g2_fill_2 FILLER_57_373 ();
 sg13g2_fill_2 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_50 ();
 sg13g2_fill_2 FILLER_58_73 ();
 sg13g2_fill_1 FILLER_58_75 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_91 ();
 sg13g2_fill_2 FILLER_58_101 ();
 sg13g2_fill_2 FILLER_58_113 ();
 sg13g2_decap_8 FILLER_58_124 ();
 sg13g2_decap_8 FILLER_58_131 ();
 sg13g2_decap_4 FILLER_58_138 ();
 sg13g2_fill_2 FILLER_58_159 ();
 sg13g2_fill_1 FILLER_58_161 ();
 sg13g2_fill_1 FILLER_58_197 ();
 sg13g2_fill_2 FILLER_58_203 ();
 sg13g2_fill_2 FILLER_58_227 ();
 sg13g2_fill_1 FILLER_58_240 ();
 sg13g2_fill_1 FILLER_58_282 ();
 sg13g2_fill_1 FILLER_58_306 ();
 sg13g2_fill_1 FILLER_58_333 ();
 sg13g2_fill_1 FILLER_58_370 ();
 sg13g2_fill_2 FILLER_58_397 ();
 sg13g2_fill_1 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_59_66 ();
 sg13g2_decap_4 FILLER_59_94 ();
 sg13g2_fill_2 FILLER_59_98 ();
 sg13g2_fill_2 FILLER_59_130 ();
 sg13g2_fill_2 FILLER_59_209 ();
 sg13g2_fill_1 FILLER_59_211 ();
 sg13g2_decap_8 FILLER_59_253 ();
 sg13g2_decap_8 FILLER_59_260 ();
 sg13g2_decap_8 FILLER_59_267 ();
 sg13g2_decap_4 FILLER_59_279 ();
 sg13g2_fill_1 FILLER_59_283 ();
 sg13g2_fill_2 FILLER_59_292 ();
 sg13g2_fill_1 FILLER_59_294 ();
 sg13g2_fill_2 FILLER_59_313 ();
 sg13g2_fill_2 FILLER_59_380 ();
 sg13g2_fill_1 FILLER_59_382 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_105 ();
 sg13g2_fill_1 FILLER_60_173 ();
 sg13g2_fill_2 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_decap_8 FILLER_60_245 ();
 sg13g2_decap_8 FILLER_60_252 ();
 sg13g2_decap_8 FILLER_60_259 ();
 sg13g2_decap_8 FILLER_60_266 ();
 sg13g2_fill_1 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_305 ();
 sg13g2_fill_1 FILLER_60_312 ();
 sg13g2_fill_1 FILLER_60_353 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_50 ();
 sg13g2_fill_2 FILLER_61_64 ();
 sg13g2_fill_2 FILLER_61_75 ();
 sg13g2_fill_2 FILLER_61_94 ();
 sg13g2_fill_1 FILLER_61_117 ();
 sg13g2_fill_2 FILLER_61_177 ();
 sg13g2_fill_2 FILLER_61_197 ();
 sg13g2_decap_8 FILLER_61_209 ();
 sg13g2_decap_8 FILLER_61_216 ();
 sg13g2_decap_8 FILLER_61_223 ();
 sg13g2_decap_8 FILLER_61_230 ();
 sg13g2_decap_8 FILLER_61_237 ();
 sg13g2_decap_8 FILLER_61_244 ();
 sg13g2_decap_4 FILLER_61_255 ();
 sg13g2_fill_1 FILLER_61_259 ();
 sg13g2_decap_8 FILLER_61_298 ();
 sg13g2_decap_8 FILLER_61_305 ();
 sg13g2_decap_4 FILLER_61_312 ();
 sg13g2_fill_2 FILLER_61_316 ();
 sg13g2_fill_2 FILLER_61_323 ();
 sg13g2_fill_1 FILLER_61_325 ();
 sg13g2_fill_1 FILLER_61_346 ();
 sg13g2_fill_2 FILLER_61_351 ();
 sg13g2_fill_2 FILLER_61_397 ();
 sg13g2_fill_1 FILLER_61_399 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_48 ();
 sg13g2_fill_1 FILLER_62_50 ();
 sg13g2_decap_4 FILLER_62_79 ();
 sg13g2_fill_1 FILLER_62_109 ();
 sg13g2_fill_1 FILLER_62_147 ();
 sg13g2_fill_1 FILLER_62_162 ();
 sg13g2_decap_4 FILLER_62_185 ();
 sg13g2_decap_8 FILLER_62_199 ();
 sg13g2_decap_8 FILLER_62_206 ();
 sg13g2_decap_8 FILLER_62_213 ();
 sg13g2_decap_4 FILLER_62_220 ();
 sg13g2_fill_1 FILLER_62_224 ();
 sg13g2_decap_4 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_296 ();
 sg13g2_fill_1 FILLER_62_298 ();
 sg13g2_fill_2 FILLER_62_325 ();
 sg13g2_fill_2 FILLER_62_348 ();
 sg13g2_fill_1 FILLER_62_350 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_2 ();
 sg13g2_fill_2 FILLER_63_29 ();
 sg13g2_decap_4 FILLER_63_39 ();
 sg13g2_fill_2 FILLER_63_43 ();
 sg13g2_fill_1 FILLER_63_63 ();
 sg13g2_fill_1 FILLER_63_73 ();
 sg13g2_fill_2 FILLER_63_110 ();
 sg13g2_fill_1 FILLER_63_135 ();
 sg13g2_fill_2 FILLER_63_162 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_fill_2 FILLER_63_196 ();
 sg13g2_fill_1 FILLER_63_250 ();
 sg13g2_fill_2 FILLER_63_342 ();
 sg13g2_fill_1 FILLER_63_344 ();
 sg13g2_fill_2 FILLER_63_380 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_36 ();
 sg13g2_fill_1 FILLER_64_40 ();
 sg13g2_fill_2 FILLER_64_52 ();
 sg13g2_fill_2 FILLER_64_63 ();
 sg13g2_fill_1 FILLER_64_105 ();
 sg13g2_fill_2 FILLER_64_181 ();
 sg13g2_fill_1 FILLER_64_183 ();
 sg13g2_fill_1 FILLER_64_192 ();
 sg13g2_fill_1 FILLER_64_233 ();
 sg13g2_fill_2 FILLER_64_247 ();
 sg13g2_fill_1 FILLER_64_249 ();
 sg13g2_fill_2 FILLER_64_257 ();
 sg13g2_fill_1 FILLER_64_281 ();
 sg13g2_decap_4 FILLER_64_311 ();
 sg13g2_fill_2 FILLER_64_398 ();
 sg13g2_decap_4 FILLER_65_26 ();
 sg13g2_fill_2 FILLER_65_30 ();
 sg13g2_fill_2 FILLER_65_64 ();
 sg13g2_fill_2 FILLER_65_82 ();
 sg13g2_fill_1 FILLER_65_175 ();
 sg13g2_fill_1 FILLER_65_191 ();
 sg13g2_fill_2 FILLER_65_197 ();
 sg13g2_fill_1 FILLER_65_229 ();
 sg13g2_fill_2 FILLER_65_238 ();
 sg13g2_fill_1 FILLER_65_249 ();
 sg13g2_fill_2 FILLER_65_254 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_fill_2 FILLER_65_274 ();
 sg13g2_fill_1 FILLER_65_276 ();
 sg13g2_fill_1 FILLER_65_282 ();
 sg13g2_decap_4 FILLER_65_292 ();
 sg13g2_fill_1 FILLER_65_296 ();
 sg13g2_fill_2 FILLER_65_309 ();
 sg13g2_fill_1 FILLER_65_311 ();
 sg13g2_fill_2 FILLER_65_344 ();
 sg13g2_fill_1 FILLER_65_346 ();
 sg13g2_fill_2 FILLER_65_379 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_fill_1 FILLER_66_195 ();
 sg13g2_fill_2 FILLER_66_279 ();
 sg13g2_fill_2 FILLER_66_299 ();
 sg13g2_fill_2 FILLER_66_355 ();
 sg13g2_fill_1 FILLER_66_357 ();
 sg13g2_fill_2 FILLER_66_381 ();
 sg13g2_fill_1 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_56 ();
 sg13g2_fill_1 FILLER_67_58 ();
 sg13g2_fill_2 FILLER_67_64 ();
 sg13g2_fill_1 FILLER_67_66 ();
 sg13g2_fill_2 FILLER_67_101 ();
 sg13g2_fill_1 FILLER_67_116 ();
 sg13g2_fill_1 FILLER_67_125 ();
 sg13g2_fill_1 FILLER_67_130 ();
 sg13g2_fill_2 FILLER_67_185 ();
 sg13g2_fill_2 FILLER_67_199 ();
 sg13g2_fill_1 FILLER_67_201 ();
 sg13g2_decap_4 FILLER_67_231 ();
 sg13g2_fill_2 FILLER_67_257 ();
 sg13g2_fill_1 FILLER_67_259 ();
 sg13g2_fill_2 FILLER_67_292 ();
 sg13g2_decap_4 FILLER_67_306 ();
 sg13g2_fill_2 FILLER_67_320 ();
 sg13g2_fill_1 FILLER_67_348 ();
 sg13g2_fill_2 FILLER_67_358 ();
 sg13g2_fill_2 FILLER_67_397 ();
 sg13g2_fill_1 FILLER_67_399 ();
 sg13g2_fill_1 FILLER_68_44 ();
 sg13g2_fill_2 FILLER_68_53 ();
 sg13g2_fill_2 FILLER_68_67 ();
 sg13g2_fill_2 FILLER_68_78 ();
 sg13g2_fill_2 FILLER_68_93 ();
 sg13g2_fill_2 FILLER_68_103 ();
 sg13g2_fill_1 FILLER_68_194 ();
 sg13g2_decap_8 FILLER_68_212 ();
 sg13g2_decap_4 FILLER_68_219 ();
 sg13g2_decap_8 FILLER_68_228 ();
 sg13g2_decap_8 FILLER_68_235 ();
 sg13g2_decap_8 FILLER_68_242 ();
 sg13g2_decap_4 FILLER_68_249 ();
 sg13g2_fill_2 FILLER_68_261 ();
 sg13g2_decap_4 FILLER_68_266 ();
 sg13g2_fill_1 FILLER_68_305 ();
 sg13g2_fill_1 FILLER_68_311 ();
 sg13g2_fill_1 FILLER_68_325 ();
 sg13g2_fill_2 FILLER_68_345 ();
 sg13g2_fill_2 FILLER_68_356 ();
 sg13g2_fill_1 FILLER_68_358 ();
 sg13g2_fill_1 FILLER_68_385 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_2 ();
 sg13g2_decap_8 FILLER_69_16 ();
 sg13g2_decap_8 FILLER_69_23 ();
 sg13g2_fill_1 FILLER_69_53 ();
 sg13g2_fill_2 FILLER_69_68 ();
 sg13g2_decap_4 FILLER_69_80 ();
 sg13g2_decap_4 FILLER_69_110 ();
 sg13g2_fill_1 FILLER_69_114 ();
 sg13g2_fill_2 FILLER_69_216 ();
 sg13g2_fill_1 FILLER_69_218 ();
 sg13g2_fill_2 FILLER_69_274 ();
 sg13g2_fill_1 FILLER_69_276 ();
 sg13g2_fill_1 FILLER_69_285 ();
 sg13g2_decap_4 FILLER_69_291 ();
 sg13g2_fill_2 FILLER_69_308 ();
 sg13g2_fill_1 FILLER_69_310 ();
 sg13g2_decap_4 FILLER_69_316 ();
 sg13g2_fill_1 FILLER_69_333 ();
 sg13g2_fill_2 FILLER_69_345 ();
 sg13g2_fill_2 FILLER_69_378 ();
 sg13g2_fill_1 FILLER_69_398 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_10 ();
 sg13g2_fill_2 FILLER_70_15 ();
 sg13g2_fill_1 FILLER_70_43 ();
 sg13g2_decap_4 FILLER_70_106 ();
 sg13g2_decap_4 FILLER_70_136 ();
 sg13g2_fill_2 FILLER_70_140 ();
 sg13g2_fill_2 FILLER_70_146 ();
 sg13g2_fill_1 FILLER_70_148 ();
 sg13g2_fill_2 FILLER_70_219 ();
 sg13g2_decap_4 FILLER_70_225 ();
 sg13g2_fill_1 FILLER_70_229 ();
 sg13g2_decap_8 FILLER_70_234 ();
 sg13g2_fill_2 FILLER_70_241 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_fill_2 FILLER_70_249 ();
 sg13g2_fill_1 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_282 ();
 sg13g2_decap_8 FILLER_70_289 ();
 sg13g2_decap_4 FILLER_70_296 ();
 sg13g2_fill_2 FILLER_70_300 ();
 sg13g2_fill_1 FILLER_70_328 ();
 sg13g2_fill_1 FILLER_70_347 ();
 sg13g2_fill_2 FILLER_70_356 ();
 sg13g2_fill_1 FILLER_70_358 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_fill_1 FILLER_71_40 ();
 sg13g2_fill_2 FILLER_71_88 ();
 sg13g2_fill_2 FILLER_71_103 ();
 sg13g2_decap_8 FILLER_71_113 ();
 sg13g2_fill_1 FILLER_71_120 ();
 sg13g2_decap_8 FILLER_71_125 ();
 sg13g2_decap_8 FILLER_71_132 ();
 sg13g2_decap_8 FILLER_71_139 ();
 sg13g2_decap_4 FILLER_71_146 ();
 sg13g2_fill_1 FILLER_71_150 ();
 sg13g2_fill_2 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_197 ();
 sg13g2_fill_2 FILLER_71_208 ();
 sg13g2_fill_1 FILLER_71_210 ();
 sg13g2_fill_1 FILLER_71_215 ();
 sg13g2_decap_8 FILLER_71_220 ();
 sg13g2_decap_8 FILLER_71_227 ();
 sg13g2_decap_4 FILLER_71_234 ();
 sg13g2_fill_2 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_291 ();
 sg13g2_fill_1 FILLER_71_362 ();
 sg13g2_fill_1 FILLER_71_377 ();
 sg13g2_fill_1 FILLER_72_30 ();
 sg13g2_fill_2 FILLER_72_57 ();
 sg13g2_fill_1 FILLER_72_72 ();
 sg13g2_fill_2 FILLER_72_87 ();
 sg13g2_decap_4 FILLER_72_120 ();
 sg13g2_fill_1 FILLER_72_159 ();
 sg13g2_fill_2 FILLER_72_164 ();
 sg13g2_fill_1 FILLER_72_174 ();
 sg13g2_decap_8 FILLER_72_190 ();
 sg13g2_decap_8 FILLER_72_197 ();
 sg13g2_fill_1 FILLER_72_204 ();
 sg13g2_fill_2 FILLER_72_243 ();
 sg13g2_decap_4 FILLER_72_287 ();
 sg13g2_fill_2 FILLER_72_291 ();
 sg13g2_decap_4 FILLER_72_297 ();
 sg13g2_fill_2 FILLER_72_301 ();
 sg13g2_fill_2 FILLER_72_341 ();
 sg13g2_fill_1 FILLER_72_343 ();
 sg13g2_fill_2 FILLER_72_380 ();
 sg13g2_fill_1 FILLER_72_382 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_30 ();
 sg13g2_fill_1 FILLER_73_32 ();
 sg13g2_fill_1 FILLER_73_165 ();
 sg13g2_decap_8 FILLER_73_174 ();
 sg13g2_decap_4 FILLER_73_181 ();
 sg13g2_decap_8 FILLER_73_194 ();
 sg13g2_fill_2 FILLER_73_201 ();
 sg13g2_decap_4 FILLER_73_208 ();
 sg13g2_fill_2 FILLER_73_212 ();
 sg13g2_decap_4 FILLER_73_222 ();
 sg13g2_decap_8 FILLER_73_275 ();
 sg13g2_decap_4 FILLER_73_282 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_1 FILLER_73_312 ();
 sg13g2_fill_2 FILLER_73_349 ();
 sg13g2_fill_1 FILLER_73_351 ();
 sg13g2_fill_1 FILLER_73_365 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_98 ();
 sg13g2_fill_1 FILLER_74_100 ();
 sg13g2_fill_1 FILLER_74_127 ();
 sg13g2_decap_4 FILLER_74_202 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_fill_2 FILLER_74_245 ();
 sg13g2_fill_1 FILLER_74_247 ();
 sg13g2_fill_2 FILLER_74_275 ();
 sg13g2_fill_1 FILLER_74_282 ();
 sg13g2_fill_2 FILLER_74_329 ();
 sg13g2_fill_1 FILLER_74_331 ();
 sg13g2_fill_2 FILLER_74_337 ();
 sg13g2_fill_2 FILLER_74_372 ();
 sg13g2_fill_1 FILLER_74_374 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_2 FILLER_74_398 ();
 sg13g2_fill_2 FILLER_75_31 ();
 sg13g2_fill_2 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_44 ();
 sg13g2_fill_2 FILLER_75_54 ();
 sg13g2_fill_1 FILLER_75_56 ();
 sg13g2_fill_2 FILLER_75_67 ();
 sg13g2_fill_2 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_93 ();
 sg13g2_fill_2 FILLER_75_125 ();
 sg13g2_fill_1 FILLER_75_127 ();
 sg13g2_fill_2 FILLER_75_172 ();
 sg13g2_fill_1 FILLER_75_227 ();
 sg13g2_fill_1 FILLER_75_243 ();
 sg13g2_fill_1 FILLER_75_294 ();
 sg13g2_fill_1 FILLER_75_336 ();
 sg13g2_fill_2 FILLER_75_346 ();
 sg13g2_fill_1 FILLER_75_348 ();
 sg13g2_decap_4 FILLER_75_385 ();
 sg13g2_fill_1 FILLER_75_389 ();
 sg13g2_fill_1 FILLER_75_398 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_2 ();
 sg13g2_fill_2 FILLER_76_43 ();
 sg13g2_fill_2 FILLER_76_54 ();
 sg13g2_fill_1 FILLER_76_56 ();
 sg13g2_fill_2 FILLER_76_70 ();
 sg13g2_fill_2 FILLER_76_114 ();
 sg13g2_fill_1 FILLER_76_116 ();
 sg13g2_fill_2 FILLER_76_150 ();
 sg13g2_fill_2 FILLER_76_243 ();
 sg13g2_fill_2 FILLER_76_257 ();
 sg13g2_fill_1 FILLER_76_302 ();
 sg13g2_fill_2 FILLER_76_308 ();
 sg13g2_fill_2 FILLER_76_315 ();
 sg13g2_fill_2 FILLER_76_353 ();
 sg13g2_fill_1 FILLER_76_355 ();
 sg13g2_decap_8 FILLER_76_391 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_84 ();
 sg13g2_fill_2 FILLER_77_121 ();
 sg13g2_fill_1 FILLER_77_149 ();
 sg13g2_fill_1 FILLER_77_180 ();
 sg13g2_fill_2 FILLER_77_186 ();
 sg13g2_fill_1 FILLER_77_188 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_2 FILLER_77_243 ();
 sg13g2_fill_2 FILLER_77_260 ();
 sg13g2_fill_1 FILLER_77_262 ();
 sg13g2_fill_2 FILLER_77_277 ();
 sg13g2_fill_2 FILLER_77_292 ();
 sg13g2_fill_2 FILLER_77_317 ();
 sg13g2_fill_1 FILLER_77_319 ();
 sg13g2_fill_1 FILLER_77_333 ();
 sg13g2_decap_8 FILLER_77_387 ();
 sg13g2_decap_8 FILLER_77_394 ();
 sg13g2_decap_8 FILLER_77_401 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_36 ();
 sg13g2_fill_2 FILLER_78_125 ();
 sg13g2_fill_1 FILLER_78_127 ();
 sg13g2_fill_1 FILLER_78_163 ();
 sg13g2_fill_2 FILLER_78_192 ();
 sg13g2_fill_1 FILLER_78_229 ();
 sg13g2_decap_4 FILLER_78_365 ();
 sg13g2_fill_1 FILLER_78_369 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_69 ();
 sg13g2_fill_1 FILLER_79_126 ();
 sg13g2_fill_2 FILLER_79_144 ();
 sg13g2_fill_2 FILLER_79_158 ();
 sg13g2_decap_8 FILLER_79_164 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_decap_8 FILLER_79_198 ();
 sg13g2_decap_4 FILLER_79_209 ();
 sg13g2_fill_1 FILLER_79_213 ();
 sg13g2_fill_1 FILLER_79_218 ();
 sg13g2_fill_1 FILLER_79_249 ();
 sg13g2_fill_2 FILLER_79_276 ();
 sg13g2_fill_1 FILLER_79_278 ();
 sg13g2_decap_4 FILLER_79_291 ();
 sg13g2_fill_2 FILLER_79_325 ();
 sg13g2_fill_1 FILLER_79_327 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_4 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_59 ();
 sg13g2_fill_1 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_88 ();
 sg13g2_fill_2 FILLER_80_118 ();
 sg13g2_fill_2 FILLER_80_124 ();
 sg13g2_fill_1 FILLER_80_143 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_fill_2 FILLER_80_180 ();
 sg13g2_fill_1 FILLER_80_182 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_fill_2 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_239 ();
 sg13g2_fill_2 FILLER_80_246 ();
 sg13g2_fill_2 FILLER_80_267 ();
 sg13g2_fill_1 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_274 ();
 sg13g2_decap_8 FILLER_80_287 ();
 sg13g2_decap_8 FILLER_80_294 ();
 sg13g2_decap_4 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_305 ();
 sg13g2_decap_4 FILLER_80_310 ();
 sg13g2_fill_1 FILLER_80_314 ();
 sg13g2_fill_2 FILLER_80_327 ();
 sg13g2_fill_1 FILLER_80_329 ();
 sg13g2_fill_2 FILLER_80_342 ();
 sg13g2_fill_1 FILLER_80_348 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net10;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net319;
 assign uio_oe[5] = net320;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
endmodule

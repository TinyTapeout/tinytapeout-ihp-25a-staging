module tt_um_i2c_regf (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clk_regs;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire \i2c_slave_controller.ack_recieved ;
 wire \i2c_slave_controller.addr[0] ;
 wire \i2c_slave_controller.addr[1] ;
 wire \i2c_slave_controller.addr[2] ;
 wire \i2c_slave_controller.addr[3] ;
 wire \i2c_slave_controller.addr[4] ;
 wire \i2c_slave_controller.addr[5] ;
 wire \i2c_slave_controller.addr[6] ;
 wire \i2c_slave_controller.addr[7] ;
 wire \i2c_slave_controller.counter[0] ;
 wire \i2c_slave_controller.counter[1] ;
 wire \i2c_slave_controller.counter[2] ;
 wire \i2c_slave_controller.out_regf_req ;
 wire \i2c_slave_controller.out_regf_rw ;
 wire \i2c_slave_controller.out_regf_write_data[0] ;
 wire \i2c_slave_controller.out_regf_write_data[1] ;
 wire \i2c_slave_controller.out_regf_write_data[2] ;
 wire \i2c_slave_controller.out_regf_write_data[3] ;
 wire \i2c_slave_controller.out_regf_write_data[4] ;
 wire \i2c_slave_controller.out_regf_write_data[5] ;
 wire \i2c_slave_controller.out_regf_write_data[6] ;
 wire \i2c_slave_controller.out_regf_write_data[7] ;
 wire \i2c_slave_controller.out_start ;
 wire \i2c_slave_controller.out_start_reset ;
 wire \i2c_slave_controller.out_stop ;
 wire \i2c_slave_controller.out_stop_reset ;
 wire \i2c_slave_controller.reg_sda_out ;
 wire \i2c_slave_controller.start_resetter ;
 wire \i2c_slave_controller.state[0] ;
 wire \i2c_slave_controller.state[1] ;
 wire \i2c_slave_controller.state[2] ;
 wire \i2c_slave_controller.stop_resetter ;
 wire \i2c_slave_controller.write_enable ;
 wire \reg_file.reg_array[0] ;
 wire \reg_file.reg_array[100] ;
 wire \reg_file.reg_array[101] ;
 wire \reg_file.reg_array[102] ;
 wire \reg_file.reg_array[103] ;
 wire \reg_file.reg_array[104] ;
 wire \reg_file.reg_array[105] ;
 wire \reg_file.reg_array[106] ;
 wire \reg_file.reg_array[107] ;
 wire \reg_file.reg_array[108] ;
 wire \reg_file.reg_array[109] ;
 wire \reg_file.reg_array[10] ;
 wire \reg_file.reg_array[110] ;
 wire \reg_file.reg_array[111] ;
 wire \reg_file.reg_array[112] ;
 wire \reg_file.reg_array[113] ;
 wire \reg_file.reg_array[114] ;
 wire \reg_file.reg_array[115] ;
 wire \reg_file.reg_array[116] ;
 wire \reg_file.reg_array[117] ;
 wire \reg_file.reg_array[118] ;
 wire \reg_file.reg_array[119] ;
 wire \reg_file.reg_array[11] ;
 wire \reg_file.reg_array[120] ;
 wire \reg_file.reg_array[121] ;
 wire \reg_file.reg_array[122] ;
 wire \reg_file.reg_array[123] ;
 wire \reg_file.reg_array[124] ;
 wire \reg_file.reg_array[125] ;
 wire \reg_file.reg_array[126] ;
 wire \reg_file.reg_array[127] ;
 wire \reg_file.reg_array[12] ;
 wire \reg_file.reg_array[13] ;
 wire \reg_file.reg_array[14] ;
 wire \reg_file.reg_array[15] ;
 wire \reg_file.reg_array[16] ;
 wire \reg_file.reg_array[17] ;
 wire \reg_file.reg_array[18] ;
 wire \reg_file.reg_array[19] ;
 wire \reg_file.reg_array[1] ;
 wire \reg_file.reg_array[20] ;
 wire \reg_file.reg_array[21] ;
 wire \reg_file.reg_array[22] ;
 wire \reg_file.reg_array[23] ;
 wire \reg_file.reg_array[24] ;
 wire \reg_file.reg_array[25] ;
 wire \reg_file.reg_array[26] ;
 wire \reg_file.reg_array[27] ;
 wire \reg_file.reg_array[28] ;
 wire \reg_file.reg_array[29] ;
 wire \reg_file.reg_array[2] ;
 wire \reg_file.reg_array[30] ;
 wire \reg_file.reg_array[31] ;
 wire \reg_file.reg_array[32] ;
 wire \reg_file.reg_array[33] ;
 wire \reg_file.reg_array[34] ;
 wire \reg_file.reg_array[35] ;
 wire \reg_file.reg_array[36] ;
 wire \reg_file.reg_array[37] ;
 wire \reg_file.reg_array[38] ;
 wire \reg_file.reg_array[39] ;
 wire \reg_file.reg_array[3] ;
 wire \reg_file.reg_array[40] ;
 wire \reg_file.reg_array[41] ;
 wire \reg_file.reg_array[42] ;
 wire \reg_file.reg_array[43] ;
 wire \reg_file.reg_array[44] ;
 wire \reg_file.reg_array[45] ;
 wire \reg_file.reg_array[46] ;
 wire \reg_file.reg_array[47] ;
 wire \reg_file.reg_array[48] ;
 wire \reg_file.reg_array[49] ;
 wire \reg_file.reg_array[4] ;
 wire \reg_file.reg_array[50] ;
 wire \reg_file.reg_array[51] ;
 wire \reg_file.reg_array[52] ;
 wire \reg_file.reg_array[53] ;
 wire \reg_file.reg_array[54] ;
 wire \reg_file.reg_array[55] ;
 wire \reg_file.reg_array[56] ;
 wire \reg_file.reg_array[57] ;
 wire \reg_file.reg_array[58] ;
 wire \reg_file.reg_array[59] ;
 wire \reg_file.reg_array[5] ;
 wire \reg_file.reg_array[60] ;
 wire \reg_file.reg_array[61] ;
 wire \reg_file.reg_array[62] ;
 wire \reg_file.reg_array[63] ;
 wire \reg_file.reg_array[64] ;
 wire \reg_file.reg_array[65] ;
 wire \reg_file.reg_array[66] ;
 wire \reg_file.reg_array[67] ;
 wire \reg_file.reg_array[68] ;
 wire \reg_file.reg_array[69] ;
 wire \reg_file.reg_array[6] ;
 wire \reg_file.reg_array[70] ;
 wire \reg_file.reg_array[71] ;
 wire \reg_file.reg_array[72] ;
 wire \reg_file.reg_array[73] ;
 wire \reg_file.reg_array[74] ;
 wire \reg_file.reg_array[75] ;
 wire \reg_file.reg_array[76] ;
 wire \reg_file.reg_array[77] ;
 wire \reg_file.reg_array[78] ;
 wire \reg_file.reg_array[79] ;
 wire \reg_file.reg_array[7] ;
 wire \reg_file.reg_array[80] ;
 wire \reg_file.reg_array[81] ;
 wire \reg_file.reg_array[82] ;
 wire \reg_file.reg_array[83] ;
 wire \reg_file.reg_array[84] ;
 wire \reg_file.reg_array[85] ;
 wire \reg_file.reg_array[86] ;
 wire \reg_file.reg_array[87] ;
 wire \reg_file.reg_array[88] ;
 wire \reg_file.reg_array[89] ;
 wire \reg_file.reg_array[8] ;
 wire \reg_file.reg_array[90] ;
 wire \reg_file.reg_array[91] ;
 wire \reg_file.reg_array[92] ;
 wire \reg_file.reg_array[93] ;
 wire \reg_file.reg_array[94] ;
 wire \reg_file.reg_array[95] ;
 wire \reg_file.reg_array[96] ;
 wire \reg_file.reg_array[97] ;
 wire \reg_file.reg_array[98] ;
 wire \reg_file.reg_array[99] ;
 wire \reg_file.reg_array[9] ;
 wire \reg_file.reg_pointer[0] ;
 wire \reg_file.reg_pointer[1] ;
 wire \reg_file.reg_pointer[2] ;
 wire \reg_file.reg_pointer[3] ;
 wire \reg_file.state[0] ;
 wire net12;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net1;
 wire net2;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_2_0__leaf_clk_regs;
 wire clknet_2_1__leaf_clk_regs;
 wire clknet_2_2__leaf_clk_regs;
 wire clknet_2_3__leaf_clk_regs;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;

 sg13g2_inv_1 _0834_ (.Y(_0210_),
    .A(net34));
 sg13g2_inv_1 _0835_ (.Y(_0211_),
    .A(net537));
 sg13g2_inv_1 _0836_ (.Y(_0024_),
    .A(net1));
 sg13g2_inv_1 _0837_ (.Y(_0212_),
    .A(net517));
 sg13g2_inv_1 _0838_ (.Y(_0213_),
    .A(\i2c_slave_controller.addr[0] ));
 sg13g2_inv_1 _0839_ (.Y(_0214_),
    .A(net521));
 sg13g2_inv_1 _0840_ (.Y(_0215_),
    .A(net527));
 sg13g2_inv_1 _0841_ (.Y(_0216_),
    .A(\reg_file.reg_array[72] ));
 sg13g2_inv_1 _0842_ (.Y(_0217_),
    .A(\reg_file.reg_array[73] ));
 sg13g2_inv_1 _0843_ (.Y(_0218_),
    .A(\reg_file.reg_array[74] ));
 sg13g2_inv_1 _0844_ (.Y(_0219_),
    .A(\reg_file.reg_array[75] ));
 sg13g2_inv_1 _0845_ (.Y(_0220_),
    .A(\reg_file.reg_array[76] ));
 sg13g2_inv_1 _0846_ (.Y(_0221_),
    .A(\reg_file.reg_array[77] ));
 sg13g2_inv_1 _0847_ (.Y(_0222_),
    .A(\reg_file.reg_array[78] ));
 sg13g2_inv_1 _0848_ (.Y(_0223_),
    .A(\reg_file.reg_array[79] ));
 sg13g2_inv_1 _0849_ (.Y(_0224_),
    .A(uo_out[2]));
 sg13g2_inv_1 _0850_ (.Y(_0225_),
    .A(uo_out[3]));
 sg13g2_inv_1 _0851_ (.Y(_0226_),
    .A(uo_out[4]));
 sg13g2_inv_1 _0852_ (.Y(_0227_),
    .A(_0004_));
 sg13g2_inv_1 _1490__2 (.Y(net13),
    .A(clknet_1_0__leaf_clk));
 sg13g2_nor2b_1 _0854_ (.A(\i2c_slave_controller.start_resetter ),
    .B_N(net580),
    .Y(_0023_));
 sg13g2_inv_1 _0855_ (.Y(\i2c_slave_controller.out_start_reset ),
    .A(_0023_));
 sg13g2_nor3_1 _0856_ (.A(\i2c_slave_controller.addr[1] ),
    .B(\i2c_slave_controller.addr[3] ),
    .C(\i2c_slave_controller.addr[5] ),
    .Y(_0228_));
 sg13g2_nor2b_1 _0857_ (.A(\i2c_slave_controller.addr[7] ),
    .B_N(\i2c_slave_controller.addr[6] ),
    .Y(_0229_));
 sg13g2_nand4_1 _0858_ (.B(\i2c_slave_controller.addr[4] ),
    .C(_0228_),
    .A(\i2c_slave_controller.addr[2] ),
    .Y(_0230_),
    .D(_0229_));
 sg13g2_nand3b_1 _0859_ (.B(net540),
    .C(_0001_),
    .Y(_0231_),
    .A_N(\i2c_slave_controller.state[1] ));
 sg13g2_or2_1 _0860_ (.X(_0232_),
    .B(net508),
    .A(_0230_));
 sg13g2_nor3_1 _0861_ (.A(\i2c_slave_controller.addr[0] ),
    .B(_0230_),
    .C(net508),
    .Y(_0233_));
 sg13g2_nor2_2 _0862_ (.A(net519),
    .B(net520),
    .Y(_0234_));
 sg13g2_or2_1 _0863_ (.X(_0235_),
    .B(net520),
    .A(net519));
 sg13g2_nor2_1 _0864_ (.A(_0212_),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_nand2_1 _0865_ (.Y(_0237_),
    .A(net517),
    .B(_0234_));
 sg13g2_nor3_1 _0866_ (.A(_0212_),
    .B(net508),
    .C(_0235_),
    .Y(_0238_));
 sg13g2_or3_1 _0867_ (.A(_0212_),
    .B(net508),
    .C(_0235_),
    .X(_0239_));
 sg13g2_and2_1 _0868_ (.A(_0230_),
    .B(_0238_),
    .X(_0240_));
 sg13g2_nand2b_2 _0869_ (.Y(_0241_),
    .B(\i2c_slave_controller.state[0] ),
    .A_N(net538));
 sg13g2_and3_1 _0870_ (.X(_0242_),
    .A(net540),
    .B(net537),
    .C(_0237_));
 sg13g2_nor4_2 _0871_ (.A(_0233_),
    .B(_0240_),
    .C(_0241_),
    .Y(_0243_),
    .D(_0242_));
 sg13g2_nand2_1 _0872_ (.Y(_0244_),
    .A(net539),
    .B(net540));
 sg13g2_nand3_1 _0873_ (.B(net540),
    .C(net537),
    .A(net539),
    .Y(_0245_));
 sg13g2_mux2_1 _0874_ (.A0(net36),
    .A1(net507),
    .S(_0243_),
    .X(_0047_));
 sg13g2_nor2b_1 _0875_ (.A(net540),
    .B_N(net539),
    .Y(_0246_));
 sg13g2_and2_1 _0876_ (.A(net537),
    .B(_0246_),
    .X(_0247_));
 sg13g2_nand2_1 _0877_ (.Y(_0248_),
    .A(net537),
    .B(_0246_));
 sg13g2_nand2_1 _0878_ (.Y(_0249_),
    .A(_0213_),
    .B(_0247_));
 sg13g2_nor2_1 _0879_ (.A(net539),
    .B(net540),
    .Y(_0250_));
 sg13g2_or2_2 _0880_ (.X(_0251_),
    .B(\i2c_slave_controller.state[0] ),
    .A(\i2c_slave_controller.state[1] ));
 sg13g2_nor2b_1 _0881_ (.A(net539),
    .B_N(net538),
    .Y(_0252_));
 sg13g2_nand2_2 _0882_ (.Y(_0253_),
    .A(net538),
    .B(_0250_));
 sg13g2_nand2b_1 _0883_ (.Y(_0254_),
    .B(_0251_),
    .A_N(\i2c_slave_controller.state[2] ));
 sg13g2_a22oi_1 _0884_ (.Y(_0255_),
    .B1(_0253_),
    .B2(_0254_),
    .A2(_0237_),
    .A1(net540));
 sg13g2_and2_1 _0885_ (.A(_0249_),
    .B(_0255_),
    .X(_0256_));
 sg13g2_nor2b_1 _0886_ (.A(net520),
    .B_N(net519),
    .Y(_0257_));
 sg13g2_nand2_1 _0887_ (.Y(_0258_),
    .A(\i2c_slave_controller.counter[1] ),
    .B(_0210_));
 sg13g2_a21oi_1 _0888_ (.A1(uo_out[2]),
    .A2(_0257_),
    .Y(_0259_),
    .B1(\i2c_slave_controller.counter[2] ));
 sg13g2_nand2_2 _0889_ (.Y(_0260_),
    .A(net50),
    .B(net34));
 sg13g2_nand3_1 _0890_ (.B(net520),
    .C(uo_out[3]),
    .A(net519),
    .Y(_0261_));
 sg13g2_nor2b_2 _0891_ (.A(net519),
    .B_N(net520),
    .Y(_0262_));
 sg13g2_nand2b_1 _0892_ (.Y(_0263_),
    .B(net520),
    .A_N(\i2c_slave_controller.counter[1] ));
 sg13g2_a22oi_1 _0893_ (.Y(_0264_),
    .B1(_0262_),
    .B2(uo_out[1]),
    .A2(_0234_),
    .A1(uo_out[0]));
 sg13g2_nand3_1 _0894_ (.B(_0261_),
    .C(_0264_),
    .A(_0259_),
    .Y(_0265_));
 sg13g2_nand3_1 _0895_ (.B(net520),
    .C(uo_out[7]),
    .A(net519),
    .Y(_0266_));
 sg13g2_nand2_1 _0896_ (.Y(_0267_),
    .A(uo_out[5]),
    .B(_0262_));
 sg13g2_a22oi_1 _0897_ (.Y(_0268_),
    .B1(_0257_),
    .B2(uo_out[6]),
    .A2(_0234_),
    .A1(uo_out[4]));
 sg13g2_nand4_1 _0898_ (.B(_0266_),
    .C(_0267_),
    .A(\i2c_slave_controller.counter[2] ),
    .Y(_0269_),
    .D(_0268_));
 sg13g2_and3_1 _0899_ (.X(_0270_),
    .A(_0241_),
    .B(_0265_),
    .C(_0269_));
 sg13g2_mux2_1 _0900_ (.A0(net23),
    .A1(_0270_),
    .S(_0256_),
    .X(_0046_));
 sg13g2_nand2_1 _0901_ (.Y(_0271_),
    .A(net538),
    .B(_0246_));
 sg13g2_nand4_1 _0902_ (.B(_0241_),
    .C(_0248_),
    .A(net539),
    .Y(_0272_),
    .D(_0271_));
 sg13g2_mux2_1 _0903_ (.A0(net22),
    .A1(_0256_),
    .S(_0272_),
    .X(_0045_));
 sg13g2_a21o_1 _0904_ (.A2(_0253_),
    .A1(net506),
    .B1(_0237_),
    .X(_0273_));
 sg13g2_nand2_1 _0905_ (.Y(_0274_),
    .A(net537),
    .B(_0250_));
 sg13g2_nor3_1 _0906_ (.A(_0211_),
    .B(\i2c_slave_controller.out_start ),
    .C(_0251_),
    .Y(_0275_));
 sg13g2_a221oi_1 _0907_ (.B2(_0213_),
    .C1(_0275_),
    .B1(_0247_),
    .A1(_0230_),
    .Y(_0276_),
    .A2(_0238_));
 sg13g2_nand2_1 _0908_ (.Y(_0277_),
    .A(_0211_),
    .B(_0253_));
 sg13g2_nand3_1 _0909_ (.B(_0276_),
    .C(_0277_),
    .A(_0273_),
    .Y(_0278_));
 sg13g2_nand4_1 _0910_ (.B(_0273_),
    .C(_0276_),
    .A(_0234_),
    .Y(_0279_),
    .D(_0277_));
 sg13g2_mux2_1 _0911_ (.A0(net538),
    .A1(net537),
    .S(_0251_),
    .X(_0280_));
 sg13g2_nand2b_1 _0912_ (.Y(_0281_),
    .B(_0234_),
    .A_N(\i2c_slave_controller.counter[2] ));
 sg13g2_nand3_1 _0913_ (.B(_0280_),
    .C(_0281_),
    .A(_0239_),
    .Y(_0282_));
 sg13g2_and4_1 _0914_ (.A(_0273_),
    .B(_0276_),
    .C(_0277_),
    .D(_0282_),
    .X(_0283_));
 sg13g2_a21o_1 _0915_ (.A2(_0279_),
    .A1(net33),
    .B1(_0283_),
    .X(_0044_));
 sg13g2_nand3_1 _0916_ (.B(_0260_),
    .C(_0280_),
    .A(_0235_),
    .Y(_0284_));
 sg13g2_mux2_1 _0917_ (.A0(_0284_),
    .A1(net519),
    .S(_0278_),
    .X(_0043_));
 sg13g2_and4_1 _0918_ (.A(net520),
    .B(_0273_),
    .C(_0276_),
    .D(_0280_),
    .X(_0285_));
 sg13g2_a21oi_1 _0919_ (.A1(_0210_),
    .A2(_0278_),
    .Y(_0042_),
    .B1(_0285_));
 sg13g2_a21o_1 _0920_ (.A2(_0244_),
    .A1(net538),
    .B1(_0001_),
    .X(_0286_));
 sg13g2_o21ai_1 _0921_ (.B1(_0286_),
    .Y(_0287_),
    .A1(_0236_),
    .A2(_0253_));
 sg13g2_nor2_1 _0922_ (.A(\i2c_slave_controller.ack_recieved ),
    .B(_0271_),
    .Y(_0288_));
 sg13g2_or4_2 _0923_ (.A(_0242_),
    .B(_0275_),
    .C(_0287_),
    .D(_0288_),
    .X(_0289_));
 sg13g2_nand2_1 _0924_ (.Y(_0290_),
    .A(\i2c_slave_controller.addr[0] ),
    .B(_0247_));
 sg13g2_nand3_1 _0925_ (.B(_0253_),
    .C(_0290_),
    .A(net506),
    .Y(_0291_));
 sg13g2_mux2_1 _0926_ (.A0(_0291_),
    .A1(net538),
    .S(_0289_),
    .X(_0027_));
 sg13g2_nand3_1 _0927_ (.B(_0249_),
    .C(_0253_),
    .A(_0232_),
    .Y(_0292_));
 sg13g2_mux2_1 _0928_ (.A0(_0292_),
    .A1(net539),
    .S(_0289_),
    .X(_0026_));
 sg13g2_a22oi_1 _0929_ (.Y(_0293_),
    .B1(_0251_),
    .B2(_0001_),
    .A2(_0244_),
    .A1(net538));
 sg13g2_inv_1 _0930_ (.Y(_0294_),
    .A(_0293_));
 sg13g2_nand3_1 _0931_ (.B(_0249_),
    .C(_0294_),
    .A(net506),
    .Y(_0295_));
 sg13g2_mux2_1 _0932_ (.A0(_0295_),
    .A1(net540),
    .S(_0289_),
    .X(_0025_));
 sg13g2_nor2b_1 _0933_ (.A(\i2c_slave_controller.stop_resetter ),
    .B_N(net578),
    .Y(_0022_));
 sg13g2_inv_1 _0934_ (.Y(\i2c_slave_controller.out_stop_reset ),
    .A(_0022_));
 sg13g2_nor2_2 _0935_ (.A(\i2c_slave_controller.out_regf_rw ),
    .B(\reg_file.state[0] ),
    .Y(_0296_));
 sg13g2_mux2_1 _0936_ (.A0(\reg_file.reg_pointer[0] ),
    .A1(\i2c_slave_controller.out_regf_write_data[0] ),
    .S(_0296_),
    .X(_0028_));
 sg13g2_mux2_1 _0937_ (.A0(net534),
    .A1(\i2c_slave_controller.out_regf_write_data[1] ),
    .S(_0296_),
    .X(_0029_));
 sg13g2_nand2_1 _0938_ (.Y(_0297_),
    .A(\i2c_slave_controller.out_regf_write_data[2] ),
    .B(_0296_));
 sg13g2_o21ai_1 _0939_ (.B1(_0297_),
    .Y(_0030_),
    .A1(net513),
    .A2(_0296_));
 sg13g2_nand2_1 _0940_ (.Y(_0298_),
    .A(\i2c_slave_controller.out_regf_write_data[3] ),
    .B(_0296_));
 sg13g2_o21ai_1 _0941_ (.B1(_0298_),
    .Y(_0031_),
    .A1(net516),
    .A2(_0296_));
 sg13g2_nand2_1 _0942_ (.Y(_0299_),
    .A(net21),
    .B(_0274_));
 sg13g2_o21ai_1 _0943_ (.B1(_0299_),
    .Y(_0032_),
    .A1(net1),
    .A2(_0271_));
 sg13g2_o21ai_1 _0944_ (.B1(net45),
    .Y(_0300_),
    .A1(_0237_),
    .A2(net506));
 sg13g2_nand3_1 _0945_ (.B(net517),
    .C(_0234_),
    .A(net1),
    .Y(_0301_));
 sg13g2_o21ai_1 _0946_ (.B1(_0300_),
    .Y(_0033_),
    .A1(net507),
    .A2(_0301_));
 sg13g2_nand2_1 _0947_ (.Y(_0302_),
    .A(net518),
    .B(_0262_));
 sg13g2_nor2_1 _0948_ (.A(net507),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_nor2_1 _0949_ (.A(net40),
    .B(_0303_),
    .Y(_0304_));
 sg13g2_a21oi_1 _0950_ (.A1(net567),
    .A2(_0303_),
    .Y(_0034_),
    .B1(_0304_));
 sg13g2_nand2_1 _0951_ (.Y(_0305_),
    .A(net517),
    .B(_0257_));
 sg13g2_nor2_1 _0952_ (.A(net507),
    .B(_0305_),
    .Y(_0306_));
 sg13g2_nor2_1 _0953_ (.A(net41),
    .B(_0306_),
    .Y(_0307_));
 sg13g2_a21oi_1 _0954_ (.A1(net567),
    .A2(_0306_),
    .Y(_0035_),
    .B1(_0307_));
 sg13g2_nand3_1 _0955_ (.B(\i2c_slave_controller.counter[0] ),
    .C(net517),
    .A(net519),
    .Y(_0308_));
 sg13g2_nor2_2 _0956_ (.A(net506),
    .B(_0308_),
    .Y(_0309_));
 sg13g2_nor2_1 _0957_ (.A(net44),
    .B(_0309_),
    .Y(_0310_));
 sg13g2_a21oi_1 _0958_ (.A1(net567),
    .A2(_0309_),
    .Y(_0036_),
    .B1(_0310_));
 sg13g2_nand2_1 _0959_ (.Y(_0311_),
    .A(_0212_),
    .B(_0234_));
 sg13g2_o21ai_1 _0960_ (.B1(net39),
    .Y(_0312_),
    .A1(net507),
    .A2(_0311_));
 sg13g2_nand3_1 _0961_ (.B(_0212_),
    .C(_0234_),
    .A(net1),
    .Y(_0313_));
 sg13g2_o21ai_1 _0962_ (.B1(_0312_),
    .Y(_0037_),
    .A1(net507),
    .A2(_0313_));
 sg13g2_nor3_2 _0963_ (.A(net517),
    .B(net506),
    .C(_0263_),
    .Y(_0314_));
 sg13g2_nor2_1 _0964_ (.A(net38),
    .B(_0314_),
    .Y(_0315_));
 sg13g2_a21oi_1 _0965_ (.A1(net567),
    .A2(_0314_),
    .Y(_0038_),
    .B1(_0315_));
 sg13g2_nor3_2 _0966_ (.A(net517),
    .B(net506),
    .C(_0258_),
    .Y(_0316_));
 sg13g2_nor2_1 _0967_ (.A(net43),
    .B(_0316_),
    .Y(_0317_));
 sg13g2_a21oi_1 _0968_ (.A1(net567),
    .A2(_0316_),
    .Y(_0039_),
    .B1(_0317_));
 sg13g2_nor3_2 _0969_ (.A(net517),
    .B(net506),
    .C(_0260_),
    .Y(_0318_));
 sg13g2_nor2_1 _0970_ (.A(net42),
    .B(_0318_),
    .Y(_0319_));
 sg13g2_a21oi_1 _0971_ (.A1(net567),
    .A2(_0318_),
    .Y(_0040_),
    .B1(_0319_));
 sg13g2_nand2_1 _0972_ (.Y(_0320_),
    .A(net539),
    .B(net32));
 sg13g2_nand2_1 _0973_ (.Y(_0321_),
    .A(net537),
    .B(_0244_));
 sg13g2_o21ai_1 _0974_ (.B1(_0253_),
    .Y(_0322_),
    .A1(_0252_),
    .A2(_0321_));
 sg13g2_nor2_1 _0975_ (.A(net551),
    .B(_0252_),
    .Y(_0323_));
 sg13g2_a22oi_1 _0976_ (.Y(_0041_),
    .B1(_0323_),
    .B2(_0321_),
    .A2(_0322_),
    .A1(_0320_));
 sg13g2_nand2b_1 _0977_ (.Y(_0324_),
    .B(\i2c_slave_controller.out_regf_rw ),
    .A_N(\reg_file.state[0] ));
 sg13g2_and2_1 _0978_ (.A(_0000_),
    .B(_0324_),
    .X(_0048_));
 sg13g2_nor2_1 _0979_ (.A(net536),
    .B(net535),
    .Y(_0325_));
 sg13g2_xnor2_1 _0980_ (.Y(_0326_),
    .A(net526),
    .B(net503));
 sg13g2_nor2b_1 _0981_ (.A(\i2c_slave_controller.out_regf_rw ),
    .B_N(\reg_file.state[0] ),
    .Y(_0327_));
 sg13g2_nand2b_1 _0982_ (.Y(_0328_),
    .B(\reg_file.state[0] ),
    .A_N(\i2c_slave_controller.out_regf_rw ));
 sg13g2_nor2_2 _0983_ (.A(net531),
    .B(net525),
    .Y(_0329_));
 sg13g2_or2_1 _0984_ (.X(_0330_),
    .B(net525),
    .A(net531));
 sg13g2_nand3_1 _0985_ (.B(_0004_),
    .C(_0329_),
    .A(_0003_),
    .Y(_0331_));
 sg13g2_nor4_2 _0986_ (.A(\reg_file.reg_pointer[3] ),
    .B(net479),
    .C(net497),
    .Y(_0332_),
    .D(net478));
 sg13g2_nor2_1 _0987_ (.A(\reg_file.reg_array[0] ),
    .B(net470),
    .Y(_0333_));
 sg13g2_a21oi_1 _0988_ (.A1(_0005_),
    .A2(net470),
    .Y(_0049_),
    .B1(_0333_));
 sg13g2_nor2_1 _0989_ (.A(\reg_file.reg_array[1] ),
    .B(net470),
    .Y(_0334_));
 sg13g2_a21oi_1 _0990_ (.A1(_0006_),
    .A2(net470),
    .Y(_0050_),
    .B1(_0334_));
 sg13g2_nor2_1 _0991_ (.A(\reg_file.reg_array[2] ),
    .B(net470),
    .Y(_0335_));
 sg13g2_a21oi_1 _0992_ (.A1(_0007_),
    .A2(net470),
    .Y(_0051_),
    .B1(_0335_));
 sg13g2_nor2_1 _0993_ (.A(\reg_file.reg_array[3] ),
    .B(net469),
    .Y(_0336_));
 sg13g2_a21oi_1 _0994_ (.A1(_0008_),
    .A2(net469),
    .Y(_0052_),
    .B1(_0336_));
 sg13g2_nor2_1 _0995_ (.A(\reg_file.reg_array[4] ),
    .B(net470),
    .Y(_0337_));
 sg13g2_a21oi_1 _0996_ (.A1(_0009_),
    .A2(net470),
    .Y(_0053_),
    .B1(_0337_));
 sg13g2_nor2_1 _0997_ (.A(\reg_file.reg_array[5] ),
    .B(net469),
    .Y(_0338_));
 sg13g2_a21oi_1 _0998_ (.A1(_0010_),
    .A2(net469),
    .Y(_0054_),
    .B1(_0338_));
 sg13g2_nor2_1 _0999_ (.A(\reg_file.reg_array[6] ),
    .B(net469),
    .Y(_0339_));
 sg13g2_a21oi_1 _1000_ (.A1(_0011_),
    .A2(net469),
    .Y(_0055_),
    .B1(_0339_));
 sg13g2_nor2_1 _1001_ (.A(\reg_file.reg_array[7] ),
    .B(net469),
    .Y(_0340_));
 sg13g2_a21oi_1 _1002_ (.A1(_0012_),
    .A2(net469),
    .Y(_0056_),
    .B1(_0340_));
 sg13g2_nor2b_1 _1003_ (.A(net534),
    .B_N(net536),
    .Y(_0341_));
 sg13g2_and2_1 _1004_ (.A(net511),
    .B(net495),
    .X(_0342_));
 sg13g2_o21ai_1 _1005_ (.B1(net522),
    .Y(_0343_),
    .A1(_0227_),
    .A2(_0330_));
 sg13g2_nand3_1 _1006_ (.B(_0004_),
    .C(_0329_),
    .A(net516),
    .Y(_0344_));
 sg13g2_o21ai_1 _1007_ (.B1(net516),
    .Y(_0345_),
    .A1(_0227_),
    .A2(_0330_));
 sg13g2_nand3_1 _1008_ (.B(_0004_),
    .C(_0329_),
    .A(net522),
    .Y(_0346_));
 sg13g2_a21oi_2 _1009_ (.B1(net496),
    .Y(_0347_),
    .A2(_0346_),
    .A1(_0345_));
 sg13g2_nand3_1 _1010_ (.B(_0343_),
    .C(_0344_),
    .A(net499),
    .Y(_0348_));
 sg13g2_nand3_1 _1011_ (.B(net473),
    .C(net468),
    .A(net476),
    .Y(_0349_));
 sg13g2_and4_1 _1012_ (.A(\i2c_slave_controller.out_regf_write_data[0] ),
    .B(net477),
    .C(net474),
    .D(_0347_),
    .X(_0350_));
 sg13g2_a21o_1 _1013_ (.A2(_0349_),
    .A1(\reg_file.reg_array[8] ),
    .B1(_0350_),
    .X(_0057_));
 sg13g2_and4_1 _1014_ (.A(\i2c_slave_controller.out_regf_write_data[1] ),
    .B(net477),
    .C(net474),
    .D(_0347_),
    .X(_0351_));
 sg13g2_a21o_1 _1015_ (.A2(_0349_),
    .A1(\reg_file.reg_array[9] ),
    .B1(_0351_),
    .X(_0058_));
 sg13g2_and4_1 _1016_ (.A(\i2c_slave_controller.out_regf_write_data[2] ),
    .B(net477),
    .C(net474),
    .D(net468),
    .X(_0352_));
 sg13g2_a21o_1 _1017_ (.A2(_0349_),
    .A1(\reg_file.reg_array[10] ),
    .B1(_0352_),
    .X(_0059_));
 sg13g2_and4_1 _1018_ (.A(\i2c_slave_controller.out_regf_write_data[3] ),
    .B(net476),
    .C(net473),
    .D(net468),
    .X(_0353_));
 sg13g2_a21o_1 _1019_ (.A2(_0349_),
    .A1(\reg_file.reg_array[11] ),
    .B1(_0353_),
    .X(_0060_));
 sg13g2_and4_1 _1020_ (.A(\i2c_slave_controller.out_regf_write_data[4] ),
    .B(net477),
    .C(net474),
    .D(net468),
    .X(_0354_));
 sg13g2_a21o_1 _1021_ (.A2(_0349_),
    .A1(\reg_file.reg_array[12] ),
    .B1(_0354_),
    .X(_0061_));
 sg13g2_and4_1 _1022_ (.A(\i2c_slave_controller.out_regf_write_data[5] ),
    .B(net478),
    .C(net475),
    .D(net468),
    .X(_0355_));
 sg13g2_a21o_1 _1023_ (.A2(_0349_),
    .A1(\reg_file.reg_array[13] ),
    .B1(_0355_),
    .X(_0062_));
 sg13g2_and4_1 _1024_ (.A(\i2c_slave_controller.out_regf_write_data[6] ),
    .B(net476),
    .C(net473),
    .D(net468),
    .X(_0356_));
 sg13g2_a21o_1 _1025_ (.A2(_0349_),
    .A1(\reg_file.reg_array[14] ),
    .B1(_0356_),
    .X(_0063_));
 sg13g2_and4_1 _1026_ (.A(\i2c_slave_controller.out_regf_write_data[7] ),
    .B(net476),
    .C(net473),
    .D(net468),
    .X(_0357_));
 sg13g2_a21o_1 _1027_ (.A2(_0349_),
    .A1(\reg_file.reg_array[15] ),
    .B1(_0357_),
    .X(_0064_));
 sg13g2_nor2b_1 _1028_ (.A(net536),
    .B_N(net534),
    .Y(_0358_));
 sg13g2_and2_1 _1029_ (.A(net511),
    .B(net486),
    .X(_0359_));
 sg13g2_nand4_1 _1030_ (.B(_0343_),
    .C(_0344_),
    .A(net499),
    .Y(_0360_),
    .D(_0359_));
 sg13g2_nand2_1 _1031_ (.Y(_0361_),
    .A(\reg_file.reg_array[16] ),
    .B(_0360_));
 sg13g2_a21o_2 _1032_ (.A2(_0329_),
    .A1(_0003_),
    .B1(net536),
    .X(_0362_));
 sg13g2_nor2_2 _1033_ (.A(_0005_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_nand3_1 _1034_ (.B(net513),
    .C(_0363_),
    .A(net532),
    .Y(_0364_));
 sg13g2_o21ai_1 _1035_ (.B1(_0361_),
    .Y(_0065_),
    .A1(net465),
    .A2(_0364_));
 sg13g2_nand2_1 _1036_ (.Y(_0365_),
    .A(\reg_file.reg_array[17] ),
    .B(_0360_));
 sg13g2_nor2_2 _1037_ (.A(_0006_),
    .B(_0362_),
    .Y(_0366_));
 sg13g2_nand3_1 _1038_ (.B(net513),
    .C(_0366_),
    .A(net534),
    .Y(_0367_));
 sg13g2_o21ai_1 _1039_ (.B1(_0365_),
    .Y(_0066_),
    .A1(net465),
    .A2(_0367_));
 sg13g2_nand2_1 _1040_ (.Y(_0368_),
    .A(\reg_file.reg_array[18] ),
    .B(_0360_));
 sg13g2_nor2_2 _1041_ (.A(_0007_),
    .B(_0362_),
    .Y(_0369_));
 sg13g2_nand3_1 _1042_ (.B(net513),
    .C(_0369_),
    .A(net534),
    .Y(_0370_));
 sg13g2_o21ai_1 _1043_ (.B1(_0368_),
    .Y(_0067_),
    .A1(net466),
    .A2(_0370_));
 sg13g2_nand2_1 _1044_ (.Y(_0371_),
    .A(\reg_file.reg_array[19] ),
    .B(_0360_));
 sg13g2_nor2_2 _1045_ (.A(_0008_),
    .B(_0362_),
    .Y(_0372_));
 sg13g2_nand3_1 _1046_ (.B(net511),
    .C(_0372_),
    .A(net531),
    .Y(_0373_));
 sg13g2_o21ai_1 _1047_ (.B1(_0371_),
    .Y(_0068_),
    .A1(net462),
    .A2(_0373_));
 sg13g2_nand2_1 _1048_ (.Y(_0374_),
    .A(\reg_file.reg_array[20] ),
    .B(_0360_));
 sg13g2_nor2_2 _1049_ (.A(_0009_),
    .B(_0362_),
    .Y(_0375_));
 sg13g2_nand3_1 _1050_ (.B(net513),
    .C(_0375_),
    .A(net535),
    .Y(_0376_));
 sg13g2_o21ai_1 _1051_ (.B1(_0374_),
    .Y(_0069_),
    .A1(net466),
    .A2(_0376_));
 sg13g2_nand2_1 _1052_ (.Y(_0377_),
    .A(\reg_file.reg_array[21] ),
    .B(_0360_));
 sg13g2_nor2_2 _1053_ (.A(_0010_),
    .B(_0362_),
    .Y(_0378_));
 sg13g2_nand3_1 _1054_ (.B(net511),
    .C(_0378_),
    .A(net530),
    .Y(_0379_));
 sg13g2_o21ai_1 _1055_ (.B1(_0377_),
    .Y(_0070_),
    .A1(net462),
    .A2(_0379_));
 sg13g2_nand2_1 _1056_ (.Y(_0380_),
    .A(\reg_file.reg_array[22] ),
    .B(_0360_));
 sg13g2_nor2_2 _1057_ (.A(_0011_),
    .B(_0362_),
    .Y(_0381_));
 sg13g2_nand3_1 _1058_ (.B(net511),
    .C(_0381_),
    .A(net529),
    .Y(_0382_));
 sg13g2_o21ai_1 _1059_ (.B1(_0380_),
    .Y(_0071_),
    .A1(net461),
    .A2(_0382_));
 sg13g2_nand2_1 _1060_ (.Y(_0383_),
    .A(\reg_file.reg_array[23] ),
    .B(_0360_));
 sg13g2_nor2_2 _1061_ (.A(_0012_),
    .B(_0362_),
    .Y(_0384_));
 sg13g2_nand3_1 _1062_ (.B(net511),
    .C(_0384_),
    .A(net531),
    .Y(_0385_));
 sg13g2_o21ai_1 _1063_ (.B1(_0383_),
    .Y(_0072_),
    .A1(net461),
    .A2(_0385_));
 sg13g2_and2_1 _1064_ (.A(net536),
    .B(net534),
    .X(_0386_));
 sg13g2_and2_2 _1065_ (.A(net511),
    .B(net482),
    .X(_0387_));
 sg13g2_nand2_1 _1066_ (.Y(_0388_),
    .A(net513),
    .B(net484));
 sg13g2_o21ai_1 _1067_ (.B1(\reg_file.reg_array[24] ),
    .Y(_0389_),
    .A1(net465),
    .A2(net472));
 sg13g2_nand2_1 _1068_ (.Y(_0390_),
    .A(\i2c_slave_controller.out_regf_write_data[0] ),
    .B(_0387_));
 sg13g2_o21ai_1 _1069_ (.B1(_0389_),
    .Y(_0073_),
    .A1(net465),
    .A2(_0390_));
 sg13g2_o21ai_1 _1070_ (.B1(\reg_file.reg_array[25] ),
    .Y(_0391_),
    .A1(net465),
    .A2(_0388_));
 sg13g2_nand2_1 _1071_ (.Y(_0392_),
    .A(\i2c_slave_controller.out_regf_write_data[1] ),
    .B(_0387_));
 sg13g2_o21ai_1 _1072_ (.B1(_0391_),
    .Y(_0074_),
    .A1(net465),
    .A2(_0392_));
 sg13g2_o21ai_1 _1073_ (.B1(\reg_file.reg_array[26] ),
    .Y(_0393_),
    .A1(net465),
    .A2(net471));
 sg13g2_nand2_1 _1074_ (.Y(_0394_),
    .A(\i2c_slave_controller.out_regf_write_data[2] ),
    .B(_0387_));
 sg13g2_o21ai_1 _1075_ (.B1(_0393_),
    .Y(_0075_),
    .A1(net465),
    .A2(_0394_));
 sg13g2_o21ai_1 _1076_ (.B1(\reg_file.reg_array[27] ),
    .Y(_0395_),
    .A1(net461),
    .A2(net472));
 sg13g2_nand2_1 _1077_ (.Y(_0396_),
    .A(\i2c_slave_controller.out_regf_write_data[3] ),
    .B(_0387_));
 sg13g2_o21ai_1 _1078_ (.B1(_0395_),
    .Y(_0076_),
    .A1(net461),
    .A2(_0396_));
 sg13g2_o21ai_1 _1079_ (.B1(\reg_file.reg_array[28] ),
    .Y(_0397_),
    .A1(net466),
    .A2(net471));
 sg13g2_nand2_1 _1080_ (.Y(_0398_),
    .A(\i2c_slave_controller.out_regf_write_data[4] ),
    .B(_0387_));
 sg13g2_o21ai_1 _1081_ (.B1(_0397_),
    .Y(_0077_),
    .A1(net466),
    .A2(_0398_));
 sg13g2_o21ai_1 _1082_ (.B1(\reg_file.reg_array[29] ),
    .Y(_0399_),
    .A1(net466),
    .A2(net471));
 sg13g2_nand2_1 _1083_ (.Y(_0400_),
    .A(\i2c_slave_controller.out_regf_write_data[5] ),
    .B(_0387_));
 sg13g2_o21ai_1 _1084_ (.B1(_0399_),
    .Y(_0078_),
    .A1(net466),
    .A2(_0400_));
 sg13g2_o21ai_1 _1085_ (.B1(\reg_file.reg_array[30] ),
    .Y(_0401_),
    .A1(net461),
    .A2(net472));
 sg13g2_nand2_1 _1086_ (.Y(_0402_),
    .A(\i2c_slave_controller.out_regf_write_data[6] ),
    .B(_0387_));
 sg13g2_o21ai_1 _1087_ (.B1(_0401_),
    .Y(_0079_),
    .A1(net461),
    .A2(_0402_));
 sg13g2_o21ai_1 _1088_ (.B1(\reg_file.reg_array[31] ),
    .Y(_0403_),
    .A1(net461),
    .A2(net472));
 sg13g2_nand2_1 _1089_ (.Y(_0404_),
    .A(\i2c_slave_controller.out_regf_write_data[7] ),
    .B(_0387_));
 sg13g2_o21ai_1 _1090_ (.B1(_0403_),
    .Y(_0080_),
    .A1(net461),
    .A2(_0404_));
 sg13g2_nand4_1 _1091_ (.B(net524),
    .C(net502),
    .A(net515),
    .Y(_0405_),
    .D(net498));
 sg13g2_nand2_1 _1092_ (.Y(_0406_),
    .A(\reg_file.reg_array[32] ),
    .B(_0405_));
 sg13g2_nand2b_1 _1093_ (.Y(_0407_),
    .B(_0363_),
    .A_N(net532));
 sg13g2_nand3b_1 _1094_ (.B(net479),
    .C(_0363_),
    .Y(_0408_),
    .A_N(net532));
 sg13g2_o21ai_1 _1095_ (.B1(_0406_),
    .Y(_0081_),
    .A1(net464),
    .A2(_0408_));
 sg13g2_nand2_1 _1096_ (.Y(_0409_),
    .A(\reg_file.reg_array[33] ),
    .B(_0405_));
 sg13g2_nand2b_1 _1097_ (.Y(_0410_),
    .B(_0366_),
    .A_N(net532));
 sg13g2_nand3b_1 _1098_ (.B(_0326_),
    .C(_0366_),
    .Y(_0411_),
    .A_N(net532));
 sg13g2_o21ai_1 _1099_ (.B1(_0409_),
    .Y(_0082_),
    .A1(net463),
    .A2(_0411_));
 sg13g2_nand2_1 _1100_ (.Y(_0412_),
    .A(\reg_file.reg_array[34] ),
    .B(_0405_));
 sg13g2_nand2b_1 _1101_ (.Y(_0413_),
    .B(_0369_),
    .A_N(net534));
 sg13g2_nand3b_1 _1102_ (.B(net479),
    .C(_0369_),
    .Y(_0414_),
    .A_N(net532));
 sg13g2_o21ai_1 _1103_ (.B1(_0412_),
    .Y(_0083_),
    .A1(net463),
    .A2(_0414_));
 sg13g2_nand2_1 _1104_ (.Y(_0415_),
    .A(\reg_file.reg_array[35] ),
    .B(_0405_));
 sg13g2_nand2b_1 _1105_ (.Y(_0416_),
    .B(_0372_),
    .A_N(net531));
 sg13g2_nand3b_1 _1106_ (.B(net479),
    .C(_0372_),
    .Y(_0417_),
    .A_N(net529));
 sg13g2_o21ai_1 _1107_ (.B1(_0415_),
    .Y(_0084_),
    .A1(net460),
    .A2(_0417_));
 sg13g2_nand2_1 _1108_ (.Y(_0418_),
    .A(\reg_file.reg_array[36] ),
    .B(_0405_));
 sg13g2_nand2b_1 _1109_ (.Y(_0419_),
    .B(_0375_),
    .A_N(net533));
 sg13g2_nand3b_1 _1110_ (.B(net479),
    .C(_0375_),
    .Y(_0420_),
    .A_N(net533));
 sg13g2_o21ai_1 _1111_ (.B1(_0418_),
    .Y(_0085_),
    .A1(net464),
    .A2(_0420_));
 sg13g2_nand2_1 _1112_ (.Y(_0421_),
    .A(\reg_file.reg_array[37] ),
    .B(_0405_));
 sg13g2_nand2b_1 _1113_ (.Y(_0422_),
    .B(_0378_),
    .A_N(net530));
 sg13g2_nand3b_1 _1114_ (.B(net479),
    .C(_0378_),
    .Y(_0423_),
    .A_N(net530));
 sg13g2_o21ai_1 _1115_ (.B1(_0421_),
    .Y(_0086_),
    .A1(net460),
    .A2(_0423_));
 sg13g2_nand2_1 _1116_ (.Y(_0424_),
    .A(\reg_file.reg_array[38] ),
    .B(_0405_));
 sg13g2_nand2b_1 _1117_ (.Y(_0425_),
    .B(_0381_),
    .A_N(net530));
 sg13g2_nand3b_1 _1118_ (.B(net479),
    .C(_0381_),
    .Y(_0426_),
    .A_N(net529));
 sg13g2_o21ai_1 _1119_ (.B1(_0424_),
    .Y(_0087_),
    .A1(net459),
    .A2(_0426_));
 sg13g2_nand2_1 _1120_ (.Y(_0427_),
    .A(\reg_file.reg_array[39] ),
    .B(_0405_));
 sg13g2_nand2b_1 _1121_ (.Y(_0428_),
    .B(_0384_),
    .A_N(net529));
 sg13g2_nand3b_1 _1122_ (.B(net479),
    .C(_0384_),
    .Y(_0429_),
    .A_N(net529));
 sg13g2_o21ai_1 _1123_ (.B1(_0427_),
    .Y(_0088_),
    .A1(net459),
    .A2(_0429_));
 sg13g2_and2_2 _1124_ (.A(net523),
    .B(net490),
    .X(_0430_));
 sg13g2_nand4_1 _1125_ (.B(net524),
    .C(net498),
    .A(net515),
    .Y(_0431_),
    .D(net490));
 sg13g2_nand2_1 _1126_ (.Y(_0432_),
    .A(\reg_file.reg_array[40] ),
    .B(_0431_));
 sg13g2_nand2_1 _1127_ (.Y(_0433_),
    .A(\i2c_slave_controller.out_regf_write_data[0] ),
    .B(_0430_));
 sg13g2_o21ai_1 _1128_ (.B1(_0432_),
    .Y(_0089_),
    .A1(net464),
    .A2(_0433_));
 sg13g2_nand2_1 _1129_ (.Y(_0434_),
    .A(\reg_file.reg_array[41] ),
    .B(_0431_));
 sg13g2_nand2_1 _1130_ (.Y(_0435_),
    .A(\i2c_slave_controller.out_regf_write_data[1] ),
    .B(_0430_));
 sg13g2_o21ai_1 _1131_ (.B1(_0434_),
    .Y(_0090_),
    .A1(net463),
    .A2(_0435_));
 sg13g2_nand2_1 _1132_ (.Y(_0436_),
    .A(\reg_file.reg_array[42] ),
    .B(_0431_));
 sg13g2_nand2_1 _1133_ (.Y(_0437_),
    .A(\i2c_slave_controller.out_regf_write_data[2] ),
    .B(_0430_));
 sg13g2_o21ai_1 _1134_ (.B1(_0436_),
    .Y(_0091_),
    .A1(net463),
    .A2(_0437_));
 sg13g2_nand2_1 _1135_ (.Y(_0438_),
    .A(\reg_file.reg_array[43] ),
    .B(_0431_));
 sg13g2_nand2_1 _1136_ (.Y(_0439_),
    .A(\i2c_slave_controller.out_regf_write_data[3] ),
    .B(_0430_));
 sg13g2_o21ai_1 _1137_ (.B1(_0438_),
    .Y(_0092_),
    .A1(net460),
    .A2(_0439_));
 sg13g2_nand2_1 _1138_ (.Y(_0440_),
    .A(\reg_file.reg_array[44] ),
    .B(_0431_));
 sg13g2_nand2_1 _1139_ (.Y(_0441_),
    .A(\i2c_slave_controller.out_regf_write_data[4] ),
    .B(_0430_));
 sg13g2_o21ai_1 _1140_ (.B1(_0440_),
    .Y(_0093_),
    .A1(net464),
    .A2(_0441_));
 sg13g2_nand2_1 _1141_ (.Y(_0442_),
    .A(\reg_file.reg_array[45] ),
    .B(_0431_));
 sg13g2_nand2_1 _1142_ (.Y(_0443_),
    .A(\i2c_slave_controller.out_regf_write_data[5] ),
    .B(_0430_));
 sg13g2_o21ai_1 _1143_ (.B1(_0442_),
    .Y(_0094_),
    .A1(net462),
    .A2(_0443_));
 sg13g2_nand2_1 _1144_ (.Y(_0444_),
    .A(\reg_file.reg_array[46] ),
    .B(_0431_));
 sg13g2_nand2_1 _1145_ (.Y(_0445_),
    .A(\i2c_slave_controller.out_regf_write_data[6] ),
    .B(_0430_));
 sg13g2_o21ai_1 _1146_ (.B1(_0444_),
    .Y(_0095_),
    .A1(net459),
    .A2(_0445_));
 sg13g2_nand2_1 _1147_ (.Y(_0446_),
    .A(\reg_file.reg_array[47] ),
    .B(_0431_));
 sg13g2_nand2_1 _1148_ (.Y(_0447_),
    .A(\i2c_slave_controller.out_regf_write_data[7] ),
    .B(_0430_));
 sg13g2_o21ai_1 _1149_ (.B1(_0446_),
    .Y(_0096_),
    .A1(net460),
    .A2(_0447_));
 sg13g2_nand4_1 _1150_ (.B(net524),
    .C(net498),
    .A(net515),
    .Y(_0448_),
    .D(net486));
 sg13g2_nand2_1 _1151_ (.Y(_0449_),
    .A(\reg_file.reg_array[48] ),
    .B(_0448_));
 sg13g2_nand3_1 _1152_ (.B(net527),
    .C(_0363_),
    .A(net533),
    .Y(_0450_));
 sg13g2_o21ai_1 _1153_ (.B1(_0449_),
    .Y(_0097_),
    .A1(net467),
    .A2(_0450_));
 sg13g2_nand2_1 _1154_ (.Y(_0451_),
    .A(\reg_file.reg_array[49] ),
    .B(_0448_));
 sg13g2_nand3_1 _1155_ (.B(net526),
    .C(_0366_),
    .A(net532),
    .Y(_0452_));
 sg13g2_o21ai_1 _1156_ (.B1(_0451_),
    .Y(_0098_),
    .A1(net463),
    .A2(_0452_));
 sg13g2_nand2_1 _1157_ (.Y(_0453_),
    .A(\reg_file.reg_array[50] ),
    .B(_0448_));
 sg13g2_nand3_1 _1158_ (.B(net526),
    .C(_0369_),
    .A(net532),
    .Y(_0454_));
 sg13g2_o21ai_1 _1159_ (.B1(_0453_),
    .Y(_0099_),
    .A1(net463),
    .A2(_0454_));
 sg13g2_nand2_1 _1160_ (.Y(_0455_),
    .A(\reg_file.reg_array[51] ),
    .B(_0448_));
 sg13g2_nand3_1 _1161_ (.B(net523),
    .C(_0372_),
    .A(net529),
    .Y(_0456_));
 sg13g2_o21ai_1 _1162_ (.B1(_0455_),
    .Y(_0100_),
    .A1(net459),
    .A2(_0456_));
 sg13g2_nand2_1 _1163_ (.Y(_0457_),
    .A(\reg_file.reg_array[52] ),
    .B(_0448_));
 sg13g2_nand3_1 _1164_ (.B(net526),
    .C(_0375_),
    .A(net533),
    .Y(_0458_));
 sg13g2_o21ai_1 _1165_ (.B1(_0457_),
    .Y(_0101_),
    .A1(net464),
    .A2(_0458_));
 sg13g2_nand2_1 _1166_ (.Y(_0459_),
    .A(\reg_file.reg_array[53] ),
    .B(_0448_));
 sg13g2_nand3_1 _1167_ (.B(net524),
    .C(_0378_),
    .A(net530),
    .Y(_0460_));
 sg13g2_o21ai_1 _1168_ (.B1(_0459_),
    .Y(_0102_),
    .A1(net460),
    .A2(_0460_));
 sg13g2_nand2_1 _1169_ (.Y(_0461_),
    .A(\reg_file.reg_array[54] ),
    .B(_0448_));
 sg13g2_nand3_1 _1170_ (.B(net523),
    .C(_0381_),
    .A(net529),
    .Y(_0462_));
 sg13g2_o21ai_1 _1171_ (.B1(_0461_),
    .Y(_0103_),
    .A1(net459),
    .A2(_0462_));
 sg13g2_nand2_1 _1172_ (.Y(_0463_),
    .A(\reg_file.reg_array[55] ),
    .B(_0448_));
 sg13g2_nand3_1 _1173_ (.B(net523),
    .C(_0384_),
    .A(net529),
    .Y(_0464_));
 sg13g2_o21ai_1 _1174_ (.B1(_0463_),
    .Y(_0104_),
    .A1(net460),
    .A2(_0464_));
 sg13g2_and2_2 _1175_ (.A(net523),
    .B(net480),
    .X(_0465_));
 sg13g2_nand4_1 _1176_ (.B(net524),
    .C(net498),
    .A(net515),
    .Y(_0466_),
    .D(net481));
 sg13g2_nand2_1 _1177_ (.Y(_0467_),
    .A(\reg_file.reg_array[56] ),
    .B(_0466_));
 sg13g2_nand2_1 _1178_ (.Y(_0468_),
    .A(\i2c_slave_controller.out_regf_write_data[0] ),
    .B(_0465_));
 sg13g2_o21ai_1 _1179_ (.B1(_0467_),
    .Y(_0105_),
    .A1(net464),
    .A2(_0468_));
 sg13g2_nand2_1 _1180_ (.Y(_0469_),
    .A(\reg_file.reg_array[57] ),
    .B(_0466_));
 sg13g2_nand2_1 _1181_ (.Y(_0470_),
    .A(\i2c_slave_controller.out_regf_write_data[1] ),
    .B(_0465_));
 sg13g2_o21ai_1 _1182_ (.B1(_0469_),
    .Y(_0106_),
    .A1(net463),
    .A2(_0470_));
 sg13g2_nand2_1 _1183_ (.Y(_0471_),
    .A(\reg_file.reg_array[58] ),
    .B(_0466_));
 sg13g2_nand2_1 _1184_ (.Y(_0472_),
    .A(\i2c_slave_controller.out_regf_write_data[2] ),
    .B(_0465_));
 sg13g2_o21ai_1 _1185_ (.B1(_0471_),
    .Y(_0107_),
    .A1(net463),
    .A2(_0472_));
 sg13g2_nand2_1 _1186_ (.Y(_0473_),
    .A(\reg_file.reg_array[59] ),
    .B(_0466_));
 sg13g2_nand2_1 _1187_ (.Y(_0474_),
    .A(\i2c_slave_controller.out_regf_write_data[3] ),
    .B(_0465_));
 sg13g2_o21ai_1 _1188_ (.B1(_0473_),
    .Y(_0108_),
    .A1(net459),
    .A2(_0474_));
 sg13g2_nand2_1 _1189_ (.Y(_0475_),
    .A(\reg_file.reg_array[60] ),
    .B(_0466_));
 sg13g2_nand2_1 _1190_ (.Y(_0476_),
    .A(\i2c_slave_controller.out_regf_write_data[4] ),
    .B(_0465_));
 sg13g2_o21ai_1 _1191_ (.B1(_0475_),
    .Y(_0109_),
    .A1(net464),
    .A2(_0476_));
 sg13g2_nand2_1 _1192_ (.Y(_0477_),
    .A(\reg_file.reg_array[61] ),
    .B(_0466_));
 sg13g2_nand2_1 _1193_ (.Y(_0478_),
    .A(\i2c_slave_controller.out_regf_write_data[5] ),
    .B(_0465_));
 sg13g2_o21ai_1 _1194_ (.B1(_0477_),
    .Y(_0110_),
    .A1(net460),
    .A2(_0478_));
 sg13g2_nand2_1 _1195_ (.Y(_0479_),
    .A(\reg_file.reg_array[62] ),
    .B(_0466_));
 sg13g2_nand2_1 _1196_ (.Y(_0480_),
    .A(\i2c_slave_controller.out_regf_write_data[6] ),
    .B(_0465_));
 sg13g2_o21ai_1 _1197_ (.B1(_0479_),
    .Y(_0111_),
    .A1(net459),
    .A2(_0480_));
 sg13g2_nand2_1 _1198_ (.Y(_0481_),
    .A(\reg_file.reg_array[63] ),
    .B(_0466_));
 sg13g2_nand2_1 _1199_ (.Y(_0482_),
    .A(\i2c_slave_controller.out_regf_write_data[7] ),
    .B(_0465_));
 sg13g2_o21ai_1 _1200_ (.B1(_0481_),
    .Y(_0112_),
    .A1(net459),
    .A2(_0482_));
 sg13g2_nor3_1 _1201_ (.A(net536),
    .B(_0003_),
    .C(_0330_),
    .Y(_0483_));
 sg13g2_nand4_1 _1202_ (.B(_0343_),
    .C(_0344_),
    .A(net499),
    .Y(_0484_),
    .D(_0483_));
 sg13g2_nand2_1 _1203_ (.Y(_0485_),
    .A(\reg_file.reg_array[64] ),
    .B(_0484_));
 sg13g2_nand2b_2 _1204_ (.Y(_0486_),
    .B(net468),
    .A_N(_0326_));
 sg13g2_o21ai_1 _1205_ (.B1(_0485_),
    .Y(_0113_),
    .A1(_0407_),
    .A2(_0486_));
 sg13g2_nand2_1 _1206_ (.Y(_0487_),
    .A(\reg_file.reg_array[65] ),
    .B(_0484_));
 sg13g2_o21ai_1 _1207_ (.B1(_0487_),
    .Y(_0114_),
    .A1(_0410_),
    .A2(_0486_));
 sg13g2_nand2_1 _1208_ (.Y(_0488_),
    .A(\reg_file.reg_array[66] ),
    .B(_0484_));
 sg13g2_o21ai_1 _1209_ (.B1(_0488_),
    .Y(_0115_),
    .A1(_0413_),
    .A2(_0486_));
 sg13g2_nand2_1 _1210_ (.Y(_0489_),
    .A(\reg_file.reg_array[67] ),
    .B(_0484_));
 sg13g2_o21ai_1 _1211_ (.B1(_0489_),
    .Y(_0116_),
    .A1(_0416_),
    .A2(_0486_));
 sg13g2_nand2_1 _1212_ (.Y(_0490_),
    .A(\reg_file.reg_array[68] ),
    .B(_0484_));
 sg13g2_o21ai_1 _1213_ (.B1(_0490_),
    .Y(_0117_),
    .A1(_0419_),
    .A2(_0486_));
 sg13g2_nand2_1 _1214_ (.Y(_0491_),
    .A(\reg_file.reg_array[69] ),
    .B(_0484_));
 sg13g2_o21ai_1 _1215_ (.B1(_0491_),
    .Y(_0118_),
    .A1(_0422_),
    .A2(_0486_));
 sg13g2_nand2_1 _1216_ (.Y(_0492_),
    .A(\reg_file.reg_array[70] ),
    .B(_0484_));
 sg13g2_o21ai_1 _1217_ (.B1(_0492_),
    .Y(_0119_),
    .A1(_0425_),
    .A2(_0486_));
 sg13g2_nand2_1 _1218_ (.Y(_0493_),
    .A(\reg_file.reg_array[71] ),
    .B(_0484_));
 sg13g2_o21ai_1 _1219_ (.B1(_0493_),
    .Y(_0120_),
    .A1(_0428_),
    .A2(_0486_));
 sg13g2_a21oi_1 _1220_ (.A1(_0343_),
    .A2(_0344_),
    .Y(_0494_),
    .B1(net496));
 sg13g2_nand3_1 _1221_ (.B(_0345_),
    .C(_0346_),
    .A(net499),
    .Y(_0495_));
 sg13g2_and3_2 _1222_ (.X(_0496_),
    .A(net478),
    .B(net475),
    .C(_0494_));
 sg13g2_nand4_1 _1223_ (.B(net477),
    .C(net474),
    .A(\i2c_slave_controller.out_regf_write_data[0] ),
    .Y(_0497_),
    .D(net458));
 sg13g2_o21ai_1 _1224_ (.B1(_0497_),
    .Y(_0121_),
    .A1(_0216_),
    .A2(_0496_));
 sg13g2_nand4_1 _1225_ (.B(net477),
    .C(net474),
    .A(\i2c_slave_controller.out_regf_write_data[1] ),
    .Y(_0498_),
    .D(net458));
 sg13g2_o21ai_1 _1226_ (.B1(_0498_),
    .Y(_0122_),
    .A1(_0217_),
    .A2(_0496_));
 sg13g2_nand4_1 _1227_ (.B(net477),
    .C(net474),
    .A(\i2c_slave_controller.out_regf_write_data[2] ),
    .Y(_0499_),
    .D(net458));
 sg13g2_o21ai_1 _1228_ (.B1(_0499_),
    .Y(_0123_),
    .A1(_0218_),
    .A2(_0496_));
 sg13g2_nand4_1 _1229_ (.B(net476),
    .C(net473),
    .A(\i2c_slave_controller.out_regf_write_data[3] ),
    .Y(_0500_),
    .D(net458));
 sg13g2_o21ai_1 _1230_ (.B1(_0500_),
    .Y(_0124_),
    .A1(_0219_),
    .A2(_0496_));
 sg13g2_nand4_1 _1231_ (.B(net477),
    .C(net474),
    .A(\i2c_slave_controller.out_regf_write_data[4] ),
    .Y(_0501_),
    .D(net458));
 sg13g2_o21ai_1 _1232_ (.B1(_0501_),
    .Y(_0125_),
    .A1(_0220_),
    .A2(_0496_));
 sg13g2_nand4_1 _1233_ (.B(net476),
    .C(net473),
    .A(\i2c_slave_controller.out_regf_write_data[5] ),
    .Y(_0502_),
    .D(net458));
 sg13g2_o21ai_1 _1234_ (.B1(_0502_),
    .Y(_0126_),
    .A1(_0221_),
    .A2(_0496_));
 sg13g2_nand4_1 _1235_ (.B(net476),
    .C(net473),
    .A(\i2c_slave_controller.out_regf_write_data[6] ),
    .Y(_0503_),
    .D(net458));
 sg13g2_o21ai_1 _1236_ (.B1(_0503_),
    .Y(_0127_),
    .A1(_0222_),
    .A2(_0496_));
 sg13g2_nand4_1 _1237_ (.B(net476),
    .C(net473),
    .A(\i2c_slave_controller.out_regf_write_data[7] ),
    .Y(_0504_),
    .D(net458));
 sg13g2_o21ai_1 _1238_ (.B1(_0504_),
    .Y(_0128_),
    .A1(_0223_),
    .A2(_0496_));
 sg13g2_nand4_1 _1239_ (.B(_0345_),
    .C(_0346_),
    .A(net499),
    .Y(_0505_),
    .D(_0359_));
 sg13g2_nand2_1 _1240_ (.Y(_0506_),
    .A(\reg_file.reg_array[80] ),
    .B(_0505_));
 sg13g2_o21ai_1 _1241_ (.B1(_0506_),
    .Y(_0129_),
    .A1(_0364_),
    .A2(net455));
 sg13g2_nand2_1 _1242_ (.Y(_0507_),
    .A(\reg_file.reg_array[81] ),
    .B(_0505_));
 sg13g2_o21ai_1 _1243_ (.B1(_0507_),
    .Y(_0130_),
    .A1(_0367_),
    .A2(net456));
 sg13g2_nand2_1 _1244_ (.Y(_0508_),
    .A(\reg_file.reg_array[82] ),
    .B(_0505_));
 sg13g2_o21ai_1 _1245_ (.B1(_0508_),
    .Y(_0131_),
    .A1(_0370_),
    .A2(net455));
 sg13g2_nand2_1 _1246_ (.Y(_0509_),
    .A(\reg_file.reg_array[83] ),
    .B(_0505_));
 sg13g2_o21ai_1 _1247_ (.B1(_0509_),
    .Y(_0132_),
    .A1(_0373_),
    .A2(net449));
 sg13g2_nand2_1 _1248_ (.Y(_0510_),
    .A(\reg_file.reg_array[84] ),
    .B(_0505_));
 sg13g2_o21ai_1 _1249_ (.B1(_0510_),
    .Y(_0133_),
    .A1(_0376_),
    .A2(net457));
 sg13g2_nand2_1 _1250_ (.Y(_0511_),
    .A(\reg_file.reg_array[85] ),
    .B(_0505_));
 sg13g2_o21ai_1 _1251_ (.B1(_0511_),
    .Y(_0134_),
    .A1(_0379_),
    .A2(net452));
 sg13g2_nand2_1 _1252_ (.Y(_0512_),
    .A(\reg_file.reg_array[86] ),
    .B(_0505_));
 sg13g2_o21ai_1 _1253_ (.B1(_0512_),
    .Y(_0135_),
    .A1(_0382_),
    .A2(net452));
 sg13g2_nand2_1 _1254_ (.Y(_0513_),
    .A(\reg_file.reg_array[87] ),
    .B(_0505_));
 sg13g2_o21ai_1 _1255_ (.B1(_0513_),
    .Y(_0136_),
    .A1(_0385_),
    .A2(net449));
 sg13g2_o21ai_1 _1256_ (.B1(\reg_file.reg_array[88] ),
    .Y(_0514_),
    .A1(net471),
    .A2(net455));
 sg13g2_o21ai_1 _1257_ (.B1(_0514_),
    .Y(_0137_),
    .A1(_0390_),
    .A2(net455));
 sg13g2_o21ai_1 _1258_ (.B1(\reg_file.reg_array[89] ),
    .Y(_0515_),
    .A1(net471),
    .A2(net455));
 sg13g2_o21ai_1 _1259_ (.B1(_0515_),
    .Y(_0138_),
    .A1(_0392_),
    .A2(net455));
 sg13g2_o21ai_1 _1260_ (.B1(\reg_file.reg_array[90] ),
    .Y(_0516_),
    .A1(net471),
    .A2(net455));
 sg13g2_o21ai_1 _1261_ (.B1(_0516_),
    .Y(_0139_),
    .A1(_0394_),
    .A2(net455));
 sg13g2_o21ai_1 _1262_ (.B1(\reg_file.reg_array[91] ),
    .Y(_0517_),
    .A1(net472),
    .A2(net449));
 sg13g2_o21ai_1 _1263_ (.B1(_0517_),
    .Y(_0140_),
    .A1(_0396_),
    .A2(net449));
 sg13g2_o21ai_1 _1264_ (.B1(\reg_file.reg_array[92] ),
    .Y(_0518_),
    .A1(net471),
    .A2(net453));
 sg13g2_o21ai_1 _1265_ (.B1(_0518_),
    .Y(_0141_),
    .A1(_0398_),
    .A2(net453));
 sg13g2_o21ai_1 _1266_ (.B1(\reg_file.reg_array[93] ),
    .Y(_0519_),
    .A1(net471),
    .A2(net457));
 sg13g2_o21ai_1 _1267_ (.B1(_0519_),
    .Y(_0142_),
    .A1(_0400_),
    .A2(net457));
 sg13g2_o21ai_1 _1268_ (.B1(\reg_file.reg_array[94] ),
    .Y(_0520_),
    .A1(net472),
    .A2(net449));
 sg13g2_o21ai_1 _1269_ (.B1(_0520_),
    .Y(_0143_),
    .A1(_0402_),
    .A2(net449));
 sg13g2_o21ai_1 _1270_ (.B1(\reg_file.reg_array[95] ),
    .Y(_0521_),
    .A1(net472),
    .A2(net449));
 sg13g2_o21ai_1 _1271_ (.B1(_0521_),
    .Y(_0144_),
    .A1(_0404_),
    .A2(net449));
 sg13g2_nand4_1 _1272_ (.B(net526),
    .C(net503),
    .A(net521),
    .Y(_0522_),
    .D(net498));
 sg13g2_nand2_1 _1273_ (.Y(_0523_),
    .A(\reg_file.reg_array[96] ),
    .B(_0522_));
 sg13g2_o21ai_1 _1274_ (.B1(_0523_),
    .Y(_0145_),
    .A1(_0408_),
    .A2(net454));
 sg13g2_nand2_1 _1275_ (.Y(_0524_),
    .A(\reg_file.reg_array[97] ),
    .B(_0522_));
 sg13g2_o21ai_1 _1276_ (.B1(_0524_),
    .Y(_0146_),
    .A1(_0411_),
    .A2(net456));
 sg13g2_nand2_1 _1277_ (.Y(_0525_),
    .A(\reg_file.reg_array[98] ),
    .B(_0522_));
 sg13g2_o21ai_1 _1278_ (.B1(_0525_),
    .Y(_0147_),
    .A1(_0414_),
    .A2(net454));
 sg13g2_nand2_1 _1279_ (.Y(_0526_),
    .A(\reg_file.reg_array[99] ),
    .B(_0522_));
 sg13g2_o21ai_1 _1280_ (.B1(_0526_),
    .Y(_0148_),
    .A1(_0417_),
    .A2(net451));
 sg13g2_nand2_1 _1281_ (.Y(_0527_),
    .A(\reg_file.reg_array[100] ),
    .B(_0522_));
 sg13g2_o21ai_1 _1282_ (.B1(_0527_),
    .Y(_0149_),
    .A1(_0420_),
    .A2(net453));
 sg13g2_nand2_1 _1283_ (.Y(_0528_),
    .A(\reg_file.reg_array[101] ),
    .B(_0522_));
 sg13g2_o21ai_1 _1284_ (.B1(_0528_),
    .Y(_0150_),
    .A1(_0423_),
    .A2(net451));
 sg13g2_nand2_1 _1285_ (.Y(_0529_),
    .A(\reg_file.reg_array[102] ),
    .B(_0522_));
 sg13g2_o21ai_1 _1286_ (.B1(_0529_),
    .Y(_0151_),
    .A1(_0426_),
    .A2(net450));
 sg13g2_nand2_1 _1287_ (.Y(_0530_),
    .A(\reg_file.reg_array[103] ),
    .B(_0522_));
 sg13g2_o21ai_1 _1288_ (.B1(_0530_),
    .Y(_0152_),
    .A1(_0429_),
    .A2(net450));
 sg13g2_nand4_1 _1289_ (.B(net526),
    .C(net498),
    .A(net521),
    .Y(_0531_),
    .D(net492));
 sg13g2_nand2_1 _1290_ (.Y(_0532_),
    .A(\reg_file.reg_array[104] ),
    .B(_0531_));
 sg13g2_o21ai_1 _1291_ (.B1(_0532_),
    .Y(_0153_),
    .A1(_0433_),
    .A2(net454));
 sg13g2_nand2_1 _1292_ (.Y(_0533_),
    .A(\reg_file.reg_array[105] ),
    .B(_0531_));
 sg13g2_o21ai_1 _1293_ (.B1(_0533_),
    .Y(_0154_),
    .A1(_0435_),
    .A2(net454));
 sg13g2_nand2_1 _1294_ (.Y(_0534_),
    .A(\reg_file.reg_array[106] ),
    .B(_0531_));
 sg13g2_o21ai_1 _1295_ (.B1(_0534_),
    .Y(_0155_),
    .A1(_0437_),
    .A2(net454));
 sg13g2_nand2_1 _1296_ (.Y(_0535_),
    .A(\reg_file.reg_array[107] ),
    .B(_0531_));
 sg13g2_o21ai_1 _1297_ (.B1(_0535_),
    .Y(_0156_),
    .A1(_0439_),
    .A2(net451));
 sg13g2_nand2_1 _1298_ (.Y(_0536_),
    .A(\reg_file.reg_array[108] ),
    .B(_0531_));
 sg13g2_o21ai_1 _1299_ (.B1(_0536_),
    .Y(_0157_),
    .A1(_0441_),
    .A2(net453));
 sg13g2_nand2_1 _1300_ (.Y(_0537_),
    .A(\reg_file.reg_array[109] ),
    .B(_0531_));
 sg13g2_o21ai_1 _1301_ (.B1(_0537_),
    .Y(_0158_),
    .A1(_0443_),
    .A2(net451));
 sg13g2_nand2_1 _1302_ (.Y(_0538_),
    .A(\reg_file.reg_array[110] ),
    .B(_0531_));
 sg13g2_o21ai_1 _1303_ (.B1(_0538_),
    .Y(_0159_),
    .A1(_0445_),
    .A2(net450));
 sg13g2_nand2_1 _1304_ (.Y(_0539_),
    .A(\reg_file.reg_array[111] ),
    .B(_0531_));
 sg13g2_o21ai_1 _1305_ (.B1(_0539_),
    .Y(_0160_),
    .A1(_0447_),
    .A2(net450));
 sg13g2_nand4_1 _1306_ (.B(net526),
    .C(net498),
    .A(net521),
    .Y(_0540_),
    .D(net487));
 sg13g2_nand2_1 _1307_ (.Y(_0541_),
    .A(\reg_file.reg_array[112] ),
    .B(_0540_));
 sg13g2_o21ai_1 _1308_ (.B1(_0541_),
    .Y(_0161_),
    .A1(_0450_),
    .A2(net454));
 sg13g2_nand2_1 _1309_ (.Y(_0542_),
    .A(\reg_file.reg_array[113] ),
    .B(_0540_));
 sg13g2_o21ai_1 _1310_ (.B1(_0542_),
    .Y(_0162_),
    .A1(_0452_),
    .A2(net456));
 sg13g2_nand2_1 _1311_ (.Y(_0543_),
    .A(\reg_file.reg_array[114] ),
    .B(_0540_));
 sg13g2_o21ai_1 _1312_ (.B1(_0543_),
    .Y(_0163_),
    .A1(_0454_),
    .A2(net454));
 sg13g2_nand2_1 _1313_ (.Y(_0544_),
    .A(\reg_file.reg_array[115] ),
    .B(_0540_));
 sg13g2_o21ai_1 _1314_ (.B1(_0544_),
    .Y(_0164_),
    .A1(_0456_),
    .A2(net451));
 sg13g2_nand2_1 _1315_ (.Y(_0545_),
    .A(\reg_file.reg_array[116] ),
    .B(_0540_));
 sg13g2_o21ai_1 _1316_ (.B1(_0545_),
    .Y(_0165_),
    .A1(_0458_),
    .A2(net453));
 sg13g2_nand2_1 _1317_ (.Y(_0546_),
    .A(\reg_file.reg_array[117] ),
    .B(_0540_));
 sg13g2_o21ai_1 _1318_ (.B1(_0546_),
    .Y(_0166_),
    .A1(_0460_),
    .A2(net451));
 sg13g2_nand2_1 _1319_ (.Y(_0547_),
    .A(\reg_file.reg_array[118] ),
    .B(_0540_));
 sg13g2_o21ai_1 _1320_ (.B1(_0547_),
    .Y(_0167_),
    .A1(_0462_),
    .A2(net450));
 sg13g2_nand2_1 _1321_ (.Y(_0548_),
    .A(\reg_file.reg_array[119] ),
    .B(_0540_));
 sg13g2_o21ai_1 _1322_ (.B1(_0548_),
    .Y(_0168_),
    .A1(_0464_),
    .A2(net450));
 sg13g2_nand4_1 _1323_ (.B(net526),
    .C(net498),
    .A(net521),
    .Y(_0549_),
    .D(net483));
 sg13g2_nand2_1 _1324_ (.Y(_0550_),
    .A(\reg_file.reg_array[120] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1325_ (.B1(_0550_),
    .Y(_0169_),
    .A1(_0468_),
    .A2(net453));
 sg13g2_nand2_1 _1326_ (.Y(_0551_),
    .A(\reg_file.reg_array[121] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1327_ (.B1(_0551_),
    .Y(_0170_),
    .A1(_0470_),
    .A2(net453));
 sg13g2_nand2_1 _1328_ (.Y(_0552_),
    .A(\reg_file.reg_array[122] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1329_ (.B1(_0552_),
    .Y(_0171_),
    .A1(_0472_),
    .A2(net454));
 sg13g2_nand2_1 _1330_ (.Y(_0553_),
    .A(\reg_file.reg_array[123] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1331_ (.B1(_0553_),
    .Y(_0172_),
    .A1(_0474_),
    .A2(net451));
 sg13g2_nand2_1 _1332_ (.Y(_0554_),
    .A(\reg_file.reg_array[124] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1333_ (.B1(_0554_),
    .Y(_0173_),
    .A1(_0476_),
    .A2(net453));
 sg13g2_nand2_1 _1334_ (.Y(_0555_),
    .A(\reg_file.reg_array[125] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1335_ (.B1(_0555_),
    .Y(_0174_),
    .A1(_0478_),
    .A2(net451));
 sg13g2_nand2_1 _1336_ (.Y(_0556_),
    .A(\reg_file.reg_array[126] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1337_ (.B1(_0556_),
    .Y(_0175_),
    .A1(_0480_),
    .A2(net450));
 sg13g2_nand2_1 _1338_ (.Y(_0557_),
    .A(\reg_file.reg_array[127] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1339_ (.B1(_0557_),
    .Y(_0176_),
    .A1(_0482_),
    .A2(net450));
 sg13g2_nor2_1 _1340_ (.A(uo_out[0]),
    .B(net497),
    .Y(_0558_));
 sg13g2_a22oi_1 _1341_ (.Y(_0559_),
    .B1(_0386_),
    .B2(\reg_file.reg_array[88] ),
    .A2(net493),
    .A1(\reg_file.reg_array[72] ));
 sg13g2_a221oi_1 _1342_ (.B2(\reg_file.reg_array[80] ),
    .C1(net527),
    .B1(net489),
    .A1(\reg_file.reg_array[64] ),
    .Y(_0560_),
    .A2(net505));
 sg13g2_a22oi_1 _1343_ (.Y(_0561_),
    .B1(net483),
    .B2(\reg_file.reg_array[120] ),
    .A2(net488),
    .A1(\reg_file.reg_array[112] ));
 sg13g2_a221oi_1 _1344_ (.B2(\reg_file.reg_array[104] ),
    .C1(net512),
    .B1(net494),
    .A1(\reg_file.reg_array[96] ),
    .Y(_0562_),
    .A2(net504));
 sg13g2_a22oi_1 _1345_ (.Y(_0563_),
    .B1(_0561_),
    .B2(_0562_),
    .A2(_0560_),
    .A1(_0559_));
 sg13g2_nand2_1 _1346_ (.Y(_0564_),
    .A(\reg_file.reg_array[32] ),
    .B(net504));
 sg13g2_a21oi_1 _1347_ (.A1(\reg_file.reg_array[56] ),
    .A2(net484),
    .Y(_0565_),
    .B1(net512));
 sg13g2_a22oi_1 _1348_ (.Y(_0566_),
    .B1(net487),
    .B2(\reg_file.reg_array[48] ),
    .A2(net492),
    .A1(\reg_file.reg_array[40] ));
 sg13g2_nand3_1 _1349_ (.B(_0565_),
    .C(_0566_),
    .A(_0564_),
    .Y(_0567_));
 sg13g2_a22oi_1 _1350_ (.Y(_0568_),
    .B1(net489),
    .B2(\reg_file.reg_array[16] ),
    .A2(net493),
    .A1(\reg_file.reg_array[8] ));
 sg13g2_a221oi_1 _1351_ (.B2(\reg_file.reg_array[24] ),
    .C1(net528),
    .B1(net484),
    .A1(\reg_file.reg_array[0] ),
    .Y(_0569_),
    .A2(net505));
 sg13g2_a21oi_1 _1352_ (.A1(_0568_),
    .A2(_0569_),
    .Y(_0570_),
    .B1(net522));
 sg13g2_a22oi_1 _1353_ (.Y(_0571_),
    .B1(_0567_),
    .B2(_0570_),
    .A2(_0563_),
    .A1(\reg_file.reg_pointer[3] ));
 sg13g2_a21oi_1 _1354_ (.A1(net497),
    .A2(_0571_),
    .Y(_0177_),
    .B1(_0558_));
 sg13g2_nor2_1 _1355_ (.A(uo_out[1]),
    .B(net497),
    .Y(_0572_));
 sg13g2_a22oi_1 _1356_ (.Y(_0573_),
    .B1(net494),
    .B2(\reg_file.reg_array[73] ),
    .A2(net505),
    .A1(\reg_file.reg_array[65] ));
 sg13g2_a221oi_1 _1357_ (.B2(\reg_file.reg_array[89] ),
    .C1(net528),
    .B1(net484),
    .A1(\reg_file.reg_array[81] ),
    .Y(_0574_),
    .A2(net488));
 sg13g2_a22oi_1 _1358_ (.Y(_0575_),
    .B1(net483),
    .B2(\reg_file.reg_array[121] ),
    .A2(net492),
    .A1(\reg_file.reg_array[105] ));
 sg13g2_a221oi_1 _1359_ (.B2(\reg_file.reg_array[113] ),
    .C1(net512),
    .B1(net487),
    .A1(\reg_file.reg_array[97] ),
    .Y(_0576_),
    .A2(net503));
 sg13g2_a22oi_1 _1360_ (.Y(_0577_),
    .B1(_0575_),
    .B2(_0576_),
    .A2(_0574_),
    .A1(_0573_));
 sg13g2_nand2_1 _1361_ (.Y(_0578_),
    .A(\reg_file.reg_array[49] ),
    .B(net487));
 sg13g2_a21oi_1 _1362_ (.A1(\reg_file.reg_array[57] ),
    .A2(net483),
    .Y(_0579_),
    .B1(net512));
 sg13g2_a22oi_1 _1363_ (.Y(_0580_),
    .B1(net492),
    .B2(\reg_file.reg_array[41] ),
    .A2(net503),
    .A1(\reg_file.reg_array[33] ));
 sg13g2_nand3_1 _1364_ (.B(_0579_),
    .C(_0580_),
    .A(_0578_),
    .Y(_0581_));
 sg13g2_and3_1 _1365_ (.X(_0582_),
    .A(\reg_file.reg_pointer[0] ),
    .B(net534),
    .C(\reg_file.reg_array[25] ));
 sg13g2_a221oi_1 _1366_ (.B2(\reg_file.reg_array[17] ),
    .C1(_0582_),
    .B1(net488),
    .A1(\reg_file.reg_array[9] ),
    .Y(_0583_),
    .A2(net493));
 sg13g2_a21oi_1 _1367_ (.A1(\reg_file.reg_array[1] ),
    .A2(net504),
    .Y(_0584_),
    .B1(net527));
 sg13g2_a21oi_1 _1368_ (.A1(_0583_),
    .A2(_0584_),
    .Y(_0585_),
    .B1(\reg_file.reg_pointer[3] ));
 sg13g2_a22oi_1 _1369_ (.Y(_0586_),
    .B1(_0581_),
    .B2(_0585_),
    .A2(_0577_),
    .A1(net522));
 sg13g2_a21oi_1 _1370_ (.A1(net497),
    .A2(_0586_),
    .Y(_0178_),
    .B1(_0572_));
 sg13g2_a22oi_1 _1371_ (.Y(_0587_),
    .B1(net493),
    .B2(\reg_file.reg_array[74] ),
    .A2(net504),
    .A1(\reg_file.reg_array[66] ));
 sg13g2_a221oi_1 _1372_ (.B2(\reg_file.reg_array[90] ),
    .C1(net527),
    .B1(net484),
    .A1(\reg_file.reg_array[82] ),
    .Y(_0588_),
    .A2(net488));
 sg13g2_nand2_1 _1373_ (.Y(_0589_),
    .A(_0587_),
    .B(_0588_));
 sg13g2_nand2_1 _1374_ (.Y(_0590_),
    .A(\reg_file.reg_array[106] ),
    .B(net492));
 sg13g2_a21oi_1 _1375_ (.A1(\reg_file.reg_array[114] ),
    .A2(net487),
    .Y(_0591_),
    .B1(net512));
 sg13g2_a22oi_1 _1376_ (.Y(_0592_),
    .B1(net483),
    .B2(\reg_file.reg_array[122] ),
    .A2(net503),
    .A1(\reg_file.reg_array[98] ));
 sg13g2_nand3_1 _1377_ (.B(_0591_),
    .C(_0592_),
    .A(_0590_),
    .Y(_0593_));
 sg13g2_nand3_1 _1378_ (.B(_0589_),
    .C(_0593_),
    .A(net522),
    .Y(_0594_));
 sg13g2_nand2_1 _1379_ (.Y(_0595_),
    .A(\reg_file.reg_array[58] ),
    .B(net483));
 sg13g2_a21oi_1 _1380_ (.A1(\reg_file.reg_array[50] ),
    .A2(net487),
    .Y(_0596_),
    .B1(net512));
 sg13g2_a22oi_1 _1381_ (.Y(_0597_),
    .B1(net492),
    .B2(\reg_file.reg_array[42] ),
    .A2(net503),
    .A1(\reg_file.reg_array[34] ));
 sg13g2_nand3_1 _1382_ (.B(_0596_),
    .C(_0597_),
    .A(_0595_),
    .Y(_0598_));
 sg13g2_a22oi_1 _1383_ (.Y(_0599_),
    .B1(net488),
    .B2(\reg_file.reg_array[18] ),
    .A2(net493),
    .A1(\reg_file.reg_array[10] ));
 sg13g2_a221oi_1 _1384_ (.B2(\reg_file.reg_array[26] ),
    .C1(net527),
    .B1(net484),
    .A1(\reg_file.reg_array[2] ),
    .Y(_0600_),
    .A2(net504));
 sg13g2_a21oi_1 _1385_ (.A1(_0599_),
    .A2(_0600_),
    .Y(_0601_),
    .B1(net522));
 sg13g2_a21oi_1 _1386_ (.A1(_0598_),
    .A2(_0601_),
    .Y(_0602_),
    .B1(net500));
 sg13g2_a22oi_1 _1387_ (.Y(_0179_),
    .B1(_0594_),
    .B2(_0602_),
    .A2(net500),
    .A1(_0224_));
 sg13g2_a22oi_1 _1388_ (.Y(_0603_),
    .B1(net485),
    .B2(\reg_file.reg_array[51] ),
    .A2(net490),
    .A1(\reg_file.reg_array[43] ));
 sg13g2_a221oi_1 _1389_ (.B2(\reg_file.reg_array[59] ),
    .C1(net510),
    .B1(net480),
    .A1(\reg_file.reg_array[35] ),
    .Y(_0604_),
    .A2(net501));
 sg13g2_nand2_1 _1390_ (.Y(_0605_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_nand2_1 _1391_ (.Y(_0606_),
    .A(\reg_file.reg_array[27] ),
    .B(net482));
 sg13g2_a21oi_1 _1392_ (.A1(\reg_file.reg_array[11] ),
    .A2(net495),
    .Y(_0607_),
    .B1(net525));
 sg13g2_a22oi_1 _1393_ (.Y(_0608_),
    .B1(net489),
    .B2(\reg_file.reg_array[19] ),
    .A2(net505),
    .A1(\reg_file.reg_array[3] ));
 sg13g2_nand3_1 _1394_ (.B(_0607_),
    .C(_0608_),
    .A(_0606_),
    .Y(_0609_));
 sg13g2_nand3_1 _1395_ (.B(_0605_),
    .C(_0609_),
    .A(net516),
    .Y(_0610_));
 sg13g2_nand2_1 _1396_ (.Y(_0611_),
    .A(\reg_file.reg_array[115] ),
    .B(net486));
 sg13g2_a21oi_1 _1397_ (.A1(\reg_file.reg_array[123] ),
    .A2(net481),
    .Y(_0612_),
    .B1(net510));
 sg13g2_a22oi_1 _1398_ (.Y(_0613_),
    .B1(net490),
    .B2(\reg_file.reg_array[107] ),
    .A2(net502),
    .A1(\reg_file.reg_array[99] ));
 sg13g2_nand3_1 _1399_ (.B(_0612_),
    .C(_0613_),
    .A(_0611_),
    .Y(_0614_));
 sg13g2_and3_1 _1400_ (.X(_0615_),
    .A(net536),
    .B(net531),
    .C(\reg_file.reg_array[91] ));
 sg13g2_a221oi_1 _1401_ (.B2(\reg_file.reg_array[83] ),
    .C1(_0615_),
    .B1(net486),
    .A1(\reg_file.reg_array[75] ),
    .Y(_0616_),
    .A2(net495));
 sg13g2_a21oi_1 _1402_ (.A1(\reg_file.reg_array[67] ),
    .A2(net505),
    .Y(_0617_),
    .B1(net528));
 sg13g2_a21oi_1 _1403_ (.A1(_0616_),
    .A2(_0617_),
    .Y(_0618_),
    .B1(net516));
 sg13g2_a21oi_1 _1404_ (.A1(_0614_),
    .A2(_0618_),
    .Y(_0619_),
    .B1(net499));
 sg13g2_a22oi_1 _1405_ (.Y(_0180_),
    .B1(_0610_),
    .B2(_0619_),
    .A2(net499),
    .A1(_0225_));
 sg13g2_a22oi_1 _1406_ (.Y(_0620_),
    .B1(net488),
    .B2(\reg_file.reg_array[84] ),
    .A2(net493),
    .A1(\reg_file.reg_array[76] ));
 sg13g2_a221oi_1 _1407_ (.B2(\reg_file.reg_array[92] ),
    .C1(net527),
    .B1(net484),
    .A1(\reg_file.reg_array[68] ),
    .Y(_0621_),
    .A2(net504));
 sg13g2_nand2_1 _1408_ (.Y(_0622_),
    .A(_0620_),
    .B(_0621_));
 sg13g2_nand2_1 _1409_ (.Y(_0623_),
    .A(\reg_file.reg_array[124] ),
    .B(net483));
 sg13g2_a21oi_1 _1410_ (.A1(\reg_file.reg_array[108] ),
    .A2(net492),
    .Y(_0624_),
    .B1(net512));
 sg13g2_a22oi_1 _1411_ (.Y(_0625_),
    .B1(net487),
    .B2(\reg_file.reg_array[116] ),
    .A2(net503),
    .A1(\reg_file.reg_array[100] ));
 sg13g2_nand3_1 _1412_ (.B(_0624_),
    .C(_0625_),
    .A(_0623_),
    .Y(_0626_));
 sg13g2_nand3_1 _1413_ (.B(_0622_),
    .C(_0626_),
    .A(net522),
    .Y(_0627_));
 sg13g2_nand2_1 _1414_ (.Y(_0628_),
    .A(\reg_file.reg_array[52] ),
    .B(net487));
 sg13g2_a21oi_1 _1415_ (.A1(\reg_file.reg_array[36] ),
    .A2(net503),
    .Y(_0629_),
    .B1(net512));
 sg13g2_a22oi_1 _1416_ (.Y(_0630_),
    .B1(net483),
    .B2(\reg_file.reg_array[60] ),
    .A2(net492),
    .A1(\reg_file.reg_array[44] ));
 sg13g2_nand3_1 _1417_ (.B(_0629_),
    .C(_0630_),
    .A(_0628_),
    .Y(_0631_));
 sg13g2_and3_1 _1418_ (.X(_0632_),
    .A(\reg_file.reg_pointer[0] ),
    .B(net535),
    .C(\reg_file.reg_array[28] ));
 sg13g2_a221oi_1 _1419_ (.B2(\reg_file.reg_array[20] ),
    .C1(_0632_),
    .B1(net488),
    .A1(\reg_file.reg_array[12] ),
    .Y(_0633_),
    .A2(net493));
 sg13g2_a21oi_1 _1420_ (.A1(\reg_file.reg_array[4] ),
    .A2(net504),
    .Y(_0634_),
    .B1(net528));
 sg13g2_a21oi_1 _1421_ (.A1(_0633_),
    .A2(_0634_),
    .Y(_0635_),
    .B1(net521));
 sg13g2_a21oi_1 _1422_ (.A1(_0631_),
    .A2(_0635_),
    .Y(_0636_),
    .B1(net500));
 sg13g2_a22oi_1 _1423_ (.Y(_0181_),
    .B1(_0627_),
    .B2(_0636_),
    .A2(net499),
    .A1(_0226_));
 sg13g2_nor2_1 _1424_ (.A(uo_out[5]),
    .B(net496),
    .Y(_0637_));
 sg13g2_a22oi_1 _1425_ (.Y(_0638_),
    .B1(net491),
    .B2(\reg_file.reg_array[77] ),
    .A2(net501),
    .A1(\reg_file.reg_array[69] ));
 sg13g2_a221oi_1 _1426_ (.B2(\reg_file.reg_array[93] ),
    .C1(net523),
    .B1(net481),
    .A1(\reg_file.reg_array[85] ),
    .Y(_0639_),
    .A2(net485));
 sg13g2_a22oi_1 _1427_ (.Y(_0640_),
    .B1(net481),
    .B2(\reg_file.reg_array[125] ),
    .A2(net491),
    .A1(\reg_file.reg_array[109] ));
 sg13g2_a221oi_1 _1428_ (.B2(\reg_file.reg_array[117] ),
    .C1(net510),
    .B1(net485),
    .A1(\reg_file.reg_array[101] ),
    .Y(_0641_),
    .A2(net501));
 sg13g2_a22oi_1 _1429_ (.Y(_0642_),
    .B1(_0640_),
    .B2(_0641_),
    .A2(_0639_),
    .A1(_0638_));
 sg13g2_nand2_1 _1430_ (.Y(_0643_),
    .A(\reg_file.reg_array[45] ),
    .B(net491));
 sg13g2_a21oi_1 _1431_ (.A1(\reg_file.reg_array[61] ),
    .A2(net481),
    .Y(_0644_),
    .B1(net510));
 sg13g2_a22oi_1 _1432_ (.Y(_0645_),
    .B1(net485),
    .B2(\reg_file.reg_array[53] ),
    .A2(net502),
    .A1(\reg_file.reg_array[37] ));
 sg13g2_nand3_1 _1433_ (.B(_0644_),
    .C(_0645_),
    .A(_0643_),
    .Y(_0646_));
 sg13g2_a22oi_1 _1434_ (.Y(_0647_),
    .B1(net482),
    .B2(\reg_file.reg_array[29] ),
    .A2(net493),
    .A1(\reg_file.reg_array[13] ));
 sg13g2_a221oi_1 _1435_ (.B2(\reg_file.reg_array[21] ),
    .C1(net525),
    .B1(net486),
    .A1(\reg_file.reg_array[5] ),
    .Y(_0648_),
    .A2(net502));
 sg13g2_a21oi_1 _1436_ (.A1(_0647_),
    .A2(_0648_),
    .Y(_0649_),
    .B1(net521));
 sg13g2_a22oi_1 _1437_ (.Y(_0650_),
    .B1(_0646_),
    .B2(_0649_),
    .A2(_0642_),
    .A1(net521));
 sg13g2_a21oi_1 _1438_ (.A1(net496),
    .A2(_0650_),
    .Y(_0182_),
    .B1(_0637_));
 sg13g2_nor2_1 _1439_ (.A(uo_out[6]),
    .B(net496),
    .Y(_0651_));
 sg13g2_a22oi_1 _1440_ (.Y(_0652_),
    .B1(net491),
    .B2(\reg_file.reg_array[14] ),
    .A2(net502),
    .A1(\reg_file.reg_array[6] ));
 sg13g2_a221oi_1 _1441_ (.B2(\reg_file.reg_array[30] ),
    .C1(net523),
    .B1(net480),
    .A1(\reg_file.reg_array[22] ),
    .Y(_0653_),
    .A2(net489));
 sg13g2_a22oi_1 _1442_ (.Y(_0654_),
    .B1(net480),
    .B2(\reg_file.reg_array[62] ),
    .A2(net490),
    .A1(\reg_file.reg_array[46] ));
 sg13g2_a221oi_1 _1443_ (.B2(\reg_file.reg_array[54] ),
    .C1(net510),
    .B1(net485),
    .A1(\reg_file.reg_array[38] ),
    .Y(_0655_),
    .A2(net501));
 sg13g2_a22oi_1 _1444_ (.Y(_0656_),
    .B1(_0654_),
    .B2(_0655_),
    .A2(_0653_),
    .A1(_0652_));
 sg13g2_nand2_1 _1445_ (.Y(_0657_),
    .A(\reg_file.reg_array[102] ),
    .B(net501));
 sg13g2_a21oi_1 _1446_ (.A1(\reg_file.reg_array[126] ),
    .A2(net480),
    .Y(_0658_),
    .B1(net510));
 sg13g2_a22oi_1 _1447_ (.Y(_0659_),
    .B1(net485),
    .B2(\reg_file.reg_array[118] ),
    .A2(net490),
    .A1(\reg_file.reg_array[110] ));
 sg13g2_nand3_1 _1448_ (.B(_0658_),
    .C(_0659_),
    .A(_0657_),
    .Y(_0660_));
 sg13g2_a22oi_1 _1449_ (.Y(_0661_),
    .B1(net480),
    .B2(\reg_file.reg_array[94] ),
    .A2(net501),
    .A1(\reg_file.reg_array[70] ));
 sg13g2_a221oi_1 _1450_ (.B2(\reg_file.reg_array[86] ),
    .C1(net523),
    .B1(net486),
    .A1(\reg_file.reg_array[78] ),
    .Y(_0662_),
    .A2(net491));
 sg13g2_a21oi_1 _1451_ (.A1(_0661_),
    .A2(_0662_),
    .Y(_0663_),
    .B1(net515));
 sg13g2_a22oi_1 _1452_ (.Y(_0664_),
    .B1(_0660_),
    .B2(_0663_),
    .A2(_0656_),
    .A1(net515));
 sg13g2_a21oi_1 _1453_ (.A1(net496),
    .A2(_0664_),
    .Y(_0183_),
    .B1(_0651_));
 sg13g2_nor2_1 _1454_ (.A(uo_out[7]),
    .B(net496),
    .Y(_0665_));
 sg13g2_a22oi_1 _1455_ (.Y(_0666_),
    .B1(net482),
    .B2(\reg_file.reg_array[31] ),
    .A2(net502),
    .A1(\reg_file.reg_array[7] ));
 sg13g2_a221oi_1 _1456_ (.B2(\reg_file.reg_array[23] ),
    .C1(net525),
    .B1(net489),
    .A1(\reg_file.reg_array[15] ),
    .Y(_0667_),
    .A2(net491));
 sg13g2_a22oi_1 _1457_ (.Y(_0668_),
    .B1(net480),
    .B2(\reg_file.reg_array[63] ),
    .A2(net485),
    .A1(\reg_file.reg_array[55] ));
 sg13g2_a221oi_1 _1458_ (.B2(\reg_file.reg_array[47] ),
    .C1(net510),
    .B1(net490),
    .A1(\reg_file.reg_array[39] ),
    .Y(_0669_),
    .A2(net501));
 sg13g2_a22oi_1 _1459_ (.Y(_0670_),
    .B1(_0668_),
    .B2(_0669_),
    .A2(_0667_),
    .A1(_0666_));
 sg13g2_nand2_1 _1460_ (.Y(_0671_),
    .A(\reg_file.reg_array[119] ),
    .B(net485));
 sg13g2_a21oi_1 _1461_ (.A1(\reg_file.reg_array[103] ),
    .A2(net501),
    .Y(_0672_),
    .B1(net510));
 sg13g2_a22oi_1 _1462_ (.Y(_0673_),
    .B1(net480),
    .B2(\reg_file.reg_array[127] ),
    .A2(net490),
    .A1(\reg_file.reg_array[111] ));
 sg13g2_nand3_1 _1463_ (.B(_0672_),
    .C(_0673_),
    .A(_0671_),
    .Y(_0674_));
 sg13g2_and3_1 _1464_ (.X(_0193_),
    .A(net536),
    .B(net531),
    .C(\reg_file.reg_array[95] ));
 sg13g2_a221oi_1 _1465_ (.B2(\reg_file.reg_array[87] ),
    .C1(_0193_),
    .B1(net486),
    .A1(\reg_file.reg_array[79] ),
    .Y(_0194_),
    .A2(net491));
 sg13g2_a21oi_1 _1466_ (.A1(\reg_file.reg_array[71] ),
    .A2(net502),
    .Y(_0195_),
    .B1(net525));
 sg13g2_a21oi_1 _1467_ (.A1(_0194_),
    .A2(_0195_),
    .Y(_0196_),
    .B1(net515));
 sg13g2_a22oi_1 _1468_ (.Y(_0197_),
    .B1(_0674_),
    .B2(_0196_),
    .A2(_0670_),
    .A1(net515));
 sg13g2_a21oi_1 _1469_ (.A1(net496),
    .A2(_0197_),
    .Y(_0184_),
    .B1(_0665_));
 sg13g2_nand2_1 _1470_ (.Y(_0198_),
    .A(net32),
    .B(_0239_));
 sg13g2_o21ai_1 _1471_ (.B1(_0198_),
    .Y(_0185_),
    .A1(net508),
    .A2(_0301_));
 sg13g2_nor2_1 _1472_ (.A(net509),
    .B(_0302_),
    .Y(_0199_));
 sg13g2_mux2_1 _1473_ (.A0(net29),
    .A1(net1),
    .S(_0199_),
    .X(_0186_));
 sg13g2_nor2_1 _1474_ (.A(net509),
    .B(_0305_),
    .Y(_0200_));
 sg13g2_mux2_1 _1475_ (.A0(net27),
    .A1(net1),
    .S(_0200_),
    .X(_0187_));
 sg13g2_nor2_1 _1476_ (.A(net509),
    .B(_0308_),
    .Y(_0201_));
 sg13g2_nor2_1 _1477_ (.A(net28),
    .B(_0201_),
    .Y(_0202_));
 sg13g2_a21oi_1 _1478_ (.A1(_0024_),
    .A2(_0201_),
    .Y(_0188_),
    .B1(_0202_));
 sg13g2_o21ai_1 _1479_ (.B1(net26),
    .Y(_0203_),
    .A1(net508),
    .A2(_0311_));
 sg13g2_o21ai_1 _1480_ (.B1(_0203_),
    .Y(_0189_),
    .A1(net508),
    .A2(_0313_));
 sg13g2_nor3_1 _1481_ (.A(net518),
    .B(net508),
    .C(_0263_),
    .Y(_0204_));
 sg13g2_nor2_1 _1482_ (.A(net30),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_a21oi_1 _1483_ (.A1(net567),
    .A2(_0204_),
    .Y(_0190_),
    .B1(_0205_));
 sg13g2_nor3_1 _1484_ (.A(net518),
    .B(net509),
    .C(_0258_),
    .Y(_0206_));
 sg13g2_nor2_1 _1485_ (.A(net25),
    .B(_0206_),
    .Y(_0207_));
 sg13g2_a21oi_1 _1486_ (.A1(_0024_),
    .A2(_0206_),
    .Y(_0191_),
    .B1(_0207_));
 sg13g2_nor3_1 _1487_ (.A(net518),
    .B(net509),
    .C(_0260_),
    .Y(_0208_));
 sg13g2_nor2_1 _1488_ (.A(net31),
    .B(_0208_),
    .Y(_0209_));
 sg13g2_a21oi_1 _1489_ (.A1(_0024_),
    .A2(_0208_),
    .Y(_0192_),
    .B1(_0209_));
 sg13g2_inv_1 _1491__3 (.Y(net14),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1492__4 (.Y(net15),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1493__5 (.Y(net16),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1494__6 (.Y(net17),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1495__7 (.Y(net18),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1496__8 (.Y(net19),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1497__9 (.Y(net20),
    .A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _1498_ (.CLK(net12),
    .RESET_B(net578),
    .D(net48),
    .Q_N(_0832_),
    .Q(\i2c_slave_controller.state[0] ));
 sg13g2_dfrbp_1 _1499_ (.CLK(net13),
    .RESET_B(net578),
    .D(_0026_),
    .Q_N(_0831_),
    .Q(\i2c_slave_controller.state[1] ));
 sg13g2_dfrbp_1 _1500_ (.CLK(net14),
    .RESET_B(net580),
    .D(_0027_),
    .Q_N(_0001_),
    .Q(\i2c_slave_controller.state[2] ));
 sg13g2_dfrbp_1 _1501_ (.CLK(net551),
    .RESET_B(net579),
    .D(_0028_),
    .Q_N(_0004_),
    .Q(\reg_file.reg_pointer[0] ));
 sg13g2_dfrbp_1 _1502_ (.CLK(net564),
    .RESET_B(net595),
    .D(_0029_),
    .Q_N(_0830_),
    .Q(\reg_file.reg_pointer[1] ));
 sg13g2_dfrbp_1 _1503_ (.CLK(net563),
    .RESET_B(net593),
    .D(_0030_),
    .Q_N(_0829_),
    .Q(\reg_file.reg_pointer[2] ));
 sg13g2_dfrbp_1 _1504_ (.CLK(net551),
    .RESET_B(net579),
    .D(_0031_),
    .Q_N(_0003_),
    .Q(\reg_file.reg_pointer[3] ));
 sg13g2_dfrbp_1 _1505_ (.CLK(clknet_2_1__leaf_clk_regs),
    .RESET_B(net578),
    .D(_0032_),
    .Q_N(_0828_),
    .Q(\i2c_slave_controller.ack_recieved ));
 sg13g2_dfrbp_1 _1506_ (.CLK(clknet_2_1__leaf_clk_regs),
    .RESET_B(net591),
    .D(_0033_),
    .Q_N(_0005_),
    .Q(\i2c_slave_controller.out_regf_write_data[0] ));
 sg13g2_dfrbp_1 _1507_ (.CLK(clknet_2_2__leaf_clk_regs),
    .RESET_B(net596),
    .D(_0034_),
    .Q_N(_0006_),
    .Q(\i2c_slave_controller.out_regf_write_data[1] ));
 sg13g2_dfrbp_1 _1508_ (.CLK(clknet_2_3__leaf_clk_regs),
    .RESET_B(net596),
    .D(_0035_),
    .Q_N(_0007_),
    .Q(\i2c_slave_controller.out_regf_write_data[2] ));
 sg13g2_dfrbp_1 _1509_ (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net577),
    .D(_0036_),
    .Q_N(_0008_),
    .Q(\i2c_slave_controller.out_regf_write_data[3] ));
 sg13g2_dfrbp_1 _1510_ (.CLK(clknet_2_2__leaf_clk_regs),
    .RESET_B(net592),
    .D(_0037_),
    .Q_N(_0009_),
    .Q(\i2c_slave_controller.out_regf_write_data[4] ));
 sg13g2_dfrbp_1 _1511_ (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net579),
    .D(_0038_),
    .Q_N(_0010_),
    .Q(\i2c_slave_controller.out_regf_write_data[5] ));
 sg13g2_dfrbp_1 _1512_ (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net577),
    .D(_0039_),
    .Q_N(_0011_),
    .Q(\i2c_slave_controller.out_regf_write_data[6] ));
 sg13g2_dfrbp_1 _1513_ (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net576),
    .D(_0040_),
    .Q_N(_0012_),
    .Q(\i2c_slave_controller.out_regf_write_data[7] ));
 sg13g2_dfrbp_1 _1514_ (.CLK(clknet_2_1__leaf_clk_regs),
    .RESET_B(net578),
    .D(_0041_),
    .Q_N(_0827_),
    .Q(\i2c_slave_controller.out_regf_req ));
 sg13g2_dfrbp_1 _1515_ (.CLK(net15),
    .RESET_B(net592),
    .D(net35),
    .Q_N(_0826_),
    .Q(\i2c_slave_controller.counter[0] ));
 sg13g2_dfrbp_1 _1516_ (.CLK(net16),
    .RESET_B(net592),
    .D(_0043_),
    .Q_N(_0825_),
    .Q(\i2c_slave_controller.counter[1] ));
 sg13g2_dfrbp_1 _1517_ (.CLK(net17),
    .RESET_B(net580),
    .D(_0044_),
    .Q_N(_0002_),
    .Q(\i2c_slave_controller.counter[2] ));
 sg13g2_dfrbp_1 _1518_ (.CLK(net18),
    .RESET_B(net578),
    .D(_0045_),
    .Q_N(_0824_),
    .Q(\i2c_slave_controller.write_enable ));
 sg13g2_dfrbp_1 _1519_ (.CLK(net19),
    .RESET_B(net580),
    .D(net24),
    .Q_N(_0833_),
    .Q(\i2c_slave_controller.reg_sda_out ));
 sg13g2_dfrbp_1 _1520_ (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net578),
    .D(\i2c_slave_controller.out_stop ),
    .Q_N(_0823_),
    .Q(\i2c_slave_controller.stop_resetter ));
 sg13g2_dfrbp_1 _1521_ (.CLK(net20),
    .RESET_B(net595),
    .D(net37),
    .Q_N(_0822_),
    .Q(\i2c_slave_controller.out_regf_rw ));
 sg13g2_dfrbp_1 _1522_ (.CLK(net1),
    .RESET_B(_0022_),
    .D(clknet_1_0__leaf_clk),
    .Q_N(_0821_),
    .Q(\i2c_slave_controller.out_stop ));
 sg13g2_dfrbp_1 _1523_ (.CLK(net565),
    .RESET_B(net595),
    .D(_0048_),
    .Q_N(_0000_),
    .Q(\reg_file.state[0] ));
 sg13g2_dfrbp_1 _1524_ (.CLK(clknet_2_1__leaf_clk_regs),
    .RESET_B(net580),
    .D(\i2c_slave_controller.out_start ),
    .Q_N(_0820_),
    .Q(\i2c_slave_controller.start_resetter ));
 sg13g2_dfrbp_1 _1525_ (.CLK(net567),
    .RESET_B(_0023_),
    .D(clknet_1_0__leaf_clk),
    .Q_N(_0819_),
    .Q(\i2c_slave_controller.out_start ));
 sg13g2_dfrbp_1 _1526_ (.CLK(net564),
    .RESET_B(net595),
    .D(_0049_),
    .Q_N(_0818_),
    .Q(\reg_file.reg_array[0] ));
 sg13g2_dfrbp_1 _1527_ (.CLK(net564),
    .RESET_B(net595),
    .D(_0050_),
    .Q_N(_0817_),
    .Q(\reg_file.reg_array[1] ));
 sg13g2_dfrbp_1 _1528_ (.CLK(net564),
    .RESET_B(net595),
    .D(_0051_),
    .Q_N(_0816_),
    .Q(\reg_file.reg_array[2] ));
 sg13g2_dfrbp_1 _1529_ (.CLK(net549),
    .RESET_B(net577),
    .D(_0052_),
    .Q_N(_0815_),
    .Q(\reg_file.reg_array[3] ));
 sg13g2_dfrbp_1 _1530_ (.CLK(net565),
    .RESET_B(net591),
    .D(_0053_),
    .Q_N(_0814_),
    .Q(\reg_file.reg_array[4] ));
 sg13g2_dfrbp_1 _1531_ (.CLK(net551),
    .RESET_B(net579),
    .D(_0054_),
    .Q_N(_0813_),
    .Q(\reg_file.reg_array[5] ));
 sg13g2_dfrbp_1 _1532_ (.CLK(net549),
    .RESET_B(net576),
    .D(_0055_),
    .Q_N(_0812_),
    .Q(\reg_file.reg_array[6] ));
 sg13g2_dfrbp_1 _1533_ (.CLK(net549),
    .RESET_B(net576),
    .D(_0056_),
    .Q_N(_0811_),
    .Q(\reg_file.reg_array[7] ));
 sg13g2_dfrbp_1 _1534_ (.CLK(net558),
    .RESET_B(net587),
    .D(_0057_),
    .Q_N(_0810_),
    .Q(\reg_file.reg_array[8] ));
 sg13g2_dfrbp_1 _1535_ (.CLK(net562),
    .RESET_B(net593),
    .D(_0058_),
    .Q_N(_0809_),
    .Q(\reg_file.reg_array[9] ));
 sg13g2_dfrbp_1 _1536_ (.CLK(net562),
    .RESET_B(net593),
    .D(_0059_),
    .Q_N(_0808_),
    .Q(\reg_file.reg_array[10] ));
 sg13g2_dfrbp_1 _1537_ (.CLK(net550),
    .RESET_B(net577),
    .D(_0060_),
    .Q_N(_0807_),
    .Q(\reg_file.reg_array[11] ));
 sg13g2_dfrbp_1 _1538_ (.CLK(net565),
    .RESET_B(net591),
    .D(_0061_),
    .Q_N(_0806_),
    .Q(\reg_file.reg_array[12] ));
 sg13g2_dfrbp_1 _1539_ (.CLK(net547),
    .RESET_B(net574),
    .D(_0062_),
    .Q_N(_0805_),
    .Q(\reg_file.reg_array[13] ));
 sg13g2_dfrbp_1 _1540_ (.CLK(net550),
    .RESET_B(net577),
    .D(_0063_),
    .Q_N(_0804_),
    .Q(\reg_file.reg_array[14] ));
 sg13g2_dfrbp_1 _1541_ (.CLK(net544),
    .RESET_B(net571),
    .D(_0064_),
    .Q_N(_0803_),
    .Q(\reg_file.reg_array[15] ));
 sg13g2_dfrbp_1 _1542_ (.CLK(net558),
    .RESET_B(net587),
    .D(_0065_),
    .Q_N(_0802_),
    .Q(\reg_file.reg_array[16] ));
 sg13g2_dfrbp_1 _1543_ (.CLK(net563),
    .RESET_B(net594),
    .D(_0066_),
    .Q_N(_0801_),
    .Q(\reg_file.reg_array[17] ));
 sg13g2_dfrbp_1 _1544_ (.CLK(net563),
    .RESET_B(net594),
    .D(_0067_),
    .Q_N(_0800_),
    .Q(\reg_file.reg_array[18] ));
 sg13g2_dfrbp_1 _1545_ (.CLK(net549),
    .RESET_B(net577),
    .D(_0068_),
    .Q_N(_0799_),
    .Q(\reg_file.reg_array[19] ));
 sg13g2_dfrbp_1 _1546_ (.CLK(net565),
    .RESET_B(net591),
    .D(_0069_),
    .Q_N(_0798_),
    .Q(\reg_file.reg_array[20] ));
 sg13g2_dfrbp_1 _1547_ (.CLK(net547),
    .RESET_B(net574),
    .D(_0070_),
    .Q_N(_0797_),
    .Q(\reg_file.reg_array[21] ));
 sg13g2_dfrbp_1 _1548_ (.CLK(net543),
    .RESET_B(net570),
    .D(_0071_),
    .Q_N(_0796_),
    .Q(\reg_file.reg_array[22] ));
 sg13g2_dfrbp_1 _1549_ (.CLK(net543),
    .RESET_B(net570),
    .D(_0072_),
    .Q_N(_0795_),
    .Q(\reg_file.reg_array[23] ));
 sg13g2_dfrbp_1 _1550_ (.CLK(net562),
    .RESET_B(net593),
    .D(_0073_),
    .Q_N(_0794_),
    .Q(\reg_file.reg_array[24] ));
 sg13g2_dfrbp_1 _1551_ (.CLK(net562),
    .RESET_B(net593),
    .D(_0074_),
    .Q_N(_0793_),
    .Q(\reg_file.reg_array[25] ));
 sg13g2_dfrbp_1 _1552_ (.CLK(net562),
    .RESET_B(net593),
    .D(_0075_),
    .Q_N(_0792_),
    .Q(\reg_file.reg_array[26] ));
 sg13g2_dfrbp_1 _1553_ (.CLK(net550),
    .RESET_B(net576),
    .D(_0076_),
    .Q_N(_0791_),
    .Q(\reg_file.reg_array[27] ));
 sg13g2_dfrbp_1 _1554_ (.CLK(net565),
    .RESET_B(net591),
    .D(_0077_),
    .Q_N(_0790_),
    .Q(\reg_file.reg_array[28] ));
 sg13g2_dfrbp_1 _1555_ (.CLK(net561),
    .RESET_B(net584),
    .D(_0078_),
    .Q_N(_0789_),
    .Q(\reg_file.reg_array[29] ));
 sg13g2_dfrbp_1 _1556_ (.CLK(net543),
    .RESET_B(net570),
    .D(_0079_),
    .Q_N(_0788_),
    .Q(\reg_file.reg_array[30] ));
 sg13g2_dfrbp_1 _1557_ (.CLK(net549),
    .RESET_B(net576),
    .D(_0080_),
    .Q_N(_0787_),
    .Q(\reg_file.reg_array[31] ));
 sg13g2_dfrbp_1 _1558_ (.CLK(net559),
    .RESET_B(net587),
    .D(_0081_),
    .Q_N(_0786_),
    .Q(\reg_file.reg_array[32] ));
 sg13g2_dfrbp_1 _1559_ (.CLK(net557),
    .RESET_B(net586),
    .D(_0082_),
    .Q_N(_0785_),
    .Q(\reg_file.reg_array[33] ));
 sg13g2_dfrbp_1 _1560_ (.CLK(net556),
    .RESET_B(net585),
    .D(_0083_),
    .Q_N(_0784_),
    .Q(\reg_file.reg_array[34] ));
 sg13g2_dfrbp_1 _1561_ (.CLK(net546),
    .RESET_B(net573),
    .D(_0084_),
    .Q_N(_0783_),
    .Q(\reg_file.reg_array[35] ));
 sg13g2_dfrbp_1 _1562_ (.CLK(net553),
    .RESET_B(net582),
    .D(_0085_),
    .Q_N(_0782_),
    .Q(\reg_file.reg_array[36] ));
 sg13g2_dfrbp_1 _1563_ (.CLK(net548),
    .RESET_B(net575),
    .D(_0086_),
    .Q_N(_0781_),
    .Q(\reg_file.reg_array[37] ));
 sg13g2_dfrbp_1 _1564_ (.CLK(net542),
    .RESET_B(net569),
    .D(_0087_),
    .Q_N(_0780_),
    .Q(\reg_file.reg_array[38] ));
 sg13g2_dfrbp_1 _1565_ (.CLK(net542),
    .RESET_B(net569),
    .D(_0088_),
    .Q_N(_0779_),
    .Q(\reg_file.reg_array[39] ));
 sg13g2_dfrbp_1 _1566_ (.CLK(net556),
    .RESET_B(net585),
    .D(_0089_),
    .Q_N(_0778_),
    .Q(\reg_file.reg_array[40] ));
 sg13g2_dfrbp_1 _1567_ (.CLK(net556),
    .RESET_B(net585),
    .D(_0090_),
    .Q_N(_0777_),
    .Q(\reg_file.reg_array[41] ));
 sg13g2_dfrbp_1 _1568_ (.CLK(net556),
    .RESET_B(net585),
    .D(_0091_),
    .Q_N(_0776_),
    .Q(\reg_file.reg_array[42] ));
 sg13g2_dfrbp_1 _1569_ (.CLK(net542),
    .RESET_B(net569),
    .D(_0092_),
    .Q_N(_0775_),
    .Q(\reg_file.reg_array[43] ));
 sg13g2_dfrbp_1 _1570_ (.CLK(net553),
    .RESET_B(net582),
    .D(_0093_),
    .Q_N(_0774_),
    .Q(\reg_file.reg_array[44] ));
 sg13g2_dfrbp_1 _1571_ (.CLK(net548),
    .RESET_B(net573),
    .D(_0094_),
    .Q_N(_0773_),
    .Q(\reg_file.reg_array[45] ));
 sg13g2_dfrbp_1 _1572_ (.CLK(net541),
    .RESET_B(net568),
    .D(_0095_),
    .Q_N(_0772_),
    .Q(\reg_file.reg_array[46] ));
 sg13g2_dfrbp_1 _1573_ (.CLK(net541),
    .RESET_B(net568),
    .D(_0096_),
    .Q_N(_0771_),
    .Q(\reg_file.reg_array[47] ));
 sg13g2_dfrbp_1 _1574_ (.CLK(net556),
    .RESET_B(net585),
    .D(_0097_),
    .Q_N(_0770_),
    .Q(\reg_file.reg_array[48] ));
 sg13g2_dfrbp_1 _1575_ (.CLK(net557),
    .RESET_B(net586),
    .D(_0098_),
    .Q_N(_0769_),
    .Q(\reg_file.reg_array[49] ));
 sg13g2_dfrbp_1 _1576_ (.CLK(net557),
    .RESET_B(net586),
    .D(_0099_),
    .Q_N(_0768_),
    .Q(\reg_file.reg_array[50] ));
 sg13g2_dfrbp_1 _1577_ (.CLK(net542),
    .RESET_B(net569),
    .D(_0100_),
    .Q_N(_0767_),
    .Q(\reg_file.reg_array[51] ));
 sg13g2_dfrbp_1 _1578_ (.CLK(net554),
    .RESET_B(net583),
    .D(_0101_),
    .Q_N(_0766_),
    .Q(\reg_file.reg_array[52] ));
 sg13g2_dfrbp_1 _1579_ (.CLK(net546),
    .RESET_B(net575),
    .D(_0102_),
    .Q_N(_0765_),
    .Q(\reg_file.reg_array[53] ));
 sg13g2_dfrbp_1 _1580_ (.CLK(net541),
    .RESET_B(net568),
    .D(_0103_),
    .Q_N(_0764_),
    .Q(\reg_file.reg_array[54] ));
 sg13g2_dfrbp_1 _1581_ (.CLK(net543),
    .RESET_B(net570),
    .D(_0104_),
    .Q_N(_0763_),
    .Q(\reg_file.reg_array[55] ));
 sg13g2_dfrbp_1 _1582_ (.CLK(net555),
    .RESET_B(net584),
    .D(_0105_),
    .Q_N(_0762_),
    .Q(\reg_file.reg_array[56] ));
 sg13g2_dfrbp_1 _1583_ (.CLK(net553),
    .RESET_B(net582),
    .D(_0106_),
    .Q_N(_0761_),
    .Q(\reg_file.reg_array[57] ));
 sg13g2_dfrbp_1 _1584_ (.CLK(net554),
    .RESET_B(net583),
    .D(_0107_),
    .Q_N(_0760_),
    .Q(\reg_file.reg_array[58] ));
 sg13g2_dfrbp_1 _1585_ (.CLK(net542),
    .RESET_B(net569),
    .D(_0108_),
    .Q_N(_0759_),
    .Q(\reg_file.reg_array[59] ));
 sg13g2_dfrbp_1 _1586_ (.CLK(net553),
    .RESET_B(net582),
    .D(_0109_),
    .Q_N(_0758_),
    .Q(\reg_file.reg_array[60] ));
 sg13g2_dfrbp_1 _1587_ (.CLK(net548),
    .RESET_B(net575),
    .D(_0110_),
    .Q_N(_0757_),
    .Q(\reg_file.reg_array[61] ));
 sg13g2_dfrbp_1 _1588_ (.CLK(net541),
    .RESET_B(net568),
    .D(_0111_),
    .Q_N(_0756_),
    .Q(\reg_file.reg_array[62] ));
 sg13g2_dfrbp_1 _1589_ (.CLK(net543),
    .RESET_B(net570),
    .D(_0112_),
    .Q_N(_0755_),
    .Q(\reg_file.reg_array[63] ));
 sg13g2_dfrbp_1 _1590_ (.CLK(net559),
    .RESET_B(net588),
    .D(_0113_),
    .Q_N(_0754_),
    .Q(\reg_file.reg_array[64] ));
 sg13g2_dfrbp_1 _1591_ (.CLK(net558),
    .RESET_B(net587),
    .D(_0114_),
    .Q_N(_0753_),
    .Q(\reg_file.reg_array[65] ));
 sg13g2_dfrbp_1 _1592_ (.CLK(net558),
    .RESET_B(net588),
    .D(_0115_),
    .Q_N(_0752_),
    .Q(\reg_file.reg_array[66] ));
 sg13g2_dfrbp_1 _1593_ (.CLK(net551),
    .RESET_B(net579),
    .D(_0116_),
    .Q_N(_0751_),
    .Q(\reg_file.reg_array[67] ));
 sg13g2_dfrbp_1 _1594_ (.CLK(net555),
    .RESET_B(net584),
    .D(_0117_),
    .Q_N(_0750_),
    .Q(\reg_file.reg_array[68] ));
 sg13g2_dfrbp_1 _1595_ (.CLK(net547),
    .RESET_B(net574),
    .D(_0118_),
    .Q_N(_0749_),
    .Q(\reg_file.reg_array[69] ));
 sg13g2_dfrbp_1 _1596_ (.CLK(net544),
    .RESET_B(net571),
    .D(_0119_),
    .Q_N(_0748_),
    .Q(\reg_file.reg_array[70] ));
 sg13g2_dfrbp_1 _1597_ (.CLK(net544),
    .RESET_B(net571),
    .D(_0120_),
    .Q_N(_0747_),
    .Q(\reg_file.reg_array[71] ));
 sg13g2_dfrbp_1 _1598_ (.CLK(net558),
    .RESET_B(net587),
    .D(_0121_),
    .Q_N(_0746_),
    .Q(\reg_file.reg_array[72] ));
 sg13g2_dfrbp_1 _1599_ (.CLK(net555),
    .RESET_B(net584),
    .D(_0122_),
    .Q_N(_0745_),
    .Q(\reg_file.reg_array[73] ));
 sg13g2_dfrbp_1 _1600_ (.CLK(net562),
    .RESET_B(net593),
    .D(_0123_),
    .Q_N(_0744_),
    .Q(\reg_file.reg_array[74] ));
 sg13g2_dfrbp_1 _1601_ (.CLK(net551),
    .RESET_B(net579),
    .D(_0124_),
    .Q_N(_0743_),
    .Q(\reg_file.reg_array[75] ));
 sg13g2_dfrbp_1 _1602_ (.CLK(net555),
    .RESET_B(net584),
    .D(_0125_),
    .Q_N(_0742_),
    .Q(\reg_file.reg_array[76] ));
 sg13g2_dfrbp_1 _1603_ (.CLK(net547),
    .RESET_B(net574),
    .D(_0126_),
    .Q_N(_0741_),
    .Q(\reg_file.reg_array[77] ));
 sg13g2_dfrbp_1 _1604_ (.CLK(net547),
    .RESET_B(net574),
    .D(_0127_),
    .Q_N(_0740_),
    .Q(\reg_file.reg_array[78] ));
 sg13g2_dfrbp_1 _1605_ (.CLK(net547),
    .RESET_B(net574),
    .D(_0128_),
    .Q_N(_0739_),
    .Q(\reg_file.reg_array[79] ));
 sg13g2_dfrbp_1 _1606_ (.CLK(net558),
    .RESET_B(net587),
    .D(_0129_),
    .Q_N(_0738_),
    .Q(\reg_file.reg_array[80] ));
 sg13g2_dfrbp_1 _1607_ (.CLK(net563),
    .RESET_B(net594),
    .D(_0130_),
    .Q_N(_0737_),
    .Q(\reg_file.reg_array[81] ));
 sg13g2_dfrbp_1 _1608_ (.CLK(net563),
    .RESET_B(net594),
    .D(_0131_),
    .Q_N(_0736_),
    .Q(\reg_file.reg_array[82] ));
 sg13g2_dfrbp_1 _1609_ (.CLK(net550),
    .RESET_B(net577),
    .D(_0132_),
    .Q_N(_0735_),
    .Q(\reg_file.reg_array[83] ));
 sg13g2_dfrbp_1 _1610_ (.CLK(net565),
    .RESET_B(net591),
    .D(_0133_),
    .Q_N(_0734_),
    .Q(\reg_file.reg_array[84] ));
 sg13g2_dfrbp_1 _1611_ (.CLK(net547),
    .RESET_B(net574),
    .D(_0134_),
    .Q_N(_0733_),
    .Q(\reg_file.reg_array[85] ));
 sg13g2_dfrbp_1 _1612_ (.CLK(net544),
    .RESET_B(net571),
    .D(_0135_),
    .Q_N(_0732_),
    .Q(\reg_file.reg_array[86] ));
 sg13g2_dfrbp_1 _1613_ (.CLK(net549),
    .RESET_B(net576),
    .D(_0136_),
    .Q_N(_0731_),
    .Q(\reg_file.reg_array[87] ));
 sg13g2_dfrbp_1 _1614_ (.CLK(net558),
    .RESET_B(net587),
    .D(_0137_),
    .Q_N(_0730_),
    .Q(\reg_file.reg_array[88] ));
 sg13g2_dfrbp_1 _1615_ (.CLK(net562),
    .RESET_B(net593),
    .D(_0138_),
    .Q_N(_0729_),
    .Q(\reg_file.reg_array[89] ));
 sg13g2_dfrbp_1 _1616_ (.CLK(net562),
    .RESET_B(net594),
    .D(_0139_),
    .Q_N(_0728_),
    .Q(\reg_file.reg_array[90] ));
 sg13g2_dfrbp_1 _1617_ (.CLK(net549),
    .RESET_B(net576),
    .D(_0140_),
    .Q_N(_0727_),
    .Q(\reg_file.reg_array[91] ));
 sg13g2_dfrbp_1 _1618_ (.CLK(net555),
    .RESET_B(net584),
    .D(_0141_),
    .Q_N(_0726_),
    .Q(\reg_file.reg_array[92] ));
 sg13g2_dfrbp_1 _1619_ (.CLK(net561),
    .RESET_B(net590),
    .D(_0142_),
    .Q_N(_0725_),
    .Q(\reg_file.reg_array[93] ));
 sg13g2_dfrbp_1 _1620_ (.CLK(net543),
    .RESET_B(net570),
    .D(_0143_),
    .Q_N(_0724_),
    .Q(\reg_file.reg_array[94] ));
 sg13g2_dfrbp_1 _1621_ (.CLK(net549),
    .RESET_B(net576),
    .D(_0144_),
    .Q_N(_0723_),
    .Q(\reg_file.reg_array[95] ));
 sg13g2_dfrbp_1 _1622_ (.CLK(net559),
    .RESET_B(net588),
    .D(_0145_),
    .Q_N(_0722_),
    .Q(\reg_file.reg_array[96] ));
 sg13g2_dfrbp_1 _1623_ (.CLK(net557),
    .RESET_B(net586),
    .D(_0146_),
    .Q_N(_0721_),
    .Q(\reg_file.reg_array[97] ));
 sg13g2_dfrbp_1 _1624_ (.CLK(net556),
    .RESET_B(net585),
    .D(_0147_),
    .Q_N(_0720_),
    .Q(\reg_file.reg_array[98] ));
 sg13g2_dfrbp_1 _1625_ (.CLK(net546),
    .RESET_B(net573),
    .D(_0148_),
    .Q_N(_0719_),
    .Q(\reg_file.reg_array[99] ));
 sg13g2_dfrbp_1 _1626_ (.CLK(net553),
    .RESET_B(net582),
    .D(_0149_),
    .Q_N(_0718_),
    .Q(\reg_file.reg_array[100] ));
 sg13g2_dfrbp_1 _1627_ (.CLK(net546),
    .RESET_B(net573),
    .D(_0150_),
    .Q_N(_0717_),
    .Q(\reg_file.reg_array[101] ));
 sg13g2_dfrbp_1 _1628_ (.CLK(net542),
    .RESET_B(net569),
    .D(_0151_),
    .Q_N(_0716_),
    .Q(\reg_file.reg_array[102] ));
 sg13g2_dfrbp_1 _1629_ (.CLK(net544),
    .RESET_B(net571),
    .D(_0152_),
    .Q_N(_0715_),
    .Q(\reg_file.reg_array[103] ));
 sg13g2_dfrbp_1 _1630_ (.CLK(net558),
    .RESET_B(net587),
    .D(_0153_),
    .Q_N(_0714_),
    .Q(\reg_file.reg_array[104] ));
 sg13g2_dfrbp_1 _1631_ (.CLK(net556),
    .RESET_B(net585),
    .D(_0154_),
    .Q_N(_0713_),
    .Q(\reg_file.reg_array[105] ));
 sg13g2_dfrbp_1 _1632_ (.CLK(net556),
    .RESET_B(net585),
    .D(_0155_),
    .Q_N(_0712_),
    .Q(\reg_file.reg_array[106] ));
 sg13g2_dfrbp_1 _1633_ (.CLK(net546),
    .RESET_B(net573),
    .D(_0156_),
    .Q_N(_0711_),
    .Q(\reg_file.reg_array[107] ));
 sg13g2_dfrbp_1 _1634_ (.CLK(net553),
    .RESET_B(net582),
    .D(_0157_),
    .Q_N(_0710_),
    .Q(\reg_file.reg_array[108] ));
 sg13g2_dfrbp_1 _1635_ (.CLK(net548),
    .RESET_B(net574),
    .D(_0158_),
    .Q_N(_0709_),
    .Q(\reg_file.reg_array[109] ));
 sg13g2_dfrbp_1 _1636_ (.CLK(net541),
    .RESET_B(net568),
    .D(_0159_),
    .Q_N(_0708_),
    .Q(\reg_file.reg_array[110] ));
 sg13g2_dfrbp_1 _1637_ (.CLK(net541),
    .RESET_B(net568),
    .D(_0160_),
    .Q_N(_0707_),
    .Q(\reg_file.reg_array[111] ));
 sg13g2_dfrbp_1 _1638_ (.CLK(net559),
    .RESET_B(net588),
    .D(_0161_),
    .Q_N(_0706_),
    .Q(\reg_file.reg_array[112] ));
 sg13g2_dfrbp_1 _1639_ (.CLK(net557),
    .RESET_B(net586),
    .D(_0162_),
    .Q_N(_0705_),
    .Q(\reg_file.reg_array[113] ));
 sg13g2_dfrbp_1 _1640_ (.CLK(net557),
    .RESET_B(net586),
    .D(_0163_),
    .Q_N(_0704_),
    .Q(\reg_file.reg_array[114] ));
 sg13g2_dfrbp_1 _1641_ (.CLK(net546),
    .RESET_B(net573),
    .D(_0164_),
    .Q_N(_0703_),
    .Q(\reg_file.reg_array[115] ));
 sg13g2_dfrbp_1 _1642_ (.CLK(net554),
    .RESET_B(net583),
    .D(_0165_),
    .Q_N(_0702_),
    .Q(\reg_file.reg_array[116] ));
 sg13g2_dfrbp_1 _1643_ (.CLK(net546),
    .RESET_B(net573),
    .D(_0166_),
    .Q_N(_0701_),
    .Q(\reg_file.reg_array[117] ));
 sg13g2_dfrbp_1 _1644_ (.CLK(net541),
    .RESET_B(net568),
    .D(_0167_),
    .Q_N(_0700_),
    .Q(\reg_file.reg_array[118] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(net543),
    .RESET_B(net570),
    .D(_0168_),
    .Q_N(_0699_),
    .Q(\reg_file.reg_array[119] ));
 sg13g2_dfrbp_1 _1646_ (.CLK(net555),
    .RESET_B(net590),
    .D(_0169_),
    .Q_N(_0698_),
    .Q(\reg_file.reg_array[120] ));
 sg13g2_dfrbp_1 _1647_ (.CLK(net553),
    .RESET_B(net582),
    .D(_0170_),
    .Q_N(_0697_),
    .Q(\reg_file.reg_array[121] ));
 sg13g2_dfrbp_1 _1648_ (.CLK(net554),
    .RESET_B(net583),
    .D(_0171_),
    .Q_N(_0696_),
    .Q(\reg_file.reg_array[122] ));
 sg13g2_dfrbp_1 _1649_ (.CLK(net546),
    .RESET_B(net573),
    .D(_0172_),
    .Q_N(_0695_),
    .Q(\reg_file.reg_array[123] ));
 sg13g2_dfrbp_1 _1650_ (.CLK(net553),
    .RESET_B(net582),
    .D(_0173_),
    .Q_N(_0694_),
    .Q(\reg_file.reg_array[124] ));
 sg13g2_dfrbp_1 _1651_ (.CLK(net547),
    .RESET_B(net575),
    .D(_0174_),
    .Q_N(_0693_),
    .Q(\reg_file.reg_array[125] ));
 sg13g2_dfrbp_1 _1652_ (.CLK(net541),
    .RESET_B(net568),
    .D(_0175_),
    .Q_N(_0692_),
    .Q(\reg_file.reg_array[126] ));
 sg13g2_dfrbp_1 _1653_ (.CLK(net543),
    .RESET_B(net570),
    .D(_0176_),
    .Q_N(_0691_),
    .Q(\reg_file.reg_array[127] ));
 sg13g2_dfrbp_1 _1654_ (.CLK(net566),
    .RESET_B(net595),
    .D(_0177_),
    .Q_N(_0690_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1655_ (.CLK(net564),
    .RESET_B(net595),
    .D(_0178_),
    .Q_N(_0689_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1656_ (.CLK(net564),
    .RESET_B(net596),
    .D(_0179_),
    .Q_N(_0688_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1657_ (.CLK(net551),
    .RESET_B(net579),
    .D(_0180_),
    .Q_N(_0687_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1658_ (.CLK(net565),
    .RESET_B(net591),
    .D(_0181_),
    .Q_N(_0686_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1659_ (.CLK(net552),
    .RESET_B(net579),
    .D(_0182_),
    .Q_N(_0685_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1660_ (.CLK(net552),
    .RESET_B(net580),
    .D(_0183_),
    .Q_N(_0684_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1661_ (.CLK(net551),
    .RESET_B(net580),
    .D(_0184_),
    .Q_N(_0683_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1662_ (.CLK(clknet_2_1__leaf_clk_regs),
    .RESET_B(net592),
    .D(_0185_),
    .Q_N(_0682_),
    .Q(\i2c_slave_controller.addr[0] ));
 sg13g2_dfrbp_1 _1663_ (.CLK(clknet_2_2__leaf_clk_regs),
    .RESET_B(net596),
    .D(_0186_),
    .Q_N(_0681_),
    .Q(\i2c_slave_controller.addr[1] ));
 sg13g2_dfrbp_1 _1664_ (.CLK(clknet_2_3__leaf_clk_regs),
    .RESET_B(net592),
    .D(_0187_),
    .Q_N(_0680_),
    .Q(\i2c_slave_controller.addr[2] ));
 sg13g2_dfrbp_1 _1665_ (.CLK(clknet_2_3__leaf_clk_regs),
    .RESET_B(net596),
    .D(_0188_),
    .Q_N(_0679_),
    .Q(\i2c_slave_controller.addr[3] ));
 sg13g2_dfrbp_1 _1666_ (.CLK(clknet_2_2__leaf_clk_regs),
    .RESET_B(net591),
    .D(_0189_),
    .Q_N(_0678_),
    .Q(\i2c_slave_controller.addr[4] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(clknet_2_2__leaf_clk_regs),
    .RESET_B(net596),
    .D(_0190_),
    .Q_N(_0677_),
    .Q(\i2c_slave_controller.addr[5] ));
 sg13g2_dfrbp_1 _1668_ (.CLK(clknet_2_3__leaf_clk_regs),
    .RESET_B(net592),
    .D(_0191_),
    .Q_N(_0676_),
    .Q(\i2c_slave_controller.addr[6] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(clknet_2_3__leaf_clk_regs),
    .RESET_B(net596),
    .D(_0192_),
    .Q_N(_0675_),
    .Q(\i2c_slave_controller.addr[7] ));
 sg13g2_inv_1 _0853__1 (.Y(net12),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_i2c_regf_3 (.L_LO(net3));
 sg13g2_tielo tt_um_i2c_regf_4 (.L_LO(net4));
 sg13g2_tielo tt_um_i2c_regf_5 (.L_LO(net5));
 sg13g2_tielo tt_um_i2c_regf_6 (.L_LO(net6));
 sg13g2_tielo tt_um_i2c_regf_7 (.L_LO(net7));
 sg13g2_tielo tt_um_i2c_regf_8 (.L_LO(net8));
 sg13g2_tielo tt_um_i2c_regf_9 (.L_LO(net9));
 sg13g2_tielo tt_um_i2c_regf_10 (.L_LO(net10));
 sg13g2_tiehi tt_um_i2c_regf_11 (.L_HI(net11));
 sg13g2_buf_1 _1680_ (.A(\i2c_slave_controller.write_enable ),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1681_ (.A(\i2c_slave_controller.reg_sda_out ),
    .X(uio_out[0]));
 sg13g2_buf_1 _1682_ (.A(\i2c_slave_controller.out_start ),
    .X(uio_out[1]));
 sg13g2_buf_1 _1683_ (.A(\i2c_slave_controller.out_start_reset ),
    .X(uio_out[2]));
 sg13g2_buf_1 _1684_ (.A(\i2c_slave_controller.out_stop ),
    .X(uio_out[3]));
 sg13g2_buf_1 _1685_ (.A(\i2c_slave_controller.out_stop_reset ),
    .X(uio_out[4]));
 sg13g2_buf_2 fanout449 (.A(net452),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(net452),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_0495_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(net457),
    .X(net453));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(net456));
 sg13g2_buf_2 fanout455 (.A(net456),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(net457),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_0495_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_0494_),
    .X(net458));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(net460));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(net462));
 sg13g2_buf_2 fanout461 (.A(net462),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(net467),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(net467));
 sg13g2_buf_2 fanout465 (.A(net466),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net467),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_0348_),
    .X(net467));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(_0347_));
 sg13g2_buf_2 fanout469 (.A(_0332_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_0332_),
    .X(net470));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(net472));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(_0388_));
 sg13g2_buf_2 fanout473 (.A(net475),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_1 fanout475 (.A(_0342_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(net478),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_0331_),
    .X(net478));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(_0326_));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(net482));
 sg13g2_buf_2 fanout481 (.A(net482),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_0386_),
    .X(net482));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(net484));
 sg13g2_buf_2 fanout484 (.A(_0386_),
    .X(net484));
 sg13g2_buf_4 fanout485 (.X(net485),
    .A(net486));
 sg13g2_buf_2 fanout486 (.A(net489),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(net489));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(_0358_));
 sg13g2_buf_2 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net495));
 sg13g2_buf_2 fanout492 (.A(net494),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(net495),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_0341_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_0328_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_0328_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net500),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_0327_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(net502),
    .X(net501));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(net505));
 sg13g2_buf_2 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(net505));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(_0325_));
 sg13g2_buf_2 fanout506 (.A(_0245_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_0245_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_0231_),
    .X(net508));
 sg13g2_buf_1 fanout509 (.A(_0231_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(net514),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net514),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(net514),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_0215_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_0214_),
    .X(net515));
 sg13g2_buf_1 fanout516 (.A(_0214_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_0002_),
    .X(net517));
 sg13g2_buf_1 fanout518 (.A(_0002_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(net50),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(\i2c_slave_controller.counter[0] ),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(\reg_file.reg_pointer[3] ),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(net525),
    .X(net523));
 sg13g2_buf_1 fanout524 (.A(net525),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(net528),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(net527),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(\reg_file.reg_pointer[2] ),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(\reg_file.reg_pointer[1] ),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(net533),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(\reg_file.reg_pointer[1] ),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_1 fanout535 (.A(\reg_file.reg_pointer[1] ),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(\reg_file.reg_pointer[0] ),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_0001_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(net46),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(net49),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net47),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net545),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net545),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net545),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_1 fanout545 (.A(net566),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(net548),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net566),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(net550),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net552),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_1 fanout552 (.A(net566),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net555),
    .X(net553));
 sg13g2_buf_1 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(net561),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net560),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(net560),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net560),
    .X(net558));
 sg13g2_buf_1 fanout559 (.A(net560),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_1 fanout561 (.A(net566),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net564),
    .X(net562));
 sg13g2_buf_1 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net565),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(\i2c_slave_controller.out_regf_req ),
    .X(net566));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(_0024_));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(net572));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(net572));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(net572));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net581),
    .X(net572));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(net575));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(net575));
 sg13g2_buf_2 fanout575 (.A(net581),
    .X(net575));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(net577));
 sg13g2_buf_4 fanout577 (.X(net577),
    .A(net578));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(net581));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(net581));
 sg13g2_buf_4 fanout580 (.X(net580),
    .A(net581));
 sg13g2_buf_2 fanout581 (.A(rst_n),
    .X(net581));
 sg13g2_buf_4 fanout582 (.X(net582),
    .A(net584));
 sg13g2_buf_2 fanout583 (.A(net584),
    .X(net583));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(net590));
 sg13g2_buf_4 fanout585 (.X(net585),
    .A(net589));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(net589));
 sg13g2_buf_4 fanout587 (.X(net587),
    .A(net589));
 sg13g2_buf_2 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(rst_n),
    .X(net590));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(net597));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(net597));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(net597));
 sg13g2_buf_2 fanout594 (.A(net597),
    .X(net594));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(net596));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(net597));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(uio_in[0]),
    .X(net1));
 sg13g2_tielo tt_um_i2c_regf_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_2_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_2_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_2_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_2_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_3__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\i2c_slave_controller.ack_recieved ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold2 (.A(\i2c_slave_controller.write_enable ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold3 (.A(\i2c_slave_controller.reg_sda_out ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0046_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i2c_slave_controller.addr[6] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i2c_slave_controller.addr[4] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i2c_slave_controller.addr[2] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i2c_slave_controller.addr[3] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i2c_slave_controller.addr[1] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i2c_slave_controller.addr[5] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i2c_slave_controller.addr[7] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i2c_slave_controller.addr[0] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i2c_slave_controller.counter[2] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i2c_slave_controller.counter[0] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0042_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i2c_slave_controller.out_regf_rw ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0047_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i2c_slave_controller.out_regf_write_data[5] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i2c_slave_controller.out_regf_write_data[4] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i2c_slave_controller.out_regf_write_data[1] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i2c_slave_controller.out_regf_write_data[2] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i2c_slave_controller.out_regf_write_data[7] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i2c_slave_controller.out_regf_write_data[6] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i2c_slave_controller.out_regf_write_data[3] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i2c_slave_controller.out_regf_write_data[0] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i2c_slave_controller.state[2] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i2c_slave_controller.state[0] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0025_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i2c_slave_controller.state[1] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i2c_slave_controller.counter[1] ),
    .X(net50));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_fill_1 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_4 FILLER_7_268 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_4 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_37 ();
 sg13g2_decap_8 FILLER_8_44 ();
 sg13g2_decap_8 FILLER_8_51 ();
 sg13g2_decap_8 FILLER_8_58 ();
 sg13g2_fill_2 FILLER_8_65 ();
 sg13g2_fill_1 FILLER_8_67 ();
 sg13g2_fill_1 FILLER_8_124 ();
 sg13g2_decap_8 FILLER_8_155 ();
 sg13g2_decap_4 FILLER_8_162 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_decap_4 FILLER_8_199 ();
 sg13g2_fill_2 FILLER_8_203 ();
 sg13g2_fill_2 FILLER_8_239 ();
 sg13g2_decap_8 FILLER_8_267 ();
 sg13g2_decap_8 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_288 ();
 sg13g2_fill_1 FILLER_8_295 ();
 sg13g2_fill_1 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_4 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_62 ();
 sg13g2_decap_8 FILLER_9_97 ();
 sg13g2_fill_1 FILLER_9_104 ();
 sg13g2_fill_2 FILLER_9_158 ();
 sg13g2_fill_1 FILLER_9_160 ();
 sg13g2_decap_4 FILLER_9_196 ();
 sg13g2_decap_4 FILLER_9_226 ();
 sg13g2_decap_4 FILLER_9_234 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_decap_4 FILLER_9_264 ();
 sg13g2_fill_2 FILLER_9_268 ();
 sg13g2_fill_1 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_fill_2 FILLER_9_380 ();
 sg13g2_fill_1 FILLER_9_382 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_37 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_fill_2 FILLER_10_79 ();
 sg13g2_fill_1 FILLER_10_81 ();
 sg13g2_fill_2 FILLER_10_86 ();
 sg13g2_fill_1 FILLER_10_88 ();
 sg13g2_fill_2 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_131 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_230 ();
 sg13g2_decap_4 FILLER_10_237 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_295 ();
 sg13g2_decap_4 FILLER_10_309 ();
 sg13g2_decap_4 FILLER_10_334 ();
 sg13g2_fill_2 FILLER_10_338 ();
 sg13g2_decap_4 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_44 ();
 sg13g2_decap_8 FILLER_11_51 ();
 sg13g2_decap_4 FILLER_11_58 ();
 sg13g2_fill_1 FILLER_11_62 ();
 sg13g2_decap_4 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_92 ();
 sg13g2_decap_8 FILLER_11_99 ();
 sg13g2_fill_2 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_108 ();
 sg13g2_fill_2 FILLER_11_113 ();
 sg13g2_fill_2 FILLER_11_123 ();
 sg13g2_decap_4 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_165 ();
 sg13g2_fill_1 FILLER_11_174 ();
 sg13g2_decap_4 FILLER_11_201 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_4 FILLER_11_242 ();
 sg13g2_fill_1 FILLER_11_246 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_decap_4 FILLER_11_266 ();
 sg13g2_fill_1 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_4 FILLER_11_287 ();
 sg13g2_fill_1 FILLER_11_291 ();
 sg13g2_decap_4 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_2 FILLER_12_29 ();
 sg13g2_fill_1 FILLER_12_31 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_2 FILLER_12_86 ();
 sg13g2_decap_4 FILLER_12_124 ();
 sg13g2_fill_1 FILLER_12_132 ();
 sg13g2_decap_8 FILLER_12_143 ();
 sg13g2_decap_8 FILLER_12_150 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_decap_8 FILLER_12_163 ();
 sg13g2_decap_8 FILLER_12_185 ();
 sg13g2_decap_8 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_199 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_fill_1 FILLER_12_218 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_fill_2 FILLER_12_241 ();
 sg13g2_fill_2 FILLER_12_259 ();
 sg13g2_fill_2 FILLER_12_292 ();
 sg13g2_fill_1 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_304 ();
 sg13g2_fill_2 FILLER_12_311 ();
 sg13g2_fill_1 FILLER_12_319 ();
 sg13g2_fill_2 FILLER_12_335 ();
 sg13g2_fill_1 FILLER_12_337 ();
 sg13g2_fill_1 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_9 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_fill_1 FILLER_13_25 ();
 sg13g2_fill_2 FILLER_13_31 ();
 sg13g2_fill_1 FILLER_13_33 ();
 sg13g2_decap_8 FILLER_13_43 ();
 sg13g2_decap_4 FILLER_13_50 ();
 sg13g2_fill_1 FILLER_13_54 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_fill_2 FILLER_13_69 ();
 sg13g2_fill_1 FILLER_13_71 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_decap_8 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_106 ();
 sg13g2_fill_1 FILLER_13_108 ();
 sg13g2_fill_2 FILLER_13_119 ();
 sg13g2_decap_4 FILLER_13_286 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_decap_4 FILLER_13_322 ();
 sg13g2_decap_4 FILLER_13_334 ();
 sg13g2_fill_2 FILLER_13_338 ();
 sg13g2_fill_1 FILLER_13_347 ();
 sg13g2_fill_1 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_30 ();
 sg13g2_fill_1 FILLER_14_101 ();
 sg13g2_fill_2 FILLER_14_110 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_fill_2 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_145 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_decap_4 FILLER_14_164 ();
 sg13g2_fill_1 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_4 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_fill_2 FILLER_14_262 ();
 sg13g2_fill_2 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_fill_1 FILLER_14_324 ();
 sg13g2_decap_4 FILLER_14_338 ();
 sg13g2_fill_2 FILLER_14_362 ();
 sg13g2_fill_1 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_4 FILLER_14_377 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_fill_1 FILLER_15_25 ();
 sg13g2_decap_4 FILLER_15_44 ();
 sg13g2_fill_1 FILLER_15_48 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_4 FILLER_15_74 ();
 sg13g2_fill_2 FILLER_15_87 ();
 sg13g2_decap_8 FILLER_15_94 ();
 sg13g2_decap_4 FILLER_15_126 ();
 sg13g2_fill_1 FILLER_15_130 ();
 sg13g2_fill_2 FILLER_15_149 ();
 sg13g2_fill_1 FILLER_15_160 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_decap_4 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_195 ();
 sg13g2_decap_8 FILLER_15_202 ();
 sg13g2_fill_2 FILLER_15_209 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_1 FILLER_15_220 ();
 sg13g2_decap_4 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_251 ();
 sg13g2_fill_1 FILLER_15_270 ();
 sg13g2_fill_1 FILLER_15_281 ();
 sg13g2_fill_2 FILLER_15_295 ();
 sg13g2_fill_1 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_343 ();
 sg13g2_fill_2 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_fill_2 FILLER_15_372 ();
 sg13g2_fill_1 FILLER_15_374 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_16_61 ();
 sg13g2_fill_1 FILLER_16_73 ();
 sg13g2_fill_2 FILLER_16_107 ();
 sg13g2_fill_1 FILLER_16_109 ();
 sg13g2_decap_4 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_123 ();
 sg13g2_decap_4 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_fill_1 FILLER_16_281 ();
 sg13g2_decap_4 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_fill_1 FILLER_16_354 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_fill_1 FILLER_17_31 ();
 sg13g2_decap_8 FILLER_17_41 ();
 sg13g2_decap_4 FILLER_17_48 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_76 ();
 sg13g2_decap_8 FILLER_17_86 ();
 sg13g2_decap_4 FILLER_17_93 ();
 sg13g2_fill_2 FILLER_17_97 ();
 sg13g2_fill_2 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_118 ();
 sg13g2_decap_8 FILLER_17_124 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_174 ();
 sg13g2_fill_2 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_4 FILLER_17_209 ();
 sg13g2_fill_2 FILLER_17_233 ();
 sg13g2_fill_1 FILLER_17_235 ();
 sg13g2_decap_8 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_decap_8 FILLER_17_271 ();
 sg13g2_decap_8 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_285 ();
 sg13g2_fill_1 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_4 FILLER_17_329 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_decap_4 FILLER_17_339 ();
 sg13g2_fill_2 FILLER_17_343 ();
 sg13g2_fill_2 FILLER_17_363 ();
 sg13g2_decap_4 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_373 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_54 ();
 sg13g2_fill_1 FILLER_18_56 ();
 sg13g2_fill_2 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_156 ();
 sg13g2_fill_1 FILLER_18_158 ();
 sg13g2_fill_2 FILLER_18_164 ();
 sg13g2_fill_1 FILLER_18_166 ();
 sg13g2_decap_8 FILLER_18_181 ();
 sg13g2_decap_4 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_decap_4 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_232 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_250 ();
 sg13g2_fill_2 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_fill_2 FILLER_18_309 ();
 sg13g2_fill_1 FILLER_18_311 ();
 sg13g2_decap_4 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_346 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_4 FILLER_19_21 ();
 sg13g2_fill_2 FILLER_19_25 ();
 sg13g2_decap_4 FILLER_19_53 ();
 sg13g2_fill_1 FILLER_19_57 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_fill_2 FILLER_19_97 ();
 sg13g2_fill_1 FILLER_19_99 ();
 sg13g2_decap_8 FILLER_19_108 ();
 sg13g2_decap_4 FILLER_19_141 ();
 sg13g2_decap_4 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_162 ();
 sg13g2_decap_8 FILLER_19_204 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_decap_4 FILLER_19_281 ();
 sg13g2_decap_4 FILLER_19_311 ();
 sg13g2_fill_1 FILLER_19_327 ();
 sg13g2_fill_2 FILLER_19_333 ();
 sg13g2_fill_1 FILLER_19_335 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_348 ();
 sg13g2_fill_1 FILLER_19_350 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_19_380 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_decap_8 FILLER_20_38 ();
 sg13g2_fill_2 FILLER_20_45 ();
 sg13g2_decap_4 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_69 ();
 sg13g2_decap_8 FILLER_20_76 ();
 sg13g2_decap_4 FILLER_20_83 ();
 sg13g2_fill_2 FILLER_20_92 ();
 sg13g2_fill_1 FILLER_20_94 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_122 ();
 sg13g2_fill_2 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_decap_8 FILLER_20_176 ();
 sg13g2_decap_8 FILLER_20_183 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_4 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_283 ();
 sg13g2_decap_4 FILLER_20_317 ();
 sg13g2_fill_2 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_354 ();
 sg13g2_fill_2 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_2 FILLER_21_44 ();
 sg13g2_fill_2 FILLER_21_55 ();
 sg13g2_fill_1 FILLER_21_113 ();
 sg13g2_decap_8 FILLER_21_128 ();
 sg13g2_decap_8 FILLER_21_135 ();
 sg13g2_decap_8 FILLER_21_142 ();
 sg13g2_fill_2 FILLER_21_185 ();
 sg13g2_fill_2 FILLER_21_192 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_decap_4 FILLER_21_223 ();
 sg13g2_fill_2 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_295 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_decap_4 FILLER_21_323 ();
 sg13g2_fill_2 FILLER_21_327 ();
 sg13g2_decap_4 FILLER_21_339 ();
 sg13g2_decap_4 FILLER_21_348 ();
 sg13g2_fill_1 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_4 FILLER_21_383 ();
 sg13g2_fill_2 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_56 ();
 sg13g2_decap_4 FILLER_22_62 ();
 sg13g2_fill_2 FILLER_22_66 ();
 sg13g2_fill_2 FILLER_22_89 ();
 sg13g2_fill_2 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_99 ();
 sg13g2_fill_1 FILLER_22_110 ();
 sg13g2_decap_4 FILLER_22_156 ();
 sg13g2_fill_1 FILLER_22_160 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_fill_1 FILLER_22_180 ();
 sg13g2_decap_4 FILLER_22_207 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_237 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_decap_4 FILLER_22_323 ();
 sg13g2_fill_1 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_346 ();
 sg13g2_fill_1 FILLER_22_348 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_38 ();
 sg13g2_decap_4 FILLER_23_45 ();
 sg13g2_decap_8 FILLER_23_54 ();
 sg13g2_fill_1 FILLER_23_61 ();
 sg13g2_decap_8 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_73 ();
 sg13g2_fill_2 FILLER_23_86 ();
 sg13g2_decap_4 FILLER_23_103 ();
 sg13g2_fill_2 FILLER_23_107 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_4 FILLER_23_130 ();
 sg13g2_fill_2 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_146 ();
 sg13g2_decap_8 FILLER_23_160 ();
 sg13g2_decap_4 FILLER_23_167 ();
 sg13g2_fill_2 FILLER_23_171 ();
 sg13g2_fill_2 FILLER_23_178 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_4 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_214 ();
 sg13g2_fill_2 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_241 ();
 sg13g2_decap_8 FILLER_23_246 ();
 sg13g2_decap_4 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_decap_4 FILLER_23_263 ();
 sg13g2_fill_2 FILLER_23_267 ();
 sg13g2_fill_2 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_decap_4 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_291 ();
 sg13g2_fill_1 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_decap_4 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_104 ();
 sg13g2_decap_4 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_115 ();
 sg13g2_decap_4 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_fill_1 FILLER_24_148 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_decap_4 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_195 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_fill_2 FILLER_24_222 ();
 sg13g2_fill_1 FILLER_24_224 ();
 sg13g2_fill_2 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_267 ();
 sg13g2_fill_1 FILLER_24_269 ();
 sg13g2_decap_4 FILLER_24_278 ();
 sg13g2_decap_4 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_decap_4 FILLER_24_319 ();
 sg13g2_fill_2 FILLER_24_323 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_4 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_358 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_36 ();
 sg13g2_fill_1 FILLER_25_38 ();
 sg13g2_decap_4 FILLER_25_43 ();
 sg13g2_decap_4 FILLER_25_52 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_1 FILLER_25_89 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_fill_2 FILLER_25_134 ();
 sg13g2_fill_2 FILLER_25_141 ();
 sg13g2_fill_2 FILLER_25_148 ();
 sg13g2_fill_2 FILLER_25_157 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_fill_2 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_222 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_271 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_decap_8 FILLER_25_302 ();
 sg13g2_fill_2 FILLER_25_309 ();
 sg13g2_fill_1 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_318 ();
 sg13g2_fill_2 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_358 ();
 sg13g2_fill_2 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_fill_2 FILLER_25_377 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_39 ();
 sg13g2_fill_2 FILLER_26_50 ();
 sg13g2_fill_1 FILLER_26_52 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_decap_4 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_fill_2 FILLER_26_118 ();
 sg13g2_decap_8 FILLER_26_146 ();
 sg13g2_decap_8 FILLER_26_157 ();
 sg13g2_fill_1 FILLER_26_170 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_decap_8 FILLER_26_202 ();
 sg13g2_fill_2 FILLER_26_209 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_4 FILLER_26_301 ();
 sg13g2_fill_2 FILLER_26_305 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_fill_2 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_fill_1 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_30 ();
 sg13g2_fill_1 FILLER_27_36 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_decap_4 FILLER_27_71 ();
 sg13g2_fill_2 FILLER_27_75 ();
 sg13g2_fill_1 FILLER_27_81 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_123 ();
 sg13g2_decap_4 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_fill_2 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_decap_4 FILLER_27_277 ();
 sg13g2_decap_4 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_decap_8 FILLER_28_96 ();
 sg13g2_fill_2 FILLER_28_103 ();
 sg13g2_decap_4 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_115 ();
 sg13g2_decap_8 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_fill_1 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_237 ();
 sg13g2_fill_2 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_decap_8 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_4 FILLER_28_348 ();
 sg13g2_fill_1 FILLER_28_352 ();
 sg13g2_decap_4 FILLER_28_369 ();
 sg13g2_fill_2 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_39 ();
 sg13g2_fill_2 FILLER_29_45 ();
 sg13g2_fill_1 FILLER_29_47 ();
 sg13g2_fill_2 FILLER_29_74 ();
 sg13g2_fill_1 FILLER_29_76 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_decap_4 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_fill_1 FILLER_29_186 ();
 sg13g2_decap_4 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_275 ();
 sg13g2_decap_8 FILLER_29_282 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_decap_4 FILLER_29_318 ();
 sg13g2_fill_1 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_decap_4 FILLER_29_347 ();
 sg13g2_decap_4 FILLER_29_375 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_58 ();
 sg13g2_decap_8 FILLER_30_85 ();
 sg13g2_fill_1 FILLER_30_92 ();
 sg13g2_decap_4 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_decap_4 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_decap_8 FILLER_30_241 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_decap_4 FILLER_30_386 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_4 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_fill_2 FILLER_31_135 ();
 sg13g2_decap_4 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_176 ();
 sg13g2_decap_4 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_4 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_decap_4 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_decap_4 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_342 ();
 sg13g2_decap_4 FILLER_31_371 ();
 sg13g2_fill_1 FILLER_31_379 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_4 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_60 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_fill_1 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_fill_2 FILLER_32_152 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_204 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_4 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_decap_4 FILLER_32_319 ();
 sg13g2_fill_2 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_116 ();
 sg13g2_fill_2 FILLER_33_123 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_decap_8 FILLER_33_152 ();
 sg13g2_decap_8 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_243 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_4 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_107 ();
 sg13g2_decap_4 FILLER_34_137 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_fill_2 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_decap_8 FILLER_34_267 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_293 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_fill_2 FILLER_34_305 ();
 sg13g2_fill_1 FILLER_34_307 ();
 sg13g2_fill_2 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_378 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_185 ();
 sg13g2_fill_1 FILLER_35_198 ();
 sg13g2_fill_1 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_252 ();
 sg13g2_fill_2 FILLER_35_270 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_342 ();
 sg13g2_fill_2 FILLER_35_380 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_2 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_137 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_363 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_4 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_189 ();
 sg13g2_decap_4 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_275 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_362 ();
 sg13g2_fill_2 FILLER_37_373 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_8 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_4 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_4 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_decap_4 FILLER_38_216 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_decap_4 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_280 ();
 sg13g2_fill_1 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_379 ();
 sg13g2_fill_1 FILLER_38_381 ();
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net2;
 assign uio_oe[3] = net3;
 assign uio_oe[4] = net4;
 assign uio_oe[5] = net5;
 assign uio_oe[6] = net6;
 assign uio_oe[7] = net7;
 assign uio_out[5] = net8;
 assign uio_out[6] = net9;
 assign uio_out[7] = net10;
endmodule

module tt_um_wokwi_group_3 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire net174;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire \proj_10.net10 ;
 wire \proj_10.net11 ;
 wire \proj_10.net12 ;
 wire \proj_10.net13 ;
 wire \proj_10.net9 ;
 wire \proj_12.net10 ;
 wire \proj_12.net11 ;
 wire \proj_12.net12 ;
 wire \proj_12.net13 ;
 wire \proj_12.net18 ;
 wire \proj_12.net19 ;
 wire \proj_12.net20 ;
 wire \proj_12.net21 ;
 wire \proj_12.net22 ;
 wire \proj_12.net23 ;
 wire \proj_12.net24 ;
 wire \proj_12.net25 ;
 wire \proj_12.net26 ;
 wire \proj_12.net27 ;
 wire \proj_12.net28 ;
 wire \proj_12.net29 ;
 wire \proj_12.net9 ;
 wire \proj_13.net12 ;
 wire \proj_13.net13 ;
 wire \proj_13.net7 ;
 wire \proj_13.net8 ;
 wire \proj_14.net100 ;
 wire \proj_14.net101 ;
 wire \proj_14.net102 ;
 wire \proj_14.net104 ;
 wire \proj_14.net105 ;
 wire \proj_14.net106 ;
 wire \proj_14.net108 ;
 wire \proj_14.net11 ;
 wire \proj_14.net110 ;
 wire \proj_14.net111 ;
 wire \proj_14.net112 ;
 wire \proj_14.net114 ;
 wire \proj_14.net115 ;
 wire \proj_14.net116 ;
 wire \proj_14.net117 ;
 wire \proj_14.net119 ;
 wire \proj_14.net12 ;
 wire \proj_14.net120 ;
 wire \proj_14.net121 ;
 wire \proj_14.net122 ;
 wire \proj_14.net124 ;
 wire \proj_14.net125 ;
 wire \proj_14.net126 ;
 wire \proj_14.net127 ;
 wire \proj_14.net129 ;
 wire \proj_14.net13 ;
 wire \proj_14.net130 ;
 wire \proj_14.net131 ;
 wire \proj_14.net132 ;
 wire \proj_14.net133 ;
 wire \proj_14.net135 ;
 wire \proj_14.net136 ;
 wire \proj_14.net137 ;
 wire \proj_14.net138 ;
 wire \proj_14.net14 ;
 wire \proj_14.net140 ;
 wire \proj_14.net141 ;
 wire \proj_14.net142 ;
 wire \proj_14.net143 ;
 wire \proj_14.net145 ;
 wire \proj_14.net146 ;
 wire \proj_14.net147 ;
 wire \proj_14.net148 ;
 wire \proj_14.net15 ;
 wire \proj_14.net150 ;
 wire \proj_14.net151 ;
 wire \proj_14.net152 ;
 wire \proj_14.net153 ;
 wire \proj_14.net155 ;
 wire \proj_14.net156 ;
 wire \proj_14.net157 ;
 wire \proj_14.net158 ;
 wire \proj_14.net16 ;
 wire \proj_14.net160 ;
 wire \proj_14.net161 ;
 wire \proj_14.net162 ;
 wire \proj_14.net163 ;
 wire \proj_14.net165 ;
 wire \proj_14.net166 ;
 wire \proj_14.net167 ;
 wire \proj_14.net168 ;
 wire \proj_14.net17 ;
 wire \proj_14.net170 ;
 wire \proj_14.net171 ;
 wire \proj_14.net172 ;
 wire \proj_14.net173 ;
 wire \proj_14.net175 ;
 wire \proj_14.net176 ;
 wire \proj_14.net177 ;
 wire \proj_14.net178 ;
 wire \proj_14.net180 ;
 wire \proj_14.net181 ;
 wire \proj_14.net182 ;
 wire \proj_14.net183 ;
 wire \proj_14.net184 ;
 wire \proj_14.net185 ;
 wire \proj_14.net186 ;
 wire \proj_14.net187 ;
 wire \proj_14.net188 ;
 wire \proj_14.net189 ;
 wire \proj_14.net190 ;
 wire \proj_14.net191 ;
 wire \proj_14.net192 ;
 wire \proj_14.net193 ;
 wire \proj_14.net194 ;
 wire \proj_14.net195 ;
 wire \proj_14.net196 ;
 wire \proj_14.net197 ;
 wire \proj_14.net198 ;
 wire \proj_14.net199 ;
 wire \proj_14.net200 ;
 wire \proj_14.net201 ;
 wire \proj_14.net202 ;
 wire \proj_14.net203 ;
 wire \proj_14.net204 ;
 wire \proj_14.net205 ;
 wire \proj_14.net206 ;
 wire \proj_14.net207 ;
 wire \proj_14.net209 ;
 wire \proj_14.net210 ;
 wire \proj_14.net211 ;
 wire \proj_14.net212 ;
 wire \proj_14.net214 ;
 wire \proj_14.net215 ;
 wire \proj_14.net216 ;
 wire \proj_14.net217 ;
 wire \proj_14.net218 ;
 wire \proj_14.net219 ;
 wire \proj_14.net220 ;
 wire \proj_14.net221 ;
 wire \proj_14.net222 ;
 wire \proj_14.net223 ;
 wire \proj_14.net224 ;
 wire \proj_14.net226 ;
 wire \proj_14.net227 ;
 wire \proj_14.net228 ;
 wire \proj_14.net229 ;
 wire \proj_14.net23 ;
 wire \proj_14.net231 ;
 wire \proj_14.net232 ;
 wire \proj_14.net233 ;
 wire \proj_14.net234 ;
 wire \proj_14.net235 ;
 wire \proj_14.net236 ;
 wire \proj_14.net237 ;
 wire \proj_14.net238 ;
 wire \proj_14.net239 ;
 wire \proj_14.net240 ;
 wire \proj_14.net241 ;
 wire \proj_14.net242 ;
 wire \proj_14.net243 ;
 wire \proj_14.net244 ;
 wire \proj_14.net245 ;
 wire \proj_14.net246 ;
 wire \proj_14.net247 ;
 wire \proj_14.net248 ;
 wire \proj_14.net249 ;
 wire \proj_14.net25 ;
 wire \proj_14.net250 ;
 wire \proj_14.net251 ;
 wire \proj_14.net252 ;
 wire \proj_14.net253 ;
 wire \proj_14.net254 ;
 wire \proj_14.net255 ;
 wire \proj_14.net256 ;
 wire \proj_14.net257 ;
 wire \proj_14.net258 ;
 wire \proj_14.net259 ;
 wire \proj_14.net26 ;
 wire \proj_14.net260 ;
 wire \proj_14.net261 ;
 wire \proj_14.net262 ;
 wire \proj_14.net263 ;
 wire \proj_14.net264 ;
 wire \proj_14.net265 ;
 wire \proj_14.net266 ;
 wire \proj_14.net267 ;
 wire \proj_14.net268 ;
 wire \proj_14.net269 ;
 wire \proj_14.net27 ;
 wire \proj_14.net270 ;
 wire \proj_14.net271 ;
 wire \proj_14.net272 ;
 wire \proj_14.net273 ;
 wire \proj_14.net274 ;
 wire \proj_14.net275 ;
 wire \proj_14.net276 ;
 wire \proj_14.net277 ;
 wire \proj_14.net278 ;
 wire \proj_14.net279 ;
 wire \proj_14.net28 ;
 wire \proj_14.net280 ;
 wire \proj_14.net281 ;
 wire \proj_14.net282 ;
 wire \proj_14.net283 ;
 wire \proj_14.net284 ;
 wire \proj_14.net285 ;
 wire \proj_14.net286 ;
 wire \proj_14.net287 ;
 wire \proj_14.net288 ;
 wire \proj_14.net289 ;
 wire \proj_14.net29 ;
 wire \proj_14.net30 ;
 wire \proj_14.net31 ;
 wire \proj_14.net32 ;
 wire \proj_14.net33 ;
 wire \proj_14.net34 ;
 wire \proj_14.net36 ;
 wire \proj_14.net37 ;
 wire \proj_14.net38 ;
 wire \proj_14.net39 ;
 wire \proj_14.net40 ;
 wire \proj_14.net41 ;
 wire \proj_14.net42 ;
 wire \proj_14.net43 ;
 wire \proj_14.net44 ;
 wire \proj_14.net45 ;
 wire \proj_14.net46 ;
 wire \proj_14.net47 ;
 wire \proj_14.net48 ;
 wire \proj_14.net50 ;
 wire \proj_14.net51 ;
 wire \proj_14.net52 ;
 wire \proj_14.net53 ;
 wire \proj_14.net54 ;
 wire \proj_14.net55 ;
 wire \proj_14.net56 ;
 wire \proj_14.net57 ;
 wire \proj_14.net58 ;
 wire \proj_14.net59 ;
 wire \proj_14.net60 ;
 wire \proj_14.net61 ;
 wire \proj_14.net62 ;
 wire \proj_14.net63 ;
 wire \proj_14.net64 ;
 wire \proj_14.net65 ;
 wire \proj_14.net66 ;
 wire \proj_14.net67 ;
 wire \proj_14.net68 ;
 wire \proj_14.net69 ;
 wire \proj_14.net70 ;
 wire \proj_14.net71 ;
 wire \proj_14.net72 ;
 wire \proj_14.net73 ;
 wire \proj_14.net74 ;
 wire \proj_14.net75 ;
 wire \proj_14.net76 ;
 wire \proj_14.net77 ;
 wire \proj_14.net78 ;
 wire \proj_14.net79 ;
 wire \proj_14.net80 ;
 wire \proj_14.net81 ;
 wire \proj_14.net82 ;
 wire \proj_14.net83 ;
 wire \proj_14.net84 ;
 wire \proj_14.net85 ;
 wire \proj_14.net86 ;
 wire \proj_14.net87 ;
 wire \proj_14.net88 ;
 wire \proj_14.net89 ;
 wire \proj_14.net90 ;
 wire \proj_14.net91 ;
 wire \proj_14.net92 ;
 wire \proj_14.net93 ;
 wire \proj_14.net94 ;
 wire \proj_14.net95 ;
 wire \proj_14.net96 ;
 wire \proj_14.net97 ;
 wire \proj_14.net98 ;
 wire \proj_14.net99 ;
 wire \proj_15.net15 ;
 wire \proj_15.net16 ;
 wire \proj_15.net17 ;
 wire \proj_15.net18 ;
 wire \proj_15.net7 ;
 wire \proj_15.net8 ;
 wire \proj_15.net9 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__0.net9 ;
 wire \proj__1.net10 ;
 wire \proj__1.net16 ;
 wire \proj__1.net17 ;
 wire \proj__1.net18 ;
 wire \proj__1.net19 ;
 wire \proj__1.net20 ;
 wire \proj__1.net21 ;
 wire \proj__1.net22 ;
 wire \proj__1.net23 ;
 wire \proj__1.net24 ;
 wire \proj__1.net9 ;
 wire \proj__2.net10 ;
 wire \proj__2.net11 ;
 wire \proj__2.net12 ;
 wire \proj__2.net9 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net3 ;
 wire \proj__3.net4 ;
 wire \proj__3.net5 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net13 ;
 wire \proj__4.net14 ;
 wire \proj__4.net15 ;
 wire \proj__4.net16 ;
 wire \proj__4.net17 ;
 wire \proj__4.net18 ;
 wire \proj__5.net10 ;
 wire \proj__5.net11 ;
 wire \proj__5.net12 ;
 wire \proj__5.net9 ;
 wire \proj__6.net10 ;
 wire \proj__6.net9 ;
 wire \proj__7.net14 ;
 wire \proj__7.net15 ;
 wire \proj__7.net5 ;
 wire \proj__7.net6 ;
 wire \proj__7.net7 ;
 wire \proj__7.net8 ;
 wire \proj__8.net7 ;
 wire \proj__9.net11 ;
 wire \proj__9.net12 ;
 wire \proj__9.net13 ;
 wire \proj__9.net14 ;
 wire \proj__9.net15 ;
 wire \proj__9.net17 ;
 wire \proj__9.net5 ;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire \proj_10.nand1/b ;
 wire net175;
 wire \proj_13.flop1/notq ;
 wire net176;
 wire \proj_13.flop2/notq ;
 wire net177;
 wire \proj_13.flop3/notq ;
 wire \proj_14.flop1/_0_ ;
 wire \proj_14.flop1/_1_ ;
 wire net63;
 wire net64;
 wire \proj_14.flop10/_0_ ;
 wire \proj_14.flop10/_1_ ;
 wire net65;
 wire net66;
 wire \proj_14.flop11/_0_ ;
 wire \proj_14.flop11/_1_ ;
 wire net88;
 wire net89;
 wire \proj_14.flop12/_0_ ;
 wire \proj_14.flop12/_1_ ;
 wire net90;
 wire net91;
 wire \proj_14.flop13/_0_ ;
 wire \proj_14.flop13/_1_ ;
 wire net92;
 wire net93;
 wire \proj_14.flop14/_0_ ;
 wire \proj_14.flop14/_1_ ;
 wire net94;
 wire net95;
 wire \proj_14.flop15/_0_ ;
 wire \proj_14.flop15/_1_ ;
 wire net96;
 wire net97;
 wire \proj_14.flop16/_0_ ;
 wire \proj_14.flop16/_1_ ;
 wire net98;
 wire net99;
 wire \proj_14.flop17/_0_ ;
 wire \proj_14.flop17/_1_ ;
 wire net100;
 wire net101;
 wire \proj_14.flop18/_0_ ;
 wire \proj_14.flop18/_1_ ;
 wire net102;
 wire net103;
 wire \proj_14.flop19/_0_ ;
 wire \proj_14.flop19/_1_ ;
 wire net104;
 wire net105;
 wire \proj_14.flop2/_0_ ;
 wire \proj_14.flop2/_1_ ;
 wire net106;
 wire net107;
 wire \proj_14.flop20/_0_ ;
 wire \proj_14.flop20/_1_ ;
 wire net108;
 wire net109;
 wire \proj_14.flop21/_0_ ;
 wire \proj_14.flop21/_1_ ;
 wire net110;
 wire net111;
 wire \proj_14.flop22/_0_ ;
 wire \proj_14.flop22/_1_ ;
 wire net112;
 wire net113;
 wire \proj_14.flop23/_0_ ;
 wire \proj_14.flop23/_1_ ;
 wire net114;
 wire net115;
 wire \proj_14.flop24/_0_ ;
 wire \proj_14.flop24/_1_ ;
 wire net116;
 wire net117;
 wire \proj_14.flop25/_0_ ;
 wire \proj_14.flop25/_1_ ;
 wire net118;
 wire net119;
 wire \proj_14.flop25/notq ;
 wire \proj_14.flop26/_0_ ;
 wire \proj_14.flop26/_1_ ;
 wire net120;
 wire net121;
 wire \proj_14.flop26/notq ;
 wire \proj_14.flop27/_0_ ;
 wire \proj_14.flop27/_1_ ;
 wire net122;
 wire net123;
 wire \proj_14.flop27/q ;
 wire net178;
 wire \proj_14.flop28/notq ;
 wire \proj_14.flop29/_0_ ;
 wire \proj_14.flop29/_1_ ;
 wire net124;
 wire net125;
 wire \proj_14.flop3/_0_ ;
 wire \proj_14.flop3/_1_ ;
 wire net126;
 wire net127;
 wire \proj_14.flop30/_0_ ;
 wire \proj_14.flop30/_1_ ;
 wire net128;
 wire net129;
 wire \proj_14.flop31/_0_ ;
 wire \proj_14.flop31/_1_ ;
 wire net130;
 wire net131;
 wire \proj_14.flop31/notq ;
 wire \proj_14.flop32/_0_ ;
 wire \proj_14.flop32/_1_ ;
 wire net132;
 wire net133;
 wire \proj_14.flop32/notq ;
 wire \proj_14.flop33/_0_ ;
 wire \proj_14.flop33/_1_ ;
 wire net134;
 wire net135;
 wire \proj_14.flop33/notq ;
 wire \proj_14.flop34/_0_ ;
 wire \proj_14.flop34/_1_ ;
 wire net136;
 wire net137;
 wire \proj_14.flop34/notq ;
 wire \proj_14.flop35/_0_ ;
 wire \proj_14.flop35/_1_ ;
 wire net138;
 wire net139;
 wire \proj_14.flop35/notq ;
 wire \proj_14.flop36/_0_ ;
 wire \proj_14.flop36/_1_ ;
 wire net140;
 wire net141;
 wire \proj_14.flop36/notq ;
 wire \proj_14.flop37/_0_ ;
 wire \proj_14.flop37/_1_ ;
 wire net142;
 wire net143;
 wire \proj_14.flop37/notq ;
 wire \proj_14.flop4/_0_ ;
 wire \proj_14.flop4/_1_ ;
 wire net144;
 wire net145;
 wire net179;
 wire \proj_14.flop46/notq ;
 wire net180;
 wire \proj_14.flop47/notq ;
 wire net181;
 wire \proj_14.flop48/notq ;
 wire net182;
 wire \proj_14.flop49/notq ;
 wire \proj_14.flop5/_0_ ;
 wire \proj_14.flop5/_1_ ;
 wire net146;
 wire net147;
 wire net183;
 wire \proj_14.flop50/notq ;
 wire net184;
 wire \proj_14.flop51/notq ;
 wire net185;
 wire \proj_14.flop52/notq ;
 wire net186;
 wire \proj_14.flop53/notq ;
 wire net187;
 wire \proj_14.flop54/notq ;
 wire net188;
 wire \proj_14.flop55/notq ;
 wire net189;
 wire \proj_14.flop56/notq ;
 wire \proj_14.flop6/_0_ ;
 wire \proj_14.flop6/_1_ ;
 wire net148;
 wire net149;
 wire \proj_14.flop7/_0_ ;
 wire \proj_14.flop7/_1_ ;
 wire net150;
 wire net151;
 wire \proj_14.flop8/_0_ ;
 wire \proj_14.flop8/_1_ ;
 wire net152;
 wire net153;
 wire \proj_14.flop9/_0_ ;
 wire \proj_14.flop9/_1_ ;
 wire net154;
 wire net155;
 wire \proj__4.flop1/_0_ ;
 wire \proj__4.flop1/_1_ ;
 wire net156;
 wire net157;
 wire \proj__4.flop1/q ;
 wire \proj__4.flop1/s ;
 wire \proj__4.flop2/_0_ ;
 wire \proj__4.flop2/_1_ ;
 wire net158;
 wire net159;
 wire \proj__4.flop2/q ;
 wire \proj__4.flop2/s ;
 wire \proj__4.flop3/_0_ ;
 wire \proj__4.flop3/_1_ ;
 wire net160;
 wire net161;
 wire \proj__4.flop3/q ;
 wire \proj__4.flop3/s ;
 wire \proj__4.flop4/_0_ ;
 wire \proj__4.flop4/_1_ ;
 wire net162;
 wire net163;
 wire \proj__4.flop4/q ;
 wire \proj__4.flop4/s ;
 wire \proj__4.flop5/_0_ ;
 wire \proj__4.flop5/_1_ ;
 wire net164;
 wire net165;
 wire \proj__4.flop5/notq ;
 wire \proj__4.flop5/s ;
 wire \proj__4.flop6/_0_ ;
 wire \proj__4.flop6/_1_ ;
 wire net166;
 wire net167;
 wire \proj__4.flop6/notq ;
 wire \proj__4.flop6/s ;
 wire \proj__4.flop8/_0_ ;
 wire \proj__4.flop8/_1_ ;
 wire net168;
 wire net169;
 wire \proj__4.flop8/notq ;
 wire \proj__4.flop8/s ;
 wire \proj__4.flop9/_0_ ;
 wire \proj__4.flop9/_1_ ;
 wire net170;
 wire net171;
 wire \proj__4.flop9/notq ;
 wire \proj__4.flop9/s ;
 wire net190;
 wire net191;
 wire clk_regs;
 wire \proj__9.flop1/_0_ ;
 wire \proj__9.flop1/_1_ ;
 wire net172;
 wire net173;
 wire \proj__9.flop1/notq ;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;

 sg13g2_inv_1 _115_ (.Y(_053_),
    .A(net6));
 sg13g2_inv_1 _116_ (.Y(_054_),
    .A(net9));
 sg13g2_inv_1 _117_ (.Y(_055_),
    .A(net8));
 sg13g2_inv_1 _118_ (.Y(_056_),
    .A(\proj__0.net9 ));
 sg13g2_inv_1 _119_ (.Y(_057_),
    .A(\proj__0.net10 ));
 sg13g2_nor2b_2 _120_ (.A(net9),
    .B_N(net8),
    .Y(_058_));
 sg13g2_nor2b_1 _121_ (.A(net7),
    .B_N(net6),
    .Y(_059_));
 sg13g2_and2_2 _122_ (.A(_058_),
    .B(_059_),
    .X(_060_));
 sg13g2_nand2_2 _123_ (.Y(_061_),
    .A(net9),
    .B(net8));
 sg13g2_nor2b_1 _124_ (.A(net6),
    .B_N(net7),
    .Y(_062_));
 sg13g2_nor2_2 _125_ (.A(net6),
    .B(net7),
    .Y(_063_));
 sg13g2_a22oi_1 _126_ (.Y(_064_),
    .B1(_063_),
    .B2(_055_),
    .A2(net75),
    .A1(_054_));
 sg13g2_o21ai_1 _127_ (.B1(_064_),
    .Y(_065_),
    .A1(_053_),
    .A2(_061_));
 sg13g2_o21ai_1 _128_ (.B1(net5),
    .Y(_066_),
    .A1(_060_),
    .A2(_065_));
 sg13g2_nor2b_2 _129_ (.A(net8),
    .B_N(net9),
    .Y(_067_));
 sg13g2_and2_2 _130_ (.A(_062_),
    .B(_067_),
    .X(_068_));
 sg13g2_and2_1 _131_ (.A(net6),
    .B(net7),
    .X(_069_));
 sg13g2_and2_2 _132_ (.A(_058_),
    .B(_069_),
    .X(_070_));
 sg13g2_nand2_1 _133_ (.Y(_071_),
    .A(_058_),
    .B(_069_));
 sg13g2_and2_2 _134_ (.A(_058_),
    .B(_063_),
    .X(_072_));
 sg13g2_nand2_1 _135_ (.Y(_073_),
    .A(\proj__4.net18 ),
    .B(_072_));
 sg13g2_a22oi_1 _136_ (.Y(_074_),
    .B1(_070_),
    .B2(\proj__7.net8 ),
    .A2(_068_),
    .A1(\proj_10.net13 ));
 sg13g2_nand3_1 _137_ (.B(_073_),
    .C(_074_),
    .A(_066_),
    .Y(uo_out[7]));
 sg13g2_nor2_2 _138_ (.A(net9),
    .B(net8),
    .Y(_075_));
 sg13g2_and2_2 _139_ (.A(_063_),
    .B(_075_),
    .X(_076_));
 sg13g2_and2_1 _140_ (.A(\proj__4.net11 ),
    .B(_072_),
    .X(_077_));
 sg13g2_nand3_1 _141_ (.B(net75),
    .C(_067_),
    .A(\proj_10.net9 ),
    .Y(_000_));
 sg13g2_nor2b_2 _142_ (.A(_061_),
    .B_N(_063_),
    .Y(_001_));
 sg13g2_and2_1 _143_ (.A(_058_),
    .B(net75),
    .X(_002_));
 sg13g2_and2_1 _144_ (.A(_069_),
    .B(_075_),
    .X(_003_));
 sg13g2_a22oi_1 _145_ (.Y(_004_),
    .B1(_069_),
    .B2(_075_),
    .A2(net75),
    .A1(_058_));
 sg13g2_nor2b_1 _146_ (.A(_004_),
    .B_N(net84),
    .Y(_005_));
 sg13g2_nand3_1 _147_ (.B(net75),
    .C(_075_),
    .A(\proj__2.net9 ),
    .Y(_006_));
 sg13g2_nand3_1 _148_ (.B(_059_),
    .C(_067_),
    .A(\proj__9.net5 ),
    .Y(_007_));
 sg13g2_nor2b_2 _149_ (.A(_061_),
    .B_N(net75),
    .Y(_008_));
 sg13g2_and3_1 _150_ (.X(_009_),
    .A(\proj__8.net7 ),
    .B(_063_),
    .C(_067_));
 sg13g2_nor2b_2 _151_ (.A(_061_),
    .B_N(_069_),
    .Y(_010_));
 sg13g2_nor3_2 _152_ (.A(_053_),
    .B(net7),
    .C(_061_),
    .Y(_011_));
 sg13g2_a22oi_1 _153_ (.Y(_012_),
    .B1(_011_),
    .B2(\proj_13.net7 ),
    .A2(_010_),
    .A1(\proj_15.net7 ));
 sg13g2_nand3_1 _154_ (.B(_059_),
    .C(_075_),
    .A(\proj__1.net9 ),
    .Y(_013_));
 sg13g2_nand4_1 _155_ (.B(_006_),
    .C(_007_),
    .A(_000_),
    .Y(_014_),
    .D(_013_));
 sg13g2_nor4_1 _156_ (.A(_076_),
    .B(_077_),
    .C(_005_),
    .D(_014_),
    .Y(_015_));
 sg13g2_a22oi_1 _157_ (.Y(_016_),
    .B1(_008_),
    .B2(\proj_14.net11 ),
    .A2(_070_),
    .A1(\proj__7.net5 ));
 sg13g2_a221oi_1 _158_ (.B2(\proj_12.net9 ),
    .C1(_009_),
    .B1(_001_),
    .A1(\proj__5.net9 ),
    .Y(_017_),
    .A2(_060_));
 sg13g2_and3_1 _159_ (.X(_018_),
    .A(_012_),
    .B(_016_),
    .C(_017_));
 sg13g2_a22oi_1 _160_ (.Y(uo_out[0]),
    .B1(_015_),
    .B2(_018_),
    .A2(_076_),
    .A1(_056_));
 sg13g2_a22oi_1 _161_ (.Y(_019_),
    .B1(_070_),
    .B2(\proj__7.net6 ),
    .A2(_068_),
    .A1(net79));
 sg13g2_a22oi_1 _162_ (.Y(_020_),
    .B1(_011_),
    .B2(\proj_13.net8 ),
    .A2(_008_),
    .A1(\proj_14.net12 ));
 sg13g2_a22oi_1 _163_ (.Y(_021_),
    .B1(_010_),
    .B2(\proj_15.net8 ),
    .A2(_001_),
    .A1(\proj_12.net10 ));
 sg13g2_a21oi_1 _164_ (.A1(\proj__4.net12 ),
    .A2(_072_),
    .Y(_022_),
    .B1(_009_));
 sg13g2_nand3_1 _165_ (.B(_062_),
    .C(_075_),
    .A(\proj__2.net10 ),
    .Y(_023_));
 sg13g2_nand2b_1 _166_ (.Y(_024_),
    .B(net82),
    .A_N(_004_));
 sg13g2_and4_1 _167_ (.A(_021_),
    .B(_022_),
    .C(_023_),
    .D(_024_),
    .X(_025_));
 sg13g2_nand3_1 _168_ (.B(_020_),
    .C(_025_),
    .A(_019_),
    .Y(uo_out[1]));
 sg13g2_and2_1 _169_ (.A(\proj_12.net11 ),
    .B(_001_),
    .X(_026_));
 sg13g2_a221oi_1 _170_ (.B2(\proj__4.net13 ),
    .C1(_026_),
    .B1(_072_),
    .A1(clknet_1_0__leaf_clk),
    .Y(_027_),
    .A2(_070_));
 sg13g2_a21oi_1 _171_ (.A1(\proj_14.net13 ),
    .A2(_008_),
    .Y(_028_),
    .B1(_076_));
 sg13g2_a22oi_1 _172_ (.Y(_029_),
    .B1(_010_),
    .B2(\proj_15.net9 ),
    .A2(_002_),
    .A1(\proj__6.net9 ));
 sg13g2_nand3_1 _173_ (.B(net75),
    .C(_075_),
    .A(\proj__2.net11 ),
    .Y(_030_));
 sg13g2_a21oi_1 _174_ (.A1(net3),
    .A2(_068_),
    .Y(_031_),
    .B1(_009_));
 sg13g2_and4_1 _175_ (.A(_028_),
    .B(_029_),
    .C(_030_),
    .D(_031_),
    .X(_032_));
 sg13g2_a22oi_1 _176_ (.Y(uo_out[2]),
    .B1(_027_),
    .B2(_032_),
    .A2(_076_),
    .A1(_057_));
 sg13g2_nand2_1 _177_ (.Y(_033_),
    .A(\proj__6.net10 ),
    .B(_002_));
 sg13g2_nand2_1 _178_ (.Y(_034_),
    .A(\proj_12.net12 ),
    .B(_001_));
 sg13g2_and3_1 _179_ (.X(_035_),
    .A(\proj__2.net12 ),
    .B(net75),
    .C(_075_));
 sg13g2_a221oi_1 _180_ (.B2(\proj_14.net14 ),
    .C1(_035_),
    .B1(_008_),
    .A1(\proj__4.net14 ),
    .Y(_036_),
    .A2(_072_));
 sg13g2_nand4_1 _181_ (.B(_033_),
    .C(_034_),
    .A(_031_),
    .Y(_037_),
    .D(_036_));
 sg13g2_mux2_1 _182_ (.A0(_037_),
    .A1(\proj__0.net11 ),
    .S(_076_),
    .X(uo_out[3]));
 sg13g2_nand3b_1 _183_ (.B(_064_),
    .C(_071_),
    .Y(_038_),
    .A_N(_011_));
 sg13g2_nand2_1 _184_ (.Y(_039_),
    .A(net2),
    .B(_038_));
 sg13g2_nand2_1 _185_ (.Y(_040_),
    .A(\proj_10.net10 ),
    .B(_068_));
 sg13g2_nand2_1 _186_ (.Y(_041_),
    .A(\proj_14.net15 ),
    .B(_008_));
 sg13g2_a22oi_1 _187_ (.Y(_042_),
    .B1(_001_),
    .B2(\proj_12.net13 ),
    .A2(_060_),
    .A1(\proj__5.net10 ));
 sg13g2_a22oi_1 _188_ (.Y(_043_),
    .B1(_003_),
    .B2(\proj__3.net3 ),
    .A2(_072_),
    .A1(\proj__4.net15 ));
 sg13g2_and3_1 _189_ (.X(_044_),
    .A(_013_),
    .B(_040_),
    .C(_043_));
 sg13g2_nand4_1 _190_ (.B(_041_),
    .C(_042_),
    .A(_039_),
    .Y(uo_out[4]),
    .D(_044_));
 sg13g2_a22oi_1 _191_ (.Y(_045_),
    .B1(_072_),
    .B2(\proj__4.net16 ),
    .A2(_068_),
    .A1(\proj_10.net11 ));
 sg13g2_nand2_1 _192_ (.Y(_046_),
    .A(\proj_14.net16 ),
    .B(_008_));
 sg13g2_a22oi_1 _193_ (.Y(_047_),
    .B1(_003_),
    .B2(\proj__3.net4 ),
    .A2(_060_),
    .A1(\proj__5.net11 ));
 sg13g2_nand4_1 _194_ (.B(_045_),
    .C(_046_),
    .A(_013_),
    .Y(_048_),
    .D(_047_));
 sg13g2_a21o_2 _195_ (.A2(_038_),
    .A1(net76),
    .B1(_048_),
    .X(uo_out[5]));
 sg13g2_nand2_1 _196_ (.Y(_049_),
    .A(net4),
    .B(_065_));
 sg13g2_a22oi_1 _197_ (.Y(_050_),
    .B1(_003_),
    .B2(\proj__3.net5 ),
    .A2(_072_),
    .A1(\proj__4.net17 ));
 sg13g2_a22oi_1 _198_ (.Y(_051_),
    .B1(_070_),
    .B2(\proj__7.net7 ),
    .A2(_060_),
    .A1(\proj__5.net12 ));
 sg13g2_a22oi_1 _199_ (.Y(_052_),
    .B1(_008_),
    .B2(\proj_14.net17 ),
    .A2(_068_),
    .A1(\proj_10.net12 ));
 sg13g2_nand4_1 _200_ (.B(_050_),
    .C(_051_),
    .A(_049_),
    .Y(uo_out[6]),
    .D(_052_));
 sg13g2_tiehi \proj_13.flop1/_1__153  (.L_HI(net174));
 sg13g2_tielo \proj_14.flop10/_4__11  (.L_LO(net11));
 sg13g2_tielo \proj_14.flop11/_4__12  (.L_LO(net12));
 sg13g2_tielo \proj_14.flop12/_4__13  (.L_LO(net13));
 sg13g2_tielo \proj_14.flop13/_4__14  (.L_LO(net14));
 sg13g2_tielo \proj_14.flop14/_4__15  (.L_LO(net15));
 sg13g2_tielo \proj_14.flop15/_4__16  (.L_LO(net16));
 sg13g2_tielo \proj_14.flop16/_4__17  (.L_LO(net17));
 sg13g2_tielo \proj_14.flop17/_4__18  (.L_LO(net18));
 sg13g2_tielo \proj_14.flop18/_4__19  (.L_LO(net19));
 sg13g2_tielo \proj_14.flop19/_4__20  (.L_LO(net20));
 sg13g2_tielo \proj_14.flop2/_4__21  (.L_LO(net21));
 sg13g2_tielo \proj_14.flop20/_4__22  (.L_LO(net22));
 sg13g2_tielo \proj_14.flop21/_4__23  (.L_LO(net23));
 sg13g2_tielo \proj_14.flop22/_4__24  (.L_LO(net24));
 sg13g2_tielo \proj_14.flop23/_4__25  (.L_LO(net25));
 sg13g2_tielo \proj_14.flop24/_4__26  (.L_LO(net26));
 sg13g2_tielo \proj_14.flop25/_4__27  (.L_LO(net27));
 sg13g2_tielo \proj_14.flop26/_4__28  (.L_LO(net28));
 sg13g2_tielo \proj_14.flop27/_4__29  (.L_LO(net29));
 sg13g2_tielo \proj_14.flop29/_4__30  (.L_LO(net30));
 sg13g2_tielo \proj_14.flop3/_4__31  (.L_LO(net31));
 sg13g2_tielo \proj_14.flop30/_4__32  (.L_LO(net32));
 sg13g2_tielo \proj_14.flop32/_4__33  (.L_LO(net33));
 sg13g2_tielo \proj_14.flop33/_4__34  (.L_LO(net34));
 sg13g2_tielo \proj_14.flop34/_4__35  (.L_LO(net35));
 sg13g2_tielo \proj_14.flop35/_5__36  (.L_LO(net36));
 sg13g2_tielo \proj_14.flop36/_4__37  (.L_LO(net37));
 sg13g2_tielo \proj_14.flop37/_5__38  (.L_LO(net38));
 sg13g2_tielo \proj_14.flop4/_5__39  (.L_LO(net39));
 sg13g2_tielo \proj_14.flop5/_4__40  (.L_LO(net40));
 sg13g2_tielo \proj_14.flop6/_5__41  (.L_LO(net41));
 sg13g2_tielo \proj_14.flop7/_4__42  (.L_LO(net42));
 sg13g2_tielo \proj_14.flop8/_4__43  (.L_LO(net43));
 sg13g2_tielo \proj_14.flop9/_5__44  (.L_LO(net44));
 sg13g2_tielo \proj__9.flop1/_4__45  (.L_LO(net45));
 sg13g2_tielo tt_um_wokwi_group_3_46 (.L_LO(net46));
 sg13g2_tielo tt_um_wokwi_group_3_47 (.L_LO(net47));
 sg13g2_tielo tt_um_wokwi_group_3_48 (.L_LO(net48));
 sg13g2_tielo tt_um_wokwi_group_3_49 (.L_LO(net49));
 sg13g2_tielo tt_um_wokwi_group_3_50 (.L_LO(net50));
 sg13g2_tielo tt_um_wokwi_group_3_51 (.L_LO(net51));
 sg13g2_tielo tt_um_wokwi_group_3_52 (.L_LO(net52));
 sg13g2_tielo tt_um_wokwi_group_3_53 (.L_LO(net53));
 sg13g2_tielo tt_um_wokwi_group_3_54 (.L_LO(net54));
 sg13g2_tielo tt_um_wokwi_group_3_55 (.L_LO(net55));
 sg13g2_tielo tt_um_wokwi_group_3_56 (.L_LO(net56));
 sg13g2_tielo tt_um_wokwi_group_3_57 (.L_LO(net57));
 sg13g2_tielo tt_um_wokwi_group_3_58 (.L_LO(net58));
 sg13g2_tielo tt_um_wokwi_group_3_59 (.L_LO(net59));
 sg13g2_tielo tt_um_wokwi_group_3_60 (.L_LO(net60));
 sg13g2_tielo tt_um_wokwi_group_3_61 (.L_LO(net61));
 sg13g2_tielo \proj_14.flop1/dffsr_62  (.L_LO(net62));
 sg13g2_mux2_1 \proj_10.mux2/_0_  (.A0(net84),
    .A1(net81),
    .S(net80),
    .X(\proj_10.net9 ));
 sg13g2_nand2_1 \proj_10.nand1/_0_  (.Y(\proj_10.net10 ),
    .A(\proj_10.nand1/b ),
    .B(net77));
 sg13g2_inv_1 \proj_10.not1/_0_  (.Y(\proj_10.net12 ),
    .A(net4));
 sg13g2_inv_1 \proj_10.not2/_0_  (.Y(\proj_10.net13 ),
    .A(net5));
 sg13g2_xor2_1 \proj_10.xor1/_0_  (.B(net2),
    .A(net76),
    .X(\proj_10.net11 ));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net81),
    .B(net84),
    .X(\proj_12.net18 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(net77),
    .B(net79),
    .X(\proj_12.net20 ));
 sg13g2_and2_1 \proj_12.and4/_0_  (.A(\proj_12.net19 ),
    .B(\proj_12.net18 ),
    .X(\proj_12.net21 ));
 sg13g2_and2_1 \proj_12.and5/_0_  (.A(net76),
    .B(net2),
    .X(\proj_12.net24 ));
 sg13g2_and2_1 \proj_12.and6/_0_  (.A(\proj_12.net23 ),
    .B(\proj_12.net22 ),
    .X(\proj_12.net25 ));
 sg13g2_and2_1 \proj_12.and7/_0_  (.A(net5),
    .B(net4),
    .X(\proj_12.net28 ));
 sg13g2_and2_1 \proj_12.and8/_0_  (.A(\proj_12.net27 ),
    .B(\proj_12.net26 ),
    .X(\proj_12.net29 ));
 sg13g2_or2_1 \proj_12.or1/_0_  (.X(\proj_12.net22 ),
    .B(\proj_12.net21 ),
    .A(\proj_12.net20 ));
 sg13g2_or2_1 \proj_12.or2/_0_  (.X(\proj_12.net26 ),
    .B(\proj_12.net25 ),
    .A(\proj_12.net24 ));
 sg13g2_or2_1 \proj_12.or3/_0_  (.X(\proj_12.net13 ),
    .B(\proj_12.net29 ),
    .A(\proj_12.net28 ));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net85),
    .A(net81),
    .X(\proj_12.net9 ));
 sg13g2_xor2_1 \proj_12.xor2/_0_  (.B(net80),
    .A(net77),
    .X(\proj_12.net19 ));
 sg13g2_xor2_1 \proj_12.xor3/_0_  (.B(\proj_12.net19 ),
    .A(\proj_12.net18 ),
    .X(\proj_12.net10 ));
 sg13g2_xor2_1 \proj_12.xor4/_0_  (.B(net2),
    .A(net76),
    .X(\proj_12.net23 ));
 sg13g2_xor2_1 \proj_12.xor5/_0_  (.B(\proj_12.net23 ),
    .A(\proj_12.net22 ),
    .X(\proj_12.net11 ));
 sg13g2_xor2_1 \proj_12.xor6/_0_  (.B(net4),
    .A(net5),
    .X(\proj_12.net27 ));
 sg13g2_xor2_1 \proj_12.xor7/_0_  (.B(\proj_12.net27 ),
    .A(\proj_12.net26 ),
    .X(\proj_12.net12 ));
 sg13g2_dfrbp_1 \proj_13.flop1/_1_  (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net174),
    .D(net86),
    .Q_N(\proj_13.flop1/notq ),
    .Q(\proj_13.net12 ));
 sg13g2_tiehi \proj_13.flop2/_1__154  (.L_HI(net175));
 sg13g2_dfrbp_1 \proj_13.flop2/_1_  (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net175),
    .D(net193),
    .Q_N(\proj_13.flop2/notq ),
    .Q(\proj_13.net13 ));
 sg13g2_tiehi \proj_13.flop3/_1__155  (.L_HI(net176));
 sg13g2_dfrbp_1 \proj_13.flop3/_1_  (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net176),
    .D(net194),
    .Q_N(\proj_13.flop3/notq ),
    .Q(\proj_13.net8 ));
 sg13g2_tiehi \proj_14.flop28/_1__156  (.L_HI(net177));
 sg13g2_inv_1 \proj_13.not5/_0_  (.Y(\proj_13.net7 ),
    .A(\proj_13.net13 ));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(\proj_14.net30 ),
    .B(\proj_14.net33 ),
    .X(\proj_14.net58 ));
 sg13g2_and2_1 \proj_14.and10/_0_  (.A(\proj_14.net32 ),
    .B(\proj_14.net30 ),
    .X(\proj_14.net64 ));
 sg13g2_and2_1 \proj_14.and11/_0_  (.A(\proj_14.net40 ),
    .B(\proj_14.net43 ),
    .X(\proj_14.net68 ));
 sg13g2_and2_1 \proj_14.and12/_0_  (.A(\proj_14.net68 ),
    .B(\proj_14.net37 ),
    .X(\proj_14.net69 ));
 sg13g2_and2_1 \proj_14.and13/_0_  (.A(\proj_14.net68 ),
    .B(\proj_14.net36 ),
    .X(\proj_14.net70 ));
 sg13g2_and2_1 \proj_14.and14/_0_  (.A(\proj_14.net39 ),
    .B(\proj_14.net43 ),
    .X(\proj_14.net71 ));
 sg13g2_and2_1 \proj_14.and15/_0_  (.A(\proj_14.net71 ),
    .B(\proj_14.net37 ),
    .X(\proj_14.net72 ));
 sg13g2_and2_1 \proj_14.and16/_0_  (.A(\proj_14.net71 ),
    .B(\proj_14.net36 ),
    .X(\proj_14.net73 ));
 sg13g2_and2_1 \proj_14.and17/_0_  (.A(\proj_14.net74 ),
    .B(\proj_14.net37 ),
    .X(\proj_14.net75 ));
 sg13g2_and2_1 \proj_14.and18/_0_  (.A(\proj_14.net74 ),
    .B(\proj_14.net36 ),
    .X(\proj_14.net76 ));
 sg13g2_and2_1 \proj_14.and19/_0_  (.A(\proj_14.net42 ),
    .B(\proj_14.net39 ),
    .X(\proj_14.net77 ));
 sg13g2_and2_1 \proj_14.and2/_0_  (.A(\proj_14.net58 ),
    .B(net249),
    .X(\proj_14.net59 ));
 sg13g2_and2_1 \proj_14.and20/_0_  (.A(\proj_14.net42 ),
    .B(\proj_14.net40 ),
    .X(\proj_14.net74 ));
 sg13g2_and2_1 \proj_14.and21/_0_  (.A(\proj_14.net54 ),
    .B(\proj_14.net57 ),
    .X(\proj_14.net78 ));
 sg13g2_and2_1 \proj_14.and22/_0_  (.A(\proj_14.net78 ),
    .B(\proj_14.net51 ),
    .X(\proj_14.net79 ));
 sg13g2_and2_1 \proj_14.and23/_0_  (.A(\proj_14.net78 ),
    .B(\proj_14.net50 ),
    .X(\proj_14.net80 ));
 sg13g2_and2_1 \proj_14.and24/_0_  (.A(\proj_14.net53 ),
    .B(\proj_14.net57 ),
    .X(\proj_14.net81 ));
 sg13g2_and2_1 \proj_14.and25/_0_  (.A(\proj_14.net81 ),
    .B(\proj_14.net51 ),
    .X(\proj_14.net82 ));
 sg13g2_and2_1 \proj_14.and26/_0_  (.A(\proj_14.net81 ),
    .B(\proj_14.net50 ),
    .X(\proj_14.net83 ));
 sg13g2_and2_1 \proj_14.and27/_0_  (.A(\proj_14.net84 ),
    .B(\proj_14.net51 ),
    .X(\proj_14.net85 ));
 sg13g2_and2_1 \proj_14.and28/_0_  (.A(\proj_14.net84 ),
    .B(\proj_14.net50 ),
    .X(\proj_14.net86 ));
 sg13g2_and2_1 \proj_14.and29/_0_  (.A(\proj_14.net56 ),
    .B(\proj_14.net53 ),
    .X(\proj_14.net87 ));
 sg13g2_and2_1 \proj_14.and3/_0_  (.A(\proj_14.net58 ),
    .B(net251),
    .X(\proj_14.net60 ));
 sg13g2_and2_1 \proj_14.and30/_0_  (.A(\proj_14.net56 ),
    .B(\proj_14.net54 ),
    .X(\proj_14.net84 ));
 sg13g2_and2_1 \proj_14.and31/_0_  (.A(\proj_14.net105 ),
    .B(\proj_14.net110 ),
    .X(\proj_14.net116 ));
 sg13g2_and2_1 \proj_14.and32/_0_  (.A(\proj_14.net116 ),
    .B(\proj_14.net114 ),
    .X(\proj_14.net121 ));
 sg13g2_and2_1 \proj_14.and33/_0_  (.A(\proj_14.net121 ),
    .B(\proj_14.net119 ),
    .X(\proj_14.net126 ));
 sg13g2_and2_1 \proj_14.and34/_0_  (.A(\proj_14.net126 ),
    .B(\proj_14.net124 ),
    .X(\proj_14.net131 ));
 sg13g2_and2_1 \proj_14.and35/_0_  (.A(\proj_14.net137 ),
    .B(\proj_14.net135 ),
    .X(\proj_14.net142 ));
 sg13g2_and2_1 \proj_14.and36/_0_  (.A(\proj_14.net142 ),
    .B(\proj_14.net140 ),
    .X(\proj_14.net147 ));
 sg13g2_and2_1 \proj_14.and37/_0_  (.A(\proj_14.net147 ),
    .B(\proj_14.net145 ),
    .X(\proj_14.net152 ));
 sg13g2_and2_1 \proj_14.and38/_0_  (.A(\proj_14.net152 ),
    .B(\proj_14.net150 ),
    .X(\proj_14.net157 ));
 sg13g2_and2_1 \proj_14.and39/_0_  (.A(\proj_14.net131 ),
    .B(\proj_14.net129 ),
    .X(\proj_14.net137 ));
 sg13g2_and2_1 \proj_14.and4/_0_  (.A(\proj_14.net29 ),
    .B(\proj_14.net33 ),
    .X(\proj_14.net61 ));
 sg13g2_and2_1 \proj_14.and40/_0_  (.A(\proj_14.net157 ),
    .B(\proj_14.net155 ),
    .X(\proj_14.net162 ));
 sg13g2_and2_1 \proj_14.and41/_0_  (.A(\proj_14.net162 ),
    .B(\proj_14.net160 ),
    .X(\proj_14.net167 ));
 sg13g2_and2_1 \proj_14.and42/_0_  (.A(\proj_14.net167 ),
    .B(\proj_14.net165 ),
    .X(\proj_14.net172 ));
 sg13g2_and2_1 \proj_14.and43/_0_  (.A(\proj_14.net172 ),
    .B(\proj_14.net170 ),
    .X(\proj_14.net177 ));
 sg13g2_and2_1 \proj_14.and44/_0_  (.A(\proj_14.net193 ),
    .B(\proj_14.net192 ),
    .X(\proj_14.net194 ));
 sg13g2_and2_1 \proj_14.and45/_0_  (.A(\proj_14.net196 ),
    .B(\proj_14.net195 ),
    .X(\proj_14.net197 ));
 sg13g2_and2_1 \proj_14.and46/_0_  (.A(\proj_14.net199 ),
    .B(\proj_14.net198 ),
    .X(\proj_14.net200 ));
 sg13g2_and2_1 \proj_14.and47/_0_  (.A(\proj_14.net202 ),
    .B(\proj_14.net201 ),
    .X(\proj_14.net203 ));
 sg13g2_and2_1 \proj_14.and48/_0_  (.A(\proj_14.net203 ),
    .B(\proj_14.net200 ),
    .X(\proj_14.net204 ));
 sg13g2_and2_1 \proj_14.and49/_0_  (.A(\proj_14.net197 ),
    .B(\proj_14.net205 ),
    .X(\proj_14.net206 ));
 sg13g2_and2_1 \proj_14.and5/_0_  (.A(\proj_14.net61 ),
    .B(net247),
    .X(\proj_14.net62 ));
 sg13g2_and2_1 \proj_14.and50/_0_  (.A(\proj_14.net204 ),
    .B(\proj_14.net206 ),
    .X(\proj_14.net178 ));
 sg13g2_and2_1 \proj_14.and51/_0_  (.A(\proj_14.net59 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net234 ));
 sg13g2_and2_1 \proj_14.and52/_0_  (.A(\proj_14.net60 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net235 ));
 sg13g2_and2_1 \proj_14.and53/_0_  (.A(\proj_14.net62 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net236 ));
 sg13g2_and2_1 \proj_14.and54/_0_  (.A(\proj_14.net63 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net237 ));
 sg13g2_and2_1 \proj_14.and55/_0_  (.A(\proj_14.net65 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net238 ));
 sg13g2_and2_1 \proj_14.and57/_0_  (.A(\proj_14.net67 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net239 ));
 sg13g2_and2_1 \proj_14.and58/_0_  (.A(\proj_14.net59 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net240 ));
 sg13g2_and2_1 \proj_14.and59/_0_  (.A(\proj_14.net60 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net241 ));
 sg13g2_and2_1 \proj_14.and6/_0_  (.A(\proj_14.net61 ),
    .B(net250),
    .X(\proj_14.net63 ));
 sg13g2_and2_1 \proj_14.and60/_0_  (.A(\proj_14.net62 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net242 ));
 sg13g2_and2_1 \proj_14.and61/_0_  (.A(\proj_14.net63 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net243 ));
 sg13g2_and2_1 \proj_14.and62/_0_  (.A(\proj_14.net65 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net244 ));
 sg13g2_and2_1 \proj_14.and63/_0_  (.A(\proj_14.net66 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net245 ));
 sg13g2_and2_1 \proj_14.and64/_0_  (.A(net196),
    .B(\proj_14.net181 ),
    .X(\proj_14.net183 ));
 sg13g2_and2_1 \proj_14.and65/_0_  (.A(\proj_14.net67 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net246 ));
 sg13g2_and2_1 \proj_14.and66/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net235 ),
    .X(\proj_14.net249 ));
 sg13g2_and2_1 \proj_14.and67/_0_  (.A(\proj_14.net235 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net248 ));
 sg13g2_and2_1 \proj_14.and68/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net238 ),
    .X(\proj_14.net252 ));
 sg13g2_and2_1 \proj_14.and69/_0_  (.A(\proj_14.net238 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net254 ));
 sg13g2_and2_1 \proj_14.and7/_0_  (.A(\proj_14.net64 ),
    .B(net249),
    .X(\proj_14.net65 ));
 sg13g2_and2_1 \proj_14.and70/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net239 ),
    .X(\proj_14.net258 ));
 sg13g2_and2_1 \proj_14.and71/_0_  (.A(\proj_14.net239 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net256 ));
 sg13g2_and2_1 \proj_14.and72/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net242 ),
    .X(\proj_14.net265 ));
 sg13g2_and2_1 \proj_14.and73/_0_  (.A(\proj_14.net242 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net261 ));
 sg13g2_and2_1 \proj_14.and74/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net245 ),
    .X(\proj_14.net267 ));
 sg13g2_and2_1 \proj_14.and75/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net246 ),
    .X(\proj_14.net259 ));
 sg13g2_and2_1 \proj_14.and76/_0_  (.A(\proj_14.net246 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net269 ));
 sg13g2_and2_1 \proj_14.and77/_0_  (.A(\proj_14.net194 ),
    .B(\proj_14.net135 ),
    .X(\proj_14.net205 ));
 sg13g2_and2_1 \proj_14.and8/_0_  (.A(\proj_14.net64 ),
    .B(net248),
    .X(\proj_14.net66 ));
 sg13g2_and2_1 \proj_14.and9/_0_  (.A(net243),
    .B(net240),
    .X(\proj_14.net67 ));
 sg13g2_inv_1 \proj_14.flop1/_4_  (.Y(\proj_14.flop1/_1_ ),
    .A(net10));
 sg13g2_inv_1 \proj_14.flop1/_5_  (.Y(\proj_14.flop1/_0_ ),
    .A(net70));
 sg13g2_tielo \proj_14.flop1/dffsr_63  (.L_LO(net63));
 sg13g2_tielo \proj_14.flop10/dffsr_64  (.L_LO(net64));
 sg13g2_sdfbbp_1 \proj_14.flop1/dffsr  (.Q(\proj_14.net26 ),
    .Q_N(\proj_14.net27 ),
    .RESET_B(\proj_14.flop1/_0_ ),
    .SET_B(\proj_14.flop1/_1_ ),
    .D(\proj_14.net23 ),
    .SCE(net63),
    .SCD(net62),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop10/_4_  (.Y(\proj_14.flop10/_1_ ),
    .A(net11));
 sg13g2_inv_1 \proj_14.flop10/_5_  (.Y(\proj_14.flop10/_0_ ),
    .A(net68));
 sg13g2_tielo \proj_14.flop10/dffsr_65  (.L_LO(net65));
 sg13g2_tielo \proj_14.flop11/dffsr_66  (.L_LO(net66));
 sg13g2_sdfbbp_1 \proj_14.flop10/dffsr  (.Q(\proj_14.net105 ),
    .Q_N(\proj_14.net106 ),
    .RESET_B(\proj_14.flop10/_0_ ),
    .SET_B(\proj_14.flop10/_1_ ),
    .D(\proj_14.net102 ),
    .SCE(net65),
    .SCD(net64),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop11/_4_  (.Y(\proj_14.flop11/_1_ ),
    .A(net12));
 sg13g2_inv_1 \proj_14.flop11/_5_  (.Y(\proj_14.flop11/_0_ ),
    .A(net68));
 sg13g2_tielo \proj_14.flop11/dffsr_67  (.L_LO(net88));
 sg13g2_tielo \proj_14.flop12/dffsr_68  (.L_LO(net89));
 sg13g2_sdfbbp_1 \proj_14.flop11/dffsr  (.Q(\proj_14.net110 ),
    .Q_N(\proj_14.net111 ),
    .RESET_B(\proj_14.flop11/_0_ ),
    .SET_B(\proj_14.flop11/_1_ ),
    .D(net208),
    .SCE(net88),
    .SCD(net66),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop12/_4_  (.Y(\proj_14.flop12/_1_ ),
    .A(net13));
 sg13g2_inv_1 \proj_14.flop12/_5_  (.Y(\proj_14.flop12/_0_ ),
    .A(net67));
 sg13g2_tielo \proj_14.flop12/dffsr_69  (.L_LO(net90));
 sg13g2_tielo \proj_14.flop13/dffsr_70  (.L_LO(net91));
 sg13g2_sdfbbp_1 \proj_14.flop12/dffsr  (.Q(\proj_14.net114 ),
    .Q_N(\proj_14.net115 ),
    .RESET_B(\proj_14.flop12/_0_ ),
    .SET_B(\proj_14.flop12/_1_ ),
    .D(net206),
    .SCE(net90),
    .SCD(net89),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop13/_4_  (.Y(\proj_14.flop13/_1_ ),
    .A(net14));
 sg13g2_inv_1 \proj_14.flop13/_5_  (.Y(\proj_14.flop13/_0_ ),
    .A(net67));
 sg13g2_tielo \proj_14.flop13/dffsr_71  (.L_LO(net92));
 sg13g2_tielo \proj_14.flop14/dffsr_72  (.L_LO(net93));
 sg13g2_sdfbbp_1 \proj_14.flop13/dffsr  (.Q(\proj_14.net119 ),
    .Q_N(\proj_14.net120 ),
    .RESET_B(\proj_14.flop13/_0_ ),
    .SET_B(\proj_14.flop13/_1_ ),
    .D(net211),
    .SCE(net92),
    .SCD(net91),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop14/_4_  (.Y(\proj_14.flop14/_1_ ),
    .A(net15));
 sg13g2_inv_1 \proj_14.flop14/_5_  (.Y(\proj_14.flop14/_0_ ),
    .A(net67));
 sg13g2_tielo \proj_14.flop14/dffsr_73  (.L_LO(net94));
 sg13g2_tielo \proj_14.flop15/dffsr_74  (.L_LO(net95));
 sg13g2_sdfbbp_1 \proj_14.flop14/dffsr  (.Q(\proj_14.net124 ),
    .Q_N(\proj_14.net125 ),
    .RESET_B(\proj_14.flop14/_0_ ),
    .SET_B(\proj_14.flop14/_1_ ),
    .D(net202),
    .SCE(net94),
    .SCD(net93),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop15/_4_  (.Y(\proj_14.flop15/_1_ ),
    .A(net16));
 sg13g2_inv_1 \proj_14.flop15/_5_  (.Y(\proj_14.flop15/_0_ ),
    .A(net67));
 sg13g2_tielo \proj_14.flop15/dffsr_75  (.L_LO(net96));
 sg13g2_tielo \proj_14.flop16/dffsr_76  (.L_LO(net97));
 sg13g2_sdfbbp_1 \proj_14.flop15/dffsr  (.Q(\proj_14.net129 ),
    .Q_N(\proj_14.net130 ),
    .RESET_B(\proj_14.flop15/_0_ ),
    .SET_B(\proj_14.flop15/_1_ ),
    .D(net213),
    .SCE(net96),
    .SCD(net95),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop16/_4_  (.Y(\proj_14.flop16/_1_ ),
    .A(net17));
 sg13g2_inv_1 \proj_14.flop16/_5_  (.Y(\proj_14.flop16/_0_ ),
    .A(net68));
 sg13g2_tielo \proj_14.flop16/dffsr_77  (.L_LO(net98));
 sg13g2_tielo \proj_14.flop17/dffsr_78  (.L_LO(net99));
 sg13g2_sdfbbp_1 \proj_14.flop16/dffsr  (.Q(\proj_14.net135 ),
    .Q_N(\proj_14.net136 ),
    .RESET_B(\proj_14.flop16/_0_ ),
    .SET_B(\proj_14.flop16/_1_ ),
    .D(net221),
    .SCE(net98),
    .SCD(net97),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop17/_4_  (.Y(\proj_14.flop17/_1_ ),
    .A(net18));
 sg13g2_inv_1 \proj_14.flop17/_5_  (.Y(\proj_14.flop17/_0_ ),
    .A(net68));
 sg13g2_tielo \proj_14.flop17/dffsr_79  (.L_LO(net100));
 sg13g2_tielo \proj_14.flop18/dffsr_80  (.L_LO(net101));
 sg13g2_sdfbbp_1 \proj_14.flop17/dffsr  (.Q(\proj_14.net140 ),
    .Q_N(\proj_14.net141 ),
    .RESET_B(\proj_14.flop17/_0_ ),
    .SET_B(\proj_14.flop17/_1_ ),
    .D(net227),
    .SCE(net100),
    .SCD(net99),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop18/_4_  (.Y(\proj_14.flop18/_1_ ),
    .A(net19));
 sg13g2_inv_1 \proj_14.flop18/_5_  (.Y(\proj_14.flop18/_0_ ),
    .A(net67));
 sg13g2_tielo \proj_14.flop18/dffsr_81  (.L_LO(net102));
 sg13g2_tielo \proj_14.flop19/dffsr_82  (.L_LO(net103));
 sg13g2_sdfbbp_1 \proj_14.flop18/dffsr  (.Q(\proj_14.net145 ),
    .Q_N(\proj_14.net146 ),
    .RESET_B(\proj_14.flop18/_0_ ),
    .SET_B(\proj_14.flop18/_1_ ),
    .D(net225),
    .SCE(net102),
    .SCD(net101),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop19/_4_  (.Y(\proj_14.flop19/_1_ ),
    .A(net20));
 sg13g2_inv_1 \proj_14.flop19/_5_  (.Y(\proj_14.flop19/_0_ ),
    .A(net67));
 sg13g2_tielo \proj_14.flop19/dffsr_83  (.L_LO(net104));
 sg13g2_tielo \proj_14.flop2/dffsr_84  (.L_LO(net105));
 sg13g2_sdfbbp_1 \proj_14.flop19/dffsr  (.Q(\proj_14.net150 ),
    .Q_N(\proj_14.net151 ),
    .RESET_B(\proj_14.flop19/_0_ ),
    .SET_B(\proj_14.flop19/_1_ ),
    .D(net229),
    .SCE(net104),
    .SCD(net103),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop2/_4_  (.Y(\proj_14.flop2/_1_ ),
    .A(net21));
 sg13g2_inv_1 \proj_14.flop2/_5_  (.Y(\proj_14.flop2/_0_ ),
    .A(net70));
 sg13g2_tielo \proj_14.flop2/dffsr_85  (.L_LO(net106));
 sg13g2_tielo \proj_14.flop20/dffsr_86  (.L_LO(net107));
 sg13g2_sdfbbp_1 \proj_14.flop2/dffsr  (.Q(\proj_14.net29 ),
    .Q_N(\proj_14.net30 ),
    .RESET_B(\proj_14.flop2/_0_ ),
    .SET_B(\proj_14.flop2/_1_ ),
    .D(\proj_14.net28 ),
    .SCE(net106),
    .SCD(net105),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop20/_4_  (.Y(\proj_14.flop20/_1_ ),
    .A(net22));
 sg13g2_inv_1 \proj_14.flop20/_5_  (.Y(\proj_14.flop20/_0_ ),
    .A(net67));
 sg13g2_tielo \proj_14.flop20/dffsr_87  (.L_LO(net108));
 sg13g2_tielo \proj_14.flop21/dffsr_88  (.L_LO(net109));
 sg13g2_sdfbbp_1 \proj_14.flop20/dffsr  (.Q(\proj_14.net155 ),
    .Q_N(\proj_14.net156 ),
    .RESET_B(\proj_14.flop20/_0_ ),
    .SET_B(\proj_14.flop20/_1_ ),
    .D(net217),
    .SCE(net108),
    .SCD(net107),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop21/_4_  (.Y(\proj_14.flop21/_1_ ),
    .A(net23));
 sg13g2_inv_1 \proj_14.flop21/_5_  (.Y(\proj_14.flop21/_0_ ),
    .A(net67));
 sg13g2_tielo \proj_14.flop21/dffsr_89  (.L_LO(net110));
 sg13g2_tielo \proj_14.flop22/dffsr_90  (.L_LO(net111));
 sg13g2_sdfbbp_1 \proj_14.flop21/dffsr  (.Q(\proj_14.net160 ),
    .Q_N(\proj_14.net161 ),
    .RESET_B(\proj_14.flop21/_0_ ),
    .SET_B(\proj_14.flop21/_1_ ),
    .D(net204),
    .SCE(net110),
    .SCD(net109),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop22/_4_  (.Y(\proj_14.flop22/_1_ ),
    .A(net24));
 sg13g2_inv_1 \proj_14.flop22/_5_  (.Y(\proj_14.flop22/_0_ ),
    .A(net68));
 sg13g2_tielo \proj_14.flop22/dffsr_91  (.L_LO(net112));
 sg13g2_tielo \proj_14.flop23/dffsr_92  (.L_LO(net113));
 sg13g2_sdfbbp_1 \proj_14.flop22/dffsr  (.Q(\proj_14.net165 ),
    .Q_N(\proj_14.net166 ),
    .RESET_B(\proj_14.flop22/_0_ ),
    .SET_B(\proj_14.flop22/_1_ ),
    .D(net215),
    .SCE(net112),
    .SCD(net111),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop23/_4_  (.Y(\proj_14.flop23/_1_ ),
    .A(net25));
 sg13g2_inv_1 \proj_14.flop23/_5_  (.Y(\proj_14.flop23/_0_ ),
    .A(net68));
 sg13g2_tielo \proj_14.flop23/dffsr_93  (.L_LO(net114));
 sg13g2_tielo \proj_14.flop24/dffsr_94  (.L_LO(net115));
 sg13g2_sdfbbp_1 \proj_14.flop23/dffsr  (.Q(\proj_14.net170 ),
    .Q_N(\proj_14.net171 ),
    .RESET_B(\proj_14.flop23/_0_ ),
    .SET_B(\proj_14.flop23/_1_ ),
    .D(net223),
    .SCE(net114),
    .SCD(net113),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop24/_4_  (.Y(\proj_14.flop24/_1_ ),
    .A(net26));
 sg13g2_inv_1 \proj_14.flop24/_5_  (.Y(\proj_14.flop24/_0_ ),
    .A(net68));
 sg13g2_tielo \proj_14.flop24/dffsr_95  (.L_LO(net116));
 sg13g2_tielo \proj_14.flop25/dffsr_96  (.L_LO(net117));
 sg13g2_sdfbbp_1 \proj_14.flop24/dffsr  (.Q(\proj_14.net175 ),
    .Q_N(\proj_14.net176 ),
    .RESET_B(\proj_14.flop24/_0_ ),
    .SET_B(\proj_14.flop24/_1_ ),
    .D(net219),
    .SCE(net116),
    .SCD(net115),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop25/_4_  (.Y(\proj_14.flop25/_1_ ),
    .A(net27));
 sg13g2_inv_1 \proj_14.flop25/_5_  (.Y(\proj_14.flop25/_0_ ),
    .A(net71));
 sg13g2_tielo \proj_14.flop25/dffsr_97  (.L_LO(net118));
 sg13g2_tielo \proj_14.flop26/dffsr_98  (.L_LO(net119));
 sg13g2_sdfbbp_1 \proj_14.flop25/dffsr  (.Q(\proj_14.net180 ),
    .Q_N(\proj_14.flop25/notq ),
    .RESET_B(\proj_14.flop25/_0_ ),
    .SET_B(\proj_14.flop25/_1_ ),
    .D(\proj_14.net178 ),
    .SCE(net118),
    .SCD(net117),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop26/_4_  (.Y(\proj_14.flop26/_1_ ),
    .A(net28));
 sg13g2_inv_1 \proj_14.flop26/_5_  (.Y(\proj_14.flop26/_0_ ),
    .A(net71));
 sg13g2_tielo \proj_14.flop26/dffsr_99  (.L_LO(net120));
 sg13g2_tielo \proj_14.flop27/dffsr_100  (.L_LO(net121));
 sg13g2_sdfbbp_1 \proj_14.flop26/dffsr  (.Q(\proj_14.net181 ),
    .Q_N(\proj_14.flop26/notq ),
    .RESET_B(\proj_14.flop26/_0_ ),
    .SET_B(\proj_14.flop26/_1_ ),
    .D(net195),
    .SCE(net120),
    .SCD(net119),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop27/_4_  (.Y(\proj_14.flop27/_1_ ),
    .A(net29));
 sg13g2_inv_1 \proj_14.flop27/_5_  (.Y(\proj_14.flop27/_0_ ),
    .A(net71));
 sg13g2_tielo \proj_14.flop27/dffsr_101  (.L_LO(net122));
 sg13g2_tielo \proj_14.flop29/dffsr_102  (.L_LO(net123));
 sg13g2_sdfbbp_1 \proj_14.flop27/dffsr  (.Q(\proj_14.flop27/q ),
    .Q_N(\proj_14.net182 ),
    .RESET_B(\proj_14.flop27/_0_ ),
    .SET_B(\proj_14.flop27/_1_ ),
    .D(net198),
    .SCE(net122),
    .SCD(net121),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbp_1 \proj_14.flop28/_1_  (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net177),
    .D(\proj_14.net95 ),
    .Q_N(\proj_14.flop28/notq ),
    .Q(\proj_14.net11 ));
 sg13g2_tiehi \proj_14.flop46/_1__157  (.L_HI(net178));
 sg13g2_inv_1 \proj_14.flop29/_4_  (.Y(\proj_14.flop29/_1_ ),
    .A(net30));
 sg13g2_inv_1 \proj_14.flop29/_5_  (.Y(\proj_14.flop29/_0_ ),
    .A(net70));
 sg13g2_tielo \proj_14.flop29/dffsr_103  (.L_LO(net124));
 sg13g2_tielo \proj_14.flop3/dffsr_104  (.L_LO(net125));
 sg13g2_sdfbbp_1 \proj_14.flop29/dffsr  (.Q(\proj_14.net209 ),
    .Q_N(\proj_14.net210 ),
    .RESET_B(\proj_14.flop29/_0_ ),
    .SET_B(\proj_14.flop29/_1_ ),
    .D(net200),
    .SCE(net124),
    .SCD(net123),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop3/_4_  (.Y(\proj_14.flop3/_1_ ),
    .A(net31));
 sg13g2_inv_1 \proj_14.flop3/_5_  (.Y(\proj_14.flop3/_0_ ),
    .A(net70));
 sg13g2_tielo \proj_14.flop3/dffsr_105  (.L_LO(net126));
 sg13g2_tielo \proj_14.flop30/dffsr_106  (.L_LO(net127));
 sg13g2_sdfbbp_1 \proj_14.flop3/dffsr  (.Q(\proj_14.net32 ),
    .Q_N(\proj_14.net33 ),
    .RESET_B(\proj_14.flop3/_0_ ),
    .SET_B(\proj_14.flop3/_1_ ),
    .D(\proj_14.net31 ),
    .SCE(net126),
    .SCD(net125),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop30/_4_  (.Y(\proj_14.flop30/_1_ ),
    .A(net32));
 sg13g2_inv_1 \proj_14.flop30/_5_  (.Y(\proj_14.flop30/_0_ ),
    .A(net69));
 sg13g2_tielo \proj_14.flop30/dffsr_107  (.L_LO(net128));
 sg13g2_tielo \proj_14.flop31/dffsr_108  (.L_LO(net129));
 sg13g2_sdfbbp_1 \proj_14.flop30/dffsr  (.Q(\proj_14.net214 ),
    .Q_N(\proj_14.net215 ),
    .RESET_B(\proj_14.flop30/_0_ ),
    .SET_B(\proj_14.flop30/_1_ ),
    .D(\proj_14.net212 ),
    .SCE(net128),
    .SCD(net127),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop31/_4_  (.Y(\proj_14.flop31/_1_ ),
    .A(net69));
 sg13g2_inv_1 \proj_14.flop31/_5_  (.Y(\proj_14.flop31/_0_ ),
    .A(net69));
 sg13g2_tielo \proj_14.flop31/dffsr_109  (.L_LO(net130));
 sg13g2_tielo \proj_14.flop32/dffsr_110  (.L_LO(net131));
 sg13g2_sdfbbp_1 \proj_14.flop31/dffsr  (.Q(\proj_14.net217 ),
    .Q_N(\proj_14.flop31/notq ),
    .RESET_B(\proj_14.flop31/_0_ ),
    .SET_B(\proj_14.flop31/_1_ ),
    .D(\proj_14.net216 ),
    .SCE(net130),
    .SCD(net129),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop32/_4_  (.Y(\proj_14.flop32/_1_ ),
    .A(net33));
 sg13g2_inv_1 \proj_14.flop32/_5_  (.Y(\proj_14.flop32/_0_ ),
    .A(net69));
 sg13g2_tielo \proj_14.flop32/dffsr_111  (.L_LO(net132));
 sg13g2_tielo \proj_14.flop33/dffsr_112  (.L_LO(net133));
 sg13g2_sdfbbp_1 \proj_14.flop32/dffsr  (.Q(\proj_14.net219 ),
    .Q_N(\proj_14.flop32/notq ),
    .RESET_B(\proj_14.flop32/_0_ ),
    .SET_B(\proj_14.flop32/_1_ ),
    .D(\proj_14.net218 ),
    .SCE(net132),
    .SCD(net131),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop33/_4_  (.Y(\proj_14.flop33/_1_ ),
    .A(net34));
 sg13g2_inv_1 \proj_14.flop33/_5_  (.Y(\proj_14.flop33/_0_ ),
    .A(net69));
 sg13g2_tielo \proj_14.flop33/dffsr_113  (.L_LO(net134));
 sg13g2_tielo \proj_14.flop34/dffsr_114  (.L_LO(net135));
 sg13g2_sdfbbp_1 \proj_14.flop33/dffsr  (.Q(\proj_14.net221 ),
    .Q_N(\proj_14.flop33/notq ),
    .RESET_B(\proj_14.flop33/_0_ ),
    .SET_B(\proj_14.flop33/_1_ ),
    .D(\proj_14.net220 ),
    .SCE(net134),
    .SCD(net133),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop34/_4_  (.Y(\proj_14.flop34/_1_ ),
    .A(net35));
 sg13g2_inv_1 \proj_14.flop34/_5_  (.Y(\proj_14.flop34/_0_ ),
    .A(net69));
 sg13g2_tielo \proj_14.flop34/dffsr_115  (.L_LO(net136));
 sg13g2_tielo \proj_14.flop35/dffsr_116  (.L_LO(net137));
 sg13g2_sdfbbp_1 \proj_14.flop34/dffsr  (.Q(\proj_14.net223 ),
    .Q_N(\proj_14.flop34/notq ),
    .RESET_B(\proj_14.flop34/_0_ ),
    .SET_B(\proj_14.flop34/_1_ ),
    .D(\proj_14.net222 ),
    .SCE(net136),
    .SCD(net135),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop35/_4_  (.Y(\proj_14.flop35/_1_ ),
    .A(net69));
 sg13g2_inv_1 \proj_14.flop35/_5_  (.Y(\proj_14.flop35/_0_ ),
    .A(net36));
 sg13g2_tielo \proj_14.flop35/dffsr_117  (.L_LO(net138));
 sg13g2_tielo \proj_14.flop36/dffsr_118  (.L_LO(net139));
 sg13g2_sdfbbp_1 \proj_14.flop35/dffsr  (.Q(\proj_14.net226 ),
    .Q_N(\proj_14.flop35/notq ),
    .RESET_B(\proj_14.flop35/_0_ ),
    .SET_B(\proj_14.flop35/_1_ ),
    .D(\proj_14.net224 ),
    .SCE(net138),
    .SCD(net137),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop36/_4_  (.Y(\proj_14.flop36/_1_ ),
    .A(net37));
 sg13g2_inv_1 \proj_14.flop36/_5_  (.Y(\proj_14.flop36/_0_ ),
    .A(net70));
 sg13g2_tielo \proj_14.flop36/dffsr_119  (.L_LO(net140));
 sg13g2_tielo \proj_14.flop37/dffsr_120  (.L_LO(net141));
 sg13g2_sdfbbp_1 \proj_14.flop36/dffsr  (.Q(\proj_14.net228 ),
    .Q_N(\proj_14.flop36/notq ),
    .RESET_B(\proj_14.flop36/_0_ ),
    .SET_B(\proj_14.flop36/_1_ ),
    .D(net234),
    .SCE(net140),
    .SCD(net139),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop37/_4_  (.Y(\proj_14.flop37/_1_ ),
    .A(net71));
 sg13g2_inv_1 \proj_14.flop37/_5_  (.Y(\proj_14.flop37/_0_ ),
    .A(net38));
 sg13g2_tielo \proj_14.flop37/dffsr_121  (.L_LO(net142));
 sg13g2_tielo \proj_14.flop4/dffsr_122  (.L_LO(net143));
 sg13g2_sdfbbp_1 \proj_14.flop37/dffsr  (.Q(\proj_14.net231 ),
    .Q_N(\proj_14.flop37/notq ),
    .RESET_B(\proj_14.flop37/_0_ ),
    .SET_B(\proj_14.flop37/_1_ ),
    .D(\proj_14.net229 ),
    .SCE(net142),
    .SCD(net141),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop4/_4_  (.Y(\proj_14.flop4/_1_ ),
    .A(net70));
 sg13g2_inv_1 \proj_14.flop4/_5_  (.Y(\proj_14.flop4/_0_ ),
    .A(net39));
 sg13g2_tielo \proj_14.flop4/dffsr_123  (.L_LO(net144));
 sg13g2_tielo \proj_14.flop5/dffsr_124  (.L_LO(net145));
 sg13g2_sdfbbp_1 \proj_14.flop4/dffsr  (.Q(\proj_14.net36 ),
    .Q_N(\proj_14.net37 ),
    .RESET_B(\proj_14.flop4/_0_ ),
    .SET_B(\proj_14.flop4/_1_ ),
    .D(\proj_14.net34 ),
    .SCE(net144),
    .SCD(net143),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbp_1 \proj_14.flop46/_1_  (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net178),
    .D(\proj_14.net96 ),
    .Q_N(\proj_14.flop46/notq ),
    .Q(\proj_14.net12 ));
 sg13g2_tiehi \proj_14.flop47/_1__158  (.L_HI(net179));
 sg13g2_dfrbp_1 \proj_14.flop47/_1_  (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net179),
    .D(\proj_14.net97 ),
    .Q_N(\proj_14.flop47/notq ),
    .Q(\proj_14.net13 ));
 sg13g2_tiehi \proj_14.flop48/_1__159  (.L_HI(net180));
 sg13g2_dfrbp_1 \proj_14.flop48/_1_  (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net180),
    .D(\proj_14.net98 ),
    .Q_N(\proj_14.flop48/notq ),
    .Q(\proj_14.net14 ));
 sg13g2_tiehi \proj_14.flop49/_1__160  (.L_HI(net181));
 sg13g2_dfrbp_1 \proj_14.flop49/_1_  (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net181),
    .D(\proj_14.net99 ),
    .Q_N(\proj_14.flop49/notq ),
    .Q(\proj_14.net15 ));
 sg13g2_tiehi \proj_14.flop50/_1__161  (.L_HI(net182));
 sg13g2_inv_1 \proj_14.flop5/_4_  (.Y(\proj_14.flop5/_1_ ),
    .A(net40));
 sg13g2_inv_1 \proj_14.flop5/_5_  (.Y(\proj_14.flop5/_0_ ),
    .A(net70));
 sg13g2_tielo \proj_14.flop5/dffsr_125  (.L_LO(net146));
 sg13g2_tielo \proj_14.flop6/dffsr_126  (.L_LO(net147));
 sg13g2_sdfbbp_1 \proj_14.flop5/dffsr  (.Q(\proj_14.net39 ),
    .Q_N(\proj_14.net40 ),
    .RESET_B(\proj_14.flop5/_0_ ),
    .SET_B(\proj_14.flop5/_1_ ),
    .D(\proj_14.net38 ),
    .SCE(net146),
    .SCD(net145),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbp_1 \proj_14.flop50/_1_  (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net182),
    .D(\proj_14.net100 ),
    .Q_N(\proj_14.flop50/notq ),
    .Q(\proj_14.net16 ));
 sg13g2_tiehi \proj_14.flop51/_1__162  (.L_HI(net183));
 sg13g2_dfrbp_1 \proj_14.flop51/_1_  (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net183),
    .D(\proj_14.net101 ),
    .Q_N(\proj_14.flop51/notq ),
    .Q(\proj_14.net17 ));
 sg13g2_tiehi \proj_14.flop52/_1__163  (.L_HI(net184));
 sg13g2_dfrbp_1 \proj_14.flop52/_1_  (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net184),
    .D(net197),
    .Q_N(\proj_14.flop52/notq ),
    .Q(\proj_14.net45 ));
 sg13g2_tiehi \proj_14.flop53/_1__164  (.L_HI(net185));
 sg13g2_dfrbp_1 \proj_14.flop53/_1_  (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net185),
    .D(\proj_14.net275 ),
    .Q_N(\proj_14.flop53/notq ),
    .Q(\proj_14.net44 ));
 sg13g2_tiehi \proj_14.flop54/_1__165  (.L_HI(net186));
 sg13g2_dfrbp_1 \proj_14.flop54/_1_  (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net186),
    .D(\proj_14.net277 ),
    .Q_N(\proj_14.flop54/notq ),
    .Q(\proj_14.net46 ));
 sg13g2_tiehi \proj_14.flop55/_1__166  (.L_HI(net187));
 sg13g2_dfrbp_1 \proj_14.flop55/_1_  (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net187),
    .D(\proj_14.net280 ),
    .Q_N(\proj_14.flop55/notq ),
    .Q(\proj_14.net47 ));
 sg13g2_tiehi \proj_14.flop56/_1__167  (.L_HI(net188));
 sg13g2_dfrbp_1 \proj_14.flop56/_1_  (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net188),
    .D(\proj_14.net281 ),
    .Q_N(\proj_14.flop56/notq ),
    .Q(\proj_14.net211 ));
 sg13g2_tiehi \proj__7.flop1/_1__168  (.L_HI(net189));
 sg13g2_inv_1 \proj_14.flop6/_4_  (.Y(\proj_14.flop6/_1_ ),
    .A(net69));
 sg13g2_inv_1 \proj_14.flop6/_5_  (.Y(\proj_14.flop6/_0_ ),
    .A(net41));
 sg13g2_tielo \proj_14.flop6/dffsr_127  (.L_LO(net148));
 sg13g2_tielo \proj_14.flop7/dffsr_128  (.L_LO(net149));
 sg13g2_sdfbbp_1 \proj_14.flop6/dffsr  (.Q(\proj_14.net42 ),
    .Q_N(\proj_14.net43 ),
    .RESET_B(\proj_14.flop6/_0_ ),
    .SET_B(\proj_14.flop6/_1_ ),
    .D(\proj_14.net41 ),
    .SCE(net148),
    .SCD(net147),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop7/_4_  (.Y(\proj_14.flop7/_1_ ),
    .A(net42));
 sg13g2_inv_1 \proj_14.flop7/_5_  (.Y(\proj_14.flop7/_0_ ),
    .A(net71));
 sg13g2_tielo \proj_14.flop7/dffsr_129  (.L_LO(net150));
 sg13g2_tielo \proj_14.flop8/dffsr_130  (.L_LO(net151));
 sg13g2_sdfbbp_1 \proj_14.flop7/dffsr  (.Q(\proj_14.net50 ),
    .Q_N(\proj_14.net51 ),
    .RESET_B(\proj_14.flop7/_0_ ),
    .SET_B(\proj_14.flop7/_1_ ),
    .D(\proj_14.net48 ),
    .SCE(net150),
    .SCD(net149),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop8/_4_  (.Y(\proj_14.flop8/_1_ ),
    .A(net43));
 sg13g2_inv_1 \proj_14.flop8/_5_  (.Y(\proj_14.flop8/_0_ ),
    .A(net71));
 sg13g2_tielo \proj_14.flop8/dffsr_131  (.L_LO(net152));
 sg13g2_tielo \proj_14.flop9/dffsr_132  (.L_LO(net153));
 sg13g2_sdfbbp_1 \proj_14.flop8/dffsr  (.Q(\proj_14.net53 ),
    .Q_N(\proj_14.net54 ),
    .RESET_B(\proj_14.flop8/_0_ ),
    .SET_B(\proj_14.flop8/_1_ ),
    .D(\proj_14.net52 ),
    .SCE(net152),
    .SCD(net151),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_inv_1 \proj_14.flop9/_4_  (.Y(\proj_14.flop9/_1_ ),
    .A(net71));
 sg13g2_inv_1 \proj_14.flop9/_5_  (.Y(\proj_14.flop9/_0_ ),
    .A(net44));
 sg13g2_tielo \proj_14.flop9/dffsr_133  (.L_LO(net154));
 sg13g2_tielo \proj__4.flop1/dffsr_134  (.L_LO(net155));
 sg13g2_sdfbbp_1 \proj_14.flop9/dffsr  (.Q(\proj_14.net56 ),
    .Q_N(\proj_14.net57 ),
    .RESET_B(\proj_14.flop9/_0_ ),
    .SET_B(\proj_14.flop9/_1_ ),
    .D(\proj_14.net55 ),
    .SCE(net154),
    .SCD(net153),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_mux2_1 \proj_14.mux1/_0_  (.A0(\proj_14.net23 ),
    .A1(net231),
    .S(net74),
    .X(\proj_14.net23 ));
 sg13g2_mux2_1 \proj_14.mux10/_0_  (.A0(\proj_14.net105 ),
    .A1(net209),
    .S(net173),
    .X(\proj_14.net102 ));
 sg13g2_mux2_1 \proj_14.mux11/_0_  (.A0(\proj_14.net110 ),
    .A1(net207),
    .S(\proj_14.net105 ),
    .X(\proj_14.net108 ));
 sg13g2_mux2_1 \proj_14.mux12/_0_  (.A0(\proj_14.net114 ),
    .A1(net205),
    .S(\proj_14.net116 ),
    .X(\proj_14.net112 ));
 sg13g2_mux2_1 \proj_14.mux13/_0_  (.A0(\proj_14.net119 ),
    .A1(net210),
    .S(\proj_14.net121 ),
    .X(\proj_14.net117 ));
 sg13g2_mux2_1 \proj_14.mux14/_0_  (.A0(\proj_14.net124 ),
    .A1(net201),
    .S(\proj_14.net126 ),
    .X(\proj_14.net122 ));
 sg13g2_mux2_1 \proj_14.mux15/_0_  (.A0(\proj_14.net129 ),
    .A1(net212),
    .S(\proj_14.net131 ),
    .X(\proj_14.net127 ));
 sg13g2_mux2_1 \proj_14.mux16/_0_  (.A0(\proj_14.net135 ),
    .A1(net220),
    .S(\proj_14.net137 ),
    .X(\proj_14.net133 ));
 sg13g2_mux2_1 \proj_14.mux17/_0_  (.A0(\proj_14.net140 ),
    .A1(net226),
    .S(\proj_14.net142 ),
    .X(\proj_14.net138 ));
 sg13g2_mux2_1 \proj_14.mux18/_0_  (.A0(\proj_14.net145 ),
    .A1(net224),
    .S(\proj_14.net147 ),
    .X(\proj_14.net143 ));
 sg13g2_mux2_1 \proj_14.mux19/_0_  (.A0(\proj_14.net150 ),
    .A1(net228),
    .S(\proj_14.net152 ),
    .X(\proj_14.net148 ));
 sg13g2_mux2_1 \proj_14.mux2/_0_  (.A0(\proj_14.net28 ),
    .A1(net230),
    .S(net74),
    .X(\proj_14.net28 ));
 sg13g2_mux2_1 \proj_14.mux20/_0_  (.A0(\proj_14.net155 ),
    .A1(net216),
    .S(\proj_14.net157 ),
    .X(\proj_14.net153 ));
 sg13g2_mux2_1 \proj_14.mux21/_0_  (.A0(\proj_14.net160 ),
    .A1(net203),
    .S(\proj_14.net162 ),
    .X(\proj_14.net158 ));
 sg13g2_mux2_1 \proj_14.mux22/_0_  (.A0(\proj_14.net165 ),
    .A1(net214),
    .S(\proj_14.net167 ),
    .X(\proj_14.net163 ));
 sg13g2_mux2_1 \proj_14.mux23/_0_  (.A0(\proj_14.net170 ),
    .A1(net222),
    .S(\proj_14.net172 ),
    .X(\proj_14.net168 ));
 sg13g2_mux2_1 \proj_14.mux24/_0_  (.A0(\proj_14.net175 ),
    .A1(net218),
    .S(\proj_14.net177 ),
    .X(\proj_14.net173 ));
 sg13g2_mux2_1 \proj_14.mux25/_0_  (.A0(\proj_14.net209 ),
    .A1(net199),
    .S(net74),
    .X(\proj_14.net207 ));
 sg13g2_mux2_1 \proj_14.mux26/_0_  (.A0(\proj_14.net214 ),
    .A1(\proj_14.net233 ),
    .S(net72),
    .X(\proj_14.net212 ));
 sg13g2_mux2_1 \proj_14.mux27/_0_  (.A0(net235),
    .A1(\proj_14.net214 ),
    .S(net72),
    .X(\proj_14.net216 ));
 sg13g2_mux2_1 \proj_14.mux28/_0_  (.A0(net236),
    .A1(net235),
    .S(net72),
    .X(\proj_14.net218 ));
 sg13g2_mux2_1 \proj_14.mux29/_0_  (.A0(net238),
    .A1(net236),
    .S(net72),
    .X(\proj_14.net220 ));
 sg13g2_mux2_1 \proj_14.mux3/_0_  (.A0(\proj_14.net31 ),
    .A1(net232),
    .S(net74),
    .X(\proj_14.net31 ));
 sg13g2_mux2_1 \proj_14.mux30/_0_  (.A0(net241),
    .A1(net238),
    .S(net72),
    .X(\proj_14.net222 ));
 sg13g2_mux2_1 \proj_14.mux31/_0_  (.A0(net242),
    .A1(net241),
    .S(net73),
    .X(\proj_14.net224 ));
 sg13g2_mux2_1 \proj_14.mux32/_0_  (.A0(net233),
    .A1(\proj_14.net226 ),
    .S(net73),
    .X(\proj_14.net227 ));
 sg13g2_mux2_1 \proj_14.mux33/_0_  (.A0(net237),
    .A1(net233),
    .S(net72),
    .X(\proj_14.net229 ));
 sg13g2_mux2_1 \proj_14.mux4/_0_  (.A0(\proj_14.net34 ),
    .A1(net246),
    .S(net74),
    .X(\proj_14.net34 ));
 sg13g2_mux2_1 \proj_14.mux5/_0_  (.A0(\proj_14.net38 ),
    .A1(net240),
    .S(net72),
    .X(\proj_14.net38 ));
 sg13g2_mux2_1 \proj_14.mux6/_0_  (.A0(\proj_14.net41 ),
    .A1(net243),
    .S(net72),
    .X(\proj_14.net41 ));
 sg13g2_mux2_1 \proj_14.mux7/_0_  (.A0(\proj_14.net48 ),
    .A1(net245),
    .S(net74),
    .X(\proj_14.net48 ));
 sg13g2_mux2_1 \proj_14.mux8/_0_  (.A0(\proj_14.net52 ),
    .A1(net239),
    .S(net73),
    .X(\proj_14.net52 ));
 sg13g2_mux2_1 \proj_14.mux9/_0_  (.A0(\proj_14.net55 ),
    .A1(net244),
    .S(net73),
    .X(\proj_14.net55 ));
 sg13g2_inv_1 \proj_14.not1/_0_  (.Y(\proj_14.net132 ),
    .A(net87));
 sg13g2_inv_1 \proj_14.not10/_0_  (.Y(\proj_14.net193 ),
    .A(\proj_14.net190 ));
 sg13g2_inv_1 \proj_14.not2/_0_  (.Y(\proj_14.net202 ),
    .A(\proj_14.net184 ));
 sg13g2_inv_1 \proj_14.not3/_0_  (.Y(\proj_14.net201 ),
    .A(\proj_14.net185 ));
 sg13g2_inv_1 \proj_14.not4/_0_  (.Y(\proj_14.net198 ),
    .A(\proj_14.net187 ));
 sg13g2_inv_1 \proj_14.not5/_0_  (.Y(\proj_14.net25 ),
    .A(net87));
 sg13g2_inv_1 \proj_14.not6/_0_  (.Y(\proj_14.net199 ),
    .A(\proj_14.net186 ));
 sg13g2_inv_1 \proj_14.not7/_0_  (.Y(\proj_14.net195 ),
    .A(\proj_14.net189 ));
 sg13g2_inv_1 \proj_14.not8/_0_  (.Y(\proj_14.net196 ),
    .A(\proj_14.net188 ));
 sg13g2_inv_1 \proj_14.not9/_0_  (.Y(\proj_14.net192 ),
    .A(\proj_14.net191 ));
 sg13g2_or2_1 \proj_14.or1/_0_  (.X(\proj_14.net104 ),
    .B(\proj_14.net132 ),
    .A(\proj_14.net183 ));
 sg13g2_or2_1 \proj_14.or10/_0_  (.X(\proj_14.net96 ),
    .B(\proj_14.net60 ),
    .A(\proj_14.net89 ));
 sg13g2_or2_1 \proj_14.or11/_0_  (.X(\proj_14.net97 ),
    .B(\proj_14.net62 ),
    .A(\proj_14.net90 ));
 sg13g2_or2_1 \proj_14.or12/_0_  (.X(\proj_14.net98 ),
    .B(\proj_14.net63 ),
    .A(\proj_14.net91 ));
 sg13g2_or2_1 \proj_14.or13/_0_  (.X(\proj_14.net99 ),
    .B(\proj_14.net65 ),
    .A(\proj_14.net92 ));
 sg13g2_or2_1 \proj_14.or14/_0_  (.X(\proj_14.net100 ),
    .B(\proj_14.net66 ),
    .A(\proj_14.net93 ));
 sg13g2_or2_1 \proj_14.or15/_0_  (.X(\proj_14.net101 ),
    .B(\proj_14.net67 ),
    .A(\proj_14.net94 ));
 sg13g2_or2_1 \proj_14.or16/_0_  (.X(\proj_14.net247 ),
    .B(\proj_14.net236 ),
    .A(\proj_14.net234 ));
 sg13g2_or2_1 \proj_14.or17/_0_  (.X(\proj_14.net250 ),
    .B(\proj_14.net248 ),
    .A(\proj_14.net249 ));
 sg13g2_or2_1 \proj_14.or18/_0_  (.X(\proj_14.net255 ),
    .B(\proj_14.net254 ),
    .A(\proj_14.net252 ));
 sg13g2_or2_1 \proj_14.or19/_0_  (.X(\proj_14.net251 ),
    .B(\proj_14.net237 ),
    .A(\proj_14.net248 ));
 sg13g2_or2_1 \proj_14.or2/_0_  (.X(\proj_14.net95 ),
    .B(\proj_14.net59 ),
    .A(\proj_14.net88 ));
 sg13g2_or2_1 \proj_14.or20/_0_  (.X(\proj_14.net253 ),
    .B(\proj_14.net252 ),
    .A(\proj_14.net236 ));
 sg13g2_or2_1 \proj_14.or21/_0_  (.X(\proj_14.net257 ),
    .B(\proj_14.net254 ),
    .A(\proj_14.net256 ));
 sg13g2_or2_1 \proj_14.or22/_0_  (.X(\proj_14.net272 ),
    .B(\proj_14.net253 ),
    .A(\proj_14.net250 ));
 sg13g2_or2_1 \proj_14.or23/_0_  (.X(\proj_14.net287 ),
    .B(\proj_14.net285 ),
    .A(\proj_14.net286 ));
 sg13g2_or2_1 \proj_14.or24/_0_  (.X(\proj_14.net260 ),
    .B(\proj_14.net259 ),
    .A(\proj_14.net240 ));
 sg13g2_or2_1 \proj_14.or25/_0_  (.X(\proj_14.net262 ),
    .B(\proj_14.net261 ),
    .A(\proj_14.net240 ));
 sg13g2_or2_1 \proj_14.or26/_0_  (.X(\proj_14.net263 ),
    .B(\proj_14.net243 ),
    .A(\proj_14.net261 ));
 sg13g2_or2_1 \proj_14.or27/_0_  (.X(\proj_14.net264 ),
    .B(\proj_14.net251 ),
    .A(\proj_14.net245 ));
 sg13g2_or2_1 \proj_14.or28/_0_  (.X(\proj_14.net266 ),
    .B(\proj_14.net244 ),
    .A(\proj_14.net265 ));
 sg13g2_or2_1 \proj_14.or29/_0_  (.X(\proj_14.net268 ),
    .B(\proj_14.net244 ),
    .A(\proj_14.net267 ));
 sg13g2_or2_1 \proj_14.or3/_0_  (.X(\proj_14.net88 ),
    .B(\proj_14.net69 ),
    .A(\proj_14.net79 ));
 sg13g2_or2_1 \proj_14.or30/_0_  (.X(\proj_14.net273 ),
    .B(\proj_14.net266 ),
    .A(\proj_14.net260 ));
 sg13g2_or2_1 \proj_14.or31/_0_  (.X(\proj_14.net270 ),
    .B(\proj_14.net269 ),
    .A(\proj_14.net268 ));
 sg13g2_or2_1 \proj_14.or32/_0_  (.X(\proj_14.net271 ),
    .B(\proj_14.net256 ),
    .A(\proj_14.net258 ));
 sg13g2_or2_1 \proj_14.or33/_0_  (.X(\proj_14.net274 ),
    .B(\proj_14.net257 ),
    .A(\proj_14.net247 ));
 sg13g2_or2_1 \proj_14.or34/_0_  (.X(\proj_14.net275 ),
    .B(\proj_14.net273 ),
    .A(\proj_14.net274 ));
 sg13g2_or2_1 \proj_14.or35/_0_  (.X(\proj_14.net276 ),
    .B(\proj_14.net263 ),
    .A(\proj_14.net272 ));
 sg13g2_or2_1 \proj_14.or36/_0_  (.X(\proj_14.net277 ),
    .B(\proj_14.net270 ),
    .A(\proj_14.net276 ));
 sg13g2_or2_1 \proj_14.or37/_0_  (.X(\proj_14.net278 ),
    .B(\proj_14.net271 ),
    .A(\proj_14.net262 ));
 sg13g2_or2_1 \proj_14.or38/_0_  (.X(\proj_14.net279 ),
    .B(\proj_14.net255 ),
    .A(\proj_14.net264 ));
 sg13g2_or2_1 \proj_14.or39/_0_  (.X(\proj_14.net280 ),
    .B(\proj_14.net278 ),
    .A(\proj_14.net279 ));
 sg13g2_or2_1 \proj_14.or4/_0_  (.X(\proj_14.net89 ),
    .B(\proj_14.net70 ),
    .A(\proj_14.net80 ));
 sg13g2_or2_1 \proj_14.or40/_0_  (.X(\proj_14.net283 ),
    .B(\proj_14.net240 ),
    .A(\proj_14.net241 ));
 sg13g2_or2_1 \proj_14.or41/_0_  (.X(\proj_14.net284 ),
    .B(\proj_14.net243 ),
    .A(\proj_14.net244 ));
 sg13g2_or2_1 \proj_14.or42/_0_  (.X(\proj_14.net285 ),
    .B(\proj_14.net283 ),
    .A(\proj_14.net284 ));
 sg13g2_or2_1 \proj_14.or43/_0_  (.X(\proj_14.net286 ),
    .B(\proj_14.net259 ),
    .A(\proj_14.net258 ));
 sg13g2_or2_1 \proj_14.or44/_0_  (.X(\proj_14.net288 ),
    .B(\proj_14.net265 ),
    .A(\proj_14.net252 ));
 sg13g2_or2_1 \proj_14.or45/_0_  (.X(\proj_14.net281 ),
    .B(\proj_14.net287 ),
    .A(\proj_14.net289 ));
 sg13g2_or2_1 \proj_14.or46/_0_  (.X(\proj_14.net289 ),
    .B(\proj_14.net245 ),
    .A(\proj_14.net288 ));
 sg13g2_or2_1 \proj_14.or5/_0_  (.X(\proj_14.net90 ),
    .B(\proj_14.net72 ),
    .A(\proj_14.net82 ));
 sg13g2_or2_1 \proj_14.or6/_0_  (.X(\proj_14.net91 ),
    .B(\proj_14.net73 ),
    .A(\proj_14.net83 ));
 sg13g2_or2_1 \proj_14.or7/_0_  (.X(\proj_14.net92 ),
    .B(\proj_14.net75 ),
    .A(\proj_14.net85 ));
 sg13g2_or2_1 \proj_14.or8/_0_  (.X(\proj_14.net93 ),
    .B(\proj_14.net76 ),
    .A(\proj_14.net86 ));
 sg13g2_or2_1 \proj_14.or9/_0_  (.X(\proj_14.net94 ),
    .B(\proj_14.net77 ),
    .A(\proj_14.net87 ));
 sg13g2_xor2_1 \proj_14.xor1/_0_  (.B(net5),
    .A(\proj_14.net175 ),
    .X(\proj_14.net184 ));
 sg13g2_xor2_1 \proj_14.xor10/_0_  (.B(\proj_14.net226 ),
    .A(\proj_14.net231 ),
    .X(\proj_14.net282 ));
 sg13g2_xor2_1 \proj_14.xor11/_0_  (.B(net238),
    .A(\proj_14.net232 ),
    .X(\proj_14.net233 ));
 sg13g2_xor2_1 \proj_14.xor2/_0_  (.B(net4),
    .A(\proj_14.net170 ),
    .X(\proj_14.net185 ));
 sg13g2_xor2_1 \proj_14.xor3/_0_  (.B(net76),
    .A(\proj_14.net165 ),
    .X(\proj_14.net186 ));
 sg13g2_xor2_1 \proj_14.xor4/_0_  (.B(net2),
    .A(\proj_14.net160 ),
    .X(\proj_14.net187 ));
 sg13g2_xor2_1 \proj_14.xor5/_0_  (.B(net78),
    .A(\proj_14.net155 ),
    .X(\proj_14.net188 ));
 sg13g2_xor2_1 \proj_14.xor6/_0_  (.B(net79),
    .A(\proj_14.net150 ),
    .X(\proj_14.net189 ));
 sg13g2_xor2_1 \proj_14.xor7/_0_  (.B(net83),
    .A(\proj_14.net145 ),
    .X(\proj_14.net190 ));
 sg13g2_xor2_1 \proj_14.xor8/_0_  (.B(net86),
    .A(\proj_14.net140 ),
    .X(\proj_14.net191 ));
 sg13g2_xor2_1 \proj_14.xor9/_0_  (.B(\proj_14.net223 ),
    .A(\proj_14.net282 ),
    .X(\proj_14.net232 ));
 sg13g2_and2_1 \proj_15.and1/_0_  (.A(net80),
    .B(net84),
    .X(\proj_15.net15 ));
 sg13g2_and2_1 \proj_15.and2/_0_  (.A(\proj_15.net15 ),
    .B(net81),
    .X(\proj_15.net18 ));
 sg13g2_and2_1 \proj_15.and3/_0_  (.A(net78),
    .B(\proj_15.net7 ),
    .X(\proj_15.net17 ));
 sg13g2_or2_1 \proj_15.or1/_0_  (.X(\proj_15.net9 ),
    .B(\proj_15.net17 ),
    .A(\proj_15.net18 ));
 sg13g2_xor2_1 \proj_15.xor1/_0_  (.B(net84),
    .A(net80),
    .X(\proj_15.net7 ));
 sg13g2_xor2_1 \proj_15.xor2/_0_  (.B(\proj_15.net15 ),
    .A(net81),
    .X(\proj_15.net16 ));
 sg13g2_xor2_1 \proj_15.xor3/_0_  (.B(\proj_15.net16 ),
    .A(net78),
    .X(\proj_15.net8 ));
 sg13g2_inv_1 \proj__0.not3/_0_  (.Y(\proj__0.net10 ),
    .A(net79));
 sg13g2_inv_1 \proj__0.not4/_0_  (.Y(\proj__0.net11 ),
    .A(net77));
 sg13g2_xor2_1 \proj__0.xor1/_0_  (.B(net85),
    .A(net81),
    .X(\proj__0.net9 ));
 sg13g2_and2_1 \proj__1.and1/_0_  (.A(\proj__1.net18 ),
    .B(net84),
    .X(\proj__1.net19 ));
 sg13g2_and2_1 \proj__1.and2/_0_  (.A(\proj__1.net16 ),
    .B(net80),
    .X(\proj__1.net20 ));
 sg13g2_and2_1 \proj__1.and3/_0_  (.A(\proj__1.net10 ),
    .B(net2),
    .X(\proj__1.net21 ));
 sg13g2_and2_1 \proj__1.and4/_0_  (.A(\proj__1.net17 ),
    .B(net4),
    .X(\proj__1.net22 ));
 sg13g2_and2_1 \proj__1.and5/_0_  (.A(\proj__1.net20 ),
    .B(\proj__1.net19 ),
    .X(\proj__1.net23 ));
 sg13g2_and2_1 \proj__1.and6/_0_  (.A(\proj__1.net22 ),
    .B(\proj__1.net21 ),
    .X(\proj__1.net24 ));
 sg13g2_and2_1 \proj__1.and7/_0_  (.A(\proj__1.net24 ),
    .B(\proj__1.net23 ),
    .X(\proj__1.net9 ));
 sg13g2_inv_1 \proj__1.not1/_0_  (.Y(\proj__1.net16 ),
    .A(net78));
 sg13g2_inv_1 \proj__1.not2/_0_  (.Y(\proj__1.net17 ),
    .A(net5));
 sg13g2_inv_1 \proj__1.not3/_0_  (.Y(\proj__1.net18 ),
    .A(net83));
 sg13g2_inv_1 \proj__1.not4/_0_  (.Y(\proj__1.net10 ),
    .A(net76));
 sg13g2_inv_1 \proj__2.not1/_0_  (.Y(\proj__2.net9 ),
    .A(net85));
 sg13g2_inv_1 \proj__2.not2/_0_  (.Y(\proj__2.net10 ),
    .A(net82));
 sg13g2_inv_1 \proj__2.not3/_0_  (.Y(\proj__2.net11 ),
    .A(net79));
 sg13g2_inv_1 \proj__2.not4/_0_  (.Y(\proj__2.net12 ),
    .A(net77));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(\proj__3.net11 ),
    .B(net84),
    .X(\proj__3.net4 ));
 sg13g2_and2_1 \proj__3.and4/_0_  (.A(net81),
    .B(\proj__3.net12 ),
    .X(\proj__3.net3 ));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net11 ),
    .A(net81));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net12 ),
    .A(net84));
 sg13g2_inv_1 \proj__3.not6/_0_  (.Y(\proj__3.net5 ),
    .A(\proj__3.net13 ));
 sg13g2_or2_1 \proj__3.or4/_0_  (.X(\proj__3.net13 ),
    .B(\proj__3.net4 ),
    .A(\proj__3.net3 ));
 sg13g2_inv_1 \proj__4.flop1/_4_  (.Y(\proj__4.flop1/_1_ ),
    .A(\proj__4.flop1/s ));
 sg13g2_inv_1 \proj__4.flop1/_5_  (.Y(\proj__4.flop1/_0_ ),
    .A(net1));
 sg13g2_tielo \proj__4.flop1/dffsr_135  (.L_LO(net156));
 sg13g2_tielo \proj__4.flop2/dffsr_136  (.L_LO(net157));
 sg13g2_sdfbbp_1 \proj__4.flop1/dffsr  (.Q(\proj__4.flop1/q ),
    .Q_N(\proj__4.net11 ),
    .RESET_B(\proj__4.flop1/_0_ ),
    .SET_B(\proj__4.flop1/_1_ ),
    .D(net86),
    .SCE(net156),
    .SCD(net155),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_inv_1 \proj__4.flop2/_4_  (.Y(\proj__4.flop2/_1_ ),
    .A(\proj__4.flop2/s ));
 sg13g2_inv_1 \proj__4.flop2/_5_  (.Y(\proj__4.flop2/_0_ ),
    .A(net1));
 sg13g2_tielo \proj__4.flop2/dffsr_137  (.L_LO(net158));
 sg13g2_tielo \proj__4.flop3/dffsr_138  (.L_LO(net159));
 sg13g2_sdfbbp_1 \proj__4.flop2/dffsr  (.Q(\proj__4.flop2/q ),
    .Q_N(\proj__4.net12 ),
    .RESET_B(\proj__4.flop2/_0_ ),
    .SET_B(\proj__4.flop2/_1_ ),
    .D(net83),
    .SCE(net158),
    .SCD(net157),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 \proj__4.flop3/_4_  (.Y(\proj__4.flop3/_1_ ),
    .A(\proj__4.flop3/s ));
 sg13g2_inv_1 \proj__4.flop3/_5_  (.Y(\proj__4.flop3/_0_ ),
    .A(net87));
 sg13g2_tielo \proj__4.flop3/dffsr_139  (.L_LO(net160));
 sg13g2_tielo \proj__4.flop4/dffsr_140  (.L_LO(net161));
 sg13g2_sdfbbp_1 \proj__4.flop3/dffsr  (.Q(\proj__4.flop3/q ),
    .Q_N(\proj__4.net13 ),
    .RESET_B(\proj__4.flop3/_0_ ),
    .SET_B(\proj__4.flop3/_1_ ),
    .D(net79),
    .SCE(net160),
    .SCD(net159),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_inv_1 \proj__4.flop4/_4_  (.Y(\proj__4.flop4/_1_ ),
    .A(\proj__4.flop4/s ));
 sg13g2_inv_1 \proj__4.flop4/_5_  (.Y(\proj__4.flop4/_0_ ),
    .A(net87));
 sg13g2_tielo \proj__4.flop4/dffsr_141  (.L_LO(net162));
 sg13g2_tielo \proj__4.flop5/dffsr_142  (.L_LO(net163));
 sg13g2_sdfbbp_1 \proj__4.flop4/dffsr  (.Q(\proj__4.flop4/q ),
    .Q_N(\proj__4.net14 ),
    .RESET_B(\proj__4.flop4/_0_ ),
    .SET_B(\proj__4.flop4/_1_ ),
    .D(net77),
    .SCE(net162),
    .SCD(net161),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_inv_1 \proj__4.flop5/_4_  (.Y(\proj__4.flop5/_1_ ),
    .A(\proj__4.flop5/s ));
 sg13g2_inv_1 \proj__4.flop5/_5_  (.Y(\proj__4.flop5/_0_ ),
    .A(net87));
 sg13g2_tielo \proj__4.flop5/dffsr_143  (.L_LO(net164));
 sg13g2_tielo \proj__4.flop6/dffsr_144  (.L_LO(net165));
 sg13g2_sdfbbp_1 \proj__4.flop5/dffsr  (.Q(\proj__4.net15 ),
    .Q_N(\proj__4.flop5/notq ),
    .RESET_B(\proj__4.flop5/_0_ ),
    .SET_B(\proj__4.flop5/_1_ ),
    .D(net2),
    .SCE(net164),
    .SCD(net163),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_inv_1 \proj__4.flop6/_4_  (.Y(\proj__4.flop6/_1_ ),
    .A(\proj__4.flop6/s ));
 sg13g2_inv_1 \proj__4.flop6/_5_  (.Y(\proj__4.flop6/_0_ ),
    .A(net87));
 sg13g2_tielo \proj__4.flop6/dffsr_145  (.L_LO(net166));
 sg13g2_tielo \proj__4.flop8/dffsr_146  (.L_LO(net167));
 sg13g2_sdfbbp_1 \proj__4.flop6/dffsr  (.Q(\proj__4.net16 ),
    .Q_N(\proj__4.flop6/notq ),
    .RESET_B(\proj__4.flop6/_0_ ),
    .SET_B(\proj__4.flop6/_1_ ),
    .D(net76),
    .SCE(net166),
    .SCD(net165),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_inv_1 \proj__4.flop8/_4_  (.Y(\proj__4.flop8/_1_ ),
    .A(\proj__4.flop8/s ));
 sg13g2_inv_1 \proj__4.flop8/_5_  (.Y(\proj__4.flop8/_0_ ),
    .A(net87));
 sg13g2_tielo \proj__4.flop8/dffsr_147  (.L_LO(net168));
 sg13g2_tielo \proj__4.flop9/dffsr_148  (.L_LO(net169));
 sg13g2_sdfbbp_1 \proj__4.flop8/dffsr  (.Q(\proj__4.net17 ),
    .Q_N(\proj__4.flop8/notq ),
    .RESET_B(\proj__4.flop8/_0_ ),
    .SET_B(\proj__4.flop8/_1_ ),
    .D(net4),
    .SCE(net168),
    .SCD(net167),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_inv_1 \proj__4.flop9/_4_  (.Y(\proj__4.flop9/_1_ ),
    .A(\proj__4.flop9/s ));
 sg13g2_inv_1 \proj__4.flop9/_5_  (.Y(\proj__4.flop9/_0_ ),
    .A(net87));
 sg13g2_tielo \proj__4.flop9/dffsr_149  (.L_LO(net170));
 sg13g2_tielo \proj__9.flop1/dffsr_150  (.L_LO(net171));
 sg13g2_sdfbbp_1 \proj__4.flop9/dffsr  (.Q(\proj__4.net18 ),
    .Q_N(\proj__4.flop9/notq ),
    .RESET_B(\proj__4.flop9/_0_ ),
    .SET_B(\proj__4.flop9/_1_ ),
    .D(net5),
    .SCE(net170),
    .SCD(net169),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net82),
    .B(net85),
    .X(\proj__5.net9 ));
 sg13g2_and2_1 \proj__5.and2/_0_  (.A(net77),
    .B(net79),
    .X(\proj__5.net12 ));
 sg13g2_inv_1 \proj__5.not1/_0_  (.Y(\proj__5.net10 ),
    .A(net4));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net11 ),
    .B(net2),
    .A(net76));
 sg13g2_inv_1 \proj__6.not3/_0_  (.Y(\proj__6.net9 ),
    .A(net79));
 sg13g2_inv_1 \proj__6.not4/_0_  (.Y(\proj__6.net10 ),
    .A(net77));
 sg13g2_dfrbp_1 \proj__7.flop1/_1_  (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net189),
    .D(net5),
    .Q_N(\proj__7.net6 ),
    .Q(\proj__7.net5 ));
 sg13g2_tiehi \proj__7.flop2/_1__169  (.L_HI(net190));
 sg13g2_dfrbp_1 \proj__7.flop2/_1_  (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net190),
    .D(net192),
    .Q_N(\proj__7.net14 ),
    .Q(\proj__7.net8 ));
 sg13g2_tiehi \proj__7.flop3/_1__170  (.L_HI(net191));
 sg13g2_dfrbp_1 \proj__7.flop3/_1_  (.CLK(\proj__7.net14 ),
    .RESET_B(net191),
    .D(\proj__7.net15 ),
    .Q_N(\proj__7.net15 ),
    .Q(\proj__7.net7 ));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_and2_1 \proj__8.and1/_0_  (.A(net82),
    .B(net85),
    .X(\proj__8.net7 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(\proj__9.net11 ),
    .B(net86),
    .X(\proj__9.net12 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(net83),
    .B(\proj__9.net13 ),
    .X(\proj__9.net14 ));
 sg13g2_inv_1 \proj__9.flop1/_4_  (.Y(\proj__9.flop1/_1_ ),
    .A(net45));
 sg13g2_inv_1 \proj__9.flop1/_5_  (.Y(\proj__9.flop1/_0_ ),
    .A(\proj__9.net17 ));
 sg13g2_tielo \proj__9.flop1/dffsr_151  (.L_LO(net172));
 sg13g2_tiehi \proj_14.mux10/_0__152  (.L_HI(net173));
 sg13g2_sdfbbp_1 \proj__9.flop1/dffsr  (.Q(\proj__9.net5 ),
    .Q_N(\proj__9.flop1/notq ),
    .RESET_B(\proj__9.flop1/_0_ ),
    .SET_B(\proj__9.flop1/_1_ ),
    .D(\proj__9.net15 ),
    .SCE(net172),
    .SCD(net171),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 \proj__9.not1/_0_  (.Y(\proj__9.net11 ),
    .A(net83));
 sg13g2_inv_1 \proj__9.not2/_0_  (.Y(\proj__9.net13 ),
    .A(net86));
 sg13g2_inv_1 \proj__9.not3/_0_  (.Y(\proj__9.net17 ),
    .A(net1));
 sg13g2_or2_1 \proj__9.or1/_0_  (.X(\proj__9.net15 ),
    .B(\proj__9.net12 ),
    .A(\proj__9.net14 ));
 sg13g2_buf_2 fanout67 (.A(net68),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(\proj_14.net104 ),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(net70),
    .X(net69));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(net71));
 sg13g2_buf_2 fanout71 (.A(\proj_14.net25 ),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(net74));
 sg13g2_buf_2 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(\proj_14.net45 ));
 sg13g2_buf_2 fanout75 (.A(_062_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(net3),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(ui_in[3]),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(ui_in[3]),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(ui_in[2]),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(ui_in[2]),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(net83),
    .X(net81));
 sg13g2_buf_1 fanout82 (.A(net83),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(ui_in[1]),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(net86),
    .X(net84));
 sg13g2_buf_1 fanout85 (.A(net86),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(ui_in[0]),
    .X(net86));
 sg13g2_buf_4 fanout87 (.X(net87),
    .A(net1));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[4]));
 sg13g2_buf_1 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[6]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[7]));
 sg13g2_buf_2 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_tielo \proj_14.flop1/_4__10  (.L_LO(net10));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_1 clkload0 (.A(clknet_4_1_0_clk_regs));
 sg13g2_buf_1 clkload1 (.A(clknet_4_2_0_clk_regs));
 sg13g2_buf_1 clkload2 (.A(clknet_4_4_0_clk_regs));
 sg13g2_buf_1 clkload3 (.A(clknet_4_5_0_clk_regs));
 sg13g2_buf_1 clkload4 (.A(clknet_4_6_0_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_4_7_0_clk_regs));
 sg13g2_buf_1 clkload6 (.A(clknet_4_12_0_clk_regs));
 sg13g2_buf_1 clkload7 (.A(clknet_4_13_0_clk_regs));
 sg13g2_buf_1 clkload8 (.A(clknet_4_14_0_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_4_15_0_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\proj__7.net14 ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold2 (.A(\proj_13.net12 ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold3 (.A(\proj_13.net13 ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold4 (.A(\proj_14.net180 ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold5 (.A(\proj_14.net182 ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold6 (.A(\proj_14.net183 ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold7 (.A(\proj_14.net181 ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold8 (.A(\proj_14.net211 ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold9 (.A(\proj_14.net207 ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold10 (.A(\proj_14.net125 ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold11 (.A(\proj_14.net122 ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold12 (.A(\proj_14.net161 ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold13 (.A(\proj_14.net158 ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold14 (.A(\proj_14.net115 ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold15 (.A(\proj_14.net112 ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold16 (.A(\proj_14.net111 ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold17 (.A(\proj_14.net108 ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold18 (.A(\proj_14.net106 ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold19 (.A(\proj_14.net120 ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold20 (.A(\proj_14.net117 ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold21 (.A(\proj_14.net130 ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold22 (.A(\proj_14.net127 ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold23 (.A(\proj_14.net166 ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold24 (.A(\proj_14.net163 ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold25 (.A(\proj_14.net156 ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold26 (.A(\proj_14.net153 ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold27 (.A(\proj_14.net176 ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold28 (.A(\proj_14.net173 ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold29 (.A(\proj_14.net136 ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold30 (.A(\proj_14.net133 ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold31 (.A(\proj_14.net171 ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold32 (.A(\proj_14.net168 ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold33 (.A(\proj_14.net146 ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold34 (.A(\proj_14.net143 ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold35 (.A(\proj_14.net141 ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold36 (.A(\proj_14.net138 ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold37 (.A(\proj_14.net151 ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold38 (.A(\proj_14.net148 ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold39 (.A(\proj_14.net46 ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold40 (.A(\proj_14.net44 ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold41 (.A(\proj_14.net47 ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold42 (.A(\proj_14.net228 ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold43 (.A(\proj_14.net227 ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold44 (.A(\proj_14.net217 ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold45 (.A(\proj_14.net219 ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold46 (.A(\proj_14.net231 ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold47 (.A(\proj_14.net221 ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold48 (.A(\proj_14.net39 ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold49 (.A(\proj_14.net29 ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold50 (.A(\proj_14.net223 ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold51 (.A(\proj_14.net226 ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold52 (.A(\proj_14.net32 ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold53 (.A(\proj_14.net42 ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold54 (.A(\proj_14.net36 ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold55 (.A(\proj_14.net26 ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold56 (.A(\proj_14.net27 ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold57 (.A(\proj_14.net26 ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold58 (.A(\proj_14.net27 ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold59 (.A(\proj_14.net26 ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold60 (.A(\proj_14.net26 ),
    .X(net251));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_fill_1 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_fill_1 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_fill_1 FILLER_17_329 ();
 sg13g2_decap_4 FILLER_17_334 ();
 sg13g2_fill_1 FILLER_17_338 ();
 sg13g2_fill_1 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_fill_2 FILLER_17_403 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_82 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_99 ();
 sg13g2_decap_4 FILLER_18_106 ();
 sg13g2_decap_8 FILLER_18_113 ();
 sg13g2_decap_8 FILLER_18_120 ();
 sg13g2_decap_8 FILLER_18_127 ();
 sg13g2_decap_8 FILLER_18_134 ();
 sg13g2_decap_8 FILLER_18_141 ();
 sg13g2_decap_8 FILLER_18_148 ();
 sg13g2_decap_8 FILLER_18_155 ();
 sg13g2_decap_8 FILLER_18_162 ();
 sg13g2_decap_8 FILLER_18_169 ();
 sg13g2_decap_8 FILLER_18_176 ();
 sg13g2_decap_8 FILLER_18_183 ();
 sg13g2_decap_8 FILLER_18_195 ();
 sg13g2_decap_8 FILLER_18_202 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_decap_8 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_fill_1 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_decap_8 FILLER_18_314 ();
 sg13g2_fill_2 FILLER_18_321 ();
 sg13g2_fill_1 FILLER_18_323 ();
 sg13g2_fill_2 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_4 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_43 ();
 sg13g2_decap_8 FILLER_19_50 ();
 sg13g2_fill_1 FILLER_19_57 ();
 sg13g2_fill_2 FILLER_19_70 ();
 sg13g2_fill_1 FILLER_19_72 ();
 sg13g2_decap_8 FILLER_19_121 ();
 sg13g2_decap_8 FILLER_19_128 ();
 sg13g2_decap_8 FILLER_19_135 ();
 sg13g2_decap_8 FILLER_19_142 ();
 sg13g2_decap_8 FILLER_19_149 ();
 sg13g2_decap_8 FILLER_19_156 ();
 sg13g2_decap_8 FILLER_19_163 ();
 sg13g2_decap_8 FILLER_19_170 ();
 sg13g2_decap_8 FILLER_19_177 ();
 sg13g2_decap_8 FILLER_19_184 ();
 sg13g2_decap_8 FILLER_19_191 ();
 sg13g2_decap_8 FILLER_19_198 ();
 sg13g2_decap_8 FILLER_19_205 ();
 sg13g2_decap_8 FILLER_19_212 ();
 sg13g2_decap_8 FILLER_19_219 ();
 sg13g2_decap_8 FILLER_19_226 ();
 sg13g2_decap_8 FILLER_19_233 ();
 sg13g2_decap_4 FILLER_19_240 ();
 sg13g2_fill_1 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_357 ();
 sg13g2_decap_4 FILLER_19_379 ();
 sg13g2_fill_1 FILLER_19_383 ();
 sg13g2_fill_2 FILLER_19_398 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_127 ();
 sg13g2_fill_1 FILLER_20_129 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_4 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_fill_2 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_296 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_decap_4 FILLER_20_312 ();
 sg13g2_fill_1 FILLER_20_316 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_24 ();
 sg13g2_fill_2 FILLER_21_31 ();
 sg13g2_fill_2 FILLER_21_37 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_85 ();
 sg13g2_decap_4 FILLER_21_92 ();
 sg13g2_fill_2 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_decap_4 FILLER_21_118 ();
 sg13g2_fill_1 FILLER_21_132 ();
 sg13g2_decap_4 FILLER_21_141 ();
 sg13g2_fill_1 FILLER_21_157 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_decap_8 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_decap_8 FILLER_21_190 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_4 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_212 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_4 FILLER_21_224 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_1 FILLER_21_344 ();
 sg13g2_decap_4 FILLER_21_355 ();
 sg13g2_fill_2 FILLER_21_364 ();
 sg13g2_fill_2 FILLER_21_374 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_47 ();
 sg13g2_decap_8 FILLER_22_72 ();
 sg13g2_fill_2 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_decap_4 FILLER_22_89 ();
 sg13g2_fill_2 FILLER_22_150 ();
 sg13g2_decap_8 FILLER_22_170 ();
 sg13g2_decap_8 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_271 ();
 sg13g2_decap_4 FILLER_22_284 ();
 sg13g2_fill_2 FILLER_22_288 ();
 sg13g2_decap_4 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_303 ();
 sg13g2_fill_2 FILLER_22_310 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_11 ();
 sg13g2_decap_4 FILLER_23_20 ();
 sg13g2_fill_2 FILLER_23_24 ();
 sg13g2_decap_4 FILLER_23_33 ();
 sg13g2_fill_1 FILLER_23_37 ();
 sg13g2_fill_2 FILLER_23_60 ();
 sg13g2_fill_1 FILLER_23_62 ();
 sg13g2_fill_1 FILLER_23_101 ();
 sg13g2_fill_2 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_225 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_decap_4 FILLER_23_290 ();
 sg13g2_decap_4 FILLER_23_297 ();
 sg13g2_fill_1 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_338 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_decap_4 FILLER_24_87 ();
 sg13g2_fill_2 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_96 ();
 sg13g2_fill_2 FILLER_24_106 ();
 sg13g2_fill_2 FILLER_24_113 ();
 sg13g2_decap_4 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_decap_4 FILLER_24_148 ();
 sg13g2_fill_2 FILLER_24_152 ();
 sg13g2_decap_4 FILLER_24_157 ();
 sg13g2_fill_2 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_4 FILLER_24_175 ();
 sg13g2_decap_4 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_274 ();
 sg13g2_decap_4 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_325 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_decap_4 FILLER_24_374 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_fill_2 FILLER_24_392 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_30 ();
 sg13g2_fill_2 FILLER_25_37 ();
 sg13g2_decap_4 FILLER_25_62 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_decap_8 FILLER_25_174 ();
 sg13g2_decap_4 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_decap_4 FILLER_25_274 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_2 FILLER_25_300 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_decap_4 FILLER_25_306 ();
 sg13g2_fill_2 FILLER_25_310 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_decap_4 FILLER_25_323 ();
 sg13g2_fill_2 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_fill_2 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_72 ();
 sg13g2_fill_1 FILLER_26_118 ();
 sg13g2_decap_8 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_211 ();
 sg13g2_decap_4 FILLER_26_216 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_230 ();
 sg13g2_decap_4 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_286 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_331 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_390 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_32 ();
 sg13g2_decap_4 FILLER_27_51 ();
 sg13g2_fill_2 FILLER_27_59 ();
 sg13g2_fill_1 FILLER_27_61 ();
 sg13g2_fill_2 FILLER_27_83 ();
 sg13g2_decap_4 FILLER_27_93 ();
 sg13g2_fill_1 FILLER_27_97 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_170 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_241 ();
 sg13g2_fill_2 FILLER_27_246 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_fill_2 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_282 ();
 sg13g2_decap_4 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_318 ();
 sg13g2_decap_8 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_332 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_351 ();
 sg13g2_decap_4 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_25 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_101 ();
 sg13g2_decap_8 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_117 ();
 sg13g2_decap_8 FILLER_28_130 ();
 sg13g2_fill_2 FILLER_28_137 ();
 sg13g2_decap_4 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_fill_2 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_230 ();
 sg13g2_fill_1 FILLER_28_237 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_310 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_fill_2 FILLER_28_379 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_11 ();
 sg13g2_decap_4 FILLER_29_47 ();
 sg13g2_fill_2 FILLER_29_51 ();
 sg13g2_decap_4 FILLER_29_60 ();
 sg13g2_fill_1 FILLER_29_64 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_fill_2 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_201 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_decap_8 FILLER_29_256 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_296 ();
 sg13g2_fill_2 FILLER_29_303 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_fill_2 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_23 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_4 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_39 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_101 ();
 sg13g2_fill_2 FILLER_30_113 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_decap_4 FILLER_30_131 ();
 sg13g2_fill_2 FILLER_30_145 ();
 sg13g2_fill_1 FILLER_30_147 ();
 sg13g2_decap_4 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_decap_4 FILLER_30_179 ();
 sg13g2_decap_4 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_241 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_decap_4 FILLER_30_304 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_314 ();
 sg13g2_fill_1 FILLER_30_316 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_4 FILLER_30_329 ();
 sg13g2_decap_4 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_2 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_fill_1 FILLER_30_391 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_25 ();
 sg13g2_decap_4 FILLER_31_30 ();
 sg13g2_decap_4 FILLER_31_52 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_144 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_decap_4 FILLER_31_278 ();
 sg13g2_decap_4 FILLER_31_289 ();
 sg13g2_decap_4 FILLER_31_308 ();
 sg13g2_fill_2 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_41 ();
 sg13g2_decap_8 FILLER_32_48 ();
 sg13g2_fill_1 FILLER_32_55 ();
 sg13g2_fill_2 FILLER_32_81 ();
 sg13g2_fill_1 FILLER_32_83 ();
 sg13g2_fill_1 FILLER_32_104 ();
 sg13g2_decap_8 FILLER_32_110 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_decap_4 FILLER_32_163 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_fill_2 FILLER_32_214 ();
 sg13g2_fill_1 FILLER_32_216 ();
 sg13g2_decap_8 FILLER_32_220 ();
 sg13g2_decap_8 FILLER_32_227 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_296 ();
 sg13g2_decap_8 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_2 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_4 FILLER_32_372 ();
 sg13g2_fill_2 FILLER_32_376 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_2 FILLER_33_25 ();
 sg13g2_fill_1 FILLER_33_36 ();
 sg13g2_fill_1 FILLER_33_41 ();
 sg13g2_decap_4 FILLER_33_101 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_fill_2 FILLER_33_136 ();
 sg13g2_decap_4 FILLER_33_173 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_fill_1 FILLER_33_214 ();
 sg13g2_decap_4 FILLER_33_247 ();
 sg13g2_decap_4 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_decap_4 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_336 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_fill_2 FILLER_33_357 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_fill_2 FILLER_33_391 ();
 sg13g2_fill_1 FILLER_33_402 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_25 ();
 sg13g2_decap_8 FILLER_34_52 ();
 sg13g2_fill_1 FILLER_34_59 ();
 sg13g2_fill_1 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_111 ();
 sg13g2_decap_8 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_decap_8 FILLER_34_163 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_decap_4 FILLER_34_220 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_decap_4 FILLER_34_253 ();
 sg13g2_decap_4 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_327 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_353 ();
 sg13g2_decap_8 FILLER_34_360 ();
 sg13g2_fill_2 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_46 ();
 sg13g2_decap_8 FILLER_35_53 ();
 sg13g2_decap_8 FILLER_35_60 ();
 sg13g2_fill_1 FILLER_35_67 ();
 sg13g2_decap_8 FILLER_35_78 ();
 sg13g2_fill_1 FILLER_35_85 ();
 sg13g2_decap_4 FILLER_35_111 ();
 sg13g2_decap_8 FILLER_35_146 ();
 sg13g2_decap_8 FILLER_35_153 ();
 sg13g2_decap_8 FILLER_35_160 ();
 sg13g2_decap_8 FILLER_35_167 ();
 sg13g2_decap_8 FILLER_35_174 ();
 sg13g2_decap_8 FILLER_35_181 ();
 sg13g2_decap_8 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_decap_4 FILLER_35_252 ();
 sg13g2_fill_2 FILLER_35_256 ();
 sg13g2_decap_4 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_decap_4 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_fill_2 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_decap_4 FILLER_35_383 ();
 sg13g2_fill_2 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_4 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_130 ();
 sg13g2_decap_8 FILLER_36_135 ();
 sg13g2_decap_8 FILLER_36_142 ();
 sg13g2_decap_8 FILLER_36_149 ();
 sg13g2_decap_8 FILLER_36_156 ();
 sg13g2_decap_8 FILLER_36_163 ();
 sg13g2_decap_8 FILLER_36_170 ();
 sg13g2_decap_8 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_191 ();
 sg13g2_decap_8 FILLER_36_198 ();
 sg13g2_decap_8 FILLER_36_209 ();
 sg13g2_decap_4 FILLER_36_216 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_decap_4 FILLER_36_254 ();
 sg13g2_fill_1 FILLER_36_258 ();
 sg13g2_decap_4 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_decap_4 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_fill_1 FILLER_36_347 ();
 sg13g2_decap_4 FILLER_36_351 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_fill_2 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_fill_1 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_4 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_214 ();
 sg13g2_decap_8 FILLER_37_254 ();
 sg13g2_decap_8 FILLER_37_261 ();
 sg13g2_fill_1 FILLER_37_268 ();
 sg13g2_decap_4 FILLER_37_281 ();
 sg13g2_fill_2 FILLER_37_328 ();
 sg13g2_fill_2 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_233 ();
 sg13g2_decap_8 FILLER_38_240 ();
 sg13g2_decap_8 FILLER_38_247 ();
 sg13g2_decap_8 FILLER_38_254 ();
 sg13g2_decap_8 FILLER_38_261 ();
 sg13g2_decap_8 FILLER_38_268 ();
 sg13g2_decap_4 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_fill_1 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net46;
 assign uio_oe[1] = net47;
 assign uio_oe[2] = net48;
 assign uio_oe[3] = net49;
 assign uio_oe[4] = net50;
 assign uio_oe[5] = net51;
 assign uio_oe[6] = net52;
 assign uio_oe[7] = net53;
 assign uio_out[0] = net54;
 assign uio_out[1] = net55;
 assign uio_out[2] = net56;
 assign uio_out[3] = net57;
 assign uio_out[4] = net58;
 assign uio_out[5] = net59;
 assign uio_out[6] = net60;
 assign uio_out[7] = net61;
endmodule

module tt_um_supermic_arghunter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][9] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][9] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.i_data ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[9] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[9] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.i_data ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.i_data ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.i_data ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.i_data ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.i_data ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.i_data ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.i_data ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[9] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[0] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[10] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[11] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[12] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[13] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[14] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[15] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[16] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[17] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[18] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[1] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[2] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[3] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[4] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[5] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[6] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[7] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[8] ;
 wire \u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[9] ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.out ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.out ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.out ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.out ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.out ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.out ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.out ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.out ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.u_mux_shift.data ;
 wire \u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.u_mux_shift.sum_res ;
 wire \u_supermic_top_module.i2s_out ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][9] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][0] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][10] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][11] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][12] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][13] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][14] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][15] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][16] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][17] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][18] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][1] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][2] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][3] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][4] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][5] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][6] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][7] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][8] ;
 wire \u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][9] ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_supermic_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_supermic_top_module.u_i2s_bus.u_mux_shift.data ;
 wire \u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[0].u_ddr_to_sdr_dual.ddr_data_falling ;
 wire \u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[0].u_ddr_to_sdr_dual.ddr_data_rising ;
 wire \u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[1].u_ddr_to_sdr_dual.ddr_data_falling ;
 wire \u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[1].u_ddr_to_sdr_dual.ddr_data_rising ;
 wire \u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[2].u_ddr_to_sdr_dual.ddr_data_falling ;
 wire \u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[2].u_ddr_to_sdr_dual.ddr_data_rising ;
 wire \u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[3].u_ddr_to_sdr_dual.ddr_data_falling ;
 wire \u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[3].u_ddr_to_sdr_dual.ddr_data_rising ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net6079;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;

 sg13g2_inv_1 _10717_ (.Y(_01458_),
    .A(net5151));
 sg13g2_inv_1 _10718_ (.Y(_02332_),
    .A(net4991));
 sg13g2_inv_1 _10719_ (.Y(_02333_),
    .A(net4997));
 sg13g2_inv_1 _10720_ (.Y(_02334_),
    .A(net5005));
 sg13g2_inv_1 _10721_ (.Y(_02335_),
    .A(net5010));
 sg13g2_inv_1 _10722_ (.Y(_02336_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][0] ));
 sg13g2_inv_1 _10723_ (.Y(_02337_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][0] ));
 sg13g2_inv_1 _10724_ (.Y(_02338_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][0] ));
 sg13g2_inv_1 _10725_ (.Y(_02339_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][0] ));
 sg13g2_inv_1 _10726_ (.Y(_02340_),
    .A(_00293_));
 sg13g2_inv_1 _10727_ (.Y(_02341_),
    .A(_00294_));
 sg13g2_inv_1 _10728_ (.Y(_02342_),
    .A(_00301_));
 sg13g2_inv_1 _10729_ (.Y(_02343_),
    .A(_00308_));
 sg13g2_inv_1 _10730_ (.Y(_02344_),
    .A(_00317_));
 sg13g2_inv_1 _10731_ (.Y(_02345_),
    .A(_00333_));
 sg13g2_inv_1 _10732_ (.Y(_02346_),
    .A(_00340_));
 sg13g2_inv_1 _10733_ (.Y(_02347_),
    .A(_00349_));
 sg13g2_inv_1 _10734_ (.Y(_02348_),
    .A(_00365_));
 sg13g2_inv_1 _10735_ (.Y(_02349_),
    .A(_00372_));
 sg13g2_inv_1 _10736_ (.Y(_02350_),
    .A(_00397_));
 sg13g2_inv_1 _10737_ (.Y(_02351_),
    .A(_00404_));
 sg13g2_inv_1 _10738_ (.Y(_02352_),
    .A(_00415_));
 sg13g2_inv_1 _10739_ (.Y(_02353_),
    .A(_00420_));
 sg13g2_inv_1 _10740_ (.Y(_02354_),
    .A(_00422_));
 sg13g2_inv_1 _10741_ (.Y(_02355_),
    .A(_00429_));
 sg13g2_inv_1 _10742_ (.Y(_02356_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_inv_1 _10743_ (.Y(_02357_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_inv_1 _10744_ (.Y(_02358_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_inv_1 _10745_ (.Y(_02359_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_inv_1 _10746_ (.Y(_02360_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_inv_1 _10747_ (.Y(_02361_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_inv_1 _10748_ (.Y(_02362_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_inv_1 _10749_ (.Y(_02363_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_inv_1 _10750_ (.Y(_02364_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_inv_1 _10751_ (.Y(_02365_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_inv_1 _10752_ (.Y(_02366_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_inv_1 _10753_ (.Y(_02367_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_inv_1 _10754_ (.Y(_02368_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_inv_1 _10755_ (.Y(_02369_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_inv_1 _10756_ (.Y(_02370_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_inv_1 _10757_ (.Y(_02371_),
    .A(net4957));
 sg13g2_inv_1 _10758_ (.Y(_02372_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10759_ (.Y(_02373_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10760_ (.Y(_02374_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10761_ (.Y(_02375_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_inv_1 _10762_ (.Y(_02376_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_inv_1 _10763_ (.Y(_02377_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_inv_1 _10764_ (.Y(_02378_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_inv_1 _10765_ (.Y(_02379_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10766_ (.Y(_02380_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_inv_1 _10767_ (.Y(_02381_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_inv_1 _10768_ (.Y(_02382_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_inv_1 _10769_ (.Y(_02383_),
    .A(net4976));
 sg13g2_inv_1 _10770_ (.Y(_02384_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10771_ (.Y(_02385_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10772_ (.Y(_02386_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10773_ (.Y(_02387_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][7] ));
 sg13g2_inv_1 _10774_ (.Y(_02388_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10775_ (.Y(_02389_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_inv_1 _10776_ (.Y(_02390_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_inv_1 _10777_ (.Y(_02391_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_inv_1 _10778_ (.Y(_02392_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10779_ (.Y(_02393_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10780_ (.Y(_02394_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10781_ (.Y(_02395_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_inv_1 _10782_ (.Y(_02396_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_inv_1 _10783_ (.Y(_02397_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_inv_1 _10784_ (.Y(_02398_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_inv_1 _10785_ (.Y(_02399_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10786_ (.Y(_02400_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_inv_1 _10787_ (.Y(_02401_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_inv_1 _10788_ (.Y(_02402_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_inv_1 _10789_ (.Y(_02403_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_inv_1 _10790_ (.Y(_02404_),
    .A(net4970));
 sg13g2_inv_1 _10791_ (.Y(_02405_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10792_ (.Y(_02406_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10793_ (.Y(_02407_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10794_ (.Y(_02408_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_inv_1 _10795_ (.Y(_02409_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_inv_1 _10796_ (.Y(_02410_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_inv_1 _10797_ (.Y(_02411_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_inv_1 _10798_ (.Y(_02412_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10799_ (.Y(_02413_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10800_ (.Y(_02414_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10801_ (.Y(_02415_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10802_ (.Y(_02416_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][7] ));
 sg13g2_inv_1 _10803_ (.Y(_02417_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_inv_1 _10804_ (.Y(_02418_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_inv_1 _10805_ (.Y(_02419_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_inv_1 _10806_ (.Y(_02420_),
    .A(net4962));
 sg13g2_inv_1 _10807_ (.Y(_02421_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10808_ (.Y(_02422_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10809_ (.Y(_02423_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10810_ (.Y(_02424_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][7] ));
 sg13g2_inv_1 _10811_ (.Y(_02425_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10812_ (.Y(_02426_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10813_ (.Y(_02427_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10814_ (.Y(_02428_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10815_ (.Y(_02429_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_inv_1 _10816_ (.Y(_02430_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_inv_1 _10817_ (.Y(_02431_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_inv_1 _10818_ (.Y(_02432_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_inv_1 _10819_ (.Y(_02433_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10820_ (.Y(_02434_),
    .A(net4972));
 sg13g2_inv_1 _10821_ (.Y(_02435_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_inv_1 _10822_ (.Y(_02436_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_inv_1 _10823_ (.Y(_02437_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_inv_1 _10824_ (.Y(_02438_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10825_ (.Y(_02439_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10826_ (.Y(_02440_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10827_ (.Y(_02441_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_inv_1 _10828_ (.Y(_02442_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_inv_1 _10829_ (.Y(_02443_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_inv_1 _10830_ (.Y(_02444_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_inv_1 _10831_ (.Y(_02445_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10832_ (.Y(_02446_),
    .A(net4982));
 sg13g2_inv_1 _10833_ (.Y(_02447_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_inv_1 _10834_ (.Y(_02448_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_inv_1 _10835_ (.Y(_02449_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_inv_1 _10836_ (.Y(_02450_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_inv_1 _10837_ (.Y(_02451_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10838_ (.Y(_02452_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10839_ (.Y(_02453_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10840_ (.Y(_02454_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][7] ));
 sg13g2_inv_1 _10841_ (.Y(_02455_),
    .A(net4951));
 sg13g2_inv_1 _10842_ (.Y(_02456_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_inv_1 _10843_ (.Y(_02457_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_inv_1 _10844_ (.Y(_02458_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_inv_1 _10845_ (.Y(_02459_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_inv_1 _10846_ (.Y(_02460_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10847_ (.Y(_02461_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10848_ (.Y(_02462_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10849_ (.Y(_02463_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_inv_1 _10850_ (.Y(_02464_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_inv_1 _10851_ (.Y(_02465_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_inv_1 _10852_ (.Y(_02466_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_inv_1 _10853_ (.Y(_02467_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10854_ (.Y(_02468_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10855_ (.Y(_02469_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10856_ (.Y(_02470_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10857_ (.Y(_02471_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][7] ));
 sg13g2_inv_1 _10858_ (.Y(_02472_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10859_ (.Y(_02473_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10860_ (.Y(_02474_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10861_ (.Y(_02475_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10862_ (.Y(_02476_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][7] ));
 sg13g2_inv_1 _10863_ (.Y(_02477_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10864_ (.Y(_02478_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10865_ (.Y(_02479_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10866_ (.Y(_02480_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10867_ (.Y(_02481_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][7] ));
 sg13g2_inv_1 _10868_ (.Y(_02482_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10869_ (.Y(_02483_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10870_ (.Y(_02484_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10871_ (.Y(_02485_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10872_ (.Y(_02486_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_inv_1 _10873_ (.Y(_02487_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_inv_1 _10874_ (.Y(_02488_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_inv_1 _10875_ (.Y(_02489_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_inv_1 _10876_ (.Y(_02490_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10877_ (.Y(_02491_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10878_ (.Y(_02492_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10879_ (.Y(_02493_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10880_ (.Y(_02494_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_inv_1 _10881_ (.Y(_02495_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_inv_1 _10882_ (.Y(_02496_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_inv_1 _10883_ (.Y(_02497_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_inv_1 _10884_ (.Y(_02498_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10885_ (.Y(_02499_),
    .A(net4963));
 sg13g2_inv_1 _10886_ (.Y(_02500_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_inv_1 _10887_ (.Y(_02501_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_inv_1 _10888_ (.Y(_02502_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_inv_1 _10889_ (.Y(_02503_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][7] ));
 sg13g2_inv_1 _10890_ (.Y(_02504_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_inv_1 _10891_ (.Y(_01194_),
    .A(net5219));
 sg13g2_and2_1 _10892_ (.A(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .B(net5721),
    .X(_01807_));
 sg13g2_and2_1 _10893_ (.A(net5720),
    .B(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .X(_01806_));
 sg13g2_and2_1 _10894_ (.A(net5723),
    .B(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .X(_01805_));
 sg13g2_and2_1 _10895_ (.A(net5729),
    .B(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .X(_01804_));
 sg13g2_and2_1 _10896_ (.A(net5728),
    .B(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .X(_01803_));
 sg13g2_and2_1 _10897_ (.A(net5720),
    .B(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .X(_01802_));
 sg13g2_and2_1 _10898_ (.A(net5719),
    .B(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .X(_01801_));
 sg13g2_and2_1 _10899_ (.A(net5722),
    .B(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .X(_01800_));
 sg13g2_and2_1 _10900_ (.A(net5729),
    .B(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .X(_01799_));
 sg13g2_nand2b_1 _10901_ (.Y(_02505_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][0] ));
 sg13g2_xor2_1 _10902_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][0] ),
    .X(_00434_));
 sg13g2_nand2b_1 _10903_ (.Y(_02506_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][0] ));
 sg13g2_xor2_1 _10904_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][0] ),
    .X(_01017_));
 sg13g2_nand2b_1 _10905_ (.Y(_02507_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][0] ));
 sg13g2_xor2_1 _10906_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][0] ),
    .X(_00528_));
 sg13g2_nand2b_1 _10907_ (.Y(_02508_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][0] ));
 sg13g2_xor2_1 _10908_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][0] ),
    .X(_00453_));
 sg13g2_nand2b_1 _10909_ (.Y(_02509_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][0] ));
 sg13g2_xor2_1 _10910_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][0] ),
    .X(_00622_));
 sg13g2_nand2b_1 _10911_ (.Y(_02510_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][0] ));
 sg13g2_xor2_1 _10912_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][0] ),
    .X(_00547_));
 sg13g2_nand2b_1 _10913_ (.Y(_02511_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][0] ));
 sg13g2_xor2_1 _10914_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][0] ),
    .X(_00716_));
 sg13g2_nand2b_1 _10915_ (.Y(_02512_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][0] ));
 sg13g2_xor2_1 _10916_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][0] ),
    .X(_00641_));
 sg13g2_nand2b_1 _10917_ (.Y(_02513_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][0] ));
 sg13g2_xor2_1 _10918_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][0] ),
    .X(_00810_));
 sg13g2_nand2b_1 _10919_ (.Y(_02514_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][0] ));
 sg13g2_xor2_1 _10920_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][0] ),
    .X(_00735_));
 sg13g2_nand2b_1 _10921_ (.Y(_02515_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][0] ));
 sg13g2_xor2_1 _10922_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][0] ),
    .X(_00923_));
 sg13g2_nand2b_1 _10923_ (.Y(_02516_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][0] ));
 sg13g2_xor2_1 _10924_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][0] ),
    .X(_00998_));
 sg13g2_nand2b_1 _10925_ (.Y(_02517_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][0] ));
 sg13g2_xor2_1 _10926_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][0] ),
    .X(_00904_));
 sg13g2_nand2b_1 _10927_ (.Y(_02518_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][0] ));
 sg13g2_xor2_1 _10928_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][0] ),
    .X(_01111_));
 sg13g2_nand2b_2 _10929_ (.Y(_02519_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][0] ));
 sg13g2_xor2_1 _10930_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][0] ),
    .X(_01092_));
 sg13g2_nand2b_1 _10931_ (.Y(_02520_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][0] ));
 sg13g2_xor2_1 _10932_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[0] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][0] ),
    .X(_00829_));
 sg13g2_nor2_2 _10933_ (.A(_01458_),
    .B(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ),
    .Y(_02521_));
 sg13g2_nand2b_1 _10934_ (.Y(_02522_),
    .B(net5151),
    .A_N(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ));
 sg13g2_mux2_1 _10935_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .S(net4921),
    .X(_00234_));
 sg13g2_mux2_1 _10936_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .S(net4920),
    .X(_00245_));
 sg13g2_mux2_1 _10937_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .S(net4920),
    .X(_00248_));
 sg13g2_mux2_1 _10938_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .S(net4922),
    .X(_00249_));
 sg13g2_mux2_1 _10939_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .S(net4922),
    .X(_00250_));
 sg13g2_mux2_1 _10940_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .S(net4922),
    .X(_00251_));
 sg13g2_mux2_1 _10941_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .S(net4920),
    .X(_00252_));
 sg13g2_mux2_1 _10942_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .S(net4922),
    .X(_00253_));
 sg13g2_mux2_1 _10943_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .S(net4922),
    .X(_00254_));
 sg13g2_mux2_1 _10944_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .S(net4921),
    .X(_00224_));
 sg13g2_mux2_1 _10945_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .S(net4921),
    .X(_00225_));
 sg13g2_mux2_1 _10946_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .S(net4921),
    .X(_00226_));
 sg13g2_mux2_1 _10947_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .S(net4921),
    .X(_00227_));
 sg13g2_mux2_1 _10948_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .S(net4921),
    .X(_00228_));
 sg13g2_mux2_1 _10949_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .S(net4921),
    .X(_00229_));
 sg13g2_mux2_1 _10950_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .S(net4921),
    .X(_00230_));
 sg13g2_mux2_1 _10951_ (.A0(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .S(net4919),
    .X(_00231_));
 sg13g2_and2_1 _10952_ (.A(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .B(net4932),
    .X(_02523_));
 sg13g2_a21o_1 _10953_ (.A2(net4919),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B1(net4870),
    .X(_00232_));
 sg13g2_a21o_1 _10954_ (.A2(net4918),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B1(net4870),
    .X(_00233_));
 sg13g2_a21o_1 _10955_ (.A2(net4916),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B1(net4870),
    .X(_00235_));
 sg13g2_a21o_1 _10956_ (.A2(net4916),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .B1(net4870),
    .X(_00236_));
 sg13g2_a21o_1 _10957_ (.A2(net4913),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .B1(net4870),
    .X(_00237_));
 sg13g2_a21o_1 _10958_ (.A2(net4903),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B1(net4869),
    .X(_00238_));
 sg13g2_a21o_1 _10959_ (.A2(net4903),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B1(net4869),
    .X(_00239_));
 sg13g2_a21o_1 _10960_ (.A2(net4906),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B1(net4869),
    .X(_00240_));
 sg13g2_a21o_1 _10961_ (.A2(net4906),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B1(net4869),
    .X(_00241_));
 sg13g2_a21o_1 _10962_ (.A2(net4904),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B1(net4869),
    .X(_00242_));
 sg13g2_a21o_1 _10963_ (.A2(net4904),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B1(net4869),
    .X(_00243_));
 sg13g2_a21o_1 _10964_ (.A2(net4904),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B1(net4869),
    .X(_00244_));
 sg13g2_a21o_1 _10965_ (.A2(net4904),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B1(net4869),
    .X(_00246_));
 sg13g2_a21o_2 _10966_ (.A2(net4906),
    .A1(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B1(net4870),
    .X(_00247_));
 sg13g2_mux2_1 _10967_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .S(net4912),
    .X(_00202_));
 sg13g2_mux2_1 _10968_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .S(net4913),
    .X(_00213_));
 sg13g2_mux2_1 _10969_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .S(net4914),
    .X(_00216_));
 sg13g2_mux2_1 _10970_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .S(net4914),
    .X(_00217_));
 sg13g2_mux2_1 _10971_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .S(net4914),
    .X(_00218_));
 sg13g2_mux2_1 _10972_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .S(net4914),
    .X(_00219_));
 sg13g2_mux2_1 _10973_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .S(net4914),
    .X(_00220_));
 sg13g2_mux2_1 _10974_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .S(net4913),
    .X(_00221_));
 sg13g2_mux2_1 _10975_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .S(net4910),
    .X(_00222_));
 sg13g2_mux2_1 _10976_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .S(net4910),
    .X(_00192_));
 sg13g2_mux2_1 _10977_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .S(net4910),
    .X(_00193_));
 sg13g2_mux2_1 _10978_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .S(net4910),
    .X(_00194_));
 sg13g2_mux2_1 _10979_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .S(net4910),
    .X(_00195_));
 sg13g2_mux2_1 _10980_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .S(net4907),
    .X(_00196_));
 sg13g2_mux2_1 _10981_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .S(net4910),
    .X(_00197_));
 sg13g2_mux2_1 _10982_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .S(net4913),
    .X(_00198_));
 sg13g2_mux2_1 _10983_ (.A0(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .S(net4906),
    .X(_00199_));
 sg13g2_and2_1 _10984_ (.A(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .B(net4925),
    .X(_02524_));
 sg13g2_a21o_1 _10985_ (.A2(net4904),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B1(net4868),
    .X(_00200_));
 sg13g2_a21o_1 _10986_ (.A2(net4904),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B1(net4868),
    .X(_00201_));
 sg13g2_a21o_1 _10987_ (.A2(net4902),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B1(net4868),
    .X(_00203_));
 sg13g2_a21o_1 _10988_ (.A2(net4902),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .B1(net4867),
    .X(_00204_));
 sg13g2_a21o_1 _10989_ (.A2(net4901),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .B1(net4867),
    .X(_00205_));
 sg13g2_a21o_1 _10990_ (.A2(net4901),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B1(net4867),
    .X(_00206_));
 sg13g2_a21o_1 _10991_ (.A2(net4901),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B1(net4867),
    .X(_00207_));
 sg13g2_a21o_1 _10992_ (.A2(net4901),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B1(net4867),
    .X(_00208_));
 sg13g2_a21o_1 _10993_ (.A2(net4902),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B1(net4867),
    .X(_00209_));
 sg13g2_a21o_1 _10994_ (.A2(net4902),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B1(net4867),
    .X(_00210_));
 sg13g2_a21o_1 _10995_ (.A2(net4903),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B1(net4868),
    .X(_00211_));
 sg13g2_a21o_1 _10996_ (.A2(net4903),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B1(net4868),
    .X(_00212_));
 sg13g2_a21o_1 _10997_ (.A2(net4905),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B1(net4867),
    .X(_00214_));
 sg13g2_a21o_2 _10998_ (.A2(net4905),
    .A1(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B1(net4868),
    .X(_00215_));
 sg13g2_mux2_1 _10999_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .S(net4907),
    .X(_00170_));
 sg13g2_mux2_1 _11000_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .S(net4907),
    .X(_00181_));
 sg13g2_mux2_1 _11001_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .S(net4908),
    .X(_00184_));
 sg13g2_mux2_1 _11002_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .S(net4907),
    .X(_00185_));
 sg13g2_mux2_1 _11003_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .S(net4907),
    .X(_00186_));
 sg13g2_mux2_1 _11004_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .S(net4907),
    .X(_00187_));
 sg13g2_mux2_1 _11005_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .S(net4907),
    .X(_00188_));
 sg13g2_mux2_1 _11006_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .S(net4907),
    .X(_00189_));
 sg13g2_mux2_1 _11007_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .S(net4898),
    .X(_00190_));
 sg13g2_mux2_1 _11008_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .S(net4898),
    .X(_00160_));
 sg13g2_mux2_1 _11009_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .S(net4898),
    .X(_00161_));
 sg13g2_mux2_1 _11010_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .S(net4897),
    .X(_00162_));
 sg13g2_mux2_1 _11011_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .S(net4897),
    .X(_00163_));
 sg13g2_mux2_1 _11012_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .S(net4897),
    .X(_00164_));
 sg13g2_mux2_1 _11013_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .S(net4897),
    .X(_00165_));
 sg13g2_mux2_1 _11014_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .S(net4897),
    .X(_00166_));
 sg13g2_mux2_2 _11015_ (.A0(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .S(net4898),
    .X(_00167_));
 sg13g2_and2_1 _11016_ (.A(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .B(net4928),
    .X(_02525_));
 sg13g2_a21o_1 _11017_ (.A2(net4899),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B1(net4866),
    .X(_00168_));
 sg13g2_a21o_1 _11018_ (.A2(net4891),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B1(net4866),
    .X(_00169_));
 sg13g2_a21o_1 _11019_ (.A2(net4891),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B1(net4866),
    .X(_00171_));
 sg13g2_a21o_1 _11020_ (.A2(net4885),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .B1(net4865),
    .X(_00172_));
 sg13g2_a21o_1 _11021_ (.A2(net4882),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .B1(net4865),
    .X(_00173_));
 sg13g2_a21o_1 _11022_ (.A2(net4881),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B1(net4865),
    .X(_00174_));
 sg13g2_a21o_1 _11023_ (.A2(net4880),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B1(net4864),
    .X(_00175_));
 sg13g2_a21o_1 _11024_ (.A2(net4880),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B1(net4864),
    .X(_00176_));
 sg13g2_a21o_1 _11025_ (.A2(net4880),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B1(net4864),
    .X(_00177_));
 sg13g2_a21o_1 _11026_ (.A2(net4880),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B1(net4864),
    .X(_00178_));
 sg13g2_a21o_1 _11027_ (.A2(net4880),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B1(net4864),
    .X(_00179_));
 sg13g2_a21o_1 _11028_ (.A2(net4880),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B1(net4864),
    .X(_00180_));
 sg13g2_a21o_1 _11029_ (.A2(net4880),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B1(net4864),
    .X(_00182_));
 sg13g2_a21o_1 _11030_ (.A2(net4880),
    .A1(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B1(net4864),
    .X(_00183_));
 sg13g2_mux2_1 _11031_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .S(net4891),
    .X(_00138_));
 sg13g2_mux2_1 _11032_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .S(net4891),
    .X(_00149_));
 sg13g2_mux2_1 _11033_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .S(net4909),
    .X(_00152_));
 sg13g2_mux2_1 _11034_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .S(net4888),
    .X(_00153_));
 sg13g2_mux2_1 _11035_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .S(net4888),
    .X(_00154_));
 sg13g2_mux2_1 _11036_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .S(net4888),
    .X(_00155_));
 sg13g2_mux2_1 _11037_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .S(net4888),
    .X(_00156_));
 sg13g2_mux2_1 _11038_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .S(net4887),
    .X(_00157_));
 sg13g2_mux2_1 _11039_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .S(net4888),
    .X(_00158_));
 sg13g2_mux2_1 _11040_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .S(net4887),
    .X(_00128_));
 sg13g2_mux2_1 _11041_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .S(net4887),
    .X(_00129_));
 sg13g2_mux2_1 _11042_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .S(net4887),
    .X(_00130_));
 sg13g2_mux2_1 _11043_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .S(net4887),
    .X(_00131_));
 sg13g2_mux2_1 _11044_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .S(net4887),
    .X(_00132_));
 sg13g2_mux2_1 _11045_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .S(net4887),
    .X(_00133_));
 sg13g2_mux2_1 _11046_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .S(net4887),
    .X(_00134_));
 sg13g2_mux2_1 _11047_ (.A0(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .S(net4879),
    .X(_00135_));
 sg13g2_and2_2 _11048_ (.A(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .B(net4928),
    .X(_02526_));
 sg13g2_a21o_1 _11049_ (.A2(net4879),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B1(net4862),
    .X(_00136_));
 sg13g2_a21o_1 _11050_ (.A2(net4879),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B1(net4862),
    .X(_00137_));
 sg13g2_a21o_1 _11051_ (.A2(net4884),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B1(net4862),
    .X(_00139_));
 sg13g2_a21o_1 _11052_ (.A2(net4883),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .B1(net4862),
    .X(_00140_));
 sg13g2_a21o_1 _11053_ (.A2(net4883),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .B1(net4862),
    .X(_00141_));
 sg13g2_a21o_1 _11054_ (.A2(net4883),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B1(net4862),
    .X(_00142_));
 sg13g2_a21o_1 _11055_ (.A2(net4883),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B1(net4862),
    .X(_00143_));
 sg13g2_a21o_1 _11056_ (.A2(net4883),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B1(net4863),
    .X(_00144_));
 sg13g2_a21o_1 _11057_ (.A2(net4883),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B1(net4863),
    .X(_00145_));
 sg13g2_a21o_1 _11058_ (.A2(net4882),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B1(net4862),
    .X(_00146_));
 sg13g2_a21o_1 _11059_ (.A2(net4882),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B1(net4863),
    .X(_00147_));
 sg13g2_a21o_1 _11060_ (.A2(net4882),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B1(net4863),
    .X(_00148_));
 sg13g2_a21o_1 _11061_ (.A2(net4881),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B1(net4863),
    .X(_00150_));
 sg13g2_a21o_1 _11062_ (.A2(net4881),
    .A1(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B1(net4863),
    .X(_00151_));
 sg13g2_mux2_1 _11063_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .S(net4918),
    .X(_00106_));
 sg13g2_mux2_1 _11064_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .S(net4918),
    .X(_00117_));
 sg13g2_mux2_1 _11065_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .S(net4918),
    .X(_00120_));
 sg13g2_mux2_1 _11066_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .S(net4918),
    .X(_00121_));
 sg13g2_mux2_1 _11067_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .S(net4918),
    .X(_00122_));
 sg13g2_mux2_1 _11068_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .S(net4920),
    .X(_00123_));
 sg13g2_mux2_1 _11069_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .S(net4920),
    .X(_00124_));
 sg13g2_mux2_1 _11070_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .S(net4920),
    .X(_00125_));
 sg13g2_mux2_1 _11071_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .S(net4920),
    .X(_00126_));
 sg13g2_mux2_1 _11072_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .S(net4920),
    .X(_00096_));
 sg13g2_mux2_1 _11073_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .S(net4918),
    .X(_00097_));
 sg13g2_mux2_1 _11074_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .S(net4918),
    .X(_00098_));
 sg13g2_mux2_1 _11075_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .S(net4919),
    .X(_00099_));
 sg13g2_mux2_1 _11076_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .S(net4919),
    .X(_00100_));
 sg13g2_mux2_1 _11077_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .S(net4916),
    .X(_00101_));
 sg13g2_mux2_1 _11078_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .S(net4916),
    .X(_00102_));
 sg13g2_mux2_1 _11079_ (.A0(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .S(net4916),
    .X(_00103_));
 sg13g2_and2_1 _11080_ (.A(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .B(net4933),
    .X(_02527_));
 sg13g2_a21o_1 _11081_ (.A2(net4916),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B1(net4861),
    .X(_00104_));
 sg13g2_a21o_1 _11082_ (.A2(net4916),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B1(net4861),
    .X(_00105_));
 sg13g2_a21o_1 _11083_ (.A2(net4913),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B1(net4861),
    .X(_00107_));
 sg13g2_a21o_1 _11084_ (.A2(net4906),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .B1(net4860),
    .X(_00108_));
 sg13g2_a21o_1 _11085_ (.A2(net4903),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .B1(net4860),
    .X(_00109_));
 sg13g2_a21o_1 _11086_ (.A2(net4903),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B1(net4859),
    .X(_00110_));
 sg13g2_a21o_1 _11087_ (.A2(net4902),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B1(net4860),
    .X(_00111_));
 sg13g2_a21o_1 _11088_ (.A2(net4902),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B1(net4859),
    .X(_00112_));
 sg13g2_a21o_1 _11089_ (.A2(net4901),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B1(net4859),
    .X(_00113_));
 sg13g2_a21o_1 _11090_ (.A2(net4901),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B1(net4859),
    .X(_00114_));
 sg13g2_a21o_1 _11091_ (.A2(net4901),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B1(net4859),
    .X(_00115_));
 sg13g2_a21o_1 _11092_ (.A2(net4895),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B1(net4859),
    .X(_00116_));
 sg13g2_a21o_1 _11093_ (.A2(net4895),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B1(net4859),
    .X(_00118_));
 sg13g2_a21o_2 _11094_ (.A2(net4895),
    .A1(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B1(net4859),
    .X(_00119_));
 sg13g2_mux2_1 _11095_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .S(net4912),
    .X(_00074_));
 sg13g2_mux2_1 _11096_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .S(net4912),
    .X(_00085_));
 sg13g2_mux2_1 _11097_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .S(net4915),
    .X(_00088_));
 sg13g2_mux2_1 _11098_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .S(net4915),
    .X(_00089_));
 sg13g2_mux2_1 _11099_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .S(net4915),
    .X(_00090_));
 sg13g2_mux2_1 _11100_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .S(net4916),
    .X(_00091_));
 sg13g2_mux2_1 _11101_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .S(net4914),
    .X(_00092_));
 sg13g2_mux2_1 _11102_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .S(net4915),
    .X(_00093_));
 sg13g2_mux2_1 _11103_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .S(net4912),
    .X(_00094_));
 sg13g2_mux2_1 _11104_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .S(net4912),
    .X(_00064_));
 sg13g2_mux2_1 _11105_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .S(net4912),
    .X(_00065_));
 sg13g2_mux2_1 _11106_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .S(net4911),
    .X(_00066_));
 sg13g2_mux2_1 _11107_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .S(net4911),
    .X(_00067_));
 sg13g2_mux2_1 _11108_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .S(net4910),
    .X(_00068_));
 sg13g2_mux2_1 _11109_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .S(net4911),
    .X(_00069_));
 sg13g2_mux2_1 _11110_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .S(net4911),
    .X(_00070_));
 sg13g2_mux2_1 _11111_ (.A0(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .S(net4911),
    .X(_00071_));
 sg13g2_and2_1 _11112_ (.A(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .B(net4930),
    .X(_02528_));
 sg13g2_a21o_1 _11113_ (.A2(net4910),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B1(net4858),
    .X(_00072_));
 sg13g2_a21o_1 _11114_ (.A2(net4906),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B1(net4858),
    .X(_00073_));
 sg13g2_a21o_1 _11115_ (.A2(net4906),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B1(net4858),
    .X(_00075_));
 sg13g2_a21o_1 _11116_ (.A2(net4904),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .B1(net4858),
    .X(_00076_));
 sg13g2_a21o_1 _11117_ (.A2(net4903),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .B1(net4858),
    .X(_00077_));
 sg13g2_a21o_1 _11118_ (.A2(net4903),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B1(net4858),
    .X(_00078_));
 sg13g2_a21o_1 _11119_ (.A2(net4901),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B1(net4857),
    .X(_00079_));
 sg13g2_a21o_1 _11120_ (.A2(net4895),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B1(net4857),
    .X(_00080_));
 sg13g2_a21o_1 _11121_ (.A2(net4895),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B1(net4857),
    .X(_00081_));
 sg13g2_a21o_1 _11122_ (.A2(net4892),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B1(net4857),
    .X(_00082_));
 sg13g2_a21o_1 _11123_ (.A2(net4892),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B1(net4857),
    .X(_00083_));
 sg13g2_a21o_1 _11124_ (.A2(net4892),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B1(net4857),
    .X(_00084_));
 sg13g2_a21o_1 _11125_ (.A2(net4893),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B1(net4857),
    .X(_00086_));
 sg13g2_a21o_2 _11126_ (.A2(net4899),
    .A1(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B1(net4857),
    .X(_00087_));
 sg13g2_mux2_1 _11127_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .S(net4898),
    .X(_00042_));
 sg13g2_mux2_1 _11128_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .S(net4897),
    .X(_00053_));
 sg13g2_mux2_1 _11129_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .S(net4897),
    .X(_00056_));
 sg13g2_mux2_1 _11130_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .S(net4897),
    .X(_00057_));
 sg13g2_mux2_1 _11131_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .S(net4899),
    .X(_00058_));
 sg13g2_mux2_1 _11132_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .S(net4899),
    .X(_00059_));
 sg13g2_mux2_1 _11133_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .S(net4899),
    .X(_00060_));
 sg13g2_mux2_1 _11134_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .S(net4899),
    .X(_00061_));
 sg13g2_mux2_1 _11135_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .S(net4893),
    .X(_00062_));
 sg13g2_mux2_1 _11136_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .S(net4893),
    .X(_00032_));
 sg13g2_mux2_1 _11137_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .S(net4893),
    .X(_00033_));
 sg13g2_mux2_1 _11138_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .S(net4894),
    .X(_00034_));
 sg13g2_mux2_1 _11139_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .S(net4893),
    .X(_00035_));
 sg13g2_mux2_1 _11140_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .S(net4894),
    .X(_00036_));
 sg13g2_mux2_1 _11141_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .S(net4894),
    .X(_00037_));
 sg13g2_mux2_1 _11142_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .S(net4893),
    .X(_00038_));
 sg13g2_mux2_2 _11143_ (.A0(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .S(net4899),
    .X(_00039_));
 sg13g2_and2_1 _11144_ (.A(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .B(net4928),
    .X(_02529_));
 sg13g2_a21o_1 _11145_ (.A2(net4891),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B1(net4856),
    .X(_00040_));
 sg13g2_a21o_1 _11146_ (.A2(net4891),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B1(net4856),
    .X(_00041_));
 sg13g2_a21o_1 _11147_ (.A2(net4891),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B1(net4856),
    .X(_00043_));
 sg13g2_a21o_1 _11148_ (.A2(net4884),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .B1(net4855),
    .X(_00044_));
 sg13g2_a21o_1 _11149_ (.A2(net4884),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .B1(net4855),
    .X(_00045_));
 sg13g2_a21o_1 _11150_ (.A2(net4884),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B1(net4855),
    .X(_00046_));
 sg13g2_a21o_1 _11151_ (.A2(net4884),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B1(net4855),
    .X(_00047_));
 sg13g2_a21o_1 _11152_ (.A2(net4884),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B1(net4855),
    .X(_00048_));
 sg13g2_a21o_1 _11153_ (.A2(net4884),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B1(net4855),
    .X(_00049_));
 sg13g2_a21o_1 _11154_ (.A2(net4885),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B1(net4855),
    .X(_00050_));
 sg13g2_a21o_1 _11155_ (.A2(net4885),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B1(net4855),
    .X(_00051_));
 sg13g2_a21o_1 _11156_ (.A2(net4885),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B1(net4856),
    .X(_00052_));
 sg13g2_a21o_1 _11157_ (.A2(net4885),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B1(net4856),
    .X(_00054_));
 sg13g2_a21o_1 _11158_ (.A2(net4884),
    .A1(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B1(net4856),
    .X(_00055_));
 sg13g2_mux2_1 _11159_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .S(net4893),
    .X(_00010_));
 sg13g2_mux2_1 _11160_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .S(net4893),
    .X(_00021_));
 sg13g2_mux2_1 _11161_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .S(net4890),
    .X(_00024_));
 sg13g2_mux2_1 _11162_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .S(net4890),
    .X(_00025_));
 sg13g2_mux2_1 _11163_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .S(net4892),
    .X(_00026_));
 sg13g2_mux2_1 _11164_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .S(net4892),
    .X(_00027_));
 sg13g2_mux2_1 _11165_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .S(net4892),
    .X(_00028_));
 sg13g2_mux2_1 _11166_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .S(net4892),
    .X(_00029_));
 sg13g2_mux2_1 _11167_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .S(net4894),
    .X(_00030_));
 sg13g2_mux2_1 _11168_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .S(net4895),
    .X(_00000_));
 sg13g2_mux2_1 _11169_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .S(net4895),
    .X(_00001_));
 sg13g2_mux2_1 _11170_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .S(net4896),
    .X(_00002_));
 sg13g2_mux2_1 _11171_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .S(net4896),
    .X(_00003_));
 sg13g2_mux2_1 _11172_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .S(net4902),
    .X(_00004_));
 sg13g2_mux2_1 _11173_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .S(net4896),
    .X(_00005_));
 sg13g2_mux2_1 _11174_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .S(net4896),
    .X(_00006_));
 sg13g2_mux2_1 _11175_ (.A0(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .S(net4895),
    .X(_00007_));
 sg13g2_and2_1 _11176_ (.A(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .B(net4928),
    .X(_02530_));
 sg13g2_a21o_1 _11177_ (.A2(net4892),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B1(net4854),
    .X(_00008_));
 sg13g2_a21o_1 _11178_ (.A2(net4890),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B1(net4854),
    .X(_00009_));
 sg13g2_a21o_1 _11179_ (.A2(net4889),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B1(net4854),
    .X(_00011_));
 sg13g2_a21o_1 _11180_ (.A2(net4889),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .B1(net4854),
    .X(_00012_));
 sg13g2_a21o_1 _11181_ (.A2(net4879),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .B1(net4854),
    .X(_00013_));
 sg13g2_a21o_1 _11182_ (.A2(net4879),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B1(net4854),
    .X(_00014_));
 sg13g2_a21o_1 _11183_ (.A2(net4878),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B1(net4853),
    .X(_00015_));
 sg13g2_a21o_1 _11184_ (.A2(net4878),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B1(net4853),
    .X(_00016_));
 sg13g2_a21o_1 _11185_ (.A2(net4878),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B1(net4853),
    .X(_00017_));
 sg13g2_a21o_1 _11186_ (.A2(net4878),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B1(net4853),
    .X(_00018_));
 sg13g2_a21o_1 _11187_ (.A2(net4878),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B1(net4853),
    .X(_00019_));
 sg13g2_a21o_1 _11188_ (.A2(net4878),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B1(net4853),
    .X(_00020_));
 sg13g2_a21o_1 _11189_ (.A2(net4878),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B1(net4853),
    .X(_00022_));
 sg13g2_a21o_2 _11190_ (.A2(net4878),
    .A1(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B1(net4853),
    .X(_00023_));
 sg13g2_nor2_2 _11191_ (.A(net4989),
    .B(net4996),
    .Y(_02531_));
 sg13g2_nand2b_2 _11192_ (.Y(_02532_),
    .B(_02531_),
    .A_N(net5002));
 sg13g2_nor2b_2 _11193_ (.A(net5001),
    .B_N(net5004),
    .Y(_02533_));
 sg13g2_nand2b_2 _11194_ (.Y(_02534_),
    .B(net5005),
    .A_N(net5002));
 sg13g2_nor2_1 _11195_ (.A(_02334_),
    .B(_02532_),
    .Y(_02535_));
 sg13g2_nand2_2 _11196_ (.Y(_02536_),
    .A(_02531_),
    .B(_02533_));
 sg13g2_nand2b_2 _11197_ (.Y(_02537_),
    .B(net5003),
    .A_N(net5006));
 sg13g2_nor2b_1 _11198_ (.A(net5009),
    .B_N(net5001),
    .Y(_02538_));
 sg13g2_nand2b_2 _11199_ (.Y(_02539_),
    .B(net5000),
    .A_N(net5008));
 sg13g2_and2_1 _11200_ (.A(net5004),
    .B(net5009),
    .X(_02540_));
 sg13g2_nand2_1 _11201_ (.Y(_02541_),
    .A(net5007),
    .B(_02539_));
 sg13g2_xnor2_1 _11202_ (.Y(_02542_),
    .A(net5001),
    .B(net5004));
 sg13g2_xor2_1 _11203_ (.B(net5004),
    .A(net5001),
    .X(_02543_));
 sg13g2_nor3_1 _11204_ (.A(net4984),
    .B(_02540_),
    .C(_02543_),
    .Y(_02544_));
 sg13g2_nor2b_1 _11205_ (.A(net4997),
    .B_N(net5002),
    .Y(_02545_));
 sg13g2_nand2_1 _11206_ (.Y(_02546_),
    .A(net4984),
    .B(net5002));
 sg13g2_o21ai_1 _11207_ (.B1(net4993),
    .Y(_02547_),
    .A1(_02544_),
    .A2(_02545_));
 sg13g2_and2_2 _11208_ (.A(_02536_),
    .B(_02547_),
    .X(_02548_));
 sg13g2_nand2_1 _11209_ (.Y(_02549_),
    .A(_02536_),
    .B(_02547_));
 sg13g2_or2_2 _11210_ (.X(_02550_),
    .B(net5005),
    .A(net5001));
 sg13g2_nand2b_2 _11211_ (.Y(_02551_),
    .B(net5010),
    .A_N(net5003));
 sg13g2_nand2_1 _11212_ (.Y(_02552_),
    .A(_02335_),
    .B(_02534_));
 sg13g2_o21ai_1 _11213_ (.B1(_02551_),
    .Y(_02553_),
    .A1(net5009),
    .A2(_02533_));
 sg13g2_nand2_1 _11214_ (.Y(_02554_),
    .A(_02550_),
    .B(_02553_));
 sg13g2_a21o_1 _11215_ (.A2(_02553_),
    .A1(_02550_),
    .B1(net4984),
    .X(_02555_));
 sg13g2_nand2b_2 _11216_ (.Y(_02556_),
    .B(net5006),
    .A_N(net4996));
 sg13g2_and2_1 _11217_ (.A(net4985),
    .B(_02550_),
    .X(_02557_));
 sg13g2_a221oi_1 _11218_ (.B2(net4999),
    .C1(_02557_),
    .B1(_02554_),
    .A1(_02536_),
    .Y(_02558_),
    .A2(_02547_));
 sg13g2_nand4_1 _11219_ (.B(_02549_),
    .C(_02555_),
    .A(_02546_),
    .Y(_02559_),
    .D(_02556_));
 sg13g2_nor2_1 _11220_ (.A(net5004),
    .B(_02551_),
    .Y(_02560_));
 sg13g2_nand2b_2 _11221_ (.Y(_02561_),
    .B(net4996),
    .A_N(net4989));
 sg13g2_and2_1 _11222_ (.A(net5001),
    .B(net5009),
    .X(_02562_));
 sg13g2_nand2_1 _11223_ (.Y(_02563_),
    .A(net5000),
    .B(net5008));
 sg13g2_nand2b_1 _11224_ (.Y(_02564_),
    .B(net5008),
    .A_N(net5007));
 sg13g2_nor3_1 _11225_ (.A(_02538_),
    .B(_02560_),
    .C(_02561_),
    .Y(_02565_));
 sg13g2_nor2_2 _11226_ (.A(net4997),
    .B(net5005),
    .Y(_02566_));
 sg13g2_and2_1 _11227_ (.A(net4984),
    .B(_02551_),
    .X(_02567_));
 sg13g2_nor2_2 _11228_ (.A(net4996),
    .B(net5008),
    .Y(_02568_));
 sg13g2_nand2_1 _11229_ (.Y(_02569_),
    .A(net4984),
    .B(_02534_));
 sg13g2_o21ai_1 _11230_ (.B1(net4984),
    .Y(_02570_),
    .A1(_02335_),
    .A2(_02534_));
 sg13g2_nand3_1 _11231_ (.B(_02537_),
    .C(_02563_),
    .A(net4996),
    .Y(_02571_));
 sg13g2_nand2_1 _11232_ (.Y(_02572_),
    .A(_02570_),
    .B(_02571_));
 sg13g2_a221oi_1 _11233_ (.B2(net4991),
    .C1(_02565_),
    .B1(_02572_),
    .A1(_02531_),
    .Y(_02573_),
    .A2(_02543_));
 sg13g2_nand3_1 _11234_ (.B(_02334_),
    .C(_02551_),
    .A(net4997),
    .Y(_02574_));
 sg13g2_and2_1 _11235_ (.A(net4988),
    .B(_02574_),
    .X(_02575_));
 sg13g2_nand3b_1 _11236_ (.B(net5004),
    .C(net5009),
    .Y(_02576_),
    .A_N(net4998));
 sg13g2_nand2_1 _11237_ (.Y(_02577_),
    .A(net4995),
    .B(net5000));
 sg13g2_o21ai_1 _11238_ (.B1(_02576_),
    .Y(_02578_),
    .A1(_02533_),
    .A2(_02545_));
 sg13g2_and3_1 _11239_ (.X(_02579_),
    .A(net4990),
    .B(_02574_),
    .C(_02578_));
 sg13g2_nand2b_1 _11240_ (.Y(_02580_),
    .B(_02539_),
    .A_N(_02574_));
 sg13g2_nand2_1 _11241_ (.Y(_02581_),
    .A(net5000),
    .B(net5007));
 sg13g2_o21ai_1 _11242_ (.B1(net5002),
    .Y(_02582_),
    .A1(net5004),
    .A2(net5009));
 sg13g2_nor2_1 _11243_ (.A(_02542_),
    .B(_02562_),
    .Y(_02583_));
 sg13g2_a21oi_1 _11244_ (.A1(_02574_),
    .A2(_02583_),
    .Y(_02584_),
    .B1(net4990));
 sg13g2_a22oi_1 _11245_ (.Y(_02585_),
    .B1(_02580_),
    .B2(_02584_),
    .A2(_02578_),
    .A1(_02575_));
 sg13g2_a21o_2 _11246_ (.A2(_02584_),
    .A1(_02580_),
    .B1(_02579_),
    .X(_02586_));
 sg13g2_nand2b_1 _11247_ (.Y(_02587_),
    .B(net4999),
    .A_N(net5002));
 sg13g2_o21ai_1 _11248_ (.B1(_02587_),
    .Y(_02588_),
    .A1(net4999),
    .A2(_02533_));
 sg13g2_nand3_1 _11249_ (.B(_02552_),
    .C(_02588_),
    .A(net4993),
    .Y(_02589_));
 sg13g2_nand3_1 _11250_ (.B(_02534_),
    .C(_02564_),
    .A(net4995),
    .Y(_02590_));
 sg13g2_nand2_1 _11251_ (.Y(_02591_),
    .A(_02537_),
    .B(_02568_));
 sg13g2_nand3_1 _11252_ (.B(_02590_),
    .C(_02591_),
    .A(net4986),
    .Y(_02592_));
 sg13g2_and2_1 _11253_ (.A(_02589_),
    .B(_02592_),
    .X(_02593_));
 sg13g2_nand2_2 _11254_ (.Y(_02594_),
    .A(_02589_),
    .B(_02592_));
 sg13g2_and3_2 _11255_ (.X(_02595_),
    .A(_02573_),
    .B(_02586_),
    .C(_02594_));
 sg13g2_nand2_1 _11256_ (.Y(_02596_),
    .A(net4985),
    .B(_02542_));
 sg13g2_a22oi_1 _11257_ (.Y(_02597_),
    .B1(_02568_),
    .B2(_02537_),
    .A2(_02542_),
    .A1(net4984));
 sg13g2_a21oi_1 _11258_ (.A1(_02587_),
    .A2(_02597_),
    .Y(_02598_),
    .B1(net4987));
 sg13g2_nor4_1 _11259_ (.A(net4990),
    .B(net4998),
    .C(_02540_),
    .D(_02542_),
    .Y(_02599_));
 sg13g2_nor3_2 _11260_ (.A(_02565_),
    .B(_02598_),
    .C(_02599_),
    .Y(_02600_));
 sg13g2_nor3_2 _11261_ (.A(_02585_),
    .B(_02594_),
    .C(_02600_),
    .Y(_02601_));
 sg13g2_nor3_2 _11262_ (.A(_02586_),
    .B(_02593_),
    .C(_02600_),
    .Y(_02602_));
 sg13g2_a21o_1 _11263_ (.A2(_02564_),
    .A1(net4986),
    .B1(_02531_),
    .X(_02603_));
 sg13g2_nand2_1 _11264_ (.Y(_02604_),
    .A(_02596_),
    .B(_02603_));
 sg13g2_nand3_1 _11265_ (.B(net5007),
    .C(_02539_),
    .A(net4995),
    .Y(_02605_));
 sg13g2_and4_1 _11266_ (.A(net4988),
    .B(_02556_),
    .C(_02574_),
    .D(_02605_),
    .X(_02606_));
 sg13g2_nand4_1 _11267_ (.B(_02556_),
    .C(_02574_),
    .A(net4988),
    .Y(_02607_),
    .D(_02605_));
 sg13g2_and2_1 _11268_ (.A(_02604_),
    .B(_02607_),
    .X(_02608_));
 sg13g2_nand2_2 _11269_ (.Y(_02609_),
    .A(_02604_),
    .B(_02607_));
 sg13g2_or2_1 _11270_ (.X(_02610_),
    .B(_02582_),
    .A(_02540_));
 sg13g2_a21oi_2 _11271_ (.B1(net4987),
    .Y(_02611_),
    .A2(_02610_),
    .A1(_02557_));
 sg13g2_nand2_1 _11272_ (.Y(_02612_),
    .A(_02551_),
    .B(_02581_));
 sg13g2_a221oi_1 _11273_ (.B2(net4997),
    .C1(net4987),
    .B1(_02612_),
    .A1(_02557_),
    .Y(_02613_),
    .A2(_02610_));
 sg13g2_nor2_1 _11274_ (.A(_02564_),
    .B(_02577_),
    .Y(_02614_));
 sg13g2_nor4_2 _11275_ (.A(net4988),
    .B(_02566_),
    .C(_02568_),
    .Y(_02615_),
    .D(_02614_));
 sg13g2_nor2_1 _11276_ (.A(_02613_),
    .B(_02615_),
    .Y(_02616_));
 sg13g2_or2_2 _11277_ (.X(_02617_),
    .B(_02615_),
    .A(_02613_));
 sg13g2_a21oi_1 _11278_ (.A1(net5000),
    .A2(net5008),
    .Y(_02618_),
    .B1(net4995));
 sg13g2_a21o_1 _11279_ (.A2(_02537_),
    .A1(net4995),
    .B1(_02618_),
    .X(_02619_));
 sg13g2_or3_2 _11280_ (.A(net5002),
    .B(net5006),
    .C(net5008),
    .X(_02620_));
 sg13g2_a22oi_1 _11281_ (.Y(_02621_),
    .B1(_02618_),
    .B2(_02620_),
    .A2(_02537_),
    .A1(net4995));
 sg13g2_nor2_2 _11282_ (.A(net4986),
    .B(_02621_),
    .Y(_02622_));
 sg13g2_nand2b_1 _11283_ (.Y(_02623_),
    .B(net4988),
    .A_N(_02621_));
 sg13g2_nor2b_1 _11284_ (.A(net5008),
    .B_N(net5007),
    .Y(_02624_));
 sg13g2_nand2_1 _11285_ (.Y(_02625_),
    .A(_02335_),
    .B(_02550_));
 sg13g2_nand2_1 _11286_ (.Y(_02626_),
    .A(net5010),
    .B(_02534_));
 sg13g2_nor3_1 _11287_ (.A(_02335_),
    .B(_02533_),
    .C(_02561_),
    .Y(_02627_));
 sg13g2_a21oi_1 _11288_ (.A1(_02531_),
    .A2(_02625_),
    .Y(_02628_),
    .B1(_02627_));
 sg13g2_a21o_1 _11289_ (.A2(_02625_),
    .A1(_02531_),
    .B1(_02627_),
    .X(_02629_));
 sg13g2_nor2_1 _11290_ (.A(_02622_),
    .B(_02629_),
    .Y(_02630_));
 sg13g2_and4_1 _11291_ (.A(net4990),
    .B(net4997),
    .C(net5001),
    .D(_02334_),
    .X(_02631_));
 sg13g2_nand3_1 _11292_ (.B(net5004),
    .C(net5009),
    .A(net5001),
    .Y(_02632_));
 sg13g2_a21o_1 _11293_ (.A2(_02632_),
    .A1(net4998),
    .B1(net4990),
    .X(_02633_));
 sg13g2_a21oi_2 _11294_ (.B1(net4990),
    .Y(_02634_),
    .A2(_02632_),
    .A1(net4998));
 sg13g2_nand2_1 _11295_ (.Y(_02635_),
    .A(_02569_),
    .B(_02634_));
 sg13g2_nand2_1 _11296_ (.Y(_02636_),
    .A(net4999),
    .B(_02550_));
 sg13g2_o21ai_1 _11297_ (.B1(_02550_),
    .Y(_02637_),
    .A1(net4999),
    .A2(_02582_));
 sg13g2_nand2_1 _11298_ (.Y(_02638_),
    .A(net4992),
    .B(_02637_));
 sg13g2_a22oi_1 _11299_ (.Y(_02639_),
    .B1(_02637_),
    .B2(net4993),
    .A2(_02634_),
    .A1(_02569_));
 sg13g2_nor2b_1 _11300_ (.A(_02624_),
    .B_N(_02531_),
    .Y(_02640_));
 sg13g2_xor2_1 _11301_ (.B(net5008),
    .A(net5000),
    .X(_02641_));
 sg13g2_nand2_1 _11302_ (.Y(_02642_),
    .A(net4992),
    .B(_02566_));
 sg13g2_nand3_1 _11303_ (.B(_02566_),
    .C(_02641_),
    .A(net4989),
    .Y(_02643_));
 sg13g2_a21oi_2 _11304_ (.B1(_02640_),
    .Y(_02644_),
    .A2(_02643_),
    .A1(_02633_));
 sg13g2_o21ai_1 _11305_ (.B1(net4999),
    .Y(_02645_),
    .A1(_02334_),
    .A2(_02562_));
 sg13g2_and3_1 _11306_ (.X(_02646_),
    .A(net4993),
    .B(_02597_),
    .C(_02645_));
 sg13g2_nand3_1 _11307_ (.B(_02597_),
    .C(_02645_),
    .A(net4992),
    .Y(_02647_));
 sg13g2_and3_1 _11308_ (.X(_02648_),
    .A(net4987),
    .B(_02626_),
    .C(_02636_));
 sg13g2_nand3_1 _11309_ (.B(_02626_),
    .C(_02636_),
    .A(net4986),
    .Y(_02649_));
 sg13g2_a21oi_1 _11310_ (.A1(_02647_),
    .A2(_02649_),
    .Y(_02650_),
    .B1(_02644_));
 sg13g2_a221oi_1 _11311_ (.B2(_02649_),
    .C1(_02644_),
    .B1(_02647_),
    .A1(_02635_),
    .Y(_02651_),
    .A2(_02638_));
 sg13g2_and2_1 _11312_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][0] ),
    .B(net4814),
    .X(_02652_));
 sg13g2_and3_1 _11313_ (.X(_02653_),
    .A(_02573_),
    .B(_02586_),
    .C(_02593_));
 sg13g2_nor3_2 _11314_ (.A(_02585_),
    .B(_02593_),
    .C(_02600_),
    .Y(_02654_));
 sg13g2_nand3_1 _11315_ (.B(_02556_),
    .C(_02587_),
    .A(net4992),
    .Y(_02655_));
 sg13g2_nand2_1 _11316_ (.Y(_02656_),
    .A(_02531_),
    .B(_02582_));
 sg13g2_and2_1 _11317_ (.A(_02655_),
    .B(_02656_),
    .X(_02657_));
 sg13g2_nand2_1 _11318_ (.Y(_02658_),
    .A(_02655_),
    .B(_02656_));
 sg13g2_nor2_1 _11319_ (.A(_02540_),
    .B(_02561_),
    .Y(_02659_));
 sg13g2_nor4_1 _11320_ (.A(net4990),
    .B(net4998),
    .C(_02533_),
    .D(_02538_),
    .Y(_02660_));
 sg13g2_a21o_2 _11321_ (.A2(_02659_),
    .A1(_02552_),
    .B1(_02660_),
    .X(_02661_));
 sg13g2_or2_1 _11322_ (.X(_02662_),
    .B(_02661_),
    .A(_02611_));
 sg13g2_nor3_1 _11323_ (.A(_02611_),
    .B(_02657_),
    .C(_02661_),
    .Y(_02663_));
 sg13g2_a21o_1 _11324_ (.A2(_02620_),
    .A1(_02582_),
    .B1(net4997),
    .X(_02664_));
 sg13g2_a21o_1 _11325_ (.A2(_02664_),
    .A1(_02645_),
    .B1(net4986),
    .X(_02665_));
 sg13g2_and2_2 _11326_ (.A(_02532_),
    .B(_02665_),
    .X(_02666_));
 sg13g2_nor4_2 _11327_ (.A(_02547_),
    .B(_02611_),
    .C(_02657_),
    .Y(_02667_),
    .D(_02661_));
 sg13g2_nor3_2 _11328_ (.A(_02586_),
    .B(_02594_),
    .C(_02600_),
    .Y(_02668_));
 sg13g2_nand2_1 _11329_ (.Y(_02669_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][0] ),
    .B(net4751));
 sg13g2_a221oi_1 _11330_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][0] ),
    .C1(_02652_),
    .B1(net4876),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][0] ),
    .Y(_02670_),
    .A2(net4760));
 sg13g2_a22oi_1 _11331_ (.Y(_02671_),
    .B1(net4801),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][0] ),
    .A2(net4754),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][0] ));
 sg13g2_a22oi_1 _11332_ (.Y(_02672_),
    .B1(net4763),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][0] ),
    .A2(net4766),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][0] ));
 sg13g2_a21oi_1 _11333_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][0] ),
    .A2(net4757),
    .Y(_02673_),
    .B1(net4823));
 sg13g2_and4_1 _11334_ (.A(_02669_),
    .B(_02671_),
    .C(_02672_),
    .D(_02673_),
    .X(_02674_));
 sg13g2_a22oi_1 _11335_ (.Y(_02675_),
    .B1(_02670_),
    .B2(_02674_),
    .A2(net4823),
    .A1(_02338_));
 sg13g2_nand2_1 _11336_ (.Y(_02676_),
    .A(_00290_),
    .B(net4822));
 sg13g2_and3_1 _11337_ (.X(_02677_),
    .A(_02547_),
    .B(_02635_),
    .C(_02642_));
 sg13g2_and2_1 _11338_ (.A(_02650_),
    .B(_02677_),
    .X(_02678_));
 sg13g2_nand3_1 _11339_ (.B(_02650_),
    .C(_02677_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][0] ),
    .Y(_02679_));
 sg13g2_nand2_1 _11340_ (.Y(_02680_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][0] ),
    .B(net4813));
 sg13g2_nor3_1 _11341_ (.A(_02644_),
    .B(_02646_),
    .C(_02648_),
    .Y(_02681_));
 sg13g2_and2_1 _11342_ (.A(_02677_),
    .B(_02681_),
    .X(_02682_));
 sg13g2_nand3_1 _11343_ (.B(_02677_),
    .C(_02681_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][0] ),
    .Y(_02683_));
 sg13g2_nor4_2 _11344_ (.A(_02639_),
    .B(_02644_),
    .C(_02646_),
    .Y(_02684_),
    .D(_02648_));
 sg13g2_nand2_1 _11345_ (.Y(_02685_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][0] ),
    .B(net4799));
 sg13g2_nand4_1 _11346_ (.B(_02680_),
    .C(_02683_),
    .A(_02679_),
    .Y(_02686_),
    .D(_02685_));
 sg13g2_nand2_1 _11347_ (.Y(_02687_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][0] ),
    .B(net4800));
 sg13g2_and4_2 _11348_ (.A(_02547_),
    .B(_02635_),
    .C(_02642_),
    .D(_02644_),
    .X(_02688_));
 sg13g2_nand2_1 _11349_ (.Y(_02689_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][0] ),
    .B(net4796));
 sg13g2_and3_2 _11350_ (.X(_02690_),
    .A(_02644_),
    .B(_02647_),
    .C(_02649_));
 sg13g2_nor2_1 _11351_ (.A(net5009),
    .B(_02536_),
    .Y(_02691_));
 sg13g2_a221oi_1 _11352_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][0] ),
    .C1(net4822),
    .B1(net4848),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][0] ),
    .Y(_02692_),
    .A2(net4793));
 sg13g2_nand3_1 _11353_ (.B(_02689_),
    .C(_02692_),
    .A(_02687_),
    .Y(_02693_));
 sg13g2_o21ai_1 _11354_ (.B1(_02676_),
    .Y(_02694_),
    .A1(_02686_),
    .A2(_02693_));
 sg13g2_a221oi_1 _11355_ (.B2(_02674_),
    .C1(_02694_),
    .B1(_02670_),
    .A1(_02338_),
    .Y(_02695_),
    .A2(net4823));
 sg13g2_xor2_1 _11356_ (.B(_02694_),
    .A(_02675_),
    .X(_02696_));
 sg13g2_a22oi_1 _11357_ (.Y(_02697_),
    .B1(_02665_),
    .B2(_02532_),
    .A2(_02547_),
    .A1(_02536_));
 sg13g2_and3_1 _11358_ (.X(_02698_),
    .A(_02657_),
    .B(_02662_),
    .C(_02697_));
 sg13g2_and3_1 _11359_ (.X(_02699_),
    .A(_02532_),
    .B(_02547_),
    .C(_02665_));
 sg13g2_and3_1 _11360_ (.X(_02700_),
    .A(_02657_),
    .B(_02662_),
    .C(_02699_));
 sg13g2_a22oi_1 _11361_ (.Y(_02701_),
    .B1(net4738),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][0] ),
    .A2(net4741),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][0] ));
 sg13g2_and3_1 _11362_ (.X(_02702_),
    .A(_02658_),
    .B(_02662_),
    .C(_02699_));
 sg13g2_and3_1 _11363_ (.X(_02703_),
    .A(_02658_),
    .B(_02662_),
    .C(_02697_));
 sg13g2_nor2_1 _11364_ (.A(net4984),
    .B(_02542_),
    .Y(_02704_));
 sg13g2_a21o_1 _11365_ (.A2(_02610_),
    .A1(_02567_),
    .B1(_02704_),
    .X(_02705_));
 sg13g2_nor3_1 _11366_ (.A(net4997),
    .B(_02540_),
    .C(_02543_),
    .Y(_02706_));
 sg13g2_and2_1 _11367_ (.A(_02556_),
    .B(_02562_),
    .X(_02707_));
 sg13g2_nor4_2 _11368_ (.A(net4992),
    .B(_02533_),
    .C(_02706_),
    .Y(_02708_),
    .D(_02707_));
 sg13g2_a21oi_2 _11369_ (.B1(_02708_),
    .Y(_02709_),
    .A2(_02705_),
    .A1(net4992));
 sg13g2_a21o_2 _11370_ (.A2(_02705_),
    .A1(net4992),
    .B1(_02708_),
    .X(_02710_));
 sg13g2_nand4_1 _11371_ (.B(_02546_),
    .C(_02555_),
    .A(net4986),
    .Y(_02711_),
    .D(_02556_));
 sg13g2_nor3_1 _11372_ (.A(_02334_),
    .B(_02562_),
    .C(_02568_),
    .Y(_02712_));
 sg13g2_o21ai_1 _11373_ (.B1(net4992),
    .Y(_02713_),
    .A1(_02566_),
    .A2(_02712_));
 sg13g2_nand2_2 _11374_ (.Y(_02714_),
    .A(_02711_),
    .B(_02713_));
 sg13g2_and4_1 _11375_ (.A(_02697_),
    .B(_02710_),
    .C(_02711_),
    .D(_02713_),
    .X(_02715_));
 sg13g2_and2_1 _11376_ (.A(_02663_),
    .B(_02699_),
    .X(_02716_));
 sg13g2_nor2_2 _11377_ (.A(_02549_),
    .B(_02666_),
    .Y(_02717_));
 sg13g2_nor3_1 _11378_ (.A(_02611_),
    .B(_02658_),
    .C(_02661_),
    .Y(_02718_));
 sg13g2_and2_1 _11379_ (.A(_02699_),
    .B(_02718_),
    .X(_02719_));
 sg13g2_a22oi_1 _11380_ (.Y(_02720_),
    .B1(net4735),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][0] ),
    .A2(net4807),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][0] ));
 sg13g2_and2_1 _11381_ (.A(_02701_),
    .B(_02720_),
    .X(_02721_));
 sg13g2_a22oi_1 _11382_ (.Y(_02722_),
    .B1(net4713),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][0] ),
    .A2(net4715),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][0] ));
 sg13g2_a22oi_1 _11383_ (.Y(_02723_),
    .B1(net4710),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][0] ),
    .A2(net4849),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][0] ));
 sg13g2_a22oi_1 _11384_ (.Y(_02724_),
    .B1(net4719),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][0] ),
    .A2(net4727),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][0] ));
 sg13g2_and4_1 _11385_ (.A(net4771),
    .B(_02722_),
    .C(_02723_),
    .D(_02724_),
    .X(_02725_));
 sg13g2_a22oi_1 _11386_ (.Y(_02726_),
    .B1(_02721_),
    .B2(_02725_),
    .A2(net4834),
    .A1(_00288_));
 sg13g2_nand2_1 _11387_ (.Y(_02727_),
    .A(_00289_),
    .B(net4835));
 sg13g2_nor3_1 _11388_ (.A(net4991),
    .B(net4996),
    .C(_02537_),
    .Y(_02728_));
 sg13g2_a21o_1 _11389_ (.A2(_02568_),
    .A1(net4990),
    .B1(_02728_),
    .X(_02729_));
 sg13g2_nor2_1 _11390_ (.A(_02561_),
    .B(_02620_),
    .Y(_02730_));
 sg13g2_a21oi_2 _11391_ (.B1(_02730_),
    .Y(_02731_),
    .A2(_02729_),
    .A1(_02543_));
 sg13g2_nand2b_1 _11392_ (.Y(_02732_),
    .B(_02548_),
    .A_N(_02731_));
 sg13g2_nor3_2 _11393_ (.A(_02710_),
    .B(net4726),
    .C(_02732_),
    .Y(_02733_));
 sg13g2_nor4_2 _11394_ (.A(_02548_),
    .B(_02666_),
    .C(_02710_),
    .Y(_02734_),
    .D(net4726));
 sg13g2_nor3_2 _11395_ (.A(_02709_),
    .B(_02714_),
    .C(_02732_),
    .Y(_02735_));
 sg13g2_and2_1 _11396_ (.A(_02548_),
    .B(_02731_),
    .X(_02736_));
 sg13g2_nand2_2 _11397_ (.Y(_02737_),
    .A(_02548_),
    .B(_02731_));
 sg13g2_nor3_2 _11398_ (.A(_02710_),
    .B(net4726),
    .C(_02737_),
    .Y(_02738_));
 sg13g2_nor4_1 _11399_ (.A(_02337_),
    .B(_02710_),
    .C(net4726),
    .D(_02737_),
    .Y(_02739_));
 sg13g2_a221oi_1 _11400_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][0] ),
    .C1(net4834),
    .B1(net4729),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][0] ),
    .Y(_02740_),
    .A2(net4808));
 sg13g2_and2_1 _11401_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][0] ),
    .B(net4721),
    .X(_02741_));
 sg13g2_nor3_2 _11402_ (.A(_02709_),
    .B(net4726),
    .C(_02737_),
    .Y(_02742_));
 sg13g2_nor4_1 _11403_ (.A(_02336_),
    .B(_02709_),
    .C(net4726),
    .D(_02737_),
    .Y(_02743_));
 sg13g2_and3_2 _11404_ (.X(_02744_),
    .A(_02709_),
    .B(_02714_),
    .C(_02736_));
 sg13g2_and4_1 _11405_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][0] ),
    .B(_02709_),
    .C(net4726),
    .D(_02736_),
    .X(_02745_));
 sg13g2_and3_2 _11406_ (.X(_02746_),
    .A(_02710_),
    .B(net4726),
    .C(_02736_));
 sg13g2_nor4_1 _11407_ (.A(_02739_),
    .B(_02741_),
    .C(_02743_),
    .D(_02745_),
    .Y(_02747_));
 sg13g2_a22oi_1 _11408_ (.Y(_02748_),
    .B1(net4659),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][0] ),
    .A2(net4663),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][0] ));
 sg13g2_a22oi_1 _11409_ (.Y(_02749_),
    .B1(net4650),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][0] ),
    .A2(net4665),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][0] ));
 sg13g2_nand4_1 _11410_ (.B(_02747_),
    .C(_02748_),
    .A(_02740_),
    .Y(_02750_),
    .D(_02749_));
 sg13g2_and3_2 _11411_ (.X(_02751_),
    .A(_02726_),
    .B(_02727_),
    .C(_02750_));
 sg13g2_a21oi_2 _11412_ (.B1(_02726_),
    .Y(_02752_),
    .A2(_02750_),
    .A1(_02727_));
 sg13g2_nor3_2 _11413_ (.A(_02696_),
    .B(_02751_),
    .C(_02752_),
    .Y(_02753_));
 sg13g2_o21ai_1 _11414_ (.B1(_02696_),
    .Y(_02754_),
    .A1(_02751_),
    .A2(_02752_));
 sg13g2_nand2b_1 _11415_ (.Y(_02755_),
    .B(_02754_),
    .A_N(_02753_));
 sg13g2_nor2_1 _11416_ (.A(_02556_),
    .B(_02563_),
    .Y(_02756_));
 sg13g2_nor2b_1 _11417_ (.A(_02756_),
    .B_N(_02603_),
    .Y(_02757_));
 sg13g2_nand2b_1 _11418_ (.Y(_02758_),
    .B(_02603_),
    .A_N(_02756_));
 sg13g2_a21oi_1 _11419_ (.A1(_02577_),
    .A2(_02624_),
    .Y(_02759_),
    .B1(net4986));
 sg13g2_and2_1 _11420_ (.A(_02619_),
    .B(_02759_),
    .X(_02760_));
 sg13g2_nand2_1 _11421_ (.Y(_02761_),
    .A(_02619_),
    .B(_02759_));
 sg13g2_mux2_1 _11422_ (.A0(_02539_),
    .A1(_02551_),
    .S(net4995),
    .X(_02762_));
 sg13g2_a21oi_2 _11423_ (.B1(net4988),
    .Y(_02763_),
    .A2(_02539_),
    .A1(net5007));
 sg13g2_nand2_1 _11424_ (.Y(_02764_),
    .A(_02762_),
    .B(_02763_));
 sg13g2_a22oi_1 _11425_ (.Y(_02765_),
    .B1(_02762_),
    .B2(_02763_),
    .A2(_02759_),
    .A1(_02619_));
 sg13g2_a21oi_1 _11426_ (.A1(net5000),
    .A2(net5007),
    .Y(_02766_),
    .B1(net4995));
 sg13g2_or3_1 _11427_ (.A(net4988),
    .B(_02625_),
    .C(_02766_),
    .X(_02767_));
 sg13g2_nand2b_1 _11428_ (.Y(_02768_),
    .B(net4985),
    .A_N(_02581_));
 sg13g2_nand3_1 _11429_ (.B(_02574_),
    .C(_02768_),
    .A(net5),
    .Y(_02769_));
 sg13g2_and4_2 _11430_ (.A(_02757_),
    .B(_02765_),
    .C(_02767_),
    .D(_02769_),
    .X(_02770_));
 sg13g2_nand2_1 _11431_ (.Y(_02771_),
    .A(_02758_),
    .B(_02769_));
 sg13g2_nand2b_1 _11432_ (.Y(_02772_),
    .B(_02766_),
    .A_N(_02641_));
 sg13g2_a21o_1 _11433_ (.A2(_02772_),
    .A1(_02605_),
    .B1(net4986),
    .X(_02773_));
 sg13g2_and2_1 _11434_ (.A(_02767_),
    .B(_02773_),
    .X(_02774_));
 sg13g2_nand2_2 _11435_ (.Y(_02775_),
    .A(_02771_),
    .B(_02774_));
 sg13g2_nor2_1 _11436_ (.A(net4790),
    .B(_02775_),
    .Y(_02776_));
 sg13g2_nand3b_1 _11437_ (.B(_02771_),
    .C(_02774_),
    .Y(_02777_),
    .A_N(_02770_));
 sg13g2_or2_1 _11438_ (.X(_02778_),
    .B(_02777_),
    .A(_02340_));
 sg13g2_a221oi_1 _11439_ (.B2(_02773_),
    .C1(_02760_),
    .B1(_02767_),
    .A1(_02762_),
    .Y(_02779_),
    .A2(_02763_));
 sg13g2_a221oi_1 _11440_ (.B2(_02575_),
    .C1(_02757_),
    .B1(_02768_),
    .A1(_02761_),
    .Y(_02780_),
    .A2(_02764_));
 sg13g2_nor2_2 _11441_ (.A(_02765_),
    .B(_02774_),
    .Y(_02781_));
 sg13g2_a221oi_1 _11442_ (.B2(_02773_),
    .C1(_02339_),
    .B1(_02767_),
    .A1(_02761_),
    .Y(_02782_),
    .A2(_02764_));
 sg13g2_a221oi_1 _11443_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][0] ),
    .C1(_02782_),
    .B1(net4783),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][0] ),
    .Y(_02783_),
    .A2(_02779_));
 sg13g2_and4_1 _11444_ (.A(_02758_),
    .B(_02765_),
    .C(_02767_),
    .D(_02769_),
    .X(_02784_));
 sg13g2_a22oi_1 _11445_ (.Y(_02785_),
    .B1(net4779),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][0] ),
    .A2(_02770_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][0] ));
 sg13g2_nand3_1 _11446_ (.B(_02783_),
    .C(_02785_),
    .A(_02777_),
    .Y(_02786_));
 sg13g2_nand2_1 _11447_ (.Y(_02787_),
    .A(net5),
    .B(_02614_));
 sg13g2_mux2_1 _11448_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][0] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][0] ),
    .S(net4843),
    .X(_02788_));
 sg13g2_nand3_1 _11449_ (.B(_02786_),
    .C(_02788_),
    .A(_02778_),
    .Y(_02789_));
 sg13g2_a21o_1 _11450_ (.A2(_02786_),
    .A1(_02778_),
    .B1(_02788_),
    .X(_02790_));
 sg13g2_and2_2 _11451_ (.A(_02789_),
    .B(_02790_),
    .X(_02791_));
 sg13g2_a22oi_1 _11452_ (.Y(_02792_),
    .B1(_02623_),
    .B2(_02628_),
    .A2(_02607_),
    .A1(_02604_));
 sg13g2_and2_1 _11453_ (.A(net4819),
    .B(net4774),
    .X(_02793_));
 sg13g2_nand2_1 _11454_ (.Y(_02794_),
    .A(_00291_),
    .B(net4698));
 sg13g2_a221oi_1 _11455_ (.B2(_02628_),
    .C1(_02606_),
    .B1(_02623_),
    .A1(_02596_),
    .Y(_02795_),
    .A2(_02603_));
 sg13g2_and2_1 _11456_ (.A(net4820),
    .B(_02795_),
    .X(_02796_));
 sg13g2_nand3_1 _11457_ (.B(net4820),
    .C(_02795_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][0] ),
    .Y(_02797_));
 sg13g2_o21ai_1 _11458_ (.B1(net4775),
    .Y(_02798_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][0] ),
    .A2(net4820));
 sg13g2_and2_1 _11459_ (.A(_02617_),
    .B(_02795_),
    .X(_02799_));
 sg13g2_nand3_1 _11460_ (.B(_02617_),
    .C(_02795_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][0] ),
    .Y(_02800_));
 sg13g2_nand3_1 _11461_ (.B(_02798_),
    .C(_02800_),
    .A(_02797_),
    .Y(_02801_));
 sg13g2_nor4_2 _11462_ (.A(_02608_),
    .B(net4820),
    .C(_02622_),
    .Y(_02802_),
    .D(_02629_));
 sg13g2_nand4_1 _11463_ (.B(_02609_),
    .C(_02617_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][0] ),
    .Y(_02803_),
    .D(_02630_));
 sg13g2_nor4_2 _11464_ (.A(_02613_),
    .B(_02615_),
    .C(_02622_),
    .Y(_02804_),
    .D(_02629_));
 sg13g2_and2_1 _11465_ (.A(_02609_),
    .B(_02804_),
    .X(_02805_));
 sg13g2_nand3_1 _11466_ (.B(_02609_),
    .C(_02804_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][0] ),
    .Y(_02806_));
 sg13g2_and2_1 _11467_ (.A(_02608_),
    .B(_02804_),
    .X(_02807_));
 sg13g2_nand3_1 _11468_ (.B(_02608_),
    .C(_02804_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][0] ),
    .Y(_02808_));
 sg13g2_nand2_1 _11469_ (.Y(_02809_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][0] ),
    .B(net4873));
 sg13g2_nand4_1 _11470_ (.B(_02806_),
    .C(_02808_),
    .A(_02803_),
    .Y(_02810_),
    .D(_02809_));
 sg13g2_o21ai_1 _11471_ (.B1(_02794_),
    .Y(_02811_),
    .A1(_02801_),
    .A2(_02810_));
 sg13g2_nand2_1 _11472_ (.Y(_02812_),
    .A(_02570_),
    .B(_02634_));
 sg13g2_nand4_1 _11473_ (.B(_02541_),
    .C(_02574_),
    .A(net4988),
    .Y(_02813_),
    .D(_02591_));
 sg13g2_and2_1 _11474_ (.A(_02812_),
    .B(_02813_),
    .X(_02814_));
 sg13g2_nand2_2 _11475_ (.Y(_02815_),
    .A(_02812_),
    .B(_02813_));
 sg13g2_a21o_1 _11476_ (.A2(_02556_),
    .A1(_02553_),
    .B1(net4991),
    .X(_02816_));
 sg13g2_nand3b_1 _11477_ (.B(_02571_),
    .C(net4989),
    .Y(_02817_),
    .A_N(_02568_));
 sg13g2_a21o_2 _11478_ (.A2(_02817_),
    .A1(_02816_),
    .B1(net4848),
    .X(_02818_));
 sg13g2_a21oi_1 _11479_ (.A1(net4996),
    .A2(net5000),
    .Y(_02819_),
    .B1(net5010));
 sg13g2_and2_1 _11480_ (.A(_02568_),
    .B(_02581_),
    .X(_02820_));
 sg13g2_o21ai_1 _11481_ (.B1(net4989),
    .Y(_02821_),
    .A1(_02543_),
    .A2(_02819_));
 sg13g2_or2_1 _11482_ (.X(_02822_),
    .B(_02821_),
    .A(_02820_));
 sg13g2_and2_1 _11483_ (.A(_02561_),
    .B(_02822_),
    .X(_02823_));
 sg13g2_o21ai_1 _11484_ (.B1(_02561_),
    .Y(_02824_),
    .A1(_02820_),
    .A2(_02821_));
 sg13g2_nor3_1 _11485_ (.A(_02815_),
    .B(_02818_),
    .C(_02823_),
    .Y(_02825_));
 sg13g2_and2_1 _11486_ (.A(_02815_),
    .B(_02818_),
    .X(_02826_));
 sg13g2_nand2_2 _11487_ (.Y(_02827_),
    .A(_02815_),
    .B(_02818_));
 sg13g2_and2_1 _11488_ (.A(_02818_),
    .B(_02824_),
    .X(_02828_));
 sg13g2_nand3_1 _11489_ (.B(_02818_),
    .C(_02824_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][0] ),
    .Y(_02829_));
 sg13g2_a221oi_1 _11490_ (.B2(_02817_),
    .C1(_02824_),
    .B1(_02816_),
    .A1(_02335_),
    .Y(_02830_),
    .A2(net4852));
 sg13g2_and2_2 _11491_ (.A(_02814_),
    .B(_02830_),
    .X(_02831_));
 sg13g2_nand3_1 _11492_ (.B(_02814_),
    .C(_02830_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][0] ),
    .Y(_02832_));
 sg13g2_nor3_1 _11493_ (.A(_02814_),
    .B(_02818_),
    .C(_02823_),
    .Y(_02833_));
 sg13g2_and3_2 _11494_ (.X(_02834_),
    .A(_02814_),
    .B(_02818_),
    .C(_02823_));
 sg13g2_nand4_1 _11495_ (.B(_02814_),
    .C(_02818_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][0] ),
    .Y(_02835_),
    .D(_02823_));
 sg13g2_and2_2 _11496_ (.A(_02815_),
    .B(_02830_),
    .X(_02836_));
 sg13g2_and3_1 _11497_ (.X(_02837_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][0] ),
    .B(_02815_),
    .C(_02830_));
 sg13g2_a221oi_1 _11498_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][0] ),
    .C1(_02837_),
    .B1(net4672),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][0] ),
    .Y(_02838_),
    .A2(net4685));
 sg13g2_and4_1 _11499_ (.A(_02827_),
    .B(_02829_),
    .C(_02832_),
    .D(_02835_),
    .X(_02839_));
 sg13g2_and2_1 _11500_ (.A(_00292_),
    .B(net4681),
    .X(_02840_));
 sg13g2_a21o_2 _11501_ (.A2(_02839_),
    .A1(_02838_),
    .B1(_02840_),
    .X(_02841_));
 sg13g2_xor2_1 _11502_ (.B(_02841_),
    .A(_02811_),
    .X(_02842_));
 sg13g2_nand2_1 _11503_ (.Y(_02843_),
    .A(_02791_),
    .B(_02842_));
 sg13g2_xnor2_1 _11504_ (.Y(_02844_),
    .A(_02791_),
    .B(_02842_));
 sg13g2_inv_1 _11505_ (.Y(_02845_),
    .A(_02844_));
 sg13g2_nand3b_1 _11506_ (.B(_02754_),
    .C(_02845_),
    .Y(_02846_),
    .A_N(_02753_));
 sg13g2_nand3_1 _11507_ (.B(net4820),
    .C(_02795_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][1] ),
    .Y(_02847_));
 sg13g2_and2_2 _11508_ (.A(_02617_),
    .B(net4775),
    .X(_02848_));
 sg13g2_o21ai_1 _11509_ (.B1(net4775),
    .Y(_02849_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][1] ),
    .A2(net4820));
 sg13g2_nand3_1 _11510_ (.B(_02617_),
    .C(_02795_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][1] ),
    .Y(_02850_));
 sg13g2_nand3_1 _11511_ (.B(_02849_),
    .C(_02850_),
    .A(_02847_),
    .Y(_02851_));
 sg13g2_nand4_1 _11512_ (.B(_02609_),
    .C(_02617_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][1] ),
    .Y(_02852_),
    .D(_02630_));
 sg13g2_nand3_1 _11513_ (.B(_02608_),
    .C(_02804_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][1] ),
    .Y(_02853_));
 sg13g2_nand3_1 _11514_ (.B(_02609_),
    .C(_02804_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][1] ),
    .Y(_02854_));
 sg13g2_nand2_1 _11515_ (.Y(_02855_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][1] ),
    .B(net4873));
 sg13g2_nand4_1 _11516_ (.B(_02853_),
    .C(_02854_),
    .A(_02852_),
    .Y(_02856_),
    .D(_02855_));
 sg13g2_nand2_1 _11517_ (.Y(_02857_),
    .A(_00295_),
    .B(net4698));
 sg13g2_o21ai_1 _11518_ (.B1(_02857_),
    .Y(_02858_),
    .A1(_02851_),
    .A2(_02856_));
 sg13g2_nor3_1 _11519_ (.A(_02811_),
    .B(_02841_),
    .C(_02858_),
    .Y(_02859_));
 sg13g2_or3_1 _11520_ (.A(_02811_),
    .B(_02841_),
    .C(_02858_),
    .X(_02860_));
 sg13g2_o21ai_1 _11521_ (.B1(_02858_),
    .Y(_02861_),
    .A1(_02811_),
    .A2(_02841_));
 sg13g2_a221oi_1 _11522_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][1] ),
    .C1(net4681),
    .B1(net4670),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][1] ),
    .Y(_02862_),
    .A2(net4677));
 sg13g2_a22oi_1 _11523_ (.Y(_02863_),
    .B1(net4672),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][1] ),
    .A2(net4675),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][1] ));
 sg13g2_a22oi_1 _11524_ (.Y(_02864_),
    .B1(net4668),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][1] ),
    .A2(net4685),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][1] ));
 sg13g2_and2_1 _11525_ (.A(_02863_),
    .B(_02864_),
    .X(_02865_));
 sg13g2_a22oi_1 _11526_ (.Y(_02866_),
    .B1(_02862_),
    .B2(_02865_),
    .A2(net4681),
    .A1(_00296_));
 sg13g2_and3_1 _11527_ (.X(_02867_),
    .A(_02860_),
    .B(_02861_),
    .C(_02866_));
 sg13g2_a21oi_1 _11528_ (.A1(_02860_),
    .A2(_02861_),
    .Y(_02868_),
    .B1(_02866_));
 sg13g2_nor2_2 _11529_ (.A(_02867_),
    .B(_02868_),
    .Y(_02869_));
 sg13g2_mux2_1 _11530_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][1] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][1] ),
    .S(net4843),
    .X(_02870_));
 sg13g2_nand2b_1 _11531_ (.Y(_02871_),
    .B(_02870_),
    .A_N(_02789_));
 sg13g2_xor2_1 _11532_ (.B(_02870_),
    .A(_02789_),
    .X(_02872_));
 sg13g2_nand2_1 _11533_ (.Y(_02873_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][1] ),
    .B(net4702));
 sg13g2_a22oi_1 _11534_ (.Y(_02874_),
    .B1(net4781),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][1] ),
    .A2(net4785),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][1] ));
 sg13g2_a22oi_1 _11535_ (.Y(_02875_),
    .B1(net4777),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][1] ),
    .A2(net4788),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][1] ));
 sg13g2_nand4_1 _11536_ (.B(_02873_),
    .C(_02874_),
    .A(net4706),
    .Y(_02876_),
    .D(_02875_));
 sg13g2_o21ai_1 _11537_ (.B1(_02876_),
    .Y(_02877_),
    .A1(_02341_),
    .A2(net4706));
 sg13g2_xnor2_1 _11538_ (.Y(_02878_),
    .A(_02872_),
    .B(_02877_));
 sg13g2_nor2_1 _11539_ (.A(_02843_),
    .B(_02878_),
    .Y(_02879_));
 sg13g2_xor2_1 _11540_ (.B(_02878_),
    .A(_02843_),
    .X(_02880_));
 sg13g2_xnor2_1 _11541_ (.Y(_02881_),
    .A(_02869_),
    .B(_02880_));
 sg13g2_nor2_1 _11542_ (.A(_02846_),
    .B(_02881_),
    .Y(_02882_));
 sg13g2_xor2_1 _11543_ (.B(_02881_),
    .A(_02846_),
    .X(_02883_));
 sg13g2_a22oi_1 _11544_ (.Y(_02884_),
    .B1(net4665),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][1] ),
    .A2(net4722),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][1] ));
 sg13g2_a22oi_1 _11545_ (.Y(_02885_),
    .B1(net4659),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][1] ),
    .A2(net4663),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][1] ));
 sg13g2_and2_1 _11546_ (.A(_02884_),
    .B(_02885_),
    .X(_02886_));
 sg13g2_a221oi_1 _11547_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][1] ),
    .C1(net4836),
    .B1(net4730),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][1] ),
    .Y(_02887_),
    .A2(net4809));
 sg13g2_a22oi_1 _11548_ (.Y(_02888_),
    .B1(net4655),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][1] ),
    .A2(net4657),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][1] ));
 sg13g2_nand2_1 _11549_ (.Y(_02889_),
    .A(_02887_),
    .B(_02888_));
 sg13g2_a221oi_1 _11550_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][1] ),
    .C1(_02889_),
    .B1(net4650),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][1] ),
    .Y(_02890_),
    .A2(net4653));
 sg13g2_a22oi_1 _11551_ (.Y(_02891_),
    .B1(_02886_),
    .B2(_02890_),
    .A2(net4836),
    .A1(_00300_));
 sg13g2_a22oi_1 _11552_ (.Y(_02892_),
    .B1(net4710),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][1] ),
    .A2(net4738),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][1] ));
 sg13g2_a22oi_1 _11553_ (.Y(_02893_),
    .B1(net4719),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][1] ),
    .A2(net4735),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][1] ));
 sg13g2_and2_1 _11554_ (.A(_02892_),
    .B(_02893_),
    .X(_02894_));
 sg13g2_a22oi_1 _11555_ (.Y(_02895_),
    .B1(net4713),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][1] ),
    .A2(net4727),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][1] ));
 sg13g2_a22oi_1 _11556_ (.Y(_02896_),
    .B1(net4807),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][1] ),
    .A2(net4851),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][1] ));
 sg13g2_a22oi_1 _11557_ (.Y(_02897_),
    .B1(net4717),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][1] ),
    .A2(net4741),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][1] ));
 sg13g2_and4_1 _11558_ (.A(net4769),
    .B(_02895_),
    .C(_02896_),
    .D(_02897_),
    .X(_02898_));
 sg13g2_a22oi_1 _11559_ (.Y(_02899_),
    .B1(_02894_),
    .B2(_02898_),
    .A2(net4827),
    .A1(_00299_));
 sg13g2_and2_1 _11560_ (.A(_02751_),
    .B(_02899_),
    .X(_02900_));
 sg13g2_xor2_1 _11561_ (.B(_02899_),
    .A(_02751_),
    .X(_02901_));
 sg13g2_xnor2_1 _11562_ (.Y(_02902_),
    .A(_02891_),
    .B(_02901_));
 sg13g2_and2_1 _11563_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][1] ),
    .B(net4766),
    .X(_02903_));
 sg13g2_a221oi_1 _11564_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][1] ),
    .C1(_02903_),
    .B1(net4754),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][1] ),
    .Y(_02904_),
    .A2(net4763));
 sg13g2_a221oi_1 _11565_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][1] ),
    .C1(net4823),
    .B1(net4814),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][1] ),
    .Y(_02905_),
    .A2(net4876));
 sg13g2_a22oi_1 _11566_ (.Y(_02906_),
    .B1(net4751),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][1] ),
    .A2(net4801),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][1] ));
 sg13g2_a22oi_1 _11567_ (.Y(_02907_),
    .B1(net4757),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][1] ),
    .A2(net4760),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][1] ));
 sg13g2_and3_1 _11568_ (.X(_02908_),
    .A(_02905_),
    .B(_02906_),
    .C(_02907_));
 sg13g2_a22oi_1 _11569_ (.Y(_02909_),
    .B1(_02904_),
    .B2(_02908_),
    .A2(net4824),
    .A1(_00297_));
 sg13g2_nand2_1 _11570_ (.Y(_02910_),
    .A(_02695_),
    .B(_02909_));
 sg13g2_xnor2_1 _11571_ (.Y(_02911_),
    .A(_02695_),
    .B(_02909_));
 sg13g2_a22oi_1 _11572_ (.Y(_02912_),
    .B1(net4848),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][1] ),
    .A2(net4813),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][1] ));
 sg13g2_a22oi_1 _11573_ (.Y(_02913_),
    .B1(net4793),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][1] ),
    .A2(net4799),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][1] ));
 sg13g2_nand3_1 _11574_ (.B(_02912_),
    .C(_02913_),
    .A(net4767),
    .Y(_02914_));
 sg13g2_a22oi_1 _11575_ (.Y(_02915_),
    .B1(net4796),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][1] ),
    .A2(net4748),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][1] ));
 sg13g2_a22oi_1 _11576_ (.Y(_02916_),
    .B1(net4745),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][1] ),
    .A2(net4800),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][1] ));
 sg13g2_nand2_1 _11577_ (.Y(_02917_),
    .A(_02915_),
    .B(_02916_));
 sg13g2_nand2_1 _11578_ (.Y(_02918_),
    .A(_00298_),
    .B(net4822));
 sg13g2_o21ai_1 _11579_ (.B1(_02918_),
    .Y(_02919_),
    .A1(_02914_),
    .A2(_02917_));
 sg13g2_xor2_1 _11580_ (.B(_02919_),
    .A(_02911_),
    .X(_02920_));
 sg13g2_nand2_1 _11581_ (.Y(_02921_),
    .A(_02753_),
    .B(_02920_));
 sg13g2_xnor2_1 _11582_ (.Y(_02922_),
    .A(_02753_),
    .B(_02920_));
 sg13g2_xor2_1 _11583_ (.B(_02922_),
    .A(_02902_),
    .X(_02923_));
 sg13g2_and2_1 _11584_ (.A(_02883_),
    .B(_02923_),
    .X(_02924_));
 sg13g2_nand2_1 _11585_ (.Y(_02925_),
    .A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .B(net4914));
 sg13g2_o21ai_1 _11586_ (.B1(net4929),
    .Y(_02926_),
    .A1(_02883_),
    .A2(_02923_));
 sg13g2_o21ai_1 _11587_ (.B1(_02925_),
    .Y(_00266_),
    .A1(_02924_),
    .A2(_02926_));
 sg13g2_and2_1 _11588_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][2] ),
    .B(net4730),
    .X(_02927_));
 sg13g2_a221oi_1 _11589_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][2] ),
    .C1(_02927_),
    .B1(net4655),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][2] ),
    .Y(_02928_),
    .A2(net4663));
 sg13g2_a21oi_1 _11590_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][2] ),
    .A2(net4657),
    .Y(_02929_),
    .B1(net4836));
 sg13g2_a22oi_1 _11591_ (.Y(_02930_),
    .B1(net4653),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][2] ),
    .A2(net4659),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][2] ));
 sg13g2_a22oi_1 _11592_ (.Y(_02931_),
    .B1(net4665),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][2] ),
    .A2(net4809),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][2] ));
 sg13g2_nand3_1 _11593_ (.B(_02930_),
    .C(_02931_),
    .A(_02929_),
    .Y(_02932_));
 sg13g2_a221oi_1 _11594_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][2] ),
    .C1(_02932_),
    .B1(net4650),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][2] ),
    .Y(_02933_),
    .A2(net4722));
 sg13g2_a22oi_1 _11595_ (.Y(_02934_),
    .B1(_02928_),
    .B2(_02933_),
    .A2(net4836),
    .A1(_00307_));
 sg13g2_a21oi_1 _11596_ (.A1(_02891_),
    .A2(_02901_),
    .Y(_02935_),
    .B1(_02900_));
 sg13g2_a22oi_1 _11597_ (.Y(_02936_),
    .B1(net4727),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][2] ),
    .A2(net4807),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][2] ));
 sg13g2_a22oi_1 _11598_ (.Y(_02937_),
    .B1(net4717),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][2] ),
    .A2(net4741),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][2] ));
 sg13g2_and2_1 _11599_ (.A(_02936_),
    .B(_02937_),
    .X(_02938_));
 sg13g2_a22oi_1 _11600_ (.Y(_02939_),
    .B1(net4710),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][2] ),
    .A2(net4713),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][2] ));
 sg13g2_a22oi_1 _11601_ (.Y(_02940_),
    .B1(net4738),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][2] ),
    .A2(net4851),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][2] ));
 sg13g2_a22oi_1 _11602_ (.Y(_02941_),
    .B1(net4719),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][2] ),
    .A2(net4735),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][2] ));
 sg13g2_and4_1 _11603_ (.A(net4769),
    .B(_02939_),
    .C(_02940_),
    .D(_02941_),
    .X(_02942_));
 sg13g2_a22oi_1 _11604_ (.Y(_02943_),
    .B1(_02938_),
    .B2(_02942_),
    .A2(net4827),
    .A1(_00306_));
 sg13g2_nor2b_1 _11605_ (.A(_02935_),
    .B_N(_02943_),
    .Y(_02944_));
 sg13g2_xnor2_1 _11606_ (.Y(_02945_),
    .A(_02935_),
    .B(_02943_));
 sg13g2_xnor2_1 _11607_ (.Y(_02946_),
    .A(_02934_),
    .B(_02945_));
 sg13g2_o21ai_1 _11608_ (.B1(_02921_),
    .Y(_02947_),
    .A1(_02902_),
    .A2(_02922_));
 sg13g2_o21ai_1 _11609_ (.B1(_02910_),
    .Y(_02948_),
    .A1(_02911_),
    .A2(_02919_));
 sg13g2_and2_1 _11610_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][2] ),
    .B(net4876),
    .X(_02949_));
 sg13g2_a221oi_1 _11611_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][2] ),
    .C1(_02949_),
    .B1(net4751),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][2] ),
    .Y(_02950_),
    .A2(net4760));
 sg13g2_a221oi_1 _11612_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][2] ),
    .C1(net4824),
    .B1(net4754),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][2] ),
    .Y(_02951_),
    .A2(net4814));
 sg13g2_a22oi_1 _11613_ (.Y(_02952_),
    .B1(net4757),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][2] ),
    .A2(net4763),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][2] ));
 sg13g2_a22oi_1 _11614_ (.Y(_02953_),
    .B1(net4800),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][2] ),
    .A2(net4766),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][2] ));
 sg13g2_and3_1 _11615_ (.X(_02954_),
    .A(_02951_),
    .B(_02952_),
    .C(_02953_));
 sg13g2_a22oi_1 _11616_ (.Y(_02955_),
    .B1(_02950_),
    .B2(_02954_),
    .A2(net4824),
    .A1(_00304_));
 sg13g2_nand2_1 _11617_ (.Y(_02956_),
    .A(_02948_),
    .B(_02955_));
 sg13g2_xnor2_1 _11618_ (.Y(_02957_),
    .A(_02948_),
    .B(_02955_));
 sg13g2_nand2_1 _11619_ (.Y(_02958_),
    .A(_00305_),
    .B(net4823));
 sg13g2_a22oi_1 _11620_ (.Y(_02959_),
    .B1(net4745),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][2] ),
    .A2(net4748),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][2] ));
 sg13g2_a22oi_1 _11621_ (.Y(_02960_),
    .B1(net4847),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][2] ),
    .A2(net4793),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][2] ));
 sg13g2_a22oi_1 _11622_ (.Y(_02961_),
    .B1(net4799),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][2] ),
    .A2(net4814),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][2] ));
 sg13g2_nand3_1 _11623_ (.B(_02960_),
    .C(_02961_),
    .A(net4768),
    .Y(_02962_));
 sg13g2_a22oi_1 _11624_ (.Y(_02963_),
    .B1(net4796),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][2] ),
    .A2(net4801),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][2] ));
 sg13g2_nand2_1 _11625_ (.Y(_02964_),
    .A(_02959_),
    .B(_02963_));
 sg13g2_o21ai_1 _11626_ (.B1(_02958_),
    .Y(_02965_),
    .A1(_02962_),
    .A2(_02964_));
 sg13g2_xor2_1 _11627_ (.B(_02965_),
    .A(_02957_),
    .X(_02966_));
 sg13g2_nand2_1 _11628_ (.Y(_02967_),
    .A(_02947_),
    .B(_02966_));
 sg13g2_xnor2_1 _11629_ (.Y(_02968_),
    .A(_02947_),
    .B(_02966_));
 sg13g2_xnor2_1 _11630_ (.Y(_02969_),
    .A(_02946_),
    .B(_02968_));
 sg13g2_a21oi_1 _11631_ (.A1(_02861_),
    .A2(_02866_),
    .Y(_02970_),
    .B1(_02859_));
 sg13g2_nand2_1 _11632_ (.Y(_02971_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][2] ),
    .B(_02796_));
 sg13g2_a221oi_1 _11633_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][2] ),
    .C1(net4698),
    .B1(_02848_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][2] ),
    .Y(_02972_),
    .A2(_02799_));
 sg13g2_a22oi_1 _11634_ (.Y(_02973_),
    .B1(_02807_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][2] ),
    .A2(net4873),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][2] ));
 sg13g2_a22oi_1 _11635_ (.Y(_02974_),
    .B1(_02805_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][2] ),
    .A2(net4692),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][2] ));
 sg13g2_nand4_1 _11636_ (.B(_02972_),
    .C(_02973_),
    .A(_02971_),
    .Y(_02975_),
    .D(_02974_));
 sg13g2_nand2_1 _11637_ (.Y(_02976_),
    .A(_00302_),
    .B(net4699));
 sg13g2_nand2_1 _11638_ (.Y(_02977_),
    .A(_02975_),
    .B(_02976_));
 sg13g2_nor2_1 _11639_ (.A(_02970_),
    .B(_02977_),
    .Y(_02978_));
 sg13g2_xor2_1 _11640_ (.B(_02977_),
    .A(_02970_),
    .X(_02979_));
 sg13g2_a221oi_1 _11641_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][2] ),
    .C1(net4681),
    .B1(_02834_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][2] ),
    .Y(_02980_),
    .A2(_02828_));
 sg13g2_a22oi_1 _11642_ (.Y(_02981_),
    .B1(net4668),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][2] ),
    .A2(net4685),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][2] ));
 sg13g2_a22oi_1 _11643_ (.Y(_02982_),
    .B1(net4672),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][2] ),
    .A2(_02831_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][2] ));
 sg13g2_and2_1 _11644_ (.A(_02981_),
    .B(_02982_),
    .X(_02983_));
 sg13g2_a22oi_1 _11645_ (.Y(_02984_),
    .B1(_02980_),
    .B2(_02983_),
    .A2(net4681),
    .A1(_00303_));
 sg13g2_xnor2_1 _11646_ (.Y(_02985_),
    .A(_02979_),
    .B(_02984_));
 sg13g2_a21oi_1 _11647_ (.A1(_02869_),
    .A2(_02880_),
    .Y(_02986_),
    .B1(_02879_));
 sg13g2_o21ai_1 _11648_ (.B1(_02871_),
    .Y(_02987_),
    .A1(_02872_),
    .A2(_02877_));
 sg13g2_mux2_1 _11649_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][2] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][2] ),
    .S(net4843),
    .X(_02988_));
 sg13g2_nand2_1 _11650_ (.Y(_02989_),
    .A(_02987_),
    .B(_02988_));
 sg13g2_nor2_1 _11651_ (.A(_02987_),
    .B(_02988_),
    .Y(_02990_));
 sg13g2_xnor2_1 _11652_ (.Y(_02991_),
    .A(_02987_),
    .B(_02988_));
 sg13g2_nand2_1 _11653_ (.Y(_02992_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][2] ),
    .B(net4701));
 sg13g2_a22oi_1 _11654_ (.Y(_02993_),
    .B1(net4781),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][2] ),
    .A2(net4785),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][2] ));
 sg13g2_a22oi_1 _11655_ (.Y(_02994_),
    .B1(net4777),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][2] ),
    .A2(net4788),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][2] ));
 sg13g2_nand4_1 _11656_ (.B(_02992_),
    .C(_02993_),
    .A(net4706),
    .Y(_02995_),
    .D(_02994_));
 sg13g2_o21ai_1 _11657_ (.B1(_02995_),
    .Y(_02996_),
    .A1(_02342_),
    .A2(net4706));
 sg13g2_xnor2_1 _11658_ (.Y(_02997_),
    .A(_02991_),
    .B(_02996_));
 sg13g2_or2_1 _11659_ (.X(_02998_),
    .B(_02997_),
    .A(_02986_));
 sg13g2_and2_1 _11660_ (.A(_02986_),
    .B(_02997_),
    .X(_02999_));
 sg13g2_xor2_1 _11661_ (.B(_02997_),
    .A(_02986_),
    .X(_03000_));
 sg13g2_xnor2_1 _11662_ (.Y(_03001_),
    .A(_02985_),
    .B(_03000_));
 sg13g2_o21ai_1 _11663_ (.B1(_03001_),
    .Y(_03002_),
    .A1(_02882_),
    .A2(_02924_));
 sg13g2_nor3_1 _11664_ (.A(_02882_),
    .B(_02924_),
    .C(_03001_),
    .Y(_03003_));
 sg13g2_or3_1 _11665_ (.A(_02882_),
    .B(_02924_),
    .C(_03001_),
    .X(_03004_));
 sg13g2_and2_1 _11666_ (.A(_03002_),
    .B(_03004_),
    .X(_03005_));
 sg13g2_xnor2_1 _11667_ (.Y(_03006_),
    .A(_02969_),
    .B(_03005_));
 sg13g2_mux2_1 _11668_ (.A0(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .A1(_03006_),
    .S(net4929),
    .X(_00277_));
 sg13g2_a22oi_1 _11669_ (.Y(_03007_),
    .B1(net4663),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][3] ),
    .A2(net4722),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][3] ));
 sg13g2_a22oi_1 _11670_ (.Y(_03008_),
    .B1(net4655),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][3] ),
    .A2(net4657),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][3] ));
 sg13g2_and2_1 _11671_ (.A(_03007_),
    .B(_03008_),
    .X(_03009_));
 sg13g2_a221oi_1 _11672_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][3] ),
    .C1(net4839),
    .B1(net4730),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][3] ),
    .Y(_03010_),
    .A2(net4810));
 sg13g2_a22oi_1 _11673_ (.Y(_03011_),
    .B1(net4659),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][3] ),
    .A2(net4665),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][3] ));
 sg13g2_nand2_1 _11674_ (.Y(_03012_),
    .A(_03010_),
    .B(_03011_));
 sg13g2_a221oi_1 _11675_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][3] ),
    .C1(_03012_),
    .B1(net4650),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][3] ),
    .Y(_03013_),
    .A2(net4653));
 sg13g2_a22oi_1 _11676_ (.Y(_03014_),
    .B1(_03009_),
    .B2(_03013_),
    .A2(net4839),
    .A1(_00314_));
 sg13g2_a21oi_1 _11677_ (.A1(_02934_),
    .A2(_02945_),
    .Y(_03015_),
    .B1(_02944_));
 sg13g2_a22oi_1 _11678_ (.Y(_03016_),
    .B1(net4807),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][3] ),
    .A2(net4851),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][3] ));
 sg13g2_a22oi_1 _11679_ (.Y(_03017_),
    .B1(net4710),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][3] ),
    .A2(net4741),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][3] ));
 sg13g2_and2_1 _11680_ (.A(_03016_),
    .B(_03017_),
    .X(_03018_));
 sg13g2_a22oi_1 _11681_ (.Y(_03019_),
    .B1(net4713),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][3] ),
    .A2(net4735),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][3] ));
 sg13g2_a22oi_1 _11682_ (.Y(_03020_),
    .B1(net4719),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][3] ),
    .A2(net4738),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][3] ));
 sg13g2_a22oi_1 _11683_ (.Y(_03021_),
    .B1(net4717),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][3] ),
    .A2(net4727),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][3] ));
 sg13g2_and4_1 _11684_ (.A(net4769),
    .B(_03019_),
    .C(_03020_),
    .D(_03021_),
    .X(_03022_));
 sg13g2_a22oi_1 _11685_ (.Y(_03023_),
    .B1(_03018_),
    .B2(_03022_),
    .A2(net4833),
    .A1(_00313_));
 sg13g2_nor2b_1 _11686_ (.A(_03015_),
    .B_N(_03023_),
    .Y(_03024_));
 sg13g2_xnor2_1 _11687_ (.Y(_03025_),
    .A(_03015_),
    .B(_03023_));
 sg13g2_xnor2_1 _11688_ (.Y(_03026_),
    .A(_03014_),
    .B(_03025_));
 sg13g2_o21ai_1 _11689_ (.B1(_02967_),
    .Y(_03027_),
    .A1(_02946_),
    .A2(_02968_));
 sg13g2_o21ai_1 _11690_ (.B1(_02956_),
    .Y(_03028_),
    .A1(_02957_),
    .A2(_02965_));
 sg13g2_and2_1 _11691_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][3] ),
    .B(net4755),
    .X(_03029_));
 sg13g2_a221oi_1 _11692_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][3] ),
    .C1(_03029_),
    .B1(net4749),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][3] ),
    .Y(_03030_),
    .A2(net4758));
 sg13g2_a221oi_1 _11693_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][3] ),
    .C1(net4824),
    .B1(net4801),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][3] ),
    .Y(_03031_),
    .A2(net4815));
 sg13g2_a22oi_1 _11694_ (.Y(_03032_),
    .B1(net4761),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][3] ),
    .A2(net4764),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][3] ));
 sg13g2_a22oi_1 _11695_ (.Y(_03033_),
    .B1(net4752),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][3] ),
    .A2(net4874),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][3] ));
 sg13g2_and3_1 _11696_ (.X(_03034_),
    .A(_03031_),
    .B(_03032_),
    .C(_03033_));
 sg13g2_a22oi_1 _11697_ (.Y(_03035_),
    .B1(_03030_),
    .B2(_03034_),
    .A2(net4824),
    .A1(_00311_));
 sg13g2_nand2_1 _11698_ (.Y(_03036_),
    .A(_03028_),
    .B(_03035_));
 sg13g2_xnor2_1 _11699_ (.Y(_03037_),
    .A(_03028_),
    .B(_03035_));
 sg13g2_nand2_1 _11700_ (.Y(_03038_),
    .A(_00312_),
    .B(net4823));
 sg13g2_a22oi_1 _11701_ (.Y(_03039_),
    .B1(net4847),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][3] ),
    .A2(net4797),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][3] ));
 sg13g2_a22oi_1 _11702_ (.Y(_03040_),
    .B1(net4803),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][3] ),
    .A2(net4815),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][3] ));
 sg13g2_nand2_1 _11703_ (.Y(_03041_),
    .A(_03039_),
    .B(_03040_));
 sg13g2_a22oi_1 _11704_ (.Y(_03042_),
    .B1(net4794),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][3] ),
    .A2(net4746),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][3] ));
 sg13g2_a22oi_1 _11705_ (.Y(_03043_),
    .B1(net4791),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][3] ),
    .A2(net4743),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][3] ));
 sg13g2_nand3_1 _11706_ (.B(_03042_),
    .C(_03043_),
    .A(net4768),
    .Y(_03044_));
 sg13g2_o21ai_1 _11707_ (.B1(_03038_),
    .Y(_03045_),
    .A1(_03041_),
    .A2(_03044_));
 sg13g2_xor2_1 _11708_ (.B(_03045_),
    .A(_03037_),
    .X(_03046_));
 sg13g2_nand2_1 _11709_ (.Y(_03047_),
    .A(_03027_),
    .B(_03046_));
 sg13g2_xnor2_1 _11710_ (.Y(_03048_),
    .A(_03027_),
    .B(_03046_));
 sg13g2_xor2_1 _11711_ (.B(_03048_),
    .A(_03026_),
    .X(_03049_));
 sg13g2_a21oi_1 _11712_ (.A1(_02979_),
    .A2(_02984_),
    .Y(_03050_),
    .B1(_02978_));
 sg13g2_o21ai_1 _11713_ (.B1(net4775),
    .Y(_03051_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][3] ),
    .A2(net4821));
 sg13g2_a22oi_1 _11714_ (.Y(_03052_),
    .B1(_02799_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][3] ),
    .A2(_02796_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][3] ));
 sg13g2_a22oi_1 _11715_ (.Y(_03053_),
    .B1(_02807_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][3] ),
    .A2(_02805_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][3] ));
 sg13g2_a22oi_1 _11716_ (.Y(_03054_),
    .B1(net4692),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][3] ),
    .A2(net4873),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][3] ));
 sg13g2_nand4_1 _11717_ (.B(_03052_),
    .C(_03053_),
    .A(_03051_),
    .Y(_03055_),
    .D(_03054_));
 sg13g2_nand2_1 _11718_ (.Y(_03056_),
    .A(_00309_),
    .B(net4699));
 sg13g2_nand2_1 _11719_ (.Y(_03057_),
    .A(_03055_),
    .B(_03056_));
 sg13g2_nor2_1 _11720_ (.A(_03050_),
    .B(_03057_),
    .Y(_03058_));
 sg13g2_xor2_1 _11721_ (.B(_03057_),
    .A(_03050_),
    .X(_03059_));
 sg13g2_a221oi_1 _11722_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][3] ),
    .C1(net4682),
    .B1(net4670),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][3] ),
    .Y(_03060_),
    .A2(net4677));
 sg13g2_a22oi_1 _11723_ (.Y(_03061_),
    .B1(_02836_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][3] ),
    .A2(net4673),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][3] ));
 sg13g2_a22oi_1 _11724_ (.Y(_03062_),
    .B1(_02831_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][3] ),
    .A2(net4685),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][3] ));
 sg13g2_and2_1 _11725_ (.A(_03061_),
    .B(_03062_),
    .X(_03063_));
 sg13g2_a22oi_1 _11726_ (.Y(_03064_),
    .B1(_03060_),
    .B2(_03063_),
    .A2(net4681),
    .A1(_00310_));
 sg13g2_xnor2_1 _11727_ (.Y(_03065_),
    .A(_03059_),
    .B(_03064_));
 sg13g2_o21ai_1 _11728_ (.B1(_02998_),
    .Y(_03066_),
    .A1(_02985_),
    .A2(_02999_));
 sg13g2_o21ai_1 _11729_ (.B1(_02989_),
    .Y(_03067_),
    .A1(_02990_),
    .A2(_02996_));
 sg13g2_mux2_1 _11730_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][3] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][3] ),
    .S(net4843),
    .X(_03068_));
 sg13g2_nand2_1 _11731_ (.Y(_03069_),
    .A(_03067_),
    .B(_03068_));
 sg13g2_nor2_1 _11732_ (.A(_03067_),
    .B(_03068_),
    .Y(_03070_));
 sg13g2_xor2_1 _11733_ (.B(_03068_),
    .A(_03067_),
    .X(_03071_));
 sg13g2_nand2_1 _11734_ (.Y(_03072_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][3] ),
    .B(net4781));
 sg13g2_a22oi_1 _11735_ (.Y(_03073_),
    .B1(net4702),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][3] ),
    .A2(net4785),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][3] ));
 sg13g2_a22oi_1 _11736_ (.Y(_03074_),
    .B1(net4777),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][3] ),
    .A2(net4788),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][3] ));
 sg13g2_nand4_1 _11737_ (.B(_03072_),
    .C(_03073_),
    .A(net4706),
    .Y(_03075_),
    .D(_03074_));
 sg13g2_o21ai_1 _11738_ (.B1(_03075_),
    .Y(_03076_),
    .A1(_02343_),
    .A2(net4706));
 sg13g2_xnor2_1 _11739_ (.Y(_03077_),
    .A(_03071_),
    .B(_03076_));
 sg13g2_nand2_1 _11740_ (.Y(_03078_),
    .A(_03066_),
    .B(_03077_));
 sg13g2_nor2_1 _11741_ (.A(_03066_),
    .B(_03077_),
    .Y(_03079_));
 sg13g2_xor2_1 _11742_ (.B(_03077_),
    .A(_03066_),
    .X(_03080_));
 sg13g2_xnor2_1 _11743_ (.Y(_03081_),
    .A(_03065_),
    .B(_03080_));
 sg13g2_o21ai_1 _11744_ (.B1(_03002_),
    .Y(_03082_),
    .A1(_02969_),
    .A2(_03003_));
 sg13g2_and2_1 _11745_ (.A(_03081_),
    .B(_03082_),
    .X(_03083_));
 sg13g2_xor2_1 _11746_ (.B(_03082_),
    .A(_03081_),
    .X(_03084_));
 sg13g2_o21ai_1 _11747_ (.B1(net4929),
    .Y(_03085_),
    .A1(_03049_),
    .A2(_03084_));
 sg13g2_a21oi_1 _11748_ (.A1(_03049_),
    .A2(_03084_),
    .Y(_03086_),
    .B1(_03085_));
 sg13g2_a21o_1 _11749_ (.A2(net4914),
    .A1(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .B1(_03086_),
    .X(_00280_));
 sg13g2_a22oi_1 _11750_ (.Y(_03087_),
    .B1(net4649),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][4] ),
    .A2(net4652),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][4] ));
 sg13g2_and2_1 _11751_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][4] ),
    .B(net4810),
    .X(_03088_));
 sg13g2_a221oi_1 _11752_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][4] ),
    .C1(_03088_),
    .B1(net4658),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][4] ),
    .Y(_03089_),
    .A2(net4662));
 sg13g2_a21oi_1 _11753_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][4] ),
    .A2(net4723),
    .Y(_03090_),
    .B1(net4839));
 sg13g2_a22oi_1 _11754_ (.Y(_03091_),
    .B1(net4664),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][4] ),
    .A2(net4732),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][4] ));
 sg13g2_nand3_1 _11755_ (.B(_03090_),
    .C(_03091_),
    .A(_03087_),
    .Y(_03092_));
 sg13g2_a221oi_1 _11756_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][4] ),
    .C1(_03092_),
    .B1(net4654),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][4] ),
    .Y(_03093_),
    .A2(net4656));
 sg13g2_a22oi_1 _11757_ (.Y(_03094_),
    .B1(_03089_),
    .B2(_03093_),
    .A2(net4839),
    .A1(_00323_));
 sg13g2_a22oi_1 _11758_ (.Y(_03095_),
    .B1(net4733),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][4] ),
    .A2(net4737),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][4] ));
 sg13g2_a22oi_1 _11759_ (.Y(_03096_),
    .B1(net4734),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][4] ),
    .A2(net4740),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][4] ));
 sg13g2_and2_1 _11760_ (.A(_03095_),
    .B(_03096_),
    .X(_03097_));
 sg13g2_a22oi_1 _11761_ (.Y(_03098_),
    .B1(net4712),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][4] ),
    .A2(net4715),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][4] ));
 sg13g2_a22oi_1 _11762_ (.Y(_03099_),
    .B1(net4725),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][4] ),
    .A2(net4849),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][4] ));
 sg13g2_a22oi_1 _11763_ (.Y(_03100_),
    .B1(net4709),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][4] ),
    .A2(net4808),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][4] ));
 sg13g2_and4_1 _11764_ (.A(net4771),
    .B(_03098_),
    .C(_03099_),
    .D(_03100_),
    .X(_03101_));
 sg13g2_a22oi_1 _11765_ (.Y(_03102_),
    .B1(_03097_),
    .B2(_03101_),
    .A2(net4834),
    .A1(_00322_));
 sg13g2_a21oi_2 _11766_ (.B1(_03024_),
    .Y(_03103_),
    .A2(_03025_),
    .A1(_03014_));
 sg13g2_nor2b_1 _11767_ (.A(_03103_),
    .B_N(_03102_),
    .Y(_03104_));
 sg13g2_xnor2_1 _11768_ (.Y(_03105_),
    .A(_03102_),
    .B(_03103_));
 sg13g2_xnor2_1 _11769_ (.Y(_03106_),
    .A(_03094_),
    .B(_03105_));
 sg13g2_o21ai_1 _11770_ (.B1(_03047_),
    .Y(_03107_),
    .A1(_03026_),
    .A2(_03048_));
 sg13g2_o21ai_1 _11771_ (.B1(_03036_),
    .Y(_03108_),
    .A1(_03037_),
    .A2(_03045_));
 sg13g2_and2_1 _11772_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][4] ),
    .B(net4758),
    .X(_03109_));
 sg13g2_a221oi_1 _11773_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][4] ),
    .C1(_03109_),
    .B1(net4752),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][4] ),
    .Y(_03110_),
    .A2(net4761));
 sg13g2_a221oi_1 _11774_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][4] ),
    .C1(net4828),
    .B1(net4815),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][4] ),
    .Y(_03111_),
    .A2(net4764));
 sg13g2_a22oi_1 _11775_ (.Y(_03112_),
    .B1(net4806),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][4] ),
    .A2(net4874),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][4] ));
 sg13g2_a22oi_1 _11776_ (.Y(_03113_),
    .B1(net4749),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][4] ),
    .A2(net4755),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][4] ));
 sg13g2_and3_1 _11777_ (.X(_03114_),
    .A(_03111_),
    .B(_03112_),
    .C(_03113_));
 sg13g2_a22oi_1 _11778_ (.Y(_03115_),
    .B1(_03110_),
    .B2(_03114_),
    .A2(net4828),
    .A1(_00320_));
 sg13g2_nand2_1 _11779_ (.Y(_03116_),
    .A(_03108_),
    .B(_03115_));
 sg13g2_xnor2_1 _11780_ (.Y(_03117_),
    .A(_03108_),
    .B(_03115_));
 sg13g2_a22oi_1 _11781_ (.Y(_03118_),
    .B1(net4847),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][4] ),
    .A2(net4791),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][4] ));
 sg13g2_a22oi_1 _11782_ (.Y(_03119_),
    .B1(net4794),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][4] ),
    .A2(net4743),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][4] ));
 sg13g2_a22oi_1 _11783_ (.Y(_03120_),
    .B1(net4797),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][4] ),
    .A2(net4746),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][4] ));
 sg13g2_a22oi_1 _11784_ (.Y(_03121_),
    .B1(net4803),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][4] ),
    .A2(net4815),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][4] ));
 sg13g2_nand2_1 _11785_ (.Y(_03122_),
    .A(_03120_),
    .B(_03121_));
 sg13g2_nand3_1 _11786_ (.B(_03118_),
    .C(_03119_),
    .A(net4768),
    .Y(_03123_));
 sg13g2_nand2_1 _11787_ (.Y(_03124_),
    .A(_00321_),
    .B(net4829));
 sg13g2_o21ai_1 _11788_ (.B1(_03124_),
    .Y(_03125_),
    .A1(_03122_),
    .A2(_03123_));
 sg13g2_xor2_1 _11789_ (.B(_03125_),
    .A(_03117_),
    .X(_03126_));
 sg13g2_nand2_1 _11790_ (.Y(_03127_),
    .A(_03107_),
    .B(_03126_));
 sg13g2_xnor2_1 _11791_ (.Y(_03128_),
    .A(_03107_),
    .B(_03126_));
 sg13g2_xnor2_1 _11792_ (.Y(_03129_),
    .A(_03106_),
    .B(_03128_));
 sg13g2_a21oi_1 _11793_ (.A1(_03059_),
    .A2(_03064_),
    .Y(_03130_),
    .B1(_03058_));
 sg13g2_nand2_1 _11794_ (.Y(_03131_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][4] ),
    .B(net4696));
 sg13g2_a221oi_1 _11795_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][4] ),
    .C1(net4698),
    .B1(_02848_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][4] ),
    .Y(_03132_),
    .A2(net4694));
 sg13g2_a22oi_1 _11796_ (.Y(_03133_),
    .B1(net4692),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][4] ),
    .A2(net4873),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][4] ));
 sg13g2_a22oi_1 _11797_ (.Y(_03134_),
    .B1(net4688),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][4] ),
    .A2(net4690),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][4] ));
 sg13g2_nand4_1 _11798_ (.B(_03132_),
    .C(_03133_),
    .A(_03131_),
    .Y(_03135_),
    .D(_03134_));
 sg13g2_nand2_1 _11799_ (.Y(_03136_),
    .A(_00318_),
    .B(net4699));
 sg13g2_nand2_2 _11800_ (.Y(_03137_),
    .A(_03135_),
    .B(_03136_));
 sg13g2_nor2_1 _11801_ (.A(_03130_),
    .B(_03137_),
    .Y(_03138_));
 sg13g2_xor2_1 _11802_ (.B(_03137_),
    .A(_03130_),
    .X(_03139_));
 sg13g2_a221oi_1 _11803_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][4] ),
    .C1(net4682),
    .B1(net4670),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][4] ),
    .Y(_03140_),
    .A2(net4677));
 sg13g2_a22oi_1 _11804_ (.Y(_03141_),
    .B1(net4675),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][4] ),
    .A2(net4685),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][4] ));
 sg13g2_a22oi_1 _11805_ (.Y(_03142_),
    .B1(net4668),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][4] ),
    .A2(net4672),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][4] ));
 sg13g2_and2_1 _11806_ (.A(_03141_),
    .B(_03142_),
    .X(_03143_));
 sg13g2_a22oi_1 _11807_ (.Y(_03144_),
    .B1(_03140_),
    .B2(_03143_),
    .A2(net4682),
    .A1(_00319_));
 sg13g2_xnor2_1 _11808_ (.Y(_03145_),
    .A(_03139_),
    .B(_03144_));
 sg13g2_o21ai_1 _11809_ (.B1(_03078_),
    .Y(_03146_),
    .A1(_03065_),
    .A2(_03079_));
 sg13g2_o21ai_1 _11810_ (.B1(_03069_),
    .Y(_03147_),
    .A1(_03070_),
    .A2(_03076_));
 sg13g2_mux2_1 _11811_ (.A0(_00316_),
    .A1(_00315_),
    .S(net4843),
    .X(_03148_));
 sg13g2_nand2b_1 _11812_ (.Y(_03149_),
    .B(_03147_),
    .A_N(_03148_));
 sg13g2_xor2_1 _11813_ (.B(_03148_),
    .A(_03147_),
    .X(_03150_));
 sg13g2_nand2_1 _11814_ (.Y(_03151_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][4] ),
    .B(net4781));
 sg13g2_a22oi_1 _11815_ (.Y(_03152_),
    .B1(net4702),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][4] ),
    .A2(net4785),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][4] ));
 sg13g2_a22oi_1 _11816_ (.Y(_03153_),
    .B1(net4777),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][4] ),
    .A2(net4788),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][4] ));
 sg13g2_nand4_1 _11817_ (.B(_03151_),
    .C(_03152_),
    .A(net4707),
    .Y(_03154_),
    .D(_03153_));
 sg13g2_o21ai_1 _11818_ (.B1(_03154_),
    .Y(_03155_),
    .A1(_02344_),
    .A2(net4707));
 sg13g2_xor2_1 _11819_ (.B(_03155_),
    .A(_03150_),
    .X(_03156_));
 sg13g2_nand2_1 _11820_ (.Y(_03157_),
    .A(_03146_),
    .B(_03156_));
 sg13g2_nor2_1 _11821_ (.A(_03146_),
    .B(_03156_),
    .Y(_03158_));
 sg13g2_xor2_1 _11822_ (.B(_03156_),
    .A(_03146_),
    .X(_03159_));
 sg13g2_xnor2_1 _11823_ (.Y(_03160_),
    .A(_03145_),
    .B(_03159_));
 sg13g2_a21oi_2 _11824_ (.B1(_03083_),
    .Y(_03161_),
    .A2(_03084_),
    .A1(_03049_));
 sg13g2_nand2b_1 _11825_ (.Y(_03162_),
    .B(_03160_),
    .A_N(_03161_));
 sg13g2_nor2b_1 _11826_ (.A(_03160_),
    .B_N(_03161_),
    .Y(_03163_));
 sg13g2_xor2_1 _11827_ (.B(_03161_),
    .A(_03160_),
    .X(_03164_));
 sg13g2_xnor2_1 _11828_ (.Y(_03165_),
    .A(_03129_),
    .B(_03164_));
 sg13g2_nor2_1 _11829_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .B(net4931),
    .Y(_03166_));
 sg13g2_a21oi_1 _11830_ (.A1(net4931),
    .A2(_03165_),
    .Y(_00281_),
    .B1(_03166_));
 sg13g2_a22oi_1 _11831_ (.Y(_03167_),
    .B1(net4656),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][5] ),
    .A2(net4661),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][5] ));
 sg13g2_a22oi_1 _11832_ (.Y(_03168_),
    .B1(net4660),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][5] ),
    .A2(net4723),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][5] ));
 sg13g2_and2_1 _11833_ (.A(_03167_),
    .B(_03168_),
    .X(_03169_));
 sg13g2_a221oi_1 _11834_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][5] ),
    .C1(net4838),
    .B1(net4731),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][5] ),
    .Y(_03170_),
    .A2(net4810));
 sg13g2_a22oi_1 _11835_ (.Y(_03171_),
    .B1(_02742_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][5] ),
    .A2(net4666),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][5] ));
 sg13g2_nand2_1 _11836_ (.Y(_03172_),
    .A(_03170_),
    .B(_03171_));
 sg13g2_a221oi_1 _11837_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][5] ),
    .C1(_03172_),
    .B1(net4651),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][5] ),
    .Y(_03173_),
    .A2(_02744_));
 sg13g2_a22oi_1 _11838_ (.Y(_03174_),
    .B1(_03169_),
    .B2(_03173_),
    .A2(net4838),
    .A1(_00332_));
 sg13g2_a22oi_1 _11839_ (.Y(_03175_),
    .B1(net4712),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][5] ),
    .A2(net4850),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][5] ));
 sg13g2_a22oi_1 _11840_ (.Y(_03176_),
    .B1(net4715),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][5] ),
    .A2(net4737),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][5] ));
 sg13g2_a22oi_1 _11841_ (.Y(_03177_),
    .B1(net4720),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][5] ),
    .A2(net4734),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][5] ));
 sg13g2_a22oi_1 _11842_ (.Y(_03178_),
    .B1(net4728),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][5] ),
    .A2(net4740),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][5] ));
 sg13g2_and2_1 _11843_ (.A(_03177_),
    .B(_03178_),
    .X(_03179_));
 sg13g2_a22oi_1 _11844_ (.Y(_03180_),
    .B1(net4709),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][5] ),
    .A2(net4808),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][5] ));
 sg13g2_and4_1 _11845_ (.A(net4771),
    .B(_03175_),
    .C(_03176_),
    .D(_03180_),
    .X(_03181_));
 sg13g2_a22oi_1 _11846_ (.Y(_03182_),
    .B1(_03179_),
    .B2(_03181_),
    .A2(net4834),
    .A1(_00331_));
 sg13g2_a21oi_2 _11847_ (.B1(_03104_),
    .Y(_03183_),
    .A2(_03105_),
    .A1(_03094_));
 sg13g2_nor2b_1 _11848_ (.A(_03183_),
    .B_N(_03182_),
    .Y(_03184_));
 sg13g2_xnor2_1 _11849_ (.Y(_03185_),
    .A(_03182_),
    .B(_03183_));
 sg13g2_xnor2_1 _11850_ (.Y(_03186_),
    .A(_03174_),
    .B(_03185_));
 sg13g2_o21ai_1 _11851_ (.B1(_03127_),
    .Y(_03187_),
    .A1(_03106_),
    .A2(_03128_));
 sg13g2_o21ai_1 _11852_ (.B1(_03116_),
    .Y(_03188_),
    .A1(_03117_),
    .A2(_03125_));
 sg13g2_and2_1 _11853_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][5] ),
    .B(net4764),
    .X(_03189_));
 sg13g2_a221oi_1 _11854_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][5] ),
    .C1(_03189_),
    .B1(net4749),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][5] ),
    .Y(_03190_),
    .A2(net4761));
 sg13g2_a221oi_1 _11855_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][5] ),
    .C1(net4828),
    .B1(net4752),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][5] ),
    .Y(_03191_),
    .A2(net4815));
 sg13g2_a22oi_1 _11856_ (.Y(_03192_),
    .B1(net4803),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][5] ),
    .A2(net4874),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][5] ));
 sg13g2_a22oi_1 _11857_ (.Y(_03193_),
    .B1(net4755),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][5] ),
    .A2(net4758),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][5] ));
 sg13g2_and3_1 _11858_ (.X(_03194_),
    .A(_03191_),
    .B(_03192_),
    .C(_03193_));
 sg13g2_a22oi_1 _11859_ (.Y(_03195_),
    .B1(_03190_),
    .B2(_03194_),
    .A2(net4828),
    .A1(_00329_));
 sg13g2_nand2_1 _11860_ (.Y(_03196_),
    .A(_03188_),
    .B(_03195_));
 sg13g2_xnor2_1 _11861_ (.Y(_03197_),
    .A(_03188_),
    .B(_03195_));
 sg13g2_a22oi_1 _11862_ (.Y(_03198_),
    .B1(net4746),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][5] ),
    .A2(net4815),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][5] ));
 sg13g2_a22oi_1 _11863_ (.Y(_03199_),
    .B1(net4794),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][5] ),
    .A2(net4803),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][5] ));
 sg13g2_nand2_1 _11864_ (.Y(_03200_),
    .A(_03198_),
    .B(_03199_));
 sg13g2_a22oi_1 _11865_ (.Y(_03201_),
    .B1(net4846),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][5] ),
    .A2(net4797),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][5] ));
 sg13g2_a22oi_1 _11866_ (.Y(_03202_),
    .B1(net4791),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][5] ),
    .A2(net4743),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][5] ));
 sg13g2_nand3_1 _11867_ (.B(_03201_),
    .C(_03202_),
    .A(net4767),
    .Y(_03203_));
 sg13g2_nand2_1 _11868_ (.Y(_03204_),
    .A(_00330_),
    .B(net4827));
 sg13g2_o21ai_1 _11869_ (.B1(_03204_),
    .Y(_03205_),
    .A1(_03200_),
    .A2(_03203_));
 sg13g2_xor2_1 _11870_ (.B(_03205_),
    .A(_03197_),
    .X(_03206_));
 sg13g2_nand2_1 _11871_ (.Y(_03207_),
    .A(_03187_),
    .B(_03206_));
 sg13g2_xnor2_1 _11872_ (.Y(_03208_),
    .A(_03187_),
    .B(_03206_));
 sg13g2_xnor2_1 _11873_ (.Y(_03209_),
    .A(_03186_),
    .B(_03208_));
 sg13g2_a21oi_1 _11874_ (.A1(_03139_),
    .A2(_03144_),
    .Y(_03210_),
    .B1(_03138_));
 sg13g2_o21ai_1 _11875_ (.B1(net4774),
    .Y(_03211_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][5] ),
    .A2(net4821));
 sg13g2_a22oi_1 _11876_ (.Y(_03212_),
    .B1(net4693),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][5] ),
    .A2(net4695),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][5] ));
 sg13g2_a22oi_1 _11877_ (.Y(_03213_),
    .B1(net4688),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][5] ),
    .A2(net4691),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][5] ));
 sg13g2_a22oi_1 _11878_ (.Y(_03214_),
    .B1(net4690),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][5] ),
    .A2(net4872),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][5] ));
 sg13g2_nand4_1 _11879_ (.B(_03212_),
    .C(_03213_),
    .A(_03211_),
    .Y(_03215_),
    .D(_03214_));
 sg13g2_nand2_1 _11880_ (.Y(_03216_),
    .A(_00327_),
    .B(net4700));
 sg13g2_nand2_2 _11881_ (.Y(_03217_),
    .A(_03215_),
    .B(_03216_));
 sg13g2_nor2_1 _11882_ (.A(_03210_),
    .B(_03217_),
    .Y(_03218_));
 sg13g2_xor2_1 _11883_ (.B(_03217_),
    .A(_03210_),
    .X(_03219_));
 sg13g2_a221oi_1 _11884_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][5] ),
    .C1(net4681),
    .B1(_02834_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][5] ),
    .Y(_03220_),
    .A2(_02828_));
 sg13g2_a22oi_1 _11885_ (.Y(_03221_),
    .B1(net4672),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][5] ),
    .A2(net4675),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][5] ));
 sg13g2_a22oi_1 _11886_ (.Y(_03222_),
    .B1(net4668),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][5] ),
    .A2(net4686),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][5] ));
 sg13g2_and2_1 _11887_ (.A(_03221_),
    .B(_03222_),
    .X(_03223_));
 sg13g2_a22oi_1 _11888_ (.Y(_03224_),
    .B1(_03220_),
    .B2(_03223_),
    .A2(net4681),
    .A1(_00328_));
 sg13g2_xnor2_1 _11889_ (.Y(_03225_),
    .A(_03219_),
    .B(_03224_));
 sg13g2_o21ai_1 _11890_ (.B1(_03157_),
    .Y(_03226_),
    .A1(_03145_),
    .A2(_03158_));
 sg13g2_o21ai_1 _11891_ (.B1(_03149_),
    .Y(_03227_),
    .A1(_03150_),
    .A2(_03155_));
 sg13g2_mux2_1 _11892_ (.A0(_00325_),
    .A1(_00324_),
    .S(net4843),
    .X(_03228_));
 sg13g2_nor2b_1 _11893_ (.A(_03228_),
    .B_N(_03227_),
    .Y(_03229_));
 sg13g2_xnor2_1 _11894_ (.Y(_03230_),
    .A(_03227_),
    .B(_03228_));
 sg13g2_and2_1 _11895_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][5] ),
    .B(net4784),
    .X(_03231_));
 sg13g2_a221oi_1 _11896_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][5] ),
    .C1(_03231_),
    .B1(net4703),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][5] ),
    .Y(_03232_),
    .A2(net4782));
 sg13g2_a221oi_1 _11897_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][5] ),
    .C1(net4648),
    .B1(net4778),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][5] ),
    .Y(_03233_),
    .A2(net4789));
 sg13g2_a22oi_1 _11898_ (.Y(_03234_),
    .B1(_03232_),
    .B2(_03233_),
    .A2(net4647),
    .A1(_00326_));
 sg13g2_xor2_1 _11899_ (.B(_03234_),
    .A(_03230_),
    .X(_03235_));
 sg13g2_nand2_1 _11900_ (.Y(_03236_),
    .A(_03226_),
    .B(_03235_));
 sg13g2_nor2_1 _11901_ (.A(_03226_),
    .B(_03235_),
    .Y(_03237_));
 sg13g2_xor2_1 _11902_ (.B(_03235_),
    .A(_03226_),
    .X(_03238_));
 sg13g2_xnor2_1 _11903_ (.Y(_03239_),
    .A(_03225_),
    .B(_03238_));
 sg13g2_o21ai_1 _11904_ (.B1(_03162_),
    .Y(_03240_),
    .A1(_03129_),
    .A2(_03163_));
 sg13g2_nand2_1 _11905_ (.Y(_03241_),
    .A(_03239_),
    .B(_03240_));
 sg13g2_xnor2_1 _11906_ (.Y(_03242_),
    .A(_03239_),
    .B(_03240_));
 sg13g2_xnor2_1 _11907_ (.Y(_03243_),
    .A(_03209_),
    .B(_03242_));
 sg13g2_nor2_1 _11908_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .B(net4931),
    .Y(_03244_));
 sg13g2_a21oi_1 _11909_ (.A1(net4931),
    .A2(_03243_),
    .Y(_00282_),
    .B1(_03244_));
 sg13g2_a22oi_1 _11910_ (.Y(_03245_),
    .B1(net4656),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][6] ),
    .A2(net4661),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][6] ));
 sg13g2_a221oi_1 _11911_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][6] ),
    .C1(net4839),
    .B1(net4731),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][6] ),
    .Y(_03246_),
    .A2(net4810));
 sg13g2_nand2_1 _11912_ (.Y(_03247_),
    .A(_03245_),
    .B(_03246_));
 sg13g2_a221oi_1 _11913_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][6] ),
    .C1(_03247_),
    .B1(net4651),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][6] ),
    .Y(_03248_),
    .A2(net4652));
 sg13g2_a22oi_1 _11914_ (.Y(_03249_),
    .B1(net4660),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][6] ),
    .A2(net4723),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][6] ));
 sg13g2_a22oi_1 _11915_ (.Y(_03250_),
    .B1(net4654),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][6] ),
    .A2(net4666),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][6] ));
 sg13g2_and2_1 _11916_ (.A(_03249_),
    .B(_03250_),
    .X(_03251_));
 sg13g2_a22oi_1 _11917_ (.Y(_03252_),
    .B1(_03248_),
    .B2(_03251_),
    .A2(net4838),
    .A1(_00339_));
 sg13g2_a21oi_1 _11918_ (.A1(_03174_),
    .A2(_03185_),
    .Y(_03253_),
    .B1(_03184_));
 sg13g2_a22oi_1 _11919_ (.Y(_03254_),
    .B1(net4710),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][6] ),
    .A2(net4735),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][6] ));
 sg13g2_a22oi_1 _11920_ (.Y(_03255_),
    .B1(net4713),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][6] ),
    .A2(net4850),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][6] ));
 sg13g2_a22oi_1 _11921_ (.Y(_03256_),
    .B1(net4716),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][6] ),
    .A2(net4739),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][6] ));
 sg13g2_a22oi_1 _11922_ (.Y(_03257_),
    .B1(net4740),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][6] ),
    .A2(net4808),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][6] ));
 sg13g2_and2_1 _11923_ (.A(_03256_),
    .B(_03257_),
    .X(_03258_));
 sg13g2_a22oi_1 _11924_ (.Y(_03259_),
    .B1(net4720),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][6] ),
    .A2(net4728),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][6] ));
 sg13g2_and4_1 _11925_ (.A(net4771),
    .B(_03254_),
    .C(_03255_),
    .D(_03259_),
    .X(_03260_));
 sg13g2_a22oi_1 _11926_ (.Y(_03261_),
    .B1(_03258_),
    .B2(_03260_),
    .A2(net4834),
    .A1(_00338_));
 sg13g2_nor2b_1 _11927_ (.A(_03253_),
    .B_N(_03261_),
    .Y(_03262_));
 sg13g2_xnor2_1 _11928_ (.Y(_03263_),
    .A(_03253_),
    .B(_03261_));
 sg13g2_xnor2_1 _11929_ (.Y(_03264_),
    .A(_03252_),
    .B(_03263_));
 sg13g2_o21ai_1 _11930_ (.B1(_03207_),
    .Y(_03265_),
    .A1(_03186_),
    .A2(_03208_));
 sg13g2_o21ai_1 _11931_ (.B1(_03196_),
    .Y(_03266_),
    .A1(_03197_),
    .A2(_03205_));
 sg13g2_nand2_1 _11932_ (.Y(_03267_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][6] ),
    .B(net4750));
 sg13g2_nand2_1 _11933_ (.Y(_03268_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][6] ),
    .B(net4758));
 sg13g2_a22oi_1 _11934_ (.Y(_03269_),
    .B1(net4875),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][6] ),
    .A2(net4765),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][6] ));
 sg13g2_a21oi_1 _11935_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][6] ),
    .A2(net4803),
    .Y(_03270_),
    .B1(net4829));
 sg13g2_a22oi_1 _11936_ (.Y(_03271_),
    .B1(net4755),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][6] ),
    .A2(net4815),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][6] ));
 sg13g2_nand4_1 _11937_ (.B(_03269_),
    .C(_03270_),
    .A(_03267_),
    .Y(_03272_),
    .D(_03271_));
 sg13g2_a221oi_1 _11938_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][6] ),
    .C1(_03272_),
    .B1(net4753),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][6] ),
    .Y(_03273_),
    .A2(net4761));
 sg13g2_a22oi_1 _11939_ (.Y(_03274_),
    .B1(_03268_),
    .B2(_03273_),
    .A2(net4829),
    .A1(_00336_));
 sg13g2_nand2_1 _11940_ (.Y(_03275_),
    .A(_03266_),
    .B(_03274_));
 sg13g2_xnor2_1 _11941_ (.Y(_03276_),
    .A(_03266_),
    .B(_03274_));
 sg13g2_nand2_1 _11942_ (.Y(_03277_),
    .A(_00337_),
    .B(net4827));
 sg13g2_a22oi_1 _11943_ (.Y(_03278_),
    .B1(net4798),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][6] ),
    .A2(net4747),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][6] ));
 sg13g2_a22oi_1 _11944_ (.Y(_03279_),
    .B1(net4743),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][6] ),
    .A2(net4803),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][6] ));
 sg13g2_a22oi_1 _11945_ (.Y(_03280_),
    .B1(net4846),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][6] ),
    .A2(net4816),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][6] ));
 sg13g2_nand2_1 _11946_ (.Y(_03281_),
    .A(_03279_),
    .B(_03280_));
 sg13g2_a22oi_1 _11947_ (.Y(_03282_),
    .B1(net4792),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][6] ),
    .A2(net4795),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][6] ));
 sg13g2_nand3_1 _11948_ (.B(_03278_),
    .C(_03282_),
    .A(net4770),
    .Y(_03283_));
 sg13g2_o21ai_1 _11949_ (.B1(_03277_),
    .Y(_03284_),
    .A1(_03281_),
    .A2(_03283_));
 sg13g2_xor2_1 _11950_ (.B(_03284_),
    .A(_03276_),
    .X(_03285_));
 sg13g2_nand2_1 _11951_ (.Y(_03286_),
    .A(_03265_),
    .B(_03285_));
 sg13g2_xnor2_1 _11952_ (.Y(_03287_),
    .A(_03265_),
    .B(_03285_));
 sg13g2_xnor2_1 _11953_ (.Y(_03288_),
    .A(_03264_),
    .B(_03287_));
 sg13g2_a21oi_1 _11954_ (.A1(_03219_),
    .A2(_03224_),
    .Y(_03289_),
    .B1(_03218_));
 sg13g2_nand2_1 _11955_ (.Y(_03290_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][6] ),
    .B(net4696));
 sg13g2_a221oi_1 _11956_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][6] ),
    .C1(net4698),
    .B1(_02848_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][6] ),
    .Y(_03291_),
    .A2(net4694));
 sg13g2_a22oi_1 _11957_ (.Y(_03292_),
    .B1(net4690),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][6] ),
    .A2(net4871),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][6] ));
 sg13g2_a22oi_1 _11958_ (.Y(_03293_),
    .B1(net4688),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][6] ),
    .A2(net4692),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][6] ));
 sg13g2_nand4_1 _11959_ (.B(_03291_),
    .C(_03292_),
    .A(_03290_),
    .Y(_03294_),
    .D(_03293_));
 sg13g2_nand2_1 _11960_ (.Y(_03295_),
    .A(_00334_),
    .B(net4699));
 sg13g2_nand2_2 _11961_ (.Y(_03296_),
    .A(_03294_),
    .B(_03295_));
 sg13g2_nor2_1 _11962_ (.A(_03289_),
    .B(_03296_),
    .Y(_03297_));
 sg13g2_xor2_1 _11963_ (.B(_03296_),
    .A(_03289_),
    .X(_03298_));
 sg13g2_a221oi_1 _11964_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][6] ),
    .C1(net4682),
    .B1(net4670),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][6] ),
    .Y(_03299_),
    .A2(net4677));
 sg13g2_a22oi_1 _11965_ (.Y(_03300_),
    .B1(net4668),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][6] ),
    .A2(net4672),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][6] ));
 sg13g2_a22oi_1 _11966_ (.Y(_03301_),
    .B1(net4675),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][6] ),
    .A2(net4685),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][6] ));
 sg13g2_and2_1 _11967_ (.A(_03300_),
    .B(_03301_),
    .X(_03302_));
 sg13g2_a22oi_1 _11968_ (.Y(_03303_),
    .B1(_03299_),
    .B2(_03302_),
    .A2(net4682),
    .A1(_00335_));
 sg13g2_xnor2_1 _11969_ (.Y(_03304_),
    .A(_03298_),
    .B(_03303_));
 sg13g2_o21ai_1 _11970_ (.B1(_03236_),
    .Y(_03305_),
    .A1(_03225_),
    .A2(_03237_));
 sg13g2_a21oi_1 _11971_ (.A1(_03230_),
    .A2(_03234_),
    .Y(_03306_),
    .B1(_03229_));
 sg13g2_mux2_1 _11972_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][6] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][6] ),
    .S(net4843),
    .X(_03307_));
 sg13g2_nand2b_1 _11973_ (.Y(_03308_),
    .B(_03307_),
    .A_N(_03306_));
 sg13g2_xor2_1 _11974_ (.B(_03307_),
    .A(_03306_),
    .X(_03309_));
 sg13g2_nand2_1 _11975_ (.Y(_03310_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][6] ),
    .B(net4701));
 sg13g2_a22oi_1 _11976_ (.Y(_03311_),
    .B1(net4780),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][6] ),
    .A2(net4784),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][6] ));
 sg13g2_a22oi_1 _11977_ (.Y(_03312_),
    .B1(net4776),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][6] ),
    .A2(net4787),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][6] ));
 sg13g2_nand4_1 _11978_ (.B(_03310_),
    .C(_03311_),
    .A(net4705),
    .Y(_03313_),
    .D(_03312_));
 sg13g2_o21ai_1 _11979_ (.B1(_03313_),
    .Y(_03314_),
    .A1(_02345_),
    .A2(net4705));
 sg13g2_xor2_1 _11980_ (.B(_03314_),
    .A(_03309_),
    .X(_03315_));
 sg13g2_nand2_1 _11981_ (.Y(_03316_),
    .A(_03305_),
    .B(_03315_));
 sg13g2_nor2_1 _11982_ (.A(_03305_),
    .B(_03315_),
    .Y(_03317_));
 sg13g2_xor2_1 _11983_ (.B(_03315_),
    .A(_03305_),
    .X(_03318_));
 sg13g2_xnor2_1 _11984_ (.Y(_03319_),
    .A(_03304_),
    .B(_03318_));
 sg13g2_o21ai_1 _11985_ (.B1(_03241_),
    .Y(_03320_),
    .A1(_03209_),
    .A2(_03242_));
 sg13g2_nand2_1 _11986_ (.Y(_03321_),
    .A(_03319_),
    .B(_03320_));
 sg13g2_xnor2_1 _11987_ (.Y(_03322_),
    .A(_03319_),
    .B(_03320_));
 sg13g2_xnor2_1 _11988_ (.Y(_03323_),
    .A(_03288_),
    .B(_03322_));
 sg13g2_nor2_1 _11989_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .B(net4932),
    .Y(_03324_));
 sg13g2_a21oi_1 _11990_ (.A1(net4931),
    .A2(_03323_),
    .Y(_00283_),
    .B1(_03324_));
 sg13g2_a21oi_1 _11991_ (.A1(_03298_),
    .A2(_03303_),
    .Y(_03325_),
    .B1(_03297_));
 sg13g2_o21ai_1 _11992_ (.B1(net4775),
    .Y(_03326_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][7] ),
    .A2(net4819));
 sg13g2_a22oi_1 _11993_ (.Y(_03327_),
    .B1(net4693),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][7] ),
    .A2(net4695),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][7] ));
 sg13g2_a22oi_1 _11994_ (.Y(_03328_),
    .B1(net4687),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][7] ),
    .A2(net4689),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][7] ));
 sg13g2_a22oi_1 _11995_ (.Y(_03329_),
    .B1(net4691),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][7] ),
    .A2(net4871),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][7] ));
 sg13g2_nand4_1 _11996_ (.B(_03327_),
    .C(_03328_),
    .A(_03326_),
    .Y(_03330_),
    .D(_03329_));
 sg13g2_nand2_1 _11997_ (.Y(_03331_),
    .A(_00341_),
    .B(net4700));
 sg13g2_nand2_2 _11998_ (.Y(_03332_),
    .A(_03330_),
    .B(_03331_));
 sg13g2_nor2_1 _11999_ (.A(_03325_),
    .B(_03332_),
    .Y(_03333_));
 sg13g2_xor2_1 _12000_ (.B(_03332_),
    .A(_03325_),
    .X(_03334_));
 sg13g2_a22oi_1 _12001_ (.Y(_03335_),
    .B1(net4668),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][7] ),
    .A2(net4675),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][7] ));
 sg13g2_a221oi_1 _12002_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][7] ),
    .C1(net4683),
    .B1(net4670),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][7] ),
    .Y(_03336_),
    .A2(net4677));
 sg13g2_a22oi_1 _12003_ (.Y(_03337_),
    .B1(net4673),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][7] ),
    .A2(net4686),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][7] ));
 sg13g2_and2_1 _12004_ (.A(_03335_),
    .B(_03337_),
    .X(_03338_));
 sg13g2_a22oi_1 _12005_ (.Y(_03339_),
    .B1(_03336_),
    .B2(_03338_),
    .A2(net4683),
    .A1(_00342_));
 sg13g2_xnor2_1 _12006_ (.Y(_03340_),
    .A(_03334_),
    .B(_03339_));
 sg13g2_o21ai_1 _12007_ (.B1(_03316_),
    .Y(_03341_),
    .A1(_03304_),
    .A2(_03317_));
 sg13g2_o21ai_1 _12008_ (.B1(_03308_),
    .Y(_03342_),
    .A1(_03309_),
    .A2(_03314_));
 sg13g2_mux2_1 _12009_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][7] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][7] ),
    .S(net4843),
    .X(_03343_));
 sg13g2_nand2_1 _12010_ (.Y(_03344_),
    .A(_03342_),
    .B(_03343_));
 sg13g2_xnor2_1 _12011_ (.Y(_03345_),
    .A(_03342_),
    .B(_03343_));
 sg13g2_nand2_1 _12012_ (.Y(_03346_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][7] ),
    .B(net4780));
 sg13g2_a22oi_1 _12013_ (.Y(_03347_),
    .B1(net4701),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][7] ),
    .A2(net4784),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][7] ));
 sg13g2_a22oi_1 _12014_ (.Y(_03348_),
    .B1(net4776),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][7] ),
    .A2(net4787),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][7] ));
 sg13g2_nand4_1 _12015_ (.B(_03346_),
    .C(_03347_),
    .A(net4705),
    .Y(_03349_),
    .D(_03348_));
 sg13g2_o21ai_1 _12016_ (.B1(_03349_),
    .Y(_03350_),
    .A1(_02346_),
    .A2(net4705));
 sg13g2_xnor2_1 _12017_ (.Y(_03351_),
    .A(_03345_),
    .B(_03350_));
 sg13g2_nand2b_1 _12018_ (.Y(_03352_),
    .B(_03341_),
    .A_N(_03351_));
 sg13g2_nor2b_1 _12019_ (.A(_03341_),
    .B_N(_03351_),
    .Y(_03353_));
 sg13g2_xnor2_1 _12020_ (.Y(_03354_),
    .A(_03341_),
    .B(_03351_));
 sg13g2_xnor2_1 _12021_ (.Y(_03355_),
    .A(_03340_),
    .B(_03354_));
 sg13g2_o21ai_1 _12022_ (.B1(_03321_),
    .Y(_03356_),
    .A1(_03288_),
    .A2(_03322_));
 sg13g2_and2_1 _12023_ (.A(_03355_),
    .B(_03356_),
    .X(_03357_));
 sg13g2_xor2_1 _12024_ (.B(_03356_),
    .A(_03355_),
    .X(_03358_));
 sg13g2_and2_1 _12025_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][7] ),
    .B(net4810),
    .X(_03359_));
 sg13g2_a221oi_1 _12026_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][7] ),
    .C1(_03359_),
    .B1(_02744_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][7] ),
    .Y(_03360_),
    .A2(net4661));
 sg13g2_a21oi_1 _12027_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][7] ),
    .A2(net4654),
    .Y(_03361_),
    .B1(net4838));
 sg13g2_a22oi_1 _12028_ (.Y(_03362_),
    .B1(net4660),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][7] ),
    .A2(net4731),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][7] ));
 sg13g2_a22oi_1 _12029_ (.Y(_03363_),
    .B1(net4666),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][7] ),
    .A2(net4723),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][7] ));
 sg13g2_nand3_1 _12030_ (.B(_03362_),
    .C(_03363_),
    .A(_03361_),
    .Y(_03364_));
 sg13g2_a221oi_1 _12031_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][7] ),
    .C1(_03364_),
    .B1(net4649),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][7] ),
    .Y(_03365_),
    .A2(net4656));
 sg13g2_a22oi_1 _12032_ (.Y(_03366_),
    .B1(_03360_),
    .B2(_03365_),
    .A2(net4838),
    .A1(_00346_));
 sg13g2_nand2_1 _12033_ (.Y(_03367_),
    .A(_00345_),
    .B(net4836));
 sg13g2_a22oi_1 _12034_ (.Y(_03368_),
    .B1(net4716),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][7] ),
    .A2(net4728),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][7] ));
 sg13g2_a22oi_1 _12035_ (.Y(_03369_),
    .B1(net4736),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][7] ),
    .A2(net4849),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][7] ));
 sg13g2_a22oi_1 _12036_ (.Y(_03370_),
    .B1(net4741),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][7] ),
    .A2(net4809),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][7] ));
 sg13g2_nand2_1 _12037_ (.Y(_03371_),
    .A(_03369_),
    .B(_03370_));
 sg13g2_a22oi_1 _12038_ (.Y(_03372_),
    .B1(net4714),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][7] ),
    .A2(net4737),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][7] ));
 sg13g2_a22oi_1 _12039_ (.Y(_03373_),
    .B1(net4711),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][7] ),
    .A2(net4720),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][7] ));
 sg13g2_nand4_1 _12040_ (.B(_03368_),
    .C(_03372_),
    .A(net4771),
    .Y(_03374_),
    .D(_03373_));
 sg13g2_o21ai_1 _12041_ (.B1(_03367_),
    .Y(_03375_),
    .A1(_03371_),
    .A2(_03374_));
 sg13g2_a21oi_1 _12042_ (.A1(_03252_),
    .A2(_03263_),
    .Y(_03376_),
    .B1(_03262_));
 sg13g2_nor2_1 _12043_ (.A(_03375_),
    .B(_03376_),
    .Y(_03377_));
 sg13g2_xor2_1 _12044_ (.B(_03376_),
    .A(_03375_),
    .X(_03378_));
 sg13g2_xnor2_1 _12045_ (.Y(_03379_),
    .A(_03366_),
    .B(_03378_));
 sg13g2_o21ai_1 _12046_ (.B1(_03286_),
    .Y(_03380_),
    .A1(_03264_),
    .A2(_03287_));
 sg13g2_o21ai_1 _12047_ (.B1(_03275_),
    .Y(_03381_),
    .A1(_03276_),
    .A2(_03284_));
 sg13g2_and2_1 _12048_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][7] ),
    .B(net4805),
    .X(_03382_));
 sg13g2_a221oi_1 _12049_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][7] ),
    .C1(_03382_),
    .B1(net4750),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][7] ),
    .Y(_03383_),
    .A2(net4756));
 sg13g2_a221oi_1 _12050_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][7] ),
    .C1(net4830),
    .B1(net4817),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][7] ),
    .Y(_03384_),
    .A2(net4765));
 sg13g2_a22oi_1 _12051_ (.Y(_03385_),
    .B1(net4875),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][7] ),
    .A2(net4762),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][7] ));
 sg13g2_a22oi_1 _12052_ (.Y(_03386_),
    .B1(net4753),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][7] ),
    .A2(net4759),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][7] ));
 sg13g2_and3_1 _12053_ (.X(_03387_),
    .A(_03384_),
    .B(_03385_),
    .C(_03386_));
 sg13g2_a22oi_1 _12054_ (.Y(_03388_),
    .B1(_03383_),
    .B2(_03387_),
    .A2(net4832),
    .A1(_00343_));
 sg13g2_nand2_1 _12055_ (.Y(_03389_),
    .A(_03381_),
    .B(_03388_));
 sg13g2_xnor2_1 _12056_ (.Y(_03390_),
    .A(_03381_),
    .B(_03388_));
 sg13g2_nand2_1 _12057_ (.Y(_03391_),
    .A(_00344_),
    .B(net4827));
 sg13g2_a22oi_1 _12058_ (.Y(_03392_),
    .B1(net4846),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][7] ),
    .A2(net4798),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][7] ));
 sg13g2_a22oi_1 _12059_ (.Y(_03393_),
    .B1(net4791),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][7] ),
    .A2(net4816),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][7] ));
 sg13g2_nand3_1 _12060_ (.B(_03392_),
    .C(_03393_),
    .A(net4770),
    .Y(_03394_));
 sg13g2_a22oi_1 _12061_ (.Y(_03395_),
    .B1(net4744),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][7] ),
    .A2(net4747),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][7] ));
 sg13g2_a22oi_1 _12062_ (.Y(_03396_),
    .B1(net4795),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][7] ),
    .A2(net4804),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][7] ));
 sg13g2_nand2_1 _12063_ (.Y(_03397_),
    .A(_03395_),
    .B(_03396_));
 sg13g2_o21ai_1 _12064_ (.B1(_03391_),
    .Y(_03398_),
    .A1(_03394_),
    .A2(_03397_));
 sg13g2_xor2_1 _12065_ (.B(_03398_),
    .A(_03390_),
    .X(_03399_));
 sg13g2_nand2_1 _12066_ (.Y(_03400_),
    .A(_03380_),
    .B(_03399_));
 sg13g2_xnor2_1 _12067_ (.Y(_03401_),
    .A(_03380_),
    .B(_03399_));
 sg13g2_xor2_1 _12068_ (.B(_03401_),
    .A(_03379_),
    .X(_03402_));
 sg13g2_xnor2_1 _12069_ (.Y(_03403_),
    .A(_03358_),
    .B(_03402_));
 sg13g2_nor2_1 _12070_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .B(net4931),
    .Y(_03404_));
 sg13g2_a21oi_1 _12071_ (.A1(net4931),
    .A2(_03403_),
    .Y(_00284_),
    .B1(_03404_));
 sg13g2_a22oi_1 _12072_ (.Y(_03405_),
    .B1(net4664),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][8] ),
    .A2(net4723),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][8] ));
 sg13g2_a22oi_1 _12073_ (.Y(_03406_),
    .B1(net4658),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][8] ),
    .A2(net4661),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][8] ));
 sg13g2_and2_1 _12074_ (.A(_03405_),
    .B(_03406_),
    .X(_03407_));
 sg13g2_a221oi_1 _12075_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][8] ),
    .C1(net4838),
    .B1(net4731),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][8] ),
    .Y(_03408_),
    .A2(net4810));
 sg13g2_a22oi_1 _12076_ (.Y(_03409_),
    .B1(net4654),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][8] ),
    .A2(net4656),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][8] ));
 sg13g2_nand2_1 _12077_ (.Y(_03410_),
    .A(_03408_),
    .B(_03409_));
 sg13g2_a221oi_1 _12078_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][8] ),
    .C1(_03410_),
    .B1(net4651),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][8] ),
    .Y(_03411_),
    .A2(net4652));
 sg13g2_a22oi_1 _12079_ (.Y(_03412_),
    .B1(_03407_),
    .B2(_03411_),
    .A2(net4838),
    .A1(_00355_));
 sg13g2_a21oi_1 _12080_ (.A1(_03366_),
    .A2(_03378_),
    .Y(_03413_),
    .B1(_03377_));
 sg13g2_a22oi_1 _12081_ (.Y(_03414_),
    .B1(net4734),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][8] ),
    .A2(net4809),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][8] ));
 sg13g2_a22oi_1 _12082_ (.Y(_03415_),
    .B1(net4709),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][8] ),
    .A2(net4716),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][8] ));
 sg13g2_a22oi_1 _12083_ (.Y(_03416_),
    .B1(net4721),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][8] ),
    .A2(net4849),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][8] ));
 sg13g2_and2_1 _12084_ (.A(_03415_),
    .B(_03416_),
    .X(_03417_));
 sg13g2_a22oi_1 _12085_ (.Y(_03418_),
    .B1(net4712),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][8] ),
    .A2(net4737),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][8] ));
 sg13g2_a22oi_1 _12086_ (.Y(_03419_),
    .B1(net4728),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][8] ),
    .A2(net4742),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][8] ));
 sg13g2_and4_1 _12087_ (.A(net4771),
    .B(_03414_),
    .C(_03418_),
    .D(_03419_),
    .X(_03420_));
 sg13g2_a22oi_1 _12088_ (.Y(_03421_),
    .B1(_03417_),
    .B2(_03420_),
    .A2(net4837),
    .A1(_00354_));
 sg13g2_nor2b_1 _12089_ (.A(_03413_),
    .B_N(_03421_),
    .Y(_03422_));
 sg13g2_xnor2_1 _12090_ (.Y(_03423_),
    .A(_03413_),
    .B(_03421_));
 sg13g2_xnor2_1 _12091_ (.Y(_03424_),
    .A(_03412_),
    .B(_03423_));
 sg13g2_o21ai_1 _12092_ (.B1(_03400_),
    .Y(_03425_),
    .A1(_03379_),
    .A2(_03401_));
 sg13g2_o21ai_1 _12093_ (.B1(_03389_),
    .Y(_03426_),
    .A1(_03390_),
    .A2(_03398_));
 sg13g2_and2_1 _12094_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][8] ),
    .B(net4875),
    .X(_03427_));
 sg13g2_a221oi_1 _12095_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][8] ),
    .C1(_03427_),
    .B1(net4756),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][8] ),
    .Y(_03428_),
    .A2(net4765));
 sg13g2_a221oi_1 _12096_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][8] ),
    .C1(net4830),
    .B1(net4817),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][8] ),
    .Y(_03429_),
    .A2(net4759));
 sg13g2_a22oi_1 _12097_ (.Y(_03430_),
    .B1(net4750),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][8] ),
    .A2(net4762),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][8] ));
 sg13g2_a22oi_1 _12098_ (.Y(_03431_),
    .B1(net4805),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][8] ),
    .A2(net4753),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][8] ));
 sg13g2_and3_1 _12099_ (.X(_03432_),
    .A(_03429_),
    .B(_03430_),
    .C(_03431_));
 sg13g2_a22oi_1 _12100_ (.Y(_03433_),
    .B1(_03428_),
    .B2(_03432_),
    .A2(net4830),
    .A1(_00352_));
 sg13g2_nand2_1 _12101_ (.Y(_03434_),
    .A(_03426_),
    .B(_03433_));
 sg13g2_xnor2_1 _12102_ (.Y(_03435_),
    .A(_03426_),
    .B(_03433_));
 sg13g2_a22oi_1 _12103_ (.Y(_03436_),
    .B1(net4798),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][8] ),
    .A2(net4816),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][8] ));
 sg13g2_a22oi_1 _12104_ (.Y(_03437_),
    .B1(net4846),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][8] ),
    .A2(net4804),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][8] ));
 sg13g2_nand2_1 _12105_ (.Y(_03438_),
    .A(_03436_),
    .B(_03437_));
 sg13g2_a22oi_1 _12106_ (.Y(_03439_),
    .B1(net4744),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][8] ),
    .A2(net4747),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][8] ));
 sg13g2_a22oi_1 _12107_ (.Y(_03440_),
    .B1(net4792),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][8] ),
    .A2(net4795),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][8] ));
 sg13g2_nand3_1 _12108_ (.B(_03439_),
    .C(_03440_),
    .A(net4770),
    .Y(_03441_));
 sg13g2_nand2_1 _12109_ (.Y(_03442_),
    .A(_00353_),
    .B(net4827));
 sg13g2_o21ai_1 _12110_ (.B1(_03442_),
    .Y(_03443_),
    .A1(_03438_),
    .A2(_03441_));
 sg13g2_xor2_1 _12111_ (.B(_03443_),
    .A(_03435_),
    .X(_03444_));
 sg13g2_nand2_1 _12112_ (.Y(_03445_),
    .A(_03425_),
    .B(_03444_));
 sg13g2_xnor2_1 _12113_ (.Y(_03446_),
    .A(_03425_),
    .B(_03444_));
 sg13g2_xnor2_1 _12114_ (.Y(_03447_),
    .A(_03424_),
    .B(_03446_));
 sg13g2_a21o_1 _12115_ (.A2(_03402_),
    .A1(_03358_),
    .B1(_03357_),
    .X(_03448_));
 sg13g2_a21oi_2 _12116_ (.B1(_03333_),
    .Y(_03449_),
    .A2(_03339_),
    .A1(_03334_));
 sg13g2_o21ai_1 _12117_ (.B1(net4775),
    .Y(_03450_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][8] ),
    .A2(net4819));
 sg13g2_a22oi_1 _12118_ (.Y(_03451_),
    .B1(net4693),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][8] ),
    .A2(net4695),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][8] ));
 sg13g2_a22oi_1 _12119_ (.Y(_03452_),
    .B1(net4689),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][8] ),
    .A2(net4871),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][8] ));
 sg13g2_a22oi_1 _12120_ (.Y(_03453_),
    .B1(net4687),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][8] ),
    .A2(net4691),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][8] ));
 sg13g2_nand4_1 _12121_ (.B(_03451_),
    .C(_03452_),
    .A(_03450_),
    .Y(_03454_),
    .D(_03453_));
 sg13g2_nand2_1 _12122_ (.Y(_03455_),
    .A(_00350_),
    .B(net4697));
 sg13g2_nand2_2 _12123_ (.Y(_03456_),
    .A(_03454_),
    .B(_03455_));
 sg13g2_nor2_1 _12124_ (.A(_03449_),
    .B(_03456_),
    .Y(_03457_));
 sg13g2_xor2_1 _12125_ (.B(_03456_),
    .A(_03449_),
    .X(_03458_));
 sg13g2_a221oi_1 _12126_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][8] ),
    .C1(net4680),
    .B1(net4669),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][8] ),
    .Y(_03459_),
    .A2(net4676));
 sg13g2_a22oi_1 _12127_ (.Y(_03460_),
    .B1(net4667),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][8] ),
    .A2(net4684),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][8] ));
 sg13g2_a22oi_1 _12128_ (.Y(_03461_),
    .B1(net4671),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][8] ),
    .A2(net4674),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][8] ));
 sg13g2_and2_1 _12129_ (.A(_03460_),
    .B(_03461_),
    .X(_03462_));
 sg13g2_a22oi_1 _12130_ (.Y(_03463_),
    .B1(_03459_),
    .B2(_03462_),
    .A2(net4680),
    .A1(_00351_));
 sg13g2_xnor2_1 _12131_ (.Y(_03464_),
    .A(_03458_),
    .B(_03463_));
 sg13g2_o21ai_1 _12132_ (.B1(_03352_),
    .Y(_03465_),
    .A1(_03340_),
    .A2(_03353_));
 sg13g2_o21ai_1 _12133_ (.B1(_03344_),
    .Y(_03466_),
    .A1(_03345_),
    .A2(_03350_));
 sg13g2_mux2_1 _12134_ (.A0(_00348_),
    .A1(_00347_),
    .S(net4845),
    .X(_03467_));
 sg13g2_nand2b_1 _12135_ (.Y(_03468_),
    .B(_03466_),
    .A_N(_03467_));
 sg13g2_xor2_1 _12136_ (.B(_03467_),
    .A(_03466_),
    .X(_03469_));
 sg13g2_nand2_1 _12137_ (.Y(_03470_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][8] ),
    .B(net4780));
 sg13g2_a22oi_1 _12138_ (.Y(_03471_),
    .B1(net4701),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][8] ),
    .A2(net4784),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][8] ));
 sg13g2_a22oi_1 _12139_ (.Y(_03472_),
    .B1(net4776),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][8] ),
    .A2(net4787),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][8] ));
 sg13g2_nand4_1 _12140_ (.B(_03470_),
    .C(_03471_),
    .A(net4705),
    .Y(_03473_),
    .D(_03472_));
 sg13g2_o21ai_1 _12141_ (.B1(_03473_),
    .Y(_03474_),
    .A1(_02347_),
    .A2(net4705));
 sg13g2_xor2_1 _12142_ (.B(_03474_),
    .A(_03469_),
    .X(_03475_));
 sg13g2_nand2_1 _12143_ (.Y(_03476_),
    .A(_03465_),
    .B(_03475_));
 sg13g2_nor2_1 _12144_ (.A(_03465_),
    .B(_03475_),
    .Y(_03477_));
 sg13g2_xor2_1 _12145_ (.B(_03475_),
    .A(_03465_),
    .X(_03478_));
 sg13g2_xnor2_1 _12146_ (.Y(_03479_),
    .A(_03464_),
    .B(_03478_));
 sg13g2_nand2_1 _12147_ (.Y(_03480_),
    .A(_03448_),
    .B(_03479_));
 sg13g2_xnor2_1 _12148_ (.Y(_03481_),
    .A(_03448_),
    .B(_03479_));
 sg13g2_xnor2_1 _12149_ (.Y(_03482_),
    .A(_03447_),
    .B(_03481_));
 sg13g2_nor2_1 _12150_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .B(net4931),
    .Y(_03483_));
 sg13g2_a21oi_1 _12151_ (.A1(net4930),
    .A2(_03482_),
    .Y(_00285_),
    .B1(_03483_));
 sg13g2_a22oi_1 _12152_ (.Y(_03484_),
    .B1(_02742_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][9] ),
    .A2(net4661),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][9] ));
 sg13g2_a22oi_1 _12153_ (.Y(_03485_),
    .B1(_02738_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][9] ),
    .A2(net4664),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][9] ));
 sg13g2_and2_1 _12154_ (.A(_03484_),
    .B(_03485_),
    .X(_03486_));
 sg13g2_a221oi_1 _12155_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][9] ),
    .C1(net4839),
    .B1(net4731),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][9] ),
    .Y(_03487_),
    .A2(net4810));
 sg13g2_a22oi_1 _12156_ (.Y(_03488_),
    .B1(net4658),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][9] ),
    .A2(net4724),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][9] ));
 sg13g2_nand2_1 _12157_ (.Y(_03489_),
    .A(_03487_),
    .B(_03488_));
 sg13g2_a221oi_1 _12158_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][9] ),
    .C1(_03489_),
    .B1(net4649),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][9] ),
    .Y(_03490_),
    .A2(_02744_));
 sg13g2_a22oi_1 _12159_ (.Y(_03491_),
    .B1(_03486_),
    .B2(_03490_),
    .A2(net4838),
    .A1(_00364_));
 sg13g2_a21oi_1 _12160_ (.A1(_03412_),
    .A2(_03423_),
    .Y(_03492_),
    .B1(_03422_));
 sg13g2_a22oi_1 _12161_ (.Y(_03493_),
    .B1(net4729),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][9] ),
    .A2(net4809),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][9] ));
 sg13g2_a22oi_1 _12162_ (.Y(_03494_),
    .B1(net4734),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][9] ),
    .A2(net4737),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][9] ));
 sg13g2_and2_1 _12163_ (.A(_03493_),
    .B(_03494_),
    .X(_03495_));
 sg13g2_a22oi_1 _12164_ (.Y(_03496_),
    .B1(net4712),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][9] ),
    .A2(net4720),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][9] ));
 sg13g2_a22oi_1 _12165_ (.Y(_03497_),
    .B1(net4740),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][9] ),
    .A2(net4850),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][9] ));
 sg13g2_a22oi_1 _12166_ (.Y(_03498_),
    .B1(net4709),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][9] ),
    .A2(net4715),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][9] ));
 sg13g2_and4_1 _12167_ (.A(net4771),
    .B(_03496_),
    .C(_03497_),
    .D(_03498_),
    .X(_03499_));
 sg13g2_a22oi_1 _12168_ (.Y(_03500_),
    .B1(_03495_),
    .B2(_03499_),
    .A2(net4837),
    .A1(_00363_));
 sg13g2_nor2b_1 _12169_ (.A(_03492_),
    .B_N(_03500_),
    .Y(_03501_));
 sg13g2_xnor2_1 _12170_ (.Y(_03502_),
    .A(_03492_),
    .B(_03500_));
 sg13g2_xnor2_1 _12171_ (.Y(_03503_),
    .A(_03491_),
    .B(_03502_));
 sg13g2_o21ai_1 _12172_ (.B1(_03445_),
    .Y(_03504_),
    .A1(_03424_),
    .A2(_03446_));
 sg13g2_o21ai_1 _12173_ (.B1(_03434_),
    .Y(_03505_),
    .A1(_03435_),
    .A2(_03443_));
 sg13g2_and2_1 _12174_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][9] ),
    .B(net4875),
    .X(_03506_));
 sg13g2_a221oi_1 _12175_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][9] ),
    .C1(_03506_),
    .B1(net4805),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][9] ),
    .Y(_03507_),
    .A2(net4753));
 sg13g2_a221oi_1 _12176_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][9] ),
    .C1(net4831),
    .B1(net4756),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][9] ),
    .Y(_03508_),
    .A2(net4817));
 sg13g2_a22oi_1 _12177_ (.Y(_03509_),
    .B1(net4759),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][9] ),
    .A2(net4764),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][9] ));
 sg13g2_a22oi_1 _12178_ (.Y(_03510_),
    .B1(net4749),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][9] ),
    .A2(net4762),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][9] ));
 sg13g2_and3_1 _12179_ (.X(_03511_),
    .A(_03508_),
    .B(_03509_),
    .C(_03510_));
 sg13g2_a22oi_1 _12180_ (.Y(_03512_),
    .B1(_03507_),
    .B2(_03511_),
    .A2(net4830),
    .A1(_00361_));
 sg13g2_nand2_1 _12181_ (.Y(_03513_),
    .A(_03505_),
    .B(_03512_));
 sg13g2_xnor2_1 _12182_ (.Y(_03514_),
    .A(_03505_),
    .B(_03512_));
 sg13g2_a22oi_1 _12183_ (.Y(_03515_),
    .B1(net4792),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][9] ),
    .A2(net4816),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][9] ));
 sg13g2_a22oi_1 _12184_ (.Y(_03516_),
    .B1(net4846),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][9] ),
    .A2(net4798),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][9] ));
 sg13g2_nand3_1 _12185_ (.B(_03515_),
    .C(_03516_),
    .A(net4770),
    .Y(_03517_));
 sg13g2_a22oi_1 _12186_ (.Y(_03518_),
    .B1(net4744),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][9] ),
    .A2(net4747),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][9] ));
 sg13g2_a22oi_1 _12187_ (.Y(_03519_),
    .B1(net4795),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][9] ),
    .A2(net4804),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][9] ));
 sg13g2_nand2_1 _12188_ (.Y(_03520_),
    .A(_03518_),
    .B(_03519_));
 sg13g2_nand2_1 _12189_ (.Y(_03521_),
    .A(_00362_),
    .B(net4832));
 sg13g2_o21ai_1 _12190_ (.B1(_03521_),
    .Y(_03522_),
    .A1(_03517_),
    .A2(_03520_));
 sg13g2_xor2_1 _12191_ (.B(_03522_),
    .A(_03514_),
    .X(_03523_));
 sg13g2_nand2_1 _12192_ (.Y(_03524_),
    .A(_03504_),
    .B(_03523_));
 sg13g2_xnor2_1 _12193_ (.Y(_03525_),
    .A(_03504_),
    .B(_03523_));
 sg13g2_xnor2_1 _12194_ (.Y(_03526_),
    .A(_03503_),
    .B(_03525_));
 sg13g2_o21ai_1 _12195_ (.B1(_03480_),
    .Y(_03527_),
    .A1(_03447_),
    .A2(_03481_));
 sg13g2_a21oi_2 _12196_ (.B1(_03457_),
    .Y(_03528_),
    .A2(_03463_),
    .A1(_03458_));
 sg13g2_o21ai_1 _12197_ (.B1(net4774),
    .Y(_03529_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][9] ),
    .A2(net4819));
 sg13g2_a22oi_1 _12198_ (.Y(_03530_),
    .B1(net4693),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][9] ),
    .A2(net4695),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][9] ));
 sg13g2_a22oi_1 _12199_ (.Y(_03531_),
    .B1(net4687),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][9] ),
    .A2(net4691),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][9] ));
 sg13g2_a22oi_1 _12200_ (.Y(_03532_),
    .B1(net4689),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][9] ),
    .A2(net4871),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][9] ));
 sg13g2_nand4_1 _12201_ (.B(_03530_),
    .C(_03531_),
    .A(_03529_),
    .Y(_03533_),
    .D(_03532_));
 sg13g2_nand2_1 _12202_ (.Y(_03534_),
    .A(_00359_),
    .B(net4697));
 sg13g2_nand2_2 _12203_ (.Y(_03535_),
    .A(_03533_),
    .B(_03534_));
 sg13g2_nor2_1 _12204_ (.A(_03528_),
    .B(_03535_),
    .Y(_03536_));
 sg13g2_xor2_1 _12205_ (.B(_03535_),
    .A(_03528_),
    .X(_03537_));
 sg13g2_a221oi_1 _12206_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][9] ),
    .C1(net4680),
    .B1(net4669),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][9] ),
    .Y(_03538_),
    .A2(net4676));
 sg13g2_a22oi_1 _12207_ (.Y(_03539_),
    .B1(net4674),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][9] ),
    .A2(net4684),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][9] ));
 sg13g2_a22oi_1 _12208_ (.Y(_03540_),
    .B1(net4667),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][9] ),
    .A2(net4671),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][9] ));
 sg13g2_and2_1 _12209_ (.A(_03539_),
    .B(_03540_),
    .X(_03541_));
 sg13g2_a22oi_1 _12210_ (.Y(_03542_),
    .B1(_03538_),
    .B2(_03541_),
    .A2(net4680),
    .A1(_00360_));
 sg13g2_xnor2_1 _12211_ (.Y(_03543_),
    .A(_03537_),
    .B(_03542_));
 sg13g2_o21ai_1 _12212_ (.B1(_03476_),
    .Y(_03544_),
    .A1(_03464_),
    .A2(_03477_));
 sg13g2_o21ai_1 _12213_ (.B1(_03468_),
    .Y(_03545_),
    .A1(_03469_),
    .A2(_03474_));
 sg13g2_mux2_1 _12214_ (.A0(_00357_),
    .A1(_00356_),
    .S(net4845),
    .X(_03546_));
 sg13g2_nor2b_1 _12215_ (.A(_03546_),
    .B_N(_03545_),
    .Y(_03547_));
 sg13g2_xnor2_1 _12216_ (.Y(_03548_),
    .A(_03545_),
    .B(_03546_));
 sg13g2_and2_1 _12217_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][9] ),
    .B(net4785),
    .X(_03549_));
 sg13g2_a221oi_1 _12218_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][9] ),
    .C1(_03549_),
    .B1(net4701),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][9] ),
    .Y(_03550_),
    .A2(net4780));
 sg13g2_a221oi_1 _12219_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][9] ),
    .C1(net4647),
    .B1(net4776),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][9] ),
    .Y(_03551_),
    .A2(net4788));
 sg13g2_a22oi_1 _12220_ (.Y(_03552_),
    .B1(_03550_),
    .B2(_03551_),
    .A2(net4647),
    .A1(_00358_));
 sg13g2_xor2_1 _12221_ (.B(_03552_),
    .A(_03548_),
    .X(_03553_));
 sg13g2_nand2_1 _12222_ (.Y(_03554_),
    .A(_03544_),
    .B(_03553_));
 sg13g2_nor2_1 _12223_ (.A(_03544_),
    .B(_03553_),
    .Y(_03555_));
 sg13g2_xor2_1 _12224_ (.B(_03553_),
    .A(_03544_),
    .X(_03556_));
 sg13g2_xnor2_1 _12225_ (.Y(_03557_),
    .A(_03543_),
    .B(_03556_));
 sg13g2_nand2_1 _12226_ (.Y(_03558_),
    .A(_03527_),
    .B(_03557_));
 sg13g2_xnor2_1 _12227_ (.Y(_03559_),
    .A(_03527_),
    .B(_03557_));
 sg13g2_xnor2_1 _12228_ (.Y(_03560_),
    .A(_03526_),
    .B(_03559_));
 sg13g2_nor2_1 _12229_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .B(net4929),
    .Y(_03561_));
 sg13g2_a21oi_1 _12230_ (.A1(net4929),
    .A2(_03560_),
    .Y(_00286_),
    .B1(_03561_));
 sg13g2_and2_1 _12231_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][10] ),
    .B(_02738_),
    .X(_03562_));
 sg13g2_a221oi_1 _12232_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][10] ),
    .C1(_03562_),
    .B1(_02742_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][10] ),
    .Y(_03563_),
    .A2(net4662));
 sg13g2_a21oi_1 _12233_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][10] ),
    .A2(net4664),
    .Y(_03564_),
    .B1(net4841));
 sg13g2_a22oi_1 _12234_ (.Y(_03565_),
    .B1(net4652),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][10] ),
    .A2(net4731),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][10] ));
 sg13g2_a22oi_1 _12235_ (.Y(_03566_),
    .B1(net4649),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][10] ),
    .A2(net4811),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][10] ));
 sg13g2_nand3_1 _12236_ (.B(_03565_),
    .C(_03566_),
    .A(_03564_),
    .Y(_03567_));
 sg13g2_a221oi_1 _12237_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][10] ),
    .C1(_03567_),
    .B1(net4658),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][10] ),
    .Y(_03568_),
    .A2(net4724));
 sg13g2_a22oi_1 _12238_ (.Y(_03569_),
    .B1(_03563_),
    .B2(_03568_),
    .A2(net4841),
    .A1(_00371_));
 sg13g2_a21oi_1 _12239_ (.A1(_03491_),
    .A2(_03502_),
    .Y(_03570_),
    .B1(_03501_));
 sg13g2_a22oi_1 _12240_ (.Y(_03571_),
    .B1(net4808),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][10] ),
    .A2(net4850),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][10] ));
 sg13g2_a22oi_1 _12241_ (.Y(_03572_),
    .B1(net4710),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][10] ),
    .A2(net4716),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][10] ));
 sg13g2_and2_1 _12242_ (.A(_03571_),
    .B(_03572_),
    .X(_03573_));
 sg13g2_a22oi_1 _12243_ (.Y(_03574_),
    .B1(net4713),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][10] ),
    .A2(net4738),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][10] ));
 sg13g2_a22oi_1 _12244_ (.Y(_03575_),
    .B1(net4720),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][10] ),
    .A2(net4735),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][10] ));
 sg13g2_a22oi_1 _12245_ (.Y(_03576_),
    .B1(net4728),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][10] ),
    .A2(net4741),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][10] ));
 sg13g2_and4_1 _12246_ (.A(net4771),
    .B(_03574_),
    .C(_03575_),
    .D(_03576_),
    .X(_03577_));
 sg13g2_a22oi_1 _12247_ (.Y(_03578_),
    .B1(_03573_),
    .B2(_03577_),
    .A2(net4836),
    .A1(_00370_));
 sg13g2_nor2b_1 _12248_ (.A(_03570_),
    .B_N(_03578_),
    .Y(_03579_));
 sg13g2_xnor2_1 _12249_ (.Y(_03580_),
    .A(_03570_),
    .B(_03578_));
 sg13g2_xnor2_1 _12250_ (.Y(_03581_),
    .A(_03569_),
    .B(_03580_));
 sg13g2_o21ai_1 _12251_ (.B1(_03524_),
    .Y(_03582_),
    .A1(_03503_),
    .A2(_03525_));
 sg13g2_o21ai_1 _12252_ (.B1(_03513_),
    .Y(_03583_),
    .A1(_03514_),
    .A2(_03522_));
 sg13g2_and2_1 _12253_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][10] ),
    .B(net4765),
    .X(_03584_));
 sg13g2_a221oi_1 _12254_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][10] ),
    .C1(_03584_),
    .B1(net4752),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][10] ),
    .Y(_03585_),
    .A2(net4759));
 sg13g2_a221oi_1 _12255_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][10] ),
    .C1(net4830),
    .B1(net4817),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][10] ),
    .Y(_03586_),
    .A2(net4874));
 sg13g2_a22oi_1 _12256_ (.Y(_03587_),
    .B1(net4749),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][10] ),
    .A2(net4762),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][10] ));
 sg13g2_a22oi_1 _12257_ (.Y(_03588_),
    .B1(net4805),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][10] ),
    .A2(net4756),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][10] ));
 sg13g2_and3_1 _12258_ (.X(_03589_),
    .A(_03586_),
    .B(_03587_),
    .C(_03588_));
 sg13g2_a22oi_1 _12259_ (.Y(_03590_),
    .B1(_03585_),
    .B2(_03589_),
    .A2(net4831),
    .A1(_00368_));
 sg13g2_nand2_1 _12260_ (.Y(_03591_),
    .A(_03583_),
    .B(_03590_));
 sg13g2_xnor2_1 _12261_ (.Y(_03592_),
    .A(_03583_),
    .B(_03590_));
 sg13g2_nand2_1 _12262_ (.Y(_03593_),
    .A(_00369_),
    .B(net4832));
 sg13g2_a22oi_1 _12263_ (.Y(_03594_),
    .B1(net4847),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][10] ),
    .A2(net4744),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][10] ));
 sg13g2_a22oi_1 _12264_ (.Y(_03595_),
    .B1(net4804),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][10] ),
    .A2(net4816),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][10] ));
 sg13g2_nand2_1 _12265_ (.Y(_03596_),
    .A(_03594_),
    .B(_03595_));
 sg13g2_a22oi_1 _12266_ (.Y(_03597_),
    .B1(net4797),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][10] ),
    .A2(net4746),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][10] ));
 sg13g2_a22oi_1 _12267_ (.Y(_03598_),
    .B1(net4792),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][10] ),
    .A2(net4794),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][10] ));
 sg13g2_nand3_1 _12268_ (.B(_03597_),
    .C(_03598_),
    .A(net4769),
    .Y(_03599_));
 sg13g2_o21ai_1 _12269_ (.B1(_03593_),
    .Y(_03600_),
    .A1(_03596_),
    .A2(_03599_));
 sg13g2_xor2_1 _12270_ (.B(_03600_),
    .A(_03592_),
    .X(_03601_));
 sg13g2_nand2_1 _12271_ (.Y(_03602_),
    .A(_03582_),
    .B(_03601_));
 sg13g2_xnor2_1 _12272_ (.Y(_03603_),
    .A(_03582_),
    .B(_03601_));
 sg13g2_xnor2_1 _12273_ (.Y(_03604_),
    .A(_03581_),
    .B(_03603_));
 sg13g2_a21oi_1 _12274_ (.A1(_03537_),
    .A2(_03542_),
    .Y(_03605_),
    .B1(_03536_));
 sg13g2_o21ai_1 _12275_ (.B1(net4774),
    .Y(_03606_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][10] ),
    .A2(net4819));
 sg13g2_a22oi_1 _12276_ (.Y(_03607_),
    .B1(net4693),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][10] ),
    .A2(net4695),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][10] ));
 sg13g2_a22oi_1 _12277_ (.Y(_03608_),
    .B1(net4689),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][10] ),
    .A2(net4691),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][10] ));
 sg13g2_a22oi_1 _12278_ (.Y(_03609_),
    .B1(net4687),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][10] ),
    .A2(net4871),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][10] ));
 sg13g2_nand4_1 _12279_ (.B(_03607_),
    .C(_03608_),
    .A(_03606_),
    .Y(_03610_),
    .D(_03609_));
 sg13g2_nand2_1 _12280_ (.Y(_03611_),
    .A(_00366_),
    .B(net4697));
 sg13g2_nand2_2 _12281_ (.Y(_03612_),
    .A(_03610_),
    .B(_03611_));
 sg13g2_nor2_1 _12282_ (.A(_03605_),
    .B(_03612_),
    .Y(_03613_));
 sg13g2_xor2_1 _12283_ (.B(_03612_),
    .A(_03605_),
    .X(_03614_));
 sg13g2_a221oi_1 _12284_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][10] ),
    .C1(net4680),
    .B1(net4674),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][10] ),
    .Y(_03615_),
    .A2(net4676));
 sg13g2_a22oi_1 _12285_ (.Y(_03616_),
    .B1(net4667),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][10] ),
    .A2(net4669),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][10] ));
 sg13g2_a22oi_1 _12286_ (.Y(_03617_),
    .B1(net4671),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][10] ),
    .A2(net4684),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][10] ));
 sg13g2_and2_1 _12287_ (.A(_03616_),
    .B(_03617_),
    .X(_03618_));
 sg13g2_a22oi_1 _12288_ (.Y(_03619_),
    .B1(_03615_),
    .B2(_03618_),
    .A2(net4679),
    .A1(_00367_));
 sg13g2_xnor2_1 _12289_ (.Y(_03620_),
    .A(_03614_),
    .B(_03619_));
 sg13g2_o21ai_1 _12290_ (.B1(_03554_),
    .Y(_03621_),
    .A1(_03543_),
    .A2(_03555_));
 sg13g2_a21oi_1 _12291_ (.A1(_03548_),
    .A2(_03552_),
    .Y(_03622_),
    .B1(_03547_));
 sg13g2_mux2_1 _12292_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][10] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][10] ),
    .S(net4844),
    .X(_03623_));
 sg13g2_nand2b_1 _12293_ (.Y(_03624_),
    .B(_03623_),
    .A_N(_03622_));
 sg13g2_xor2_1 _12294_ (.B(_03623_),
    .A(_03622_),
    .X(_03625_));
 sg13g2_nand2_1 _12295_ (.Y(_03626_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][10] ),
    .B(net4701));
 sg13g2_a22oi_1 _12296_ (.Y(_03627_),
    .B1(net4780),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][10] ),
    .A2(net4784),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][10] ));
 sg13g2_nand2_1 _12297_ (.Y(_03628_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][10] ),
    .B(net4787));
 sg13g2_nand3_1 _12298_ (.B(_03627_),
    .C(_03628_),
    .A(_03626_),
    .Y(_03629_));
 sg13g2_a221oi_1 _12299_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][10] ),
    .C1(_03629_),
    .B1(net4776),
    .A1(_02348_),
    .Y(_03630_),
    .A2(net4647));
 sg13g2_xor2_1 _12300_ (.B(_03630_),
    .A(_03625_),
    .X(_03631_));
 sg13g2_nand2_1 _12301_ (.Y(_03632_),
    .A(_03621_),
    .B(_03631_));
 sg13g2_nor2_1 _12302_ (.A(_03621_),
    .B(_03631_),
    .Y(_03633_));
 sg13g2_xor2_1 _12303_ (.B(_03631_),
    .A(_03621_),
    .X(_03634_));
 sg13g2_xnor2_1 _12304_ (.Y(_03635_),
    .A(_03620_),
    .B(_03634_));
 sg13g2_o21ai_1 _12305_ (.B1(_03558_),
    .Y(_03636_),
    .A1(_03526_),
    .A2(_03559_));
 sg13g2_nand2_1 _12306_ (.Y(_03637_),
    .A(_03635_),
    .B(_03636_));
 sg13g2_nor2_1 _12307_ (.A(_03635_),
    .B(_03636_),
    .Y(_03638_));
 sg13g2_xor2_1 _12308_ (.B(_03636_),
    .A(_03635_),
    .X(_03639_));
 sg13g2_xnor2_1 _12309_ (.Y(_03640_),
    .A(_03604_),
    .B(_03639_));
 sg13g2_mux2_1 _12310_ (.A0(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .A1(_03640_),
    .S(net4929),
    .X(_00256_));
 sg13g2_and2_1 _12311_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][11] ),
    .B(net4811),
    .X(_03641_));
 sg13g2_a21oi_1 _12312_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][11] ),
    .A2(net4732),
    .Y(_03642_),
    .B1(net4841));
 sg13g2_a22oi_1 _12313_ (.Y(_03643_),
    .B1(net4654),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][11] ),
    .A2(net4664),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][11] ));
 sg13g2_a221oi_1 _12314_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][11] ),
    .C1(_03641_),
    .B1(net4649),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][11] ),
    .Y(_03644_),
    .A2(_02738_));
 sg13g2_a22oi_1 _12315_ (.Y(_03645_),
    .B1(net4652),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][11] ),
    .A2(net4724),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][11] ));
 sg13g2_nand3_1 _12316_ (.B(_03643_),
    .C(_03645_),
    .A(_03642_),
    .Y(_03646_));
 sg13g2_a221oi_1 _12317_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][11] ),
    .C1(_03646_),
    .B1(net4658),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][11] ),
    .Y(_03647_),
    .A2(net4661));
 sg13g2_a22oi_1 _12318_ (.Y(_03648_),
    .B1(_03644_),
    .B2(_03647_),
    .A2(net4841),
    .A1(_00378_));
 sg13g2_a21oi_2 _12319_ (.B1(_03579_),
    .Y(_03649_),
    .A2(_03580_),
    .A1(_03569_));
 sg13g2_a22oi_1 _12320_ (.Y(_03650_),
    .B1(net4738),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][11] ),
    .A2(net4808),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][11] ));
 sg13g2_a22oi_1 _12321_ (.Y(_03651_),
    .B1(net4728),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][11] ),
    .A2(net4740),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][11] ));
 sg13g2_and2_1 _12322_ (.A(_03650_),
    .B(_03651_),
    .X(_03652_));
 sg13g2_a22oi_1 _12323_ (.Y(_03653_),
    .B1(net4712),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][11] ),
    .A2(net4715),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][11] ));
 sg13g2_a22oi_1 _12324_ (.Y(_03654_),
    .B1(net4734),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][11] ),
    .A2(net4849),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][11] ));
 sg13g2_a22oi_1 _12325_ (.Y(_03655_),
    .B1(net4709),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][11] ),
    .A2(net4720),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][11] ));
 sg13g2_and4_1 _12326_ (.A(net4772),
    .B(_03653_),
    .C(_03654_),
    .D(_03655_),
    .X(_03656_));
 sg13g2_a22oi_1 _12327_ (.Y(_03657_),
    .B1(_03652_),
    .B2(_03656_),
    .A2(net4834),
    .A1(_00377_));
 sg13g2_nor2b_1 _12328_ (.A(_03649_),
    .B_N(_03657_),
    .Y(_03658_));
 sg13g2_xnor2_1 _12329_ (.Y(_03659_),
    .A(_03649_),
    .B(_03657_));
 sg13g2_xnor2_1 _12330_ (.Y(_03660_),
    .A(_03648_),
    .B(_03659_));
 sg13g2_o21ai_1 _12331_ (.B1(_03602_),
    .Y(_03661_),
    .A1(_03581_),
    .A2(_03603_));
 sg13g2_o21ai_1 _12332_ (.B1(_03591_),
    .Y(_03662_),
    .A1(_03592_),
    .A2(_03600_));
 sg13g2_and2_1 _12333_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][11] ),
    .B(net4755),
    .X(_03663_));
 sg13g2_a221oi_1 _12334_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][11] ),
    .C1(_03663_),
    .B1(net4758),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][11] ),
    .Y(_03664_),
    .A2(net4764));
 sg13g2_a221oi_1 _12335_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][11] ),
    .C1(net4831),
    .B1(net4817),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][11] ),
    .Y(_03665_),
    .A2(net4761));
 sg13g2_a22oi_1 _12336_ (.Y(_03666_),
    .B1(net4752),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][11] ),
    .A2(net4874),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][11] ));
 sg13g2_a22oi_1 _12337_ (.Y(_03667_),
    .B1(net4750),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][11] ),
    .A2(net4804),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][11] ));
 sg13g2_and3_1 _12338_ (.X(_03668_),
    .A(_03665_),
    .B(_03666_),
    .C(_03667_));
 sg13g2_a22oi_1 _12339_ (.Y(_03669_),
    .B1(_03664_),
    .B2(_03668_),
    .A2(net4830),
    .A1(_00375_));
 sg13g2_nand2_1 _12340_ (.Y(_03670_),
    .A(_03662_),
    .B(_03669_));
 sg13g2_xnor2_1 _12341_ (.Y(_03671_),
    .A(_03662_),
    .B(_03669_));
 sg13g2_a22oi_1 _12342_ (.Y(_03672_),
    .B1(net4746),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][11] ),
    .A2(net4816),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][11] ));
 sg13g2_a22oi_1 _12343_ (.Y(_03673_),
    .B1(net4794),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][11] ),
    .A2(net4804),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][11] ));
 sg13g2_nand2_1 _12344_ (.Y(_03674_),
    .A(_03672_),
    .B(_03673_));
 sg13g2_a22oi_1 _12345_ (.Y(_03675_),
    .B1(net4846),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][11] ),
    .A2(net4797),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][11] ));
 sg13g2_a22oi_1 _12346_ (.Y(_03676_),
    .B1(net4791),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][11] ),
    .A2(net4743),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][11] ));
 sg13g2_nand3_1 _12347_ (.B(_03675_),
    .C(_03676_),
    .A(net4769),
    .Y(_03677_));
 sg13g2_nand2_1 _12348_ (.Y(_03678_),
    .A(_00376_),
    .B(net4832));
 sg13g2_o21ai_1 _12349_ (.B1(_03678_),
    .Y(_03679_),
    .A1(_03674_),
    .A2(_03677_));
 sg13g2_xor2_1 _12350_ (.B(_03679_),
    .A(_03671_),
    .X(_03680_));
 sg13g2_nand2_1 _12351_ (.Y(_03681_),
    .A(_03661_),
    .B(_03680_));
 sg13g2_xnor2_1 _12352_ (.Y(_03682_),
    .A(_03661_),
    .B(_03680_));
 sg13g2_xnor2_1 _12353_ (.Y(_03683_),
    .A(_03660_),
    .B(_03682_));
 sg13g2_a21oi_1 _12354_ (.A1(_03614_),
    .A2(_03619_),
    .Y(_03684_),
    .B1(_03613_));
 sg13g2_nand2_1 _12355_ (.Y(_03685_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][11] ),
    .B(net4696));
 sg13g2_a221oi_1 _12356_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][11] ),
    .C1(net4698),
    .B1(_02848_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][11] ),
    .Y(_03686_),
    .A2(net4694));
 sg13g2_a22oi_1 _12357_ (.Y(_03687_),
    .B1(net4688),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][11] ),
    .A2(net4692),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][11] ));
 sg13g2_a22oi_1 _12358_ (.Y(_03688_),
    .B1(net4690),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][11] ),
    .A2(net4872),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][11] ));
 sg13g2_nand4_1 _12359_ (.B(_03686_),
    .C(_03687_),
    .A(_03685_),
    .Y(_03689_),
    .D(_03688_));
 sg13g2_nand2_1 _12360_ (.Y(_03690_),
    .A(_00373_),
    .B(net4697));
 sg13g2_nand2_1 _12361_ (.Y(_03691_),
    .A(_03689_),
    .B(_03690_));
 sg13g2_nor2_1 _12362_ (.A(_03684_),
    .B(_03691_),
    .Y(_03692_));
 sg13g2_xor2_1 _12363_ (.B(_03691_),
    .A(_03684_),
    .X(_03693_));
 sg13g2_a221oi_1 _12364_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][11] ),
    .C1(net4679),
    .B1(net4669),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][11] ),
    .Y(_03694_),
    .A2(net4676));
 sg13g2_a22oi_1 _12365_ (.Y(_03695_),
    .B1(net4667),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][11] ),
    .A2(net4671),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][11] ));
 sg13g2_a22oi_1 _12366_ (.Y(_03696_),
    .B1(net4674),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][11] ),
    .A2(net4684),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][11] ));
 sg13g2_and2_1 _12367_ (.A(_03695_),
    .B(_03696_),
    .X(_03697_));
 sg13g2_a22oi_1 _12368_ (.Y(_03698_),
    .B1(_03694_),
    .B2(_03697_),
    .A2(net4679),
    .A1(_00374_));
 sg13g2_xnor2_1 _12369_ (.Y(_03699_),
    .A(_03693_),
    .B(_03698_));
 sg13g2_o21ai_1 _12370_ (.B1(_03632_),
    .Y(_03700_),
    .A1(_03620_),
    .A2(_03633_));
 sg13g2_o21ai_1 _12371_ (.B1(_03624_),
    .Y(_03701_),
    .A1(_03625_),
    .A2(_03630_));
 sg13g2_mux2_1 _12372_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][11] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][11] ),
    .S(net4844),
    .X(_03702_));
 sg13g2_nand2_1 _12373_ (.Y(_03703_),
    .A(_03701_),
    .B(_03702_));
 sg13g2_nor2_1 _12374_ (.A(_03701_),
    .B(_03702_),
    .Y(_03704_));
 sg13g2_xor2_1 _12375_ (.B(_03702_),
    .A(_03701_),
    .X(_03705_));
 sg13g2_nand2_1 _12376_ (.Y(_03706_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][11] ),
    .B(net4701));
 sg13g2_a22oi_1 _12377_ (.Y(_03707_),
    .B1(net4780),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][11] ),
    .A2(net4784),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][11] ));
 sg13g2_a22oi_1 _12378_ (.Y(_03708_),
    .B1(net4776),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][11] ),
    .A2(net4787),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][11] ));
 sg13g2_nand4_1 _12379_ (.B(_03706_),
    .C(_03707_),
    .A(net4705),
    .Y(_03709_),
    .D(_03708_));
 sg13g2_o21ai_1 _12380_ (.B1(_03709_),
    .Y(_03710_),
    .A1(_02349_),
    .A2(net4705));
 sg13g2_xnor2_1 _12381_ (.Y(_03711_),
    .A(_03705_),
    .B(_03710_));
 sg13g2_nand2_1 _12382_ (.Y(_03712_),
    .A(_03700_),
    .B(_03711_));
 sg13g2_nor2_1 _12383_ (.A(_03700_),
    .B(_03711_),
    .Y(_03713_));
 sg13g2_xor2_1 _12384_ (.B(_03711_),
    .A(_03700_),
    .X(_03714_));
 sg13g2_xnor2_1 _12385_ (.Y(_03715_),
    .A(_03699_),
    .B(_03714_));
 sg13g2_o21ai_1 _12386_ (.B1(_03637_),
    .Y(_03716_),
    .A1(_03604_),
    .A2(_03638_));
 sg13g2_nand2_1 _12387_ (.Y(_03717_),
    .A(_03715_),
    .B(_03716_));
 sg13g2_nor2_1 _12388_ (.A(_03715_),
    .B(_03716_),
    .Y(_03718_));
 sg13g2_xor2_1 _12389_ (.B(_03716_),
    .A(_03715_),
    .X(_03719_));
 sg13g2_xnor2_1 _12390_ (.Y(_03720_),
    .A(_03683_),
    .B(_03719_));
 sg13g2_mux2_1 _12391_ (.A0(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .A1(_03720_),
    .S(net4930),
    .X(_00257_));
 sg13g2_and2_1 _12392_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][12] ),
    .B(net4723),
    .X(_03721_));
 sg13g2_a22oi_1 _12393_ (.Y(_03722_),
    .B1(net4661),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][12] ),
    .A2(net4664),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][12] ));
 sg13g2_a221oi_1 _12394_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][12] ),
    .C1(_03721_),
    .B1(net4649),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][12] ),
    .Y(_03723_),
    .A2(net4658));
 sg13g2_a21oi_1 _12395_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][12] ),
    .A2(net4652),
    .Y(_03724_),
    .B1(net4840));
 sg13g2_a22oi_1 _12396_ (.Y(_03725_),
    .B1(net4654),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][12] ),
    .A2(net4731),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][12] ));
 sg13g2_nand3_1 _12397_ (.B(_03724_),
    .C(_03725_),
    .A(_03722_),
    .Y(_03726_));
 sg13g2_a221oi_1 _12398_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][12] ),
    .C1(_03726_),
    .B1(net4656),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][12] ),
    .Y(_03727_),
    .A2(net4810));
 sg13g2_a22oi_1 _12399_ (.Y(_03728_),
    .B1(_03723_),
    .B2(_03727_),
    .A2(net4840),
    .A1(_00387_));
 sg13g2_a21oi_1 _12400_ (.A1(_03648_),
    .A2(_03659_),
    .Y(_03729_),
    .B1(_03658_));
 sg13g2_a22oi_1 _12401_ (.Y(_03730_),
    .B1(net4728),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][12] ),
    .A2(net4809),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][12] ));
 sg13g2_a22oi_1 _12402_ (.Y(_03731_),
    .B1(net4709),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][12] ),
    .A2(net4720),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][12] ));
 sg13g2_and2_1 _12403_ (.A(_03730_),
    .B(_03731_),
    .X(_03732_));
 sg13g2_a22oi_1 _12404_ (.Y(_03733_),
    .B1(net4712),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][12] ),
    .A2(net4715),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][12] ));
 sg13g2_a22oi_1 _12405_ (.Y(_03734_),
    .B1(net4734),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][12] ),
    .A2(net4740),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][12] ));
 sg13g2_a22oi_1 _12406_ (.Y(_03735_),
    .B1(net4737),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][12] ),
    .A2(net4849),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][12] ));
 sg13g2_and4_1 _12407_ (.A(net4772),
    .B(_03733_),
    .C(_03734_),
    .D(_03735_),
    .X(_03736_));
 sg13g2_a22oi_1 _12408_ (.Y(_03737_),
    .B1(_03732_),
    .B2(_03736_),
    .A2(net4835),
    .A1(_00386_));
 sg13g2_nor2b_1 _12409_ (.A(_03729_),
    .B_N(_03737_),
    .Y(_03738_));
 sg13g2_xnor2_1 _12410_ (.Y(_03739_),
    .A(_03729_),
    .B(_03737_));
 sg13g2_xnor2_1 _12411_ (.Y(_03740_),
    .A(_03728_),
    .B(_03739_));
 sg13g2_o21ai_1 _12412_ (.B1(_03681_),
    .Y(_03741_),
    .A1(_03660_),
    .A2(_03682_));
 sg13g2_o21ai_1 _12413_ (.B1(_03670_),
    .Y(_03742_),
    .A1(_03671_),
    .A2(_03679_));
 sg13g2_and2_1 _12414_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][12] ),
    .B(net4764),
    .X(_03743_));
 sg13g2_a221oi_1 _12415_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][12] ),
    .C1(_03743_),
    .B1(net4758),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][12] ),
    .Y(_03744_),
    .A2(net4761));
 sg13g2_a221oi_1 _12416_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][12] ),
    .C1(net4830),
    .B1(net4752),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][12] ),
    .Y(_03745_),
    .A2(net4817));
 sg13g2_a22oi_1 _12417_ (.Y(_03746_),
    .B1(net4805),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][12] ),
    .A2(net4874),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][12] ));
 sg13g2_a22oi_1 _12418_ (.Y(_03747_),
    .B1(net4749),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][12] ),
    .A2(net4755),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][12] ));
 sg13g2_and3_1 _12419_ (.X(_03748_),
    .A(_03745_),
    .B(_03746_),
    .C(_03747_));
 sg13g2_a22oi_1 _12420_ (.Y(_03749_),
    .B1(_03744_),
    .B2(_03748_),
    .A2(net4830),
    .A1(_00384_));
 sg13g2_nand2_1 _12421_ (.Y(_03750_),
    .A(_03742_),
    .B(_03749_));
 sg13g2_xnor2_1 _12422_ (.Y(_03751_),
    .A(_03742_),
    .B(_03749_));
 sg13g2_a22oi_1 _12423_ (.Y(_03752_),
    .B1(net4846),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][12] ),
    .A2(net4816),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][12] ));
 sg13g2_a22oi_1 _12424_ (.Y(_03753_),
    .B1(net4791),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][12] ),
    .A2(net4797),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][12] ));
 sg13g2_nand3_1 _12425_ (.B(_03752_),
    .C(_03753_),
    .A(net4769),
    .Y(_03754_));
 sg13g2_a22oi_1 _12426_ (.Y(_03755_),
    .B1(net4794),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][12] ),
    .A2(net4743),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][12] ));
 sg13g2_a22oi_1 _12427_ (.Y(_03756_),
    .B1(net4746),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][12] ),
    .A2(net4804),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][12] ));
 sg13g2_nand2_1 _12428_ (.Y(_03757_),
    .A(_03755_),
    .B(_03756_));
 sg13g2_nand2_1 _12429_ (.Y(_03758_),
    .A(_00385_),
    .B(net4832));
 sg13g2_o21ai_1 _12430_ (.B1(_03758_),
    .Y(_03759_),
    .A1(_03754_),
    .A2(_03757_));
 sg13g2_xor2_1 _12431_ (.B(_03759_),
    .A(_03751_),
    .X(_03760_));
 sg13g2_nand2_1 _12432_ (.Y(_03761_),
    .A(_03741_),
    .B(_03760_));
 sg13g2_xnor2_1 _12433_ (.Y(_03762_),
    .A(_03741_),
    .B(_03760_));
 sg13g2_xnor2_1 _12434_ (.Y(_03763_),
    .A(_03740_),
    .B(_03762_));
 sg13g2_a21oi_1 _12435_ (.A1(_03693_),
    .A2(_03698_),
    .Y(_03764_),
    .B1(_03692_));
 sg13g2_o21ai_1 _12436_ (.B1(net4774),
    .Y(_03765_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][12] ),
    .A2(net4819));
 sg13g2_a22oi_1 _12437_ (.Y(_03766_),
    .B1(net4693),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][12] ),
    .A2(net4695),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][12] ));
 sg13g2_a22oi_1 _12438_ (.Y(_03767_),
    .B1(net4691),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][12] ),
    .A2(net4871),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][12] ));
 sg13g2_a22oi_1 _12439_ (.Y(_03768_),
    .B1(net4687),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][12] ),
    .A2(net4689),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][12] ));
 sg13g2_nand4_1 _12440_ (.B(_03766_),
    .C(_03767_),
    .A(_03765_),
    .Y(_03769_),
    .D(_03768_));
 sg13g2_nand2_1 _12441_ (.Y(_03770_),
    .A(_00382_),
    .B(net4697));
 sg13g2_nand2_1 _12442_ (.Y(_03771_),
    .A(_03769_),
    .B(_03770_));
 sg13g2_nor2_1 _12443_ (.A(_03764_),
    .B(_03771_),
    .Y(_03772_));
 sg13g2_xor2_1 _12444_ (.B(_03771_),
    .A(_03764_),
    .X(_03773_));
 sg13g2_a221oi_1 _12445_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][12] ),
    .C1(net4678),
    .B1(net4671),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][12] ),
    .Y(_03774_),
    .A2(net4676));
 sg13g2_a22oi_1 _12446_ (.Y(_03775_),
    .B1(net4669),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][12] ),
    .A2(net4684),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][12] ));
 sg13g2_a22oi_1 _12447_ (.Y(_03776_),
    .B1(net4667),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][12] ),
    .A2(net4674),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][12] ));
 sg13g2_and2_1 _12448_ (.A(_03775_),
    .B(_03776_),
    .X(_03777_));
 sg13g2_a22oi_1 _12449_ (.Y(_03778_),
    .B1(_03774_),
    .B2(_03777_),
    .A2(net4678),
    .A1(_00383_));
 sg13g2_xnor2_1 _12450_ (.Y(_03779_),
    .A(_03773_),
    .B(_03778_));
 sg13g2_o21ai_1 _12451_ (.B1(_03712_),
    .Y(_03780_),
    .A1(_03699_),
    .A2(_03713_));
 sg13g2_o21ai_1 _12452_ (.B1(_03703_),
    .Y(_03781_),
    .A1(_03704_),
    .A2(_03710_));
 sg13g2_mux2_1 _12453_ (.A0(_00380_),
    .A1(_00379_),
    .S(net4845),
    .X(_03782_));
 sg13g2_nor2b_1 _12454_ (.A(_03782_),
    .B_N(_03781_),
    .Y(_03783_));
 sg13g2_nand2b_1 _12455_ (.Y(_03784_),
    .B(_03782_),
    .A_N(_03781_));
 sg13g2_xor2_1 _12456_ (.B(_03782_),
    .A(_03781_),
    .X(_03785_));
 sg13g2_and2_1 _12457_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][12] ),
    .B(net4786),
    .X(_03786_));
 sg13g2_a221oi_1 _12458_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][12] ),
    .C1(_03786_),
    .B1(net4704),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][12] ),
    .Y(_03787_),
    .A2(net4782));
 sg13g2_a221oi_1 _12459_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][12] ),
    .C1(net4648),
    .B1(net4778),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][12] ),
    .Y(_03788_),
    .A2(net4789));
 sg13g2_a22oi_1 _12460_ (.Y(_03789_),
    .B1(_03787_),
    .B2(_03788_),
    .A2(net4648),
    .A1(_00381_));
 sg13g2_xnor2_1 _12461_ (.Y(_03790_),
    .A(_03785_),
    .B(_03789_));
 sg13g2_nand2_1 _12462_ (.Y(_03791_),
    .A(_03780_),
    .B(_03790_));
 sg13g2_nor2_1 _12463_ (.A(_03780_),
    .B(_03790_),
    .Y(_03792_));
 sg13g2_xor2_1 _12464_ (.B(_03790_),
    .A(_03780_),
    .X(_03793_));
 sg13g2_xnor2_1 _12465_ (.Y(_03794_),
    .A(_03779_),
    .B(_03793_));
 sg13g2_o21ai_1 _12466_ (.B1(_03717_),
    .Y(_03795_),
    .A1(_03683_),
    .A2(_03718_));
 sg13g2_nand2_1 _12467_ (.Y(_03796_),
    .A(_03794_),
    .B(_03795_));
 sg13g2_nor2_1 _12468_ (.A(_03794_),
    .B(_03795_),
    .Y(_03797_));
 sg13g2_xor2_1 _12469_ (.B(_03795_),
    .A(_03794_),
    .X(_03798_));
 sg13g2_xnor2_1 _12470_ (.Y(_03799_),
    .A(_03763_),
    .B(_03798_));
 sg13g2_mux2_1 _12471_ (.A0(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .A1(_03799_),
    .S(net4930),
    .X(_00258_));
 sg13g2_and2_1 _12472_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][13] ),
    .B(net4723),
    .X(_03800_));
 sg13g2_a221oi_1 _12473_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][13] ),
    .C1(_03800_),
    .B1(net4649),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][13] ),
    .Y(_03801_),
    .A2(net4811));
 sg13g2_a21oi_1 _12474_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][13] ),
    .A2(net4661),
    .Y(_03802_),
    .B1(net4840));
 sg13g2_a22oi_1 _12475_ (.Y(_03803_),
    .B1(net4654),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][13] ),
    .A2(net4731),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][13] ));
 sg13g2_a22oi_1 _12476_ (.Y(_03804_),
    .B1(net4656),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][13] ),
    .A2(net4664),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][13] ));
 sg13g2_nand3_1 _12477_ (.B(_03803_),
    .C(_03804_),
    .A(_03802_),
    .Y(_03805_));
 sg13g2_a221oi_1 _12478_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][13] ),
    .C1(_03805_),
    .B1(net4652),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][13] ),
    .Y(_03806_),
    .A2(net4658));
 sg13g2_a22oi_1 _12479_ (.Y(_03807_),
    .B1(_03801_),
    .B2(_03806_),
    .A2(net4840),
    .A1(_00396_));
 sg13g2_a21oi_2 _12480_ (.B1(_03738_),
    .Y(_03808_),
    .A2(_03739_),
    .A1(_03728_));
 sg13g2_a22oi_1 _12481_ (.Y(_03809_),
    .B1(net4734),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][13] ),
    .A2(net4809),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][13] ));
 sg13g2_a22oi_1 _12482_ (.Y(_03810_),
    .B1(net4709),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][13] ),
    .A2(net4849),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][13] ));
 sg13g2_and2_1 _12483_ (.A(_03809_),
    .B(_03810_),
    .X(_03811_));
 sg13g2_a22oi_1 _12484_ (.Y(_03812_),
    .B1(net4712),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][13] ),
    .A2(net4733),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][13] ));
 sg13g2_a22oi_1 _12485_ (.Y(_03813_),
    .B1(net4715),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][13] ),
    .A2(net4737),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][13] ));
 sg13g2_a22oi_1 _12486_ (.Y(_03814_),
    .B1(net4725),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][13] ),
    .A2(net4740),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][13] ));
 sg13g2_and4_1 _12487_ (.A(net4772),
    .B(_03812_),
    .C(_03813_),
    .D(_03814_),
    .X(_03815_));
 sg13g2_a22oi_1 _12488_ (.Y(_03816_),
    .B1(_03811_),
    .B2(_03815_),
    .A2(net4835),
    .A1(_00395_));
 sg13g2_nor2b_1 _12489_ (.A(_03808_),
    .B_N(_03816_),
    .Y(_03817_));
 sg13g2_xnor2_1 _12490_ (.Y(_03818_),
    .A(_03808_),
    .B(_03816_));
 sg13g2_xnor2_1 _12491_ (.Y(_03819_),
    .A(_03807_),
    .B(_03818_));
 sg13g2_o21ai_1 _12492_ (.B1(_03761_),
    .Y(_03820_),
    .A1(_03740_),
    .A2(_03762_));
 sg13g2_o21ai_1 _12493_ (.B1(_03750_),
    .Y(_03821_),
    .A1(_03751_),
    .A2(_03759_));
 sg13g2_and2_1 _12494_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][13] ),
    .B(net4755),
    .X(_03822_));
 sg13g2_a221oi_1 _12495_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][13] ),
    .C1(_03822_),
    .B1(net4749),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][13] ),
    .Y(_03823_),
    .A2(net4758));
 sg13g2_a221oi_1 _12496_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][13] ),
    .C1(net4828),
    .B1(net4817),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][13] ),
    .Y(_03824_),
    .A2(net4761));
 sg13g2_a22oi_1 _12497_ (.Y(_03825_),
    .B1(net4806),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][13] ),
    .A2(net4874),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][13] ));
 sg13g2_a22oi_1 _12498_ (.Y(_03826_),
    .B1(net4752),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][13] ),
    .A2(net4764),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][13] ));
 sg13g2_and3_1 _12499_ (.X(_03827_),
    .A(_03824_),
    .B(_03825_),
    .C(_03826_));
 sg13g2_a22oi_1 _12500_ (.Y(_03828_),
    .B1(_03823_),
    .B2(_03827_),
    .A2(net4828),
    .A1(_00393_));
 sg13g2_nand2_1 _12501_ (.Y(_03829_),
    .A(_03821_),
    .B(_03828_));
 sg13g2_xnor2_1 _12502_ (.Y(_03830_),
    .A(_03821_),
    .B(_03828_));
 sg13g2_nand2_1 _12503_ (.Y(_03831_),
    .A(_00394_),
    .B(net4829));
 sg13g2_a22oi_1 _12504_ (.Y(_03832_),
    .B1(net4846),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][13] ),
    .A2(net4791),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][13] ));
 sg13g2_a22oi_1 _12505_ (.Y(_03833_),
    .B1(net4797),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][13] ),
    .A2(net4816),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][13] ));
 sg13g2_nand3_1 _12506_ (.B(_03832_),
    .C(_03833_),
    .A(net4769),
    .Y(_03834_));
 sg13g2_a22oi_1 _12507_ (.Y(_03835_),
    .B1(net4743),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][13] ),
    .A2(net4746),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][13] ));
 sg13g2_a22oi_1 _12508_ (.Y(_03836_),
    .B1(net4794),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][13] ),
    .A2(net4804),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][13] ));
 sg13g2_nand2_1 _12509_ (.Y(_03837_),
    .A(_03835_),
    .B(_03836_));
 sg13g2_o21ai_1 _12510_ (.B1(_03831_),
    .Y(_03838_),
    .A1(_03834_),
    .A2(_03837_));
 sg13g2_xor2_1 _12511_ (.B(_03838_),
    .A(_03830_),
    .X(_03839_));
 sg13g2_nand2_1 _12512_ (.Y(_03840_),
    .A(_03820_),
    .B(_03839_));
 sg13g2_xnor2_1 _12513_ (.Y(_03841_),
    .A(_03820_),
    .B(_03839_));
 sg13g2_xnor2_1 _12514_ (.Y(_03842_),
    .A(_03819_),
    .B(_03841_));
 sg13g2_a21oi_1 _12515_ (.A1(_03773_),
    .A2(_03778_),
    .Y(_03843_),
    .B1(_03772_));
 sg13g2_o21ai_1 _12516_ (.B1(net4774),
    .Y(_03844_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][13] ),
    .A2(net4819));
 sg13g2_a22oi_1 _12517_ (.Y(_03845_),
    .B1(net4693),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][13] ),
    .A2(net4695),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][13] ));
 sg13g2_a22oi_1 _12518_ (.Y(_03846_),
    .B1(net4687),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][13] ),
    .A2(net4871),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][13] ));
 sg13g2_a22oi_1 _12519_ (.Y(_03847_),
    .B1(net4689),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][13] ),
    .A2(net4691),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][13] ));
 sg13g2_nand4_1 _12520_ (.B(_03845_),
    .C(_03846_),
    .A(_03844_),
    .Y(_03848_),
    .D(_03847_));
 sg13g2_nand2_1 _12521_ (.Y(_03849_),
    .A(_00391_),
    .B(net4697));
 sg13g2_nand2_1 _12522_ (.Y(_03850_),
    .A(_03848_),
    .B(_03849_));
 sg13g2_nor2_1 _12523_ (.A(_03843_),
    .B(_03850_),
    .Y(_03851_));
 sg13g2_xor2_1 _12524_ (.B(_03850_),
    .A(_03843_),
    .X(_03852_));
 sg13g2_a221oi_1 _12525_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][13] ),
    .C1(net4678),
    .B1(net4669),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][13] ),
    .Y(_03853_),
    .A2(net4676));
 sg13g2_a22oi_1 _12526_ (.Y(_03854_),
    .B1(net4671),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][13] ),
    .A2(net4684),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][13] ));
 sg13g2_a22oi_1 _12527_ (.Y(_03855_),
    .B1(net4667),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][13] ),
    .A2(net4674),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][13] ));
 sg13g2_and2_1 _12528_ (.A(_03854_),
    .B(_03855_),
    .X(_03856_));
 sg13g2_a22oi_1 _12529_ (.Y(_03857_),
    .B1(_03853_),
    .B2(_03856_),
    .A2(net4678),
    .A1(_00392_));
 sg13g2_xnor2_1 _12530_ (.Y(_03858_),
    .A(_03852_),
    .B(_03857_));
 sg13g2_o21ai_1 _12531_ (.B1(_03791_),
    .Y(_03859_),
    .A1(_03779_),
    .A2(_03792_));
 sg13g2_a21oi_1 _12532_ (.A1(_03784_),
    .A2(_03789_),
    .Y(_03860_),
    .B1(_03783_));
 sg13g2_mux2_1 _12533_ (.A0(_00389_),
    .A1(_00388_),
    .S(net4844),
    .X(_03861_));
 sg13g2_nor2_1 _12534_ (.A(_03860_),
    .B(_03861_),
    .Y(_03862_));
 sg13g2_xor2_1 _12535_ (.B(_03861_),
    .A(_03860_),
    .X(_03863_));
 sg13g2_and2_1 _12536_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][13] ),
    .B(net4786),
    .X(_03864_));
 sg13g2_a221oi_1 _12537_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][13] ),
    .C1(_03864_),
    .B1(net4704),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][13] ),
    .Y(_03865_),
    .A2(net4782));
 sg13g2_a221oi_1 _12538_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][13] ),
    .C1(net4648),
    .B1(net4778),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][13] ),
    .Y(_03866_),
    .A2(net4789));
 sg13g2_a22oi_1 _12539_ (.Y(_03867_),
    .B1(_03865_),
    .B2(_03866_),
    .A2(net4648),
    .A1(_00390_));
 sg13g2_xor2_1 _12540_ (.B(_03867_),
    .A(_03863_),
    .X(_03868_));
 sg13g2_nand2_1 _12541_ (.Y(_03869_),
    .A(_03859_),
    .B(_03868_));
 sg13g2_nor2_1 _12542_ (.A(_03859_),
    .B(_03868_),
    .Y(_03870_));
 sg13g2_xor2_1 _12543_ (.B(_03868_),
    .A(_03859_),
    .X(_03871_));
 sg13g2_xnor2_1 _12544_ (.Y(_03872_),
    .A(_03858_),
    .B(_03871_));
 sg13g2_o21ai_1 _12545_ (.B1(_03796_),
    .Y(_03873_),
    .A1(_03763_),
    .A2(_03797_));
 sg13g2_nand2_1 _12546_ (.Y(_03874_),
    .A(_03872_),
    .B(_03873_));
 sg13g2_nor2_1 _12547_ (.A(_03872_),
    .B(_03873_),
    .Y(_03875_));
 sg13g2_xnor2_1 _12548_ (.Y(_03876_),
    .A(_03872_),
    .B(_03873_));
 sg13g2_xnor2_1 _12549_ (.Y(_03877_),
    .A(_03842_),
    .B(_03876_));
 sg13g2_nor2_1 _12550_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .B(net4930),
    .Y(_03878_));
 sg13g2_a21oi_1 _12551_ (.A1(net4930),
    .A2(_03877_),
    .Y(_00259_),
    .B1(_03878_));
 sg13g2_a21oi_1 _12552_ (.A1(_03852_),
    .A2(_03857_),
    .Y(_03879_),
    .B1(_03851_));
 sg13g2_o21ai_1 _12553_ (.B1(net4774),
    .Y(_03880_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][14] ),
    .A2(net4819));
 sg13g2_a22oi_1 _12554_ (.Y(_03881_),
    .B1(net4693),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][14] ),
    .A2(net4695),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][14] ));
 sg13g2_a22oi_1 _12555_ (.Y(_03882_),
    .B1(net4689),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][14] ),
    .A2(net4691),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][14] ));
 sg13g2_a22oi_1 _12556_ (.Y(_03883_),
    .B1(net4687),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][14] ),
    .A2(net4871),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][14] ));
 sg13g2_nand4_1 _12557_ (.B(_03881_),
    .C(_03882_),
    .A(_03880_),
    .Y(_03884_),
    .D(_03883_));
 sg13g2_nand2_1 _12558_ (.Y(_03885_),
    .A(_00398_),
    .B(net4697));
 sg13g2_nand2_1 _12559_ (.Y(_03886_),
    .A(_03884_),
    .B(_03885_));
 sg13g2_nor2_1 _12560_ (.A(_03879_),
    .B(_03886_),
    .Y(_03887_));
 sg13g2_xor2_1 _12561_ (.B(_03886_),
    .A(_03879_),
    .X(_03888_));
 sg13g2_a221oi_1 _12562_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][14] ),
    .C1(net4678),
    .B1(net4669),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][14] ),
    .Y(_03889_),
    .A2(net4676));
 sg13g2_a22oi_1 _12563_ (.Y(_03890_),
    .B1(net4667),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][14] ),
    .A2(net4671),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][14] ));
 sg13g2_a22oi_1 _12564_ (.Y(_03891_),
    .B1(net4674),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][14] ),
    .A2(net4684),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][14] ));
 sg13g2_and2_1 _12565_ (.A(_03890_),
    .B(_03891_),
    .X(_03892_));
 sg13g2_a22oi_1 _12566_ (.Y(_03893_),
    .B1(_03889_),
    .B2(_03892_),
    .A2(net4678),
    .A1(_00399_));
 sg13g2_xnor2_1 _12567_ (.Y(_03894_),
    .A(_03888_),
    .B(_03893_));
 sg13g2_o21ai_1 _12568_ (.B1(_03869_),
    .Y(_03895_),
    .A1(_03858_),
    .A2(_03870_));
 sg13g2_a21oi_1 _12569_ (.A1(_03863_),
    .A2(_03867_),
    .Y(_03896_),
    .B1(_03862_));
 sg13g2_mux2_1 _12570_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][14] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][14] ),
    .S(net4844),
    .X(_03897_));
 sg13g2_nand2b_1 _12571_ (.Y(_03898_),
    .B(_03897_),
    .A_N(_03896_));
 sg13g2_xor2_1 _12572_ (.B(_03897_),
    .A(_03896_),
    .X(_03899_));
 sg13g2_nand2_1 _12573_ (.Y(_03900_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][14] ),
    .B(net4783));
 sg13g2_a22oi_1 _12574_ (.Y(_03901_),
    .B1(net4704),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][14] ),
    .A2(net4786),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][14] ));
 sg13g2_a22oi_1 _12575_ (.Y(_03902_),
    .B1(net4779),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][14] ),
    .A2(net4790),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][14] ));
 sg13g2_nand4_1 _12576_ (.B(_03900_),
    .C(_03901_),
    .A(net4708),
    .Y(_03903_),
    .D(_03902_));
 sg13g2_o21ai_1 _12577_ (.B1(_03903_),
    .Y(_03904_),
    .A1(_02350_),
    .A2(net4708));
 sg13g2_xor2_1 _12578_ (.B(_03904_),
    .A(_03899_),
    .X(_03905_));
 sg13g2_nand2_1 _12579_ (.Y(_03906_),
    .A(_03895_),
    .B(_03905_));
 sg13g2_nor2_1 _12580_ (.A(_03895_),
    .B(_03905_),
    .Y(_03907_));
 sg13g2_xor2_1 _12581_ (.B(_03905_),
    .A(_03895_),
    .X(_03908_));
 sg13g2_xnor2_1 _12582_ (.Y(_03909_),
    .A(_03894_),
    .B(_03908_));
 sg13g2_o21ai_1 _12583_ (.B1(_03874_),
    .Y(_03910_),
    .A1(_03842_),
    .A2(_03875_));
 sg13g2_and2_1 _12584_ (.A(_03909_),
    .B(_03910_),
    .X(_03911_));
 sg13g2_xor2_1 _12585_ (.B(_03910_),
    .A(_03909_),
    .X(_03912_));
 sg13g2_and2_1 _12586_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][14] ),
    .B(net4811),
    .X(_03913_));
 sg13g2_a221oi_1 _12587_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][14] ),
    .C1(_03913_),
    .B1(net4654),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][14] ),
    .Y(_03914_),
    .A2(net4658));
 sg13g2_a21oi_1 _12588_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][14] ),
    .A2(net4664),
    .Y(_03915_),
    .B1(net4840));
 sg13g2_a22oi_1 _12589_ (.Y(_03916_),
    .B1(net4652),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][14] ),
    .A2(net4723),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][14] ));
 sg13g2_a22oi_1 _12590_ (.Y(_03917_),
    .B1(net4656),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][14] ),
    .A2(net4732),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][14] ));
 sg13g2_nand3_1 _12591_ (.B(_03916_),
    .C(_03917_),
    .A(_03915_),
    .Y(_03918_));
 sg13g2_a221oi_1 _12592_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][14] ),
    .C1(_03918_),
    .B1(net4649),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][14] ),
    .Y(_03919_),
    .A2(net4662));
 sg13g2_a22oi_1 _12593_ (.Y(_03920_),
    .B1(_03914_),
    .B2(_03919_),
    .A2(net4840),
    .A1(_00403_));
 sg13g2_a21oi_1 _12594_ (.A1(_03807_),
    .A2(_03818_),
    .Y(_03921_),
    .B1(_03817_));
 sg13g2_a22oi_1 _12595_ (.Y(_03922_),
    .B1(net4715),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][14] ),
    .A2(net4740),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][14] ));
 sg13g2_a22oi_1 _12596_ (.Y(_03923_),
    .B1(net4709),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][14] ),
    .A2(net4725),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][14] ));
 sg13g2_and2_1 _12597_ (.A(_03922_),
    .B(_03923_),
    .X(_03924_));
 sg13g2_a22oi_1 _12598_ (.Y(_03925_),
    .B1(net4712),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][14] ),
    .A2(net4808),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][14] ));
 sg13g2_a22oi_1 _12599_ (.Y(_03926_),
    .B1(net4737),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][14] ),
    .A2(net4849),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][14] ));
 sg13g2_a22oi_1 _12600_ (.Y(_03927_),
    .B1(net4733),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][14] ),
    .A2(net4734),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][14] ));
 sg13g2_and4_1 _12601_ (.A(net4772),
    .B(_03925_),
    .C(_03926_),
    .D(_03927_),
    .X(_03928_));
 sg13g2_a22oi_1 _12602_ (.Y(_03929_),
    .B1(_03924_),
    .B2(_03928_),
    .A2(net4835),
    .A1(_00402_));
 sg13g2_nor2b_1 _12603_ (.A(_03921_),
    .B_N(_03929_),
    .Y(_03930_));
 sg13g2_xnor2_1 _12604_ (.Y(_03931_),
    .A(_03921_),
    .B(_03929_));
 sg13g2_xnor2_1 _12605_ (.Y(_03932_),
    .A(_03920_),
    .B(_03931_));
 sg13g2_o21ai_1 _12606_ (.B1(_03840_),
    .Y(_03933_),
    .A1(_03819_),
    .A2(_03841_));
 sg13g2_o21ai_1 _12607_ (.B1(_03829_),
    .Y(_03934_),
    .A1(_03830_),
    .A2(_03838_));
 sg13g2_and2_1 _12608_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][14] ),
    .B(net4755),
    .X(_03935_));
 sg13g2_a221oi_1 _12609_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][14] ),
    .C1(_03935_),
    .B1(net4758),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][14] ),
    .Y(_03936_),
    .A2(net4761));
 sg13g2_a221oi_1 _12610_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][14] ),
    .C1(net4828),
    .B1(net4818),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][14] ),
    .Y(_03937_),
    .A2(net4764));
 sg13g2_a22oi_1 _12611_ (.Y(_03938_),
    .B1(net4803),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][14] ),
    .A2(net4752),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][14] ));
 sg13g2_a22oi_1 _12612_ (.Y(_03939_),
    .B1(net4749),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][14] ),
    .A2(net4874),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][14] ));
 sg13g2_and3_1 _12613_ (.X(_03940_),
    .A(_03937_),
    .B(_03938_),
    .C(_03939_));
 sg13g2_a22oi_1 _12614_ (.Y(_03941_),
    .B1(_03936_),
    .B2(_03940_),
    .A2(net4828),
    .A1(_00400_));
 sg13g2_nand2_1 _12615_ (.Y(_03942_),
    .A(_03934_),
    .B(_03941_));
 sg13g2_xnor2_1 _12616_ (.Y(_03943_),
    .A(_03934_),
    .B(_03941_));
 sg13g2_a22oi_1 _12617_ (.Y(_03944_),
    .B1(net4743),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][14] ),
    .A2(net4746),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][14] ));
 sg13g2_a22oi_1 _12618_ (.Y(_03945_),
    .B1(net4847),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][14] ),
    .A2(net4803),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][14] ));
 sg13g2_nand2_1 _12619_ (.Y(_03946_),
    .A(_03944_),
    .B(_03945_));
 sg13g2_a22oi_1 _12620_ (.Y(_03947_),
    .B1(net4794),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][14] ),
    .A2(net4797),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][14] ));
 sg13g2_a22oi_1 _12621_ (.Y(_03948_),
    .B1(net4791),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][14] ),
    .A2(net4815),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][14] ));
 sg13g2_nand3_1 _12622_ (.B(_03947_),
    .C(_03948_),
    .A(net4768),
    .Y(_03949_));
 sg13g2_nand2_1 _12623_ (.Y(_03950_),
    .A(_00401_),
    .B(net4823));
 sg13g2_o21ai_1 _12624_ (.B1(_03950_),
    .Y(_03951_),
    .A1(_03946_),
    .A2(_03949_));
 sg13g2_xor2_1 _12625_ (.B(_03951_),
    .A(_03943_),
    .X(_03952_));
 sg13g2_nand2_1 _12626_ (.Y(_03953_),
    .A(_03933_),
    .B(_03952_));
 sg13g2_xnor2_1 _12627_ (.Y(_03954_),
    .A(_03933_),
    .B(_03952_));
 sg13g2_xor2_1 _12628_ (.B(_03954_),
    .A(_03932_),
    .X(_03955_));
 sg13g2_xnor2_1 _12629_ (.Y(_03956_),
    .A(_03912_),
    .B(_03955_));
 sg13g2_nor2_1 _12630_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .B(net4930),
    .Y(_03957_));
 sg13g2_a21oi_1 _12631_ (.A1(net4926),
    .A2(_03956_),
    .Y(_00260_),
    .B1(_03957_));
 sg13g2_and2_1 _12632_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][15] ),
    .B(net4730),
    .X(_03958_));
 sg13g2_a22oi_1 _12633_ (.Y(_03959_),
    .B1(net4659),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][15] ),
    .A2(net4722),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][15] ));
 sg13g2_a221oi_1 _12634_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][15] ),
    .C1(_03958_),
    .B1(net4650),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][15] ),
    .Y(_03960_),
    .A2(net4657));
 sg13g2_a21oi_1 _12635_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][15] ),
    .A2(net4663),
    .Y(_03961_),
    .B1(net4840));
 sg13g2_a22oi_1 _12636_ (.Y(_03962_),
    .B1(net4653),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][15] ),
    .A2(net4811),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][15] ));
 sg13g2_nand3_1 _12637_ (.B(_03961_),
    .C(_03962_),
    .A(_03959_),
    .Y(_03963_));
 sg13g2_a221oi_1 _12638_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][15] ),
    .C1(_03963_),
    .B1(net4655),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][15] ),
    .Y(_03964_),
    .A2(net4665));
 sg13g2_a22oi_1 _12639_ (.Y(_03965_),
    .B1(_03960_),
    .B2(_03964_),
    .A2(net4840),
    .A1(_00410_));
 sg13g2_a22oi_1 _12640_ (.Y(_03966_),
    .B1(net4717),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][15] ),
    .A2(net4727),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][15] ));
 sg13g2_a22oi_1 _12641_ (.Y(_03967_),
    .B1(net4719),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][15] ),
    .A2(net4851),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][15] ));
 sg13g2_a22oi_1 _12642_ (.Y(_03968_),
    .B1(net4741),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][15] ),
    .A2(net4807),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][15] ));
 sg13g2_and2_1 _12643_ (.A(_03967_),
    .B(_03968_),
    .X(_03969_));
 sg13g2_a22oi_1 _12644_ (.Y(_03970_),
    .B1(net4713),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][15] ),
    .A2(net4738),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][15] ));
 sg13g2_a22oi_1 _12645_ (.Y(_03971_),
    .B1(net4710),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][15] ),
    .A2(net4735),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][15] ));
 sg13g2_and4_1 _12646_ (.A(net4769),
    .B(_03966_),
    .C(_03970_),
    .D(_03971_),
    .X(_03972_));
 sg13g2_a22oi_1 _12647_ (.Y(_03973_),
    .B1(_03969_),
    .B2(_03972_),
    .A2(net4827),
    .A1(_00409_));
 sg13g2_a21oi_2 _12648_ (.B1(_03930_),
    .Y(_03974_),
    .A2(_03931_),
    .A1(_03920_));
 sg13g2_nor2b_1 _12649_ (.A(_03974_),
    .B_N(_03973_),
    .Y(_03975_));
 sg13g2_xnor2_1 _12650_ (.Y(_03976_),
    .A(_03973_),
    .B(_03974_));
 sg13g2_xnor2_1 _12651_ (.Y(_03977_),
    .A(_03965_),
    .B(_03976_));
 sg13g2_o21ai_1 _12652_ (.B1(_03953_),
    .Y(_03978_),
    .A1(_03932_),
    .A2(_03954_));
 sg13g2_o21ai_1 _12653_ (.B1(_03942_),
    .Y(_03979_),
    .A1(_03943_),
    .A2(_03951_));
 sg13g2_and2_1 _12654_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][15] ),
    .B(net4760),
    .X(_03980_));
 sg13g2_a221oi_1 _12655_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][15] ),
    .C1(_03980_),
    .B1(net4751),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][15] ),
    .Y(_03981_),
    .A2(net4754));
 sg13g2_a221oi_1 _12656_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][15] ),
    .C1(net4825),
    .B1(net4813),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][15] ),
    .Y(_03982_),
    .A2(net4876));
 sg13g2_a22oi_1 _12657_ (.Y(_03983_),
    .B1(net4757),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][15] ),
    .A2(net4763),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][15] ));
 sg13g2_a22oi_1 _12658_ (.Y(_03984_),
    .B1(net4800),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][15] ),
    .A2(net4766),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][15] ));
 sg13g2_and3_1 _12659_ (.X(_03985_),
    .A(_03982_),
    .B(_03983_),
    .C(_03984_));
 sg13g2_a22oi_1 _12660_ (.Y(_03986_),
    .B1(_03981_),
    .B2(_03985_),
    .A2(net4825),
    .A1(_00407_));
 sg13g2_nand2_1 _12661_ (.Y(_03987_),
    .A(_03979_),
    .B(_03986_));
 sg13g2_xnor2_1 _12662_ (.Y(_03988_),
    .A(_03979_),
    .B(_03986_));
 sg13g2_nand2_1 _12663_ (.Y(_03989_),
    .A(_00408_),
    .B(net4823));
 sg13g2_a22oi_1 _12664_ (.Y(_03990_),
    .B1(net4793),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][15] ),
    .A2(net4799),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][15] ));
 sg13g2_a22oi_1 _12665_ (.Y(_03991_),
    .B1(net4847),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][15] ),
    .A2(net4814),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][15] ));
 sg13g2_nand3_1 _12666_ (.B(_03990_),
    .C(_03991_),
    .A(net4767),
    .Y(_03992_));
 sg13g2_a22oi_1 _12667_ (.Y(_03993_),
    .B1(net4796),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][15] ),
    .A2(net4748),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][15] ));
 sg13g2_a22oi_1 _12668_ (.Y(_03994_),
    .B1(net4745),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][15] ),
    .A2(net4801),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][15] ));
 sg13g2_nand2_1 _12669_ (.Y(_03995_),
    .A(_03993_),
    .B(_03994_));
 sg13g2_o21ai_1 _12670_ (.B1(_03989_),
    .Y(_03996_),
    .A1(_03992_),
    .A2(_03995_));
 sg13g2_xor2_1 _12671_ (.B(_03996_),
    .A(_03988_),
    .X(_03997_));
 sg13g2_nand2_1 _12672_ (.Y(_03998_),
    .A(_03978_),
    .B(_03997_));
 sg13g2_xnor2_1 _12673_ (.Y(_03999_),
    .A(_03978_),
    .B(_03997_));
 sg13g2_xnor2_1 _12674_ (.Y(_04000_),
    .A(_03977_),
    .B(_03999_));
 sg13g2_a21oi_1 _12675_ (.A1(_03888_),
    .A2(_03893_),
    .Y(_04001_),
    .B1(_03887_));
 sg13g2_o21ai_1 _12676_ (.B1(net4774),
    .Y(_04002_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][15] ),
    .A2(net4821));
 sg13g2_a22oi_1 _12677_ (.Y(_04003_),
    .B1(net4694),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][15] ),
    .A2(net4696),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][15] ));
 sg13g2_a22oi_1 _12678_ (.Y(_04004_),
    .B1(net4687),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][15] ),
    .A2(net4689),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][15] ));
 sg13g2_a22oi_1 _12679_ (.Y(_04005_),
    .B1(net4692),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][15] ),
    .A2(net4872),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][15] ));
 sg13g2_nand4_1 _12680_ (.B(_04003_),
    .C(_04004_),
    .A(_04002_),
    .Y(_04006_),
    .D(_04005_));
 sg13g2_nand2_1 _12681_ (.Y(_04007_),
    .A(_00405_),
    .B(net4697));
 sg13g2_nand2_2 _12682_ (.Y(_04008_),
    .A(_04006_),
    .B(_04007_));
 sg13g2_nor2_1 _12683_ (.A(_04001_),
    .B(_04008_),
    .Y(_04009_));
 sg13g2_xor2_1 _12684_ (.B(_04008_),
    .A(_04001_),
    .X(_04010_));
 sg13g2_a221oi_1 _12685_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][15] ),
    .C1(net4678),
    .B1(net4669),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][15] ),
    .Y(_04011_),
    .A2(net4676));
 sg13g2_a22oi_1 _12686_ (.Y(_04012_),
    .B1(net4671),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][15] ),
    .A2(net4684),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][15] ));
 sg13g2_a22oi_1 _12687_ (.Y(_04013_),
    .B1(net4667),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][15] ),
    .A2(net4674),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][15] ));
 sg13g2_and2_1 _12688_ (.A(_04012_),
    .B(_04013_),
    .X(_04014_));
 sg13g2_a22oi_1 _12689_ (.Y(_04015_),
    .B1(_04011_),
    .B2(_04014_),
    .A2(net4678),
    .A1(_00406_));
 sg13g2_xnor2_1 _12690_ (.Y(_04016_),
    .A(_04010_),
    .B(_04015_));
 sg13g2_o21ai_1 _12691_ (.B1(_03906_),
    .Y(_04017_),
    .A1(_03894_),
    .A2(_03907_));
 sg13g2_o21ai_1 _12692_ (.B1(_03898_),
    .Y(_04018_),
    .A1(_03899_),
    .A2(_03904_));
 sg13g2_mux2_1 _12693_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][15] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][15] ),
    .S(net4844),
    .X(_04019_));
 sg13g2_nand2_1 _12694_ (.Y(_04020_),
    .A(_04018_),
    .B(_04019_));
 sg13g2_xnor2_1 _12695_ (.Y(_04021_),
    .A(_04018_),
    .B(_04019_));
 sg13g2_nand2_1 _12696_ (.Y(_04022_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][15] ),
    .B(net4703));
 sg13g2_a22oi_1 _12697_ (.Y(_04023_),
    .B1(net4781),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][15] ),
    .A2(net4785),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][15] ));
 sg13g2_a22oi_1 _12698_ (.Y(_04024_),
    .B1(net4777),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][15] ),
    .A2(net4787),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][15] ));
 sg13g2_nand4_1 _12699_ (.B(_04022_),
    .C(_04023_),
    .A(net4706),
    .Y(_04025_),
    .D(_04024_));
 sg13g2_o21ai_1 _12700_ (.B1(_04025_),
    .Y(_04026_),
    .A1(_02351_),
    .A2(net4707));
 sg13g2_xnor2_1 _12701_ (.Y(_04027_),
    .A(_04021_),
    .B(_04026_));
 sg13g2_nand2b_1 _12702_ (.Y(_04028_),
    .B(_04017_),
    .A_N(_04027_));
 sg13g2_nor2b_1 _12703_ (.A(_04017_),
    .B_N(_04027_),
    .Y(_04029_));
 sg13g2_xnor2_1 _12704_ (.Y(_04030_),
    .A(_04017_),
    .B(_04027_));
 sg13g2_xnor2_1 _12705_ (.Y(_04031_),
    .A(_04016_),
    .B(_04030_));
 sg13g2_a21o_1 _12706_ (.A2(_03955_),
    .A1(_03912_),
    .B1(_03911_),
    .X(_04032_));
 sg13g2_nand2_1 _12707_ (.Y(_04033_),
    .A(_04031_),
    .B(_04032_));
 sg13g2_nor2_1 _12708_ (.A(_04031_),
    .B(_04032_),
    .Y(_04034_));
 sg13g2_xor2_1 _12709_ (.B(_04032_),
    .A(_04031_),
    .X(_04035_));
 sg13g2_xnor2_1 _12710_ (.Y(_04036_),
    .A(_04000_),
    .B(_04035_));
 sg13g2_mux2_1 _12711_ (.A0(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .A1(_04036_),
    .S(net4926),
    .X(_00261_));
 sg13g2_o21ai_1 _12712_ (.B1(_04033_),
    .Y(_04037_),
    .A1(_04000_),
    .A2(_04034_));
 sg13g2_a21oi_1 _12713_ (.A1(_04010_),
    .A2(_04015_),
    .Y(_04038_),
    .B1(_04009_));
 sg13g2_o21ai_1 _12714_ (.B1(net4775),
    .Y(_04039_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][16] ),
    .A2(net4820));
 sg13g2_a22oi_1 _12715_ (.Y(_04040_),
    .B1(net4694),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][16] ),
    .A2(net4696),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][16] ));
 sg13g2_a22oi_1 _12716_ (.Y(_04041_),
    .B1(net4688),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][16] ),
    .A2(net4692),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][16] ));
 sg13g2_a22oi_1 _12717_ (.Y(_04042_),
    .B1(net4690),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][16] ),
    .A2(net4873),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][16] ));
 sg13g2_nand4_1 _12718_ (.B(_04040_),
    .C(_04041_),
    .A(_04039_),
    .Y(_04043_),
    .D(_04042_));
 sg13g2_nand2_1 _12719_ (.Y(_04044_),
    .A(_00414_),
    .B(net4698));
 sg13g2_nand2_1 _12720_ (.Y(_04045_),
    .A(_04043_),
    .B(_04044_));
 sg13g2_nor2_1 _12721_ (.A(_04038_),
    .B(_04045_),
    .Y(_04046_));
 sg13g2_xnor2_1 _12722_ (.Y(_04047_),
    .A(_04038_),
    .B(_04045_));
 sg13g2_a221oi_1 _12723_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][16] ),
    .C1(net4682),
    .B1(_02834_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][16] ),
    .Y(_04048_),
    .A2(_02828_));
 sg13g2_a22oi_1 _12724_ (.Y(_04049_),
    .B1(net4672),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][16] ),
    .A2(_02831_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][16] ));
 sg13g2_a22oi_1 _12725_ (.Y(_04050_),
    .B1(_02836_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][16] ),
    .A2(net4685),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][16] ));
 sg13g2_nand3_1 _12726_ (.B(_04049_),
    .C(_04050_),
    .A(_04048_),
    .Y(_04051_));
 sg13g2_o21ai_1 _12727_ (.B1(_04051_),
    .Y(_04052_),
    .A1(_02352_),
    .A2(_02827_));
 sg13g2_nor2_1 _12728_ (.A(_04047_),
    .B(_04052_),
    .Y(_04053_));
 sg13g2_xnor2_1 _12729_ (.Y(_04054_),
    .A(_04047_),
    .B(_04052_));
 sg13g2_o21ai_1 _12730_ (.B1(_04028_),
    .Y(_04055_),
    .A1(_04016_),
    .A2(_04029_));
 sg13g2_o21ai_1 _12731_ (.B1(_04020_),
    .Y(_04056_),
    .A1(_04021_),
    .A2(_04026_));
 sg13g2_mux2_1 _12732_ (.A0(_00412_),
    .A1(_00411_),
    .S(net4844),
    .X(_04057_));
 sg13g2_nor2b_1 _12733_ (.A(_04057_),
    .B_N(_04056_),
    .Y(_04058_));
 sg13g2_nand2b_1 _12734_ (.Y(_04059_),
    .B(_04057_),
    .A_N(_04056_));
 sg13g2_xor2_1 _12735_ (.B(_04057_),
    .A(_04056_),
    .X(_04060_));
 sg13g2_and2_1 _12736_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][16] ),
    .B(net4784),
    .X(_04061_));
 sg13g2_a221oi_1 _12737_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][16] ),
    .C1(_04061_),
    .B1(net4701),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][16] ),
    .Y(_04062_),
    .A2(net4780));
 sg13g2_a221oi_1 _12738_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][16] ),
    .C1(net4647),
    .B1(net4776),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][16] ),
    .Y(_04063_),
    .A2(net4787));
 sg13g2_a22oi_1 _12739_ (.Y(_04064_),
    .B1(_04062_),
    .B2(_04063_),
    .A2(net4647),
    .A1(_00413_));
 sg13g2_xnor2_1 _12740_ (.Y(_04065_),
    .A(_04060_),
    .B(_04064_));
 sg13g2_nand2_1 _12741_ (.Y(_04066_),
    .A(_04055_),
    .B(_04065_));
 sg13g2_nor2_1 _12742_ (.A(_04055_),
    .B(_04065_),
    .Y(_04067_));
 sg13g2_xor2_1 _12743_ (.B(_04065_),
    .A(_04055_),
    .X(_04068_));
 sg13g2_xnor2_1 _12744_ (.Y(_04069_),
    .A(_04054_),
    .B(_04068_));
 sg13g2_and2_1 _12745_ (.A(_04037_),
    .B(_04069_),
    .X(_04070_));
 sg13g2_xor2_1 _12746_ (.B(_04069_),
    .A(_04037_),
    .X(_04071_));
 sg13g2_a22oi_1 _12747_ (.Y(_04072_),
    .B1(net4655),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][16] ),
    .A2(net4665),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][16] ));
 sg13g2_and2_1 _12748_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][16] ),
    .B(net4730),
    .X(_04073_));
 sg13g2_a221oi_1 _12749_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][16] ),
    .C1(_04073_),
    .B1(net4650),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][16] ),
    .Y(_04074_),
    .A2(net4812));
 sg13g2_a21oi_1 _12750_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][16] ),
    .A2(net4722),
    .Y(_04075_),
    .B1(net4837));
 sg13g2_a22oi_1 _12751_ (.Y(_04076_),
    .B1(net4657),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][16] ),
    .A2(net4659),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][16] ));
 sg13g2_nand3_1 _12752_ (.B(_04075_),
    .C(_04076_),
    .A(_04072_),
    .Y(_04077_));
 sg13g2_a221oi_1 _12753_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][16] ),
    .C1(_04077_),
    .B1(net4653),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][16] ),
    .Y(_04078_),
    .A2(net4663));
 sg13g2_a22oi_1 _12754_ (.Y(_04079_),
    .B1(_04074_),
    .B2(_04078_),
    .A2(net4837),
    .A1(_00419_));
 sg13g2_a21oi_1 _12755_ (.A1(_03965_),
    .A2(_03976_),
    .Y(_04080_),
    .B1(_03975_));
 sg13g2_a22oi_1 _12756_ (.Y(_04081_),
    .B1(net4718),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][16] ),
    .A2(net4742),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][16] ));
 sg13g2_a22oi_1 _12757_ (.Y(_04082_),
    .B1(net4727),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][16] ),
    .A2(net4807),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][16] ));
 sg13g2_and2_1 _12758_ (.A(_04081_),
    .B(_04082_),
    .X(_04083_));
 sg13g2_a22oi_1 _12759_ (.Y(_04084_),
    .B1(net4711),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][16] ),
    .A2(net4714),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][16] ));
 sg13g2_a22oi_1 _12760_ (.Y(_04085_),
    .B1(net4739),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][16] ),
    .A2(net4851),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][16] ));
 sg13g2_a22oi_1 _12761_ (.Y(_04086_),
    .B1(net4719),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][16] ),
    .A2(net4736),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][16] ));
 sg13g2_and4_1 _12762_ (.A(net4768),
    .B(_04084_),
    .C(_04085_),
    .D(_04086_),
    .X(_04087_));
 sg13g2_a22oi_1 _12763_ (.Y(_04088_),
    .B1(_04083_),
    .B2(_04087_),
    .A2(net4827),
    .A1(_00418_));
 sg13g2_nor2b_1 _12764_ (.A(_04080_),
    .B_N(_04088_),
    .Y(_04089_));
 sg13g2_xnor2_1 _12765_ (.Y(_04090_),
    .A(_04080_),
    .B(_04088_));
 sg13g2_xnor2_1 _12766_ (.Y(_04091_),
    .A(_04079_),
    .B(_04090_));
 sg13g2_o21ai_1 _12767_ (.B1(_03998_),
    .Y(_04092_),
    .A1(_03977_),
    .A2(_03999_));
 sg13g2_nand2_1 _12768_ (.Y(_04093_),
    .A(_00417_),
    .B(net4826));
 sg13g2_a22oi_1 _12769_ (.Y(_04094_),
    .B1(net4745),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][16] ),
    .A2(net4800),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][16] ));
 sg13g2_a22oi_1 _12770_ (.Y(_04095_),
    .B1(net4848),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][16] ),
    .A2(net4799),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][16] ));
 sg13g2_nand2_1 _12771_ (.Y(_04096_),
    .A(_04094_),
    .B(_04095_));
 sg13g2_a22oi_1 _12772_ (.Y(_04097_),
    .B1(net4796),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][16] ),
    .A2(net4748),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][16] ));
 sg13g2_a22oi_1 _12773_ (.Y(_04098_),
    .B1(net4793),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][16] ),
    .A2(net4813),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][16] ));
 sg13g2_nand3_1 _12774_ (.B(_04097_),
    .C(_04098_),
    .A(net4767),
    .Y(_04099_));
 sg13g2_o21ai_1 _12775_ (.B1(_04093_),
    .Y(_04100_),
    .A1(_04096_),
    .A2(_04099_));
 sg13g2_o21ai_1 _12776_ (.B1(_03987_),
    .Y(_04101_),
    .A1(_03988_),
    .A2(_03996_));
 sg13g2_and2_1 _12777_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][16] ),
    .B(net4876),
    .X(_04102_));
 sg13g2_a221oi_1 _12778_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][16] ),
    .C1(_04102_),
    .B1(net4760),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][16] ),
    .Y(_04103_),
    .A2(net4763));
 sg13g2_a221oi_1 _12779_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][16] ),
    .C1(net4822),
    .B1(net4800),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][16] ),
    .Y(_04104_),
    .A2(net4813));
 sg13g2_a22oi_1 _12780_ (.Y(_04105_),
    .B1(net4757),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][16] ),
    .A2(net4766),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][16] ));
 sg13g2_a22oi_1 _12781_ (.Y(_04106_),
    .B1(net4751),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][16] ),
    .A2(net4754),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][16] ));
 sg13g2_and3_1 _12782_ (.X(_04107_),
    .A(_04104_),
    .B(_04105_),
    .C(_04106_));
 sg13g2_a22oi_1 _12783_ (.Y(_04108_),
    .B1(_04103_),
    .B2(_04107_),
    .A2(net4822),
    .A1(_00416_));
 sg13g2_nand2_1 _12784_ (.Y(_04109_),
    .A(_04101_),
    .B(_04108_));
 sg13g2_xnor2_1 _12785_ (.Y(_04110_),
    .A(_04101_),
    .B(_04108_));
 sg13g2_xor2_1 _12786_ (.B(_04110_),
    .A(_04100_),
    .X(_04111_));
 sg13g2_nand2_1 _12787_ (.Y(_04112_),
    .A(_04092_),
    .B(_04111_));
 sg13g2_xnor2_1 _12788_ (.Y(_04113_),
    .A(_04092_),
    .B(_04111_));
 sg13g2_xor2_1 _12789_ (.B(_04113_),
    .A(_04091_),
    .X(_04114_));
 sg13g2_xnor2_1 _12790_ (.Y(_04115_),
    .A(_04071_),
    .B(_04114_));
 sg13g2_nor2_1 _12791_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .B(net4926),
    .Y(_04116_));
 sg13g2_a21oi_1 _12792_ (.A1(net4926),
    .A2(_04115_),
    .Y(_00262_),
    .B1(_04116_));
 sg13g2_a22oi_1 _12793_ (.Y(_04117_),
    .B1(net4657),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][17] ),
    .A2(net4721),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][17] ));
 sg13g2_a22oi_1 _12794_ (.Y(_04118_),
    .B1(net4659),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][17] ),
    .A2(net4663),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][17] ));
 sg13g2_and2_1 _12795_ (.A(_04117_),
    .B(_04118_),
    .X(_04119_));
 sg13g2_a221oi_1 _12796_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][17] ),
    .C1(net4837),
    .B1(net4729),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][17] ),
    .Y(_04120_),
    .A2(net4812));
 sg13g2_a22oi_1 _12797_ (.Y(_04121_),
    .B1(net4655),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][17] ),
    .A2(net4665),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][17] ));
 sg13g2_nand2_1 _12798_ (.Y(_04122_),
    .A(_04120_),
    .B(_04121_));
 sg13g2_a221oi_1 _12799_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][17] ),
    .C1(_04122_),
    .B1(net4650),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][17] ),
    .Y(_04123_),
    .A2(net4653));
 sg13g2_a22oi_1 _12800_ (.Y(_04124_),
    .B1(_04119_),
    .B2(_04123_),
    .A2(net4837),
    .A1(_00426_));
 sg13g2_a21oi_2 _12801_ (.B1(_04089_),
    .Y(_04125_),
    .A2(_04090_),
    .A1(_04079_));
 sg13g2_a22oi_1 _12802_ (.Y(_04126_),
    .B1(net4718),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][17] ),
    .A2(net4727),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][17] ));
 sg13g2_a22oi_1 _12803_ (.Y(_04127_),
    .B1(net4736),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][17] ),
    .A2(net4852),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][17] ));
 sg13g2_a22oi_1 _12804_ (.Y(_04128_),
    .B1(net4742),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][17] ),
    .A2(net4802),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][17] ));
 sg13g2_and2_1 _12805_ (.A(_04127_),
    .B(_04128_),
    .X(_04129_));
 sg13g2_a22oi_1 _12806_ (.Y(_04130_),
    .B1(net4714),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][17] ),
    .A2(net4739),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][17] ));
 sg13g2_a22oi_1 _12807_ (.Y(_04131_),
    .B1(net4711),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][17] ),
    .A2(net4719),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][17] ));
 sg13g2_and4_1 _12808_ (.A(net4767),
    .B(_04126_),
    .C(_04130_),
    .D(_04131_),
    .X(_04132_));
 sg13g2_a22oi_1 _12809_ (.Y(_04133_),
    .B1(_04129_),
    .B2(_04132_),
    .A2(net4826),
    .A1(_00425_));
 sg13g2_nand2b_1 _12810_ (.Y(_04134_),
    .B(_04133_),
    .A_N(_04125_));
 sg13g2_xnor2_1 _12811_ (.Y(_04135_),
    .A(_04125_),
    .B(_04133_));
 sg13g2_nand2_1 _12812_ (.Y(_04136_),
    .A(_04124_),
    .B(_04135_));
 sg13g2_xnor2_1 _12813_ (.Y(_04137_),
    .A(_04124_),
    .B(_04135_));
 sg13g2_o21ai_1 _12814_ (.B1(_04112_),
    .Y(_04138_),
    .A1(_04091_),
    .A2(_04113_));
 sg13g2_o21ai_1 _12815_ (.B1(_04109_),
    .Y(_04139_),
    .A1(_04100_),
    .A2(_04110_));
 sg13g2_nand2_1 _12816_ (.Y(_04140_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][17] ),
    .B(net4757));
 sg13g2_nand2_1 _12817_ (.Y(_04141_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][17] ),
    .B(net4751));
 sg13g2_a22oi_1 _12818_ (.Y(_04142_),
    .B1(net4877),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][17] ),
    .A2(net4760),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][17] ));
 sg13g2_a21oi_1 _12819_ (.A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][17] ),
    .A2(net4766),
    .Y(_04143_),
    .B1(net4825));
 sg13g2_a22oi_1 _12820_ (.Y(_04144_),
    .B1(net4800),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][17] ),
    .A2(net4813),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][17] ));
 sg13g2_nand4_1 _12821_ (.B(_04142_),
    .C(_04143_),
    .A(_04141_),
    .Y(_04145_),
    .D(_04144_));
 sg13g2_a221oi_1 _12822_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][17] ),
    .C1(_04145_),
    .B1(net4754),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][17] ),
    .Y(_04146_),
    .A2(net4763));
 sg13g2_a22oi_1 _12823_ (.Y(_04147_),
    .B1(_04140_),
    .B2(_04146_),
    .A2(net4822),
    .A1(_00423_));
 sg13g2_nand2_1 _12824_ (.Y(_04148_),
    .A(_04139_),
    .B(_04147_));
 sg13g2_xnor2_1 _12825_ (.Y(_04149_),
    .A(_04139_),
    .B(_04147_));
 sg13g2_nand2_1 _12826_ (.Y(_04150_),
    .A(_00424_),
    .B(net4826));
 sg13g2_a22oi_1 _12827_ (.Y(_04151_),
    .B1(net4796),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][17] ),
    .A2(net4745),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][17] ));
 sg13g2_a22oi_1 _12828_ (.Y(_04152_),
    .B1(net4848),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][17] ),
    .A2(net4799),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][17] ));
 sg13g2_a22oi_1 _12829_ (.Y(_04153_),
    .B1(net4793),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][17] ),
    .A2(net4814),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][17] ));
 sg13g2_nand3_1 _12830_ (.B(_04152_),
    .C(_04153_),
    .A(net4767),
    .Y(_04154_));
 sg13g2_a22oi_1 _12831_ (.Y(_04155_),
    .B1(net4748),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][17] ),
    .A2(net4802),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][17] ));
 sg13g2_nand2_1 _12832_ (.Y(_04156_),
    .A(_04151_),
    .B(_04155_));
 sg13g2_o21ai_1 _12833_ (.B1(_04150_),
    .Y(_04157_),
    .A1(_04154_),
    .A2(_04156_));
 sg13g2_xor2_1 _12834_ (.B(_04157_),
    .A(_04149_),
    .X(_04158_));
 sg13g2_nand2_1 _12835_ (.Y(_04159_),
    .A(_04138_),
    .B(_04158_));
 sg13g2_xnor2_1 _12836_ (.Y(_04160_),
    .A(_04138_),
    .B(_04158_));
 sg13g2_or2_1 _12837_ (.X(_04161_),
    .B(_04160_),
    .A(_04137_));
 sg13g2_xor2_1 _12838_ (.B(_04160_),
    .A(_04137_),
    .X(_04162_));
 sg13g2_a21o_1 _12839_ (.A2(_04114_),
    .A1(_04071_),
    .B1(_04070_),
    .X(_04163_));
 sg13g2_nor2_1 _12840_ (.A(_04046_),
    .B(_04053_),
    .Y(_04164_));
 sg13g2_o21ai_1 _12841_ (.B1(_02792_),
    .Y(_04165_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][17] ),
    .A2(net4821));
 sg13g2_a22oi_1 _12842_ (.Y(_04166_),
    .B1(net4694),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][17] ),
    .A2(net4696),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][17] ));
 sg13g2_a22oi_1 _12843_ (.Y(_04167_),
    .B1(net4688),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][17] ),
    .A2(net4690),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][17] ));
 sg13g2_a22oi_1 _12844_ (.Y(_04168_),
    .B1(_02802_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][17] ),
    .A2(net4877),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][17] ));
 sg13g2_nand4_1 _12845_ (.B(_04166_),
    .C(_04167_),
    .A(_04165_),
    .Y(_04169_),
    .D(_04168_));
 sg13g2_nand2_1 _12846_ (.Y(_04170_),
    .A(_00421_),
    .B(net4698));
 sg13g2_nand2_1 _12847_ (.Y(_04171_),
    .A(_04169_),
    .B(_04170_));
 sg13g2_nor2_1 _12848_ (.A(_04164_),
    .B(_04171_),
    .Y(_04172_));
 sg13g2_xnor2_1 _12849_ (.Y(_04173_),
    .A(_04164_),
    .B(_04171_));
 sg13g2_a221oi_1 _12850_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][17] ),
    .C1(net4682),
    .B1(net4670),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][17] ),
    .Y(_04174_),
    .A2(net4677));
 sg13g2_a22oi_1 _12851_ (.Y(_04175_),
    .B1(_02836_),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][17] ),
    .A2(net4685),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][17] ));
 sg13g2_a22oi_1 _12852_ (.Y(_04176_),
    .B1(net4672),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][17] ),
    .A2(net4675),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][17] ));
 sg13g2_nand3_1 _12853_ (.B(_04175_),
    .C(_04176_),
    .A(_04174_),
    .Y(_04177_));
 sg13g2_o21ai_1 _12854_ (.B1(_04177_),
    .Y(_04178_),
    .A1(_02354_),
    .A2(_02827_));
 sg13g2_nor2_1 _12855_ (.A(_04173_),
    .B(_04178_),
    .Y(_04179_));
 sg13g2_xnor2_1 _12856_ (.Y(_04180_),
    .A(_04173_),
    .B(_04178_));
 sg13g2_o21ai_1 _12857_ (.B1(_04066_),
    .Y(_04181_),
    .A1(_04054_),
    .A2(_04067_));
 sg13g2_a21oi_1 _12858_ (.A1(_04059_),
    .A2(_04064_),
    .Y(_04182_),
    .B1(_04058_));
 sg13g2_mux2_1 _12859_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][17] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][17] ),
    .S(net4844),
    .X(_04183_));
 sg13g2_nand2b_1 _12860_ (.Y(_04184_),
    .B(_04183_),
    .A_N(_04182_));
 sg13g2_xor2_1 _12861_ (.B(_04183_),
    .A(_04182_),
    .X(_04185_));
 sg13g2_nand2_1 _12862_ (.Y(_04186_),
    .A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][17] ),
    .B(net4704));
 sg13g2_a22oi_1 _12863_ (.Y(_04187_),
    .B1(net4783),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][17] ),
    .A2(net4786),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][17] ));
 sg13g2_a22oi_1 _12864_ (.Y(_04188_),
    .B1(net4779),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][17] ),
    .A2(net4790),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][17] ));
 sg13g2_nand4_1 _12865_ (.B(_04186_),
    .C(_04187_),
    .A(net4708),
    .Y(_04189_),
    .D(_04188_));
 sg13g2_o21ai_1 _12866_ (.B1(_04189_),
    .Y(_04190_),
    .A1(_02353_),
    .A2(net4708));
 sg13g2_xor2_1 _12867_ (.B(_04190_),
    .A(_04185_),
    .X(_04191_));
 sg13g2_nand2_1 _12868_ (.Y(_04192_),
    .A(_04181_),
    .B(_04191_));
 sg13g2_nor2_1 _12869_ (.A(_04181_),
    .B(_04191_),
    .Y(_04193_));
 sg13g2_xor2_1 _12870_ (.B(_04191_),
    .A(_04181_),
    .X(_04194_));
 sg13g2_xnor2_1 _12871_ (.Y(_04195_),
    .A(_04180_),
    .B(_04194_));
 sg13g2_and2_1 _12872_ (.A(_04163_),
    .B(_04195_),
    .X(_04196_));
 sg13g2_xor2_1 _12873_ (.B(_04195_),
    .A(_04163_),
    .X(_04197_));
 sg13g2_xnor2_1 _12874_ (.Y(_04198_),
    .A(_04162_),
    .B(_04197_));
 sg13g2_nor2_1 _12875_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .B(net4926),
    .Y(_04199_));
 sg13g2_a21oi_1 _12876_ (.A1(net4926),
    .A2(_04198_),
    .Y(_00263_),
    .B1(_04199_));
 sg13g2_o21ai_1 _12877_ (.B1(_04159_),
    .Y(_04200_),
    .A1(_04137_),
    .A2(_04160_));
 sg13g2_o21ai_1 _12878_ (.B1(_04148_),
    .Y(_04201_),
    .A1(_04149_),
    .A2(_04157_));
 sg13g2_a22oi_1 _12879_ (.Y(_04202_),
    .B1(net4745),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][18] ),
    .A2(net4748),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][18] ));
 sg13g2_a22oi_1 _12880_ (.Y(_04203_),
    .B1(net4848),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][18] ),
    .A2(net4802),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][18] ));
 sg13g2_nand2_1 _12881_ (.Y(_04204_),
    .A(_04202_),
    .B(_04203_));
 sg13g2_a22oi_1 _12882_ (.Y(_04205_),
    .B1(net4796),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][18] ),
    .A2(net4799),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][18] ));
 sg13g2_a22oi_1 _12883_ (.Y(_04206_),
    .B1(net4793),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][18] ),
    .A2(net4813),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][18] ));
 sg13g2_nand3_1 _12884_ (.B(_04205_),
    .C(_04206_),
    .A(net4767),
    .Y(_04207_));
 sg13g2_nand2_1 _12885_ (.Y(_04208_),
    .A(_00431_),
    .B(net4826));
 sg13g2_o21ai_1 _12886_ (.B1(_04208_),
    .Y(_04209_),
    .A1(_04204_),
    .A2(_04207_));
 sg13g2_and2_1 _12887_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][18] ),
    .B(net4800),
    .X(_04210_));
 sg13g2_a221oi_1 _12888_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][18] ),
    .C1(_04210_),
    .B1(net4760),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][18] ),
    .Y(_04211_),
    .A2(net4766));
 sg13g2_a221oi_1 _12889_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][18] ),
    .C1(net4822),
    .B1(net4754),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][18] ),
    .Y(_04212_),
    .A2(net4813));
 sg13g2_a22oi_1 _12890_ (.Y(_04213_),
    .B1(net4757),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][18] ),
    .A2(net4876),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][18] ));
 sg13g2_a22oi_1 _12891_ (.Y(_04214_),
    .B1(net4751),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][18] ),
    .A2(net4763),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][18] ));
 sg13g2_and3_1 _12892_ (.X(_04215_),
    .A(_04212_),
    .B(_04213_),
    .C(_04214_));
 sg13g2_a22oi_1 _12893_ (.Y(_04216_),
    .B1(_04211_),
    .B2(_04215_),
    .A2(net4822),
    .A1(_00430_));
 sg13g2_nand2b_1 _12894_ (.Y(_04217_),
    .B(_04216_),
    .A_N(_04209_));
 sg13g2_xnor2_1 _12895_ (.Y(_04218_),
    .A(_04209_),
    .B(_04216_));
 sg13g2_nand2b_1 _12896_ (.Y(_04219_),
    .B(_04218_),
    .A_N(_04201_));
 sg13g2_xnor2_1 _12897_ (.Y(_04220_),
    .A(_04201_),
    .B(_04218_));
 sg13g2_a21oi_1 _12898_ (.A1(_04159_),
    .A2(_04161_),
    .Y(_04221_),
    .B1(_04220_));
 sg13g2_xnor2_1 _12899_ (.Y(_04222_),
    .A(_04200_),
    .B(_04220_));
 sg13g2_a22oi_1 _12900_ (.Y(_04223_),
    .B1(net4659),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][18] ),
    .A2(net4665),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][18] ));
 sg13g2_a22oi_1 _12901_ (.Y(_04224_),
    .B1(net4655),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][18] ),
    .A2(net4720),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][18] ));
 sg13g2_and2_1 _12902_ (.A(_04223_),
    .B(_04224_),
    .X(_04225_));
 sg13g2_a221oi_1 _12903_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][18] ),
    .C1(net4834),
    .B1(net4728),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][18] ),
    .Y(_04226_),
    .A2(net4808));
 sg13g2_a22oi_1 _12904_ (.Y(_04227_),
    .B1(net4657),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][18] ),
    .A2(net4663),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][18] ));
 sg13g2_nand2_1 _12905_ (.Y(_04228_),
    .A(_04226_),
    .B(_04227_));
 sg13g2_a221oi_1 _12906_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][18] ),
    .C1(_04228_),
    .B1(net4650),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][18] ),
    .Y(_04229_),
    .A2(net4653));
 sg13g2_a22oi_1 _12907_ (.Y(_04230_),
    .B1(_04225_),
    .B2(_04229_),
    .A2(net4834),
    .A1(_00433_));
 sg13g2_a22oi_1 _12908_ (.Y(_04231_),
    .B1(net4718),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][18] ),
    .A2(net4736),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][18] ));
 sg13g2_a22oi_1 _12909_ (.Y(_04232_),
    .B1(net4727),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][18] ),
    .A2(net4739),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][18] ));
 sg13g2_a22oi_1 _12910_ (.Y(_04233_),
    .B1(net4719),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][18] ),
    .A2(net4742),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][18] ));
 sg13g2_and2_1 _12911_ (.A(_04231_),
    .B(_04233_),
    .X(_04234_));
 sg13g2_a22oi_1 _12912_ (.Y(_04235_),
    .B1(net4711),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][18] ),
    .A2(net4714),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][18] ));
 sg13g2_a22oi_1 _12913_ (.Y(_04236_),
    .B1(net4802),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][18] ),
    .A2(net4852),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][18] ));
 sg13g2_and4_1 _12914_ (.A(net4767),
    .B(_04232_),
    .C(_04235_),
    .D(_04236_),
    .X(_04237_));
 sg13g2_a22oi_1 _12915_ (.Y(_04238_),
    .B1(_04234_),
    .B2(_04237_),
    .A2(net4826),
    .A1(_00432_));
 sg13g2_nand2_1 _12916_ (.Y(_04239_),
    .A(_04230_),
    .B(_04238_));
 sg13g2_xor2_1 _12917_ (.B(_04238_),
    .A(_04230_),
    .X(_04240_));
 sg13g2_a21oi_1 _12918_ (.A1(_04134_),
    .A2(_04136_),
    .Y(_04241_),
    .B1(_04240_));
 sg13g2_nand3_1 _12919_ (.B(_04136_),
    .C(_04240_),
    .A(_04134_),
    .Y(_04242_));
 sg13g2_nand2b_1 _12920_ (.Y(_04243_),
    .B(_04242_),
    .A_N(_04241_));
 sg13g2_xor2_1 _12921_ (.B(_04243_),
    .A(_04222_),
    .X(_04244_));
 sg13g2_nor2_1 _12922_ (.A(_04172_),
    .B(_04179_),
    .Y(_04245_));
 sg13g2_o21ai_1 _12923_ (.B1(_02792_),
    .Y(_04246_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][18] ),
    .A2(net4820));
 sg13g2_a22oi_1 _12924_ (.Y(_04247_),
    .B1(net4694),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][18] ),
    .A2(net4696),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][18] ));
 sg13g2_a22oi_1 _12925_ (.Y(_04248_),
    .B1(net4688),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][18] ),
    .A2(_02802_),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][18] ));
 sg13g2_a22oi_1 _12926_ (.Y(_04249_),
    .B1(net4690),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][18] ),
    .A2(net4873),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][18] ));
 sg13g2_nand4_1 _12927_ (.B(_04247_),
    .C(_04248_),
    .A(_04246_),
    .Y(_04250_),
    .D(_04249_));
 sg13g2_nand2_1 _12928_ (.Y(_04251_),
    .A(_00428_),
    .B(net4699));
 sg13g2_nand2_1 _12929_ (.Y(_04252_),
    .A(_04250_),
    .B(_04251_));
 sg13g2_a22oi_1 _12930_ (.Y(_04253_),
    .B1(net4670),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][18] ),
    .A2(net4677),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][18] ));
 sg13g2_a22oi_1 _12931_ (.Y(_04254_),
    .B1(net4668),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][18] ),
    .A2(net4686),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][18] ));
 sg13g2_a22oi_1 _12932_ (.Y(_04255_),
    .B1(net4673),
    .B2(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][18] ),
    .A2(net4675),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][18] ));
 sg13g2_nand4_1 _12933_ (.B(_04253_),
    .C(_04254_),
    .A(_02827_),
    .Y(_04256_),
    .D(_04255_));
 sg13g2_o21ai_1 _12934_ (.B1(_04256_),
    .Y(_04257_),
    .A1(_02355_),
    .A2(_02827_));
 sg13g2_xor2_1 _12935_ (.B(_04257_),
    .A(_04252_),
    .X(_04258_));
 sg13g2_nand2_1 _12936_ (.Y(_04259_),
    .A(_04245_),
    .B(_04258_));
 sg13g2_xnor2_1 _12937_ (.Y(_04260_),
    .A(_04245_),
    .B(_04258_));
 sg13g2_o21ai_1 _12938_ (.B1(_04192_),
    .Y(_04261_),
    .A1(_04180_),
    .A2(_04193_));
 sg13g2_o21ai_1 _12939_ (.B1(_04184_),
    .Y(_04262_),
    .A1(_04185_),
    .A2(_04190_));
 sg13g2_and2_1 _12940_ (.A(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][18] ),
    .B(net4784),
    .X(_04263_));
 sg13g2_a221oi_1 _12941_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][18] ),
    .C1(_04263_),
    .B1(net4702),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][18] ),
    .Y(_04264_),
    .A2(net4780));
 sg13g2_a221oi_1 _12942_ (.B2(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][18] ),
    .C1(net4647),
    .B1(net4776),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][18] ),
    .Y(_04265_),
    .A2(net4787));
 sg13g2_a22oi_1 _12943_ (.Y(_04266_),
    .B1(_04264_),
    .B2(_04265_),
    .A2(net4647),
    .A1(_00427_));
 sg13g2_mux2_1 _12944_ (.A0(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][18] ),
    .A1(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][18] ),
    .S(net4844),
    .X(_04267_));
 sg13g2_nor2_1 _12945_ (.A(_04266_),
    .B(_04267_),
    .Y(_04268_));
 sg13g2_xor2_1 _12946_ (.B(_04267_),
    .A(_04266_),
    .X(_04269_));
 sg13g2_xnor2_1 _12947_ (.Y(_04270_),
    .A(_04262_),
    .B(_04269_));
 sg13g2_nor2b_1 _12948_ (.A(_04270_),
    .B_N(_04261_),
    .Y(_04271_));
 sg13g2_xor2_1 _12949_ (.B(_04270_),
    .A(_04261_),
    .X(_04272_));
 sg13g2_nor2b_1 _12950_ (.A(_04272_),
    .B_N(_04260_),
    .Y(_04273_));
 sg13g2_xor2_1 _12951_ (.B(_04272_),
    .A(_04260_),
    .X(_04274_));
 sg13g2_a21oi_1 _12952_ (.A1(_04162_),
    .A2(_04197_),
    .Y(_04275_),
    .B1(_04196_));
 sg13g2_nor2_1 _12953_ (.A(_04274_),
    .B(_04275_),
    .Y(_04276_));
 sg13g2_xor2_1 _12954_ (.B(_04275_),
    .A(_04274_),
    .X(_04277_));
 sg13g2_xnor2_1 _12955_ (.Y(_04278_),
    .A(_04244_),
    .B(_04277_));
 sg13g2_nor2_1 _12956_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B(net4926),
    .Y(_04279_));
 sg13g2_a21oi_1 _12957_ (.A1(net4926),
    .A2(_04278_),
    .Y(_00264_),
    .B1(_04279_));
 sg13g2_nor2_1 _12958_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B(net4925),
    .Y(_04280_));
 sg13g2_a21oi_2 _12959_ (.B1(_04276_),
    .Y(_04281_),
    .A2(_04277_),
    .A1(_04244_));
 sg13g2_nor2_1 _12960_ (.A(_04271_),
    .B(_04273_),
    .Y(_04282_));
 sg13g2_o21ai_1 _12961_ (.B1(_04259_),
    .Y(_04283_),
    .A1(_04252_),
    .A2(_04257_));
 sg13g2_a21oi_2 _12962_ (.B1(_04268_),
    .Y(_04284_),
    .A2(_04269_),
    .A1(_04262_));
 sg13g2_nand2_1 _12963_ (.Y(_04285_),
    .A(_04283_),
    .B(_04284_));
 sg13g2_xor2_1 _12964_ (.B(_04284_),
    .A(_04283_),
    .X(_04286_));
 sg13g2_nand2_1 _12965_ (.Y(_04287_),
    .A(_04282_),
    .B(_04286_));
 sg13g2_xnor2_1 _12966_ (.Y(_04288_),
    .A(_04282_),
    .B(_04286_));
 sg13g2_nor2b_1 _12967_ (.A(_04281_),
    .B_N(_04288_),
    .Y(_04289_));
 sg13g2_xnor2_1 _12968_ (.Y(_04290_),
    .A(_04281_),
    .B(_04288_));
 sg13g2_a21oi_1 _12969_ (.A1(_04222_),
    .A2(_04243_),
    .Y(_04291_),
    .B1(_04221_));
 sg13g2_nand4_1 _12970_ (.B(_04219_),
    .C(_04239_),
    .A(_04217_),
    .Y(_04292_),
    .D(_04242_));
 sg13g2_inv_1 _12971_ (.Y(_04293_),
    .A(_04292_));
 sg13g2_a22oi_1 _12972_ (.Y(_04294_),
    .B1(_04239_),
    .B2(_04242_),
    .A2(_04219_),
    .A1(_04217_));
 sg13g2_nor2_1 _12973_ (.A(_04293_),
    .B(_04294_),
    .Y(_04295_));
 sg13g2_xnor2_1 _12974_ (.Y(_04296_),
    .A(_04291_),
    .B(_04295_));
 sg13g2_xnor2_1 _12975_ (.Y(_04297_),
    .A(_04290_),
    .B(_04296_));
 sg13g2_a21oi_1 _12976_ (.A1(net4924),
    .A2(_04297_),
    .Y(_00265_),
    .B1(_04280_));
 sg13g2_nor2_1 _12977_ (.A(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B(net4924),
    .Y(_04298_));
 sg13g2_a21oi_1 _12978_ (.A1(_04290_),
    .A2(_04296_),
    .Y(_04299_),
    .B1(_04289_));
 sg13g2_o21ai_1 _12979_ (.B1(_04292_),
    .Y(_04300_),
    .A1(_04291_),
    .A2(_04294_));
 sg13g2_nand3_1 _12980_ (.B(_04287_),
    .C(_04300_),
    .A(_04285_),
    .Y(_04301_));
 sg13g2_a21oi_1 _12981_ (.A1(_04285_),
    .A2(_04287_),
    .Y(_04302_),
    .B1(_04300_));
 sg13g2_a21o_1 _12982_ (.A2(_04287_),
    .A1(_04285_),
    .B1(_04300_),
    .X(_04303_));
 sg13g2_nand2_1 _12983_ (.Y(_04304_),
    .A(_04301_),
    .B(_04303_));
 sg13g2_xnor2_1 _12984_ (.Y(_04305_),
    .A(_04299_),
    .B(_04304_));
 sg13g2_a21oi_1 _12985_ (.A1(net4924),
    .A2(_04305_),
    .Y(_00267_),
    .B1(_04298_));
 sg13g2_and2_1 _12986_ (.A(net4925),
    .B(_04301_),
    .X(_04306_));
 sg13g2_o21ai_1 _12987_ (.B1(_04306_),
    .Y(_04307_),
    .A1(_04299_),
    .A2(_04302_));
 sg13g2_o21ai_1 _12988_ (.B1(net4646),
    .Y(_00268_),
    .A1(_02356_),
    .A2(net4924));
 sg13g2_o21ai_1 _12989_ (.B1(net4646),
    .Y(_00269_),
    .A1(_02357_),
    .A2(net4924));
 sg13g2_o21ai_1 _12990_ (.B1(net4646),
    .Y(_00270_),
    .A1(_02358_),
    .A2(net4924));
 sg13g2_o21ai_1 _12991_ (.B1(_04307_),
    .Y(_00271_),
    .A1(_02359_),
    .A2(net4924));
 sg13g2_o21ai_1 _12992_ (.B1(_04307_),
    .Y(_00272_),
    .A1(_02360_),
    .A2(net4924));
 sg13g2_o21ai_1 _12993_ (.B1(_04307_),
    .Y(_00273_),
    .A1(_02361_),
    .A2(net4927));
 sg13g2_o21ai_1 _12994_ (.B1(net4646),
    .Y(_00274_),
    .A1(_02362_),
    .A2(net4927));
 sg13g2_o21ai_1 _12995_ (.B1(net4646),
    .Y(_00275_),
    .A1(_02363_),
    .A2(net4927));
 sg13g2_o21ai_1 _12996_ (.B1(net4646),
    .Y(_00276_),
    .A1(_02364_),
    .A2(net4927));
 sg13g2_o21ai_1 _12997_ (.B1(net4646),
    .Y(_00278_),
    .A1(_02365_),
    .A2(net4927));
 sg13g2_o21ai_1 _12998_ (.B1(net4646),
    .Y(_00279_),
    .A1(_02366_),
    .A2(net4927));
 sg13g2_nand2_1 _12999_ (.Y(_04308_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[0] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_xor2_1 _13000_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[0] ),
    .X(_01148_));
 sg13g2_nand2_1 _13001_ (.Y(_04309_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_nor2_1 _13002_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[1] ),
    .Y(_04310_));
 sg13g2_xor2_1 _13003_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[1] ),
    .X(_04311_));
 sg13g2_xnor2_1 _13004_ (.Y(_01158_),
    .A(_04308_),
    .B(_04311_));
 sg13g2_o21ai_1 _13005_ (.B1(_04309_),
    .Y(_04312_),
    .A1(_04308_),
    .A2(_04310_));
 sg13g2_xnor2_1 _13006_ (.Y(_04313_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[2] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_nor2b_1 _13007_ (.A(_04313_),
    .B_N(_04312_),
    .Y(_04314_));
 sg13g2_xnor2_1 _13008_ (.Y(_01159_),
    .A(_04312_),
    .B(_04313_));
 sg13g2_a21o_1 _13009_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[2] ),
    .B1(_04314_),
    .X(_04315_));
 sg13g2_xnor2_1 _13010_ (.Y(_04316_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[3] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_nor2b_1 _13011_ (.A(_04316_),
    .B_N(_04315_),
    .Y(_04317_));
 sg13g2_xnor2_1 _13012_ (.Y(_01160_),
    .A(_04315_),
    .B(_04316_));
 sg13g2_a21o_1 _13013_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[3] ),
    .B1(_04317_),
    .X(_04318_));
 sg13g2_xnor2_1 _13014_ (.Y(_04319_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[4] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_nor2b_1 _13015_ (.A(_04319_),
    .B_N(_04318_),
    .Y(_04320_));
 sg13g2_xnor2_1 _13016_ (.Y(_01161_),
    .A(_04318_),
    .B(_04319_));
 sg13g2_a21o_1 _13017_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[4] ),
    .B1(_04320_),
    .X(_04321_));
 sg13g2_nand2_1 _13018_ (.Y(_04322_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _13019_ (.Y(_04323_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _13020_ (.Y(_01162_),
    .A(_04321_),
    .B(_04323_));
 sg13g2_xnor2_1 _13021_ (.Y(_04324_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[6] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_o21ai_1 _13022_ (.B1(_04321_),
    .Y(_04325_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_a21oi_1 _13023_ (.A1(_04322_),
    .A2(_04325_),
    .Y(_04326_),
    .B1(_04324_));
 sg13g2_nand3_1 _13024_ (.B(_04324_),
    .C(_04325_),
    .A(_04322_),
    .Y(_04327_));
 sg13g2_nor2b_1 _13025_ (.A(_04326_),
    .B_N(_04327_),
    .Y(_01163_));
 sg13g2_a21oi_1 _13026_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[6] ),
    .Y(_04328_),
    .B1(_04326_));
 sg13g2_nand2_1 _13027_ (.Y(_04329_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_nor2_1 _13028_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[7] ),
    .Y(_04330_));
 sg13g2_xor2_1 _13029_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[7] ),
    .X(_04331_));
 sg13g2_xnor2_1 _13030_ (.Y(_01164_),
    .A(_04328_),
    .B(_04331_));
 sg13g2_o21ai_1 _13031_ (.B1(_04329_),
    .Y(_04332_),
    .A1(_04328_),
    .A2(_04330_));
 sg13g2_xnor2_1 _13032_ (.Y(_04333_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[8] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_nor2b_1 _13033_ (.A(_04333_),
    .B_N(_04332_),
    .Y(_04334_));
 sg13g2_xnor2_1 _13034_ (.Y(_01165_),
    .A(_04332_),
    .B(_04333_));
 sg13g2_a21o_1 _13035_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[8] ),
    .B1(_04334_),
    .X(_04335_));
 sg13g2_xnor2_1 _13036_ (.Y(_04336_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[9] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _13037_ (.Y(_01166_),
    .A(_04335_),
    .B(_04336_));
 sg13g2_nand2_1 _13038_ (.Y(_04337_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_nor2_1 _13039_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[10] ),
    .Y(_04338_));
 sg13g2_xor2_1 _13040_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[10] ),
    .X(_04339_));
 sg13g2_a21o_1 _13041_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[9] ),
    .B1(_04335_),
    .X(_04340_));
 sg13g2_o21ai_1 _13042_ (.B1(_04340_),
    .Y(_04341_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _13043_ (.Y(_01149_),
    .A(_04339_),
    .B(_04341_));
 sg13g2_o21ai_1 _13044_ (.B1(_04337_),
    .Y(_04342_),
    .A1(_04338_),
    .A2(_04341_));
 sg13g2_xnor2_1 _13045_ (.Y(_04343_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[11] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _13046_ (.Y(_01150_),
    .A(_04342_),
    .B(_04343_));
 sg13g2_xor2_1 _13047_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[12] ),
    .X(_04344_));
 sg13g2_a21o_1 _13048_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[11] ),
    .B1(_04342_),
    .X(_04345_));
 sg13g2_o21ai_1 _13049_ (.B1(_04345_),
    .Y(_04346_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_nand2b_1 _13050_ (.Y(_04347_),
    .B(_04344_),
    .A_N(_04346_));
 sg13g2_xnor2_1 _13051_ (.Y(_01151_),
    .A(_04344_),
    .B(_04346_));
 sg13g2_o21ai_1 _13052_ (.B1(_04347_),
    .Y(_04348_),
    .A1(_02368_),
    .A2(_02369_));
 sg13g2_xnor2_1 _13053_ (.Y(_04349_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[13] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_xnor2_1 _13054_ (.Y(_01152_),
    .A(_04348_),
    .B(_04349_));
 sg13g2_xor2_1 _13055_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[14] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[14] ),
    .X(_04350_));
 sg13g2_a21o_1 _13056_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[13] ),
    .B1(_04348_),
    .X(_04351_));
 sg13g2_o21ai_1 _13057_ (.B1(_04351_),
    .Y(_04352_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_nor2b_1 _13058_ (.A(_04352_),
    .B_N(_04350_),
    .Y(_04353_));
 sg13g2_xnor2_1 _13059_ (.Y(_01153_),
    .A(_04350_),
    .B(_04352_));
 sg13g2_a21o_1 _13060_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[14] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[14] ),
    .B1(_04353_),
    .X(_04354_));
 sg13g2_and2_1 _13061_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[15] ),
    .X(_04355_));
 sg13g2_or2_1 _13062_ (.X(_04356_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[15] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand2b_1 _13063_ (.Y(_04357_),
    .B(_04356_),
    .A_N(_04355_));
 sg13g2_xnor2_1 _13064_ (.Y(_01154_),
    .A(_04354_),
    .B(_04357_));
 sg13g2_and2_1 _13065_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[16] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[16] ),
    .X(_04358_));
 sg13g2_xor2_1 _13066_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[16] ),
    .X(_04359_));
 sg13g2_a21o_1 _13067_ (.A2(_04356_),
    .A1(_04354_),
    .B1(_04355_),
    .X(_04360_));
 sg13g2_xor2_1 _13068_ (.B(_04360_),
    .A(_04359_),
    .X(_01155_));
 sg13g2_a21o_1 _13069_ (.A2(_04360_),
    .A1(_04359_),
    .B1(_04358_),
    .X(_04361_));
 sg13g2_xnor2_1 _13070_ (.Y(_04362_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[17] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xnor2_1 _13071_ (.Y(_01156_),
    .A(_04361_),
    .B(_04362_));
 sg13g2_a21o_1 _13072_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[17] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[17] ),
    .B1(_04361_),
    .X(_04363_));
 sg13g2_o21ai_1 _13073_ (.B1(_04363_),
    .Y(_04364_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xor2_1 _13074_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[18] ),
    .X(_04365_));
 sg13g2_xnor2_1 _13075_ (.Y(_01157_),
    .A(_04364_),
    .B(_04365_));
 sg13g2_nand2b_1 _13076_ (.Y(_04366_),
    .B(net4958),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_nor2b_1 _13077_ (.A(net4958),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[1] ),
    .Y(_04367_));
 sg13g2_xnor2_1 _13078_ (.Y(_04368_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[1] ),
    .B(net4958));
 sg13g2_xnor2_1 _13079_ (.Y(_01139_),
    .A(_01186_),
    .B(_04368_));
 sg13g2_xnor2_1 _13080_ (.Y(_04369_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[2] ),
    .B(net4958));
 sg13g2_o21ai_1 _13081_ (.B1(_04366_),
    .Y(_04370_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[0] ),
    .A2(_04367_));
 sg13g2_nor2b_1 _13082_ (.A(_04370_),
    .B_N(_04369_),
    .Y(_04371_));
 sg13g2_xnor2_1 _13083_ (.Y(_01140_),
    .A(_04369_),
    .B(_04370_));
 sg13g2_a21oi_1 _13084_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[2] ),
    .A2(net4949),
    .Y(_04372_),
    .B1(_04371_));
 sg13g2_nor2_1 _13085_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4949),
    .Y(_04373_));
 sg13g2_nand2_1 _13086_ (.Y(_04374_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4949));
 sg13g2_nor2b_1 _13087_ (.A(_04373_),
    .B_N(_04374_),
    .Y(_04375_));
 sg13g2_xnor2_1 _13088_ (.Y(_01141_),
    .A(_04372_),
    .B(_04375_));
 sg13g2_xnor2_1 _13089_ (.Y(_04376_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[4] ),
    .B(net4958));
 sg13g2_o21ai_1 _13090_ (.B1(_04374_),
    .Y(_04377_),
    .A1(_04372_),
    .A2(_04373_));
 sg13g2_and2_1 _13091_ (.A(_04376_),
    .B(_04377_),
    .X(_04378_));
 sg13g2_xor2_1 _13092_ (.B(_04377_),
    .A(_04376_),
    .X(_01142_));
 sg13g2_xnor2_1 _13093_ (.Y(_04379_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[5] ),
    .B(net4957));
 sg13g2_a21oi_1 _13094_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[4] ),
    .A2(net4949),
    .Y(_04380_),
    .B1(_04378_));
 sg13g2_xnor2_1 _13095_ (.Y(_01143_),
    .A(_04379_),
    .B(_04380_));
 sg13g2_o21ai_1 _13096_ (.B1(net4949),
    .Y(_04381_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[4] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_and2_1 _13097_ (.A(_04378_),
    .B(_04379_),
    .X(_04382_));
 sg13g2_nor2b_1 _13098_ (.A(_04382_),
    .B_N(_04381_),
    .Y(_04383_));
 sg13g2_nand2_1 _13099_ (.Y(_04384_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4949));
 sg13g2_nor2_1 _13100_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4949),
    .Y(_04385_));
 sg13g2_xnor2_1 _13101_ (.Y(_04386_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4957));
 sg13g2_xnor2_1 _13102_ (.Y(_01144_),
    .A(_04383_),
    .B(_04386_));
 sg13g2_nand2b_1 _13103_ (.Y(_04387_),
    .B(net4957),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_xor2_1 _13104_ (.B(net4957),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[7] ),
    .X(_04388_));
 sg13g2_o21ai_1 _13105_ (.B1(_04384_),
    .Y(_04389_),
    .A1(_04383_),
    .A2(_04385_));
 sg13g2_xnor2_1 _13106_ (.Y(_01145_),
    .A(_04388_),
    .B(_04389_));
 sg13g2_xnor2_1 _13107_ (.Y(_04390_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[8] ),
    .B(net4957));
 sg13g2_o21ai_1 _13108_ (.B1(net4948),
    .Y(_04391_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_nand3_1 _13109_ (.B(_04386_),
    .C(_04387_),
    .A(_04382_),
    .Y(_04392_));
 sg13g2_and3_1 _13110_ (.X(_04393_),
    .A(_04381_),
    .B(_04391_),
    .C(_04392_));
 sg13g2_nand2b_1 _13111_ (.Y(_04394_),
    .B(_04390_),
    .A_N(_04393_));
 sg13g2_xnor2_1 _13112_ (.Y(_01146_),
    .A(_04390_),
    .B(_04393_));
 sg13g2_xor2_1 _13113_ (.B(net4957),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[9] ),
    .X(_04395_));
 sg13g2_o21ai_1 _13114_ (.B1(_04394_),
    .Y(_04396_),
    .A1(_02367_),
    .A2(net4957));
 sg13g2_xnor2_1 _13115_ (.Y(_01147_),
    .A(_04395_),
    .B(_04396_));
 sg13g2_o21ai_1 _13116_ (.B1(net4948),
    .Y(_04397_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[8] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_nor2_1 _13117_ (.A(_04394_),
    .B(_04395_),
    .Y(_04398_));
 sg13g2_nor2b_1 _13118_ (.A(_04398_),
    .B_N(_04397_),
    .Y(_04399_));
 sg13g2_nand2_1 _13119_ (.Y(_04400_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4948));
 sg13g2_nor2_1 _13120_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4948),
    .Y(_04401_));
 sg13g2_xnor2_1 _13121_ (.Y(_04402_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4956));
 sg13g2_xnor2_1 _13122_ (.Y(_01130_),
    .A(_04399_),
    .B(_04402_));
 sg13g2_xor2_1 _13123_ (.B(net4956),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[11] ),
    .X(_04403_));
 sg13g2_o21ai_1 _13124_ (.B1(_04400_),
    .Y(_04404_),
    .A1(_04399_),
    .A2(_04401_));
 sg13g2_xnor2_1 _13125_ (.Y(_01131_),
    .A(_04403_),
    .B(_04404_));
 sg13g2_xnor2_1 _13126_ (.Y(_04405_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[12] ),
    .B(net4954));
 sg13g2_nand2_1 _13127_ (.Y(_04406_),
    .A(_04398_),
    .B(_04402_));
 sg13g2_nor2_1 _13128_ (.A(_04403_),
    .B(_04406_),
    .Y(_04407_));
 sg13g2_o21ai_1 _13129_ (.B1(net4948),
    .Y(_04408_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[10] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_nand2_1 _13130_ (.Y(_04409_),
    .A(_04397_),
    .B(_04408_));
 sg13g2_inv_1 _13131_ (.Y(_04410_),
    .A(_04409_));
 sg13g2_o21ai_1 _13132_ (.B1(_04405_),
    .Y(_04411_),
    .A1(_04407_),
    .A2(_04409_));
 sg13g2_or3_1 _13133_ (.A(_04405_),
    .B(_04407_),
    .C(_04409_),
    .X(_04412_));
 sg13g2_and2_1 _13134_ (.A(_04411_),
    .B(_04412_),
    .X(_01132_));
 sg13g2_nand2_1 _13135_ (.Y(_04413_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[13] ),
    .B(net4948));
 sg13g2_nand2_1 _13136_ (.Y(_04414_),
    .A(_02370_),
    .B(net4954));
 sg13g2_nand2_1 _13137_ (.Y(_04415_),
    .A(_04413_),
    .B(_04414_));
 sg13g2_o21ai_1 _13138_ (.B1(_04411_),
    .Y(_04416_),
    .A1(_02368_),
    .A2(net4954));
 sg13g2_xnor2_1 _13139_ (.Y(_01133_),
    .A(_04415_),
    .B(_04416_));
 sg13g2_nor2b_1 _13140_ (.A(net4954),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[14] ),
    .Y(_04417_));
 sg13g2_xnor2_1 _13141_ (.Y(_04418_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[14] ),
    .B(net4954));
 sg13g2_o21ai_1 _13142_ (.B1(net4948),
    .Y(_04419_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[12] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_a22oi_1 _13143_ (.Y(_04420_),
    .B1(_04411_),
    .B2(_04419_),
    .A2(net4954),
    .A1(_02370_));
 sg13g2_xor2_1 _13144_ (.B(_04420_),
    .A(_04418_),
    .X(_01134_));
 sg13g2_xnor2_1 _13145_ (.Y(_04421_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[15] ),
    .B(net4954));
 sg13g2_a21oi_1 _13146_ (.A1(_04418_),
    .A2(_04420_),
    .Y(_04422_),
    .B1(_04417_));
 sg13g2_xnor2_1 _13147_ (.Y(_01135_),
    .A(_04421_),
    .B(_04422_));
 sg13g2_and4_1 _13148_ (.A(_04405_),
    .B(_04413_),
    .C(_04414_),
    .D(_04421_),
    .X(_04423_));
 sg13g2_nand3_1 _13149_ (.B(_04418_),
    .C(_04423_),
    .A(_04407_),
    .Y(_04424_));
 sg13g2_o21ai_1 _13150_ (.B1(net4948),
    .Y(_04425_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand4_1 _13151_ (.B(_04419_),
    .C(_04424_),
    .A(_04410_),
    .Y(_04426_),
    .D(_04425_));
 sg13g2_nor2b_1 _13152_ (.A(net4955),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[16] ),
    .Y(_04427_));
 sg13g2_xnor2_1 _13153_ (.Y(_04428_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[16] ),
    .B(net4955));
 sg13g2_xor2_1 _13154_ (.B(_04428_),
    .A(_04426_),
    .X(_01136_));
 sg13g2_a21o_1 _13155_ (.A2(_04428_),
    .A1(_04426_),
    .B1(_04427_),
    .X(_04429_));
 sg13g2_xor2_1 _13156_ (.B(net4955),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[17] ),
    .X(_04430_));
 sg13g2_xnor2_1 _13157_ (.Y(_01137_),
    .A(_04429_),
    .B(_04430_));
 sg13g2_nor3_1 _13158_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[17] ),
    .B(net4955),
    .C(_04429_),
    .Y(_04431_));
 sg13g2_nand3_1 _13159_ (.B(net4954),
    .C(_04429_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[17] ),
    .Y(_04432_));
 sg13g2_nor2b_1 _13160_ (.A(_04431_),
    .B_N(_04432_),
    .Y(_04433_));
 sg13g2_xnor2_1 _13161_ (.Y(_01138_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[18] ),
    .B(_04433_));
 sg13g2_nand2_1 _13162_ (.Y(_04434_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[0] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_xor2_1 _13163_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[0] ),
    .X(_00509_));
 sg13g2_nand2_1 _13164_ (.Y(_04435_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_nor2_1 _13165_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[1] ),
    .Y(_04436_));
 sg13g2_xor2_1 _13166_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[1] ),
    .X(_04437_));
 sg13g2_xnor2_1 _13167_ (.Y(_00519_),
    .A(_04434_),
    .B(_04437_));
 sg13g2_o21ai_1 _13168_ (.B1(_04435_),
    .Y(_04438_),
    .A1(_04434_),
    .A2(_04436_));
 sg13g2_xnor2_1 _13169_ (.Y(_04439_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[2] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_nor2b_1 _13170_ (.A(_04439_),
    .B_N(_04438_),
    .Y(_04440_));
 sg13g2_xnor2_1 _13171_ (.Y(_00520_),
    .A(_04438_),
    .B(_04439_));
 sg13g2_a21o_1 _13172_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[2] ),
    .B1(_04440_),
    .X(_04441_));
 sg13g2_xnor2_1 _13173_ (.Y(_04442_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[3] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_nor2b_1 _13174_ (.A(_04442_),
    .B_N(_04441_),
    .Y(_04443_));
 sg13g2_xnor2_1 _13175_ (.Y(_00521_),
    .A(_04441_),
    .B(_04442_));
 sg13g2_a21o_1 _13176_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[3] ),
    .B1(_04443_),
    .X(_04444_));
 sg13g2_xnor2_1 _13177_ (.Y(_04445_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[4] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_nor2b_1 _13178_ (.A(_04445_),
    .B_N(_04444_),
    .Y(_04446_));
 sg13g2_xnor2_1 _13179_ (.Y(_00522_),
    .A(_04444_),
    .B(_04445_));
 sg13g2_a21o_1 _13180_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[4] ),
    .B1(_04446_),
    .X(_04447_));
 sg13g2_nand2_1 _13181_ (.Y(_04448_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[5] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_xnor2_1 _13182_ (.Y(_04449_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[5] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_xnor2_1 _13183_ (.Y(_00523_),
    .A(_04447_),
    .B(_04449_));
 sg13g2_xnor2_1 _13184_ (.Y(_04450_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[6] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_o21ai_1 _13185_ (.B1(_04447_),
    .Y(_04451_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_a21oi_1 _13186_ (.A1(_04448_),
    .A2(_04451_),
    .Y(_04452_),
    .B1(_04450_));
 sg13g2_nand3_1 _13187_ (.B(_04450_),
    .C(_04451_),
    .A(_04448_),
    .Y(_04453_));
 sg13g2_nor2b_1 _13188_ (.A(_04452_),
    .B_N(_04453_),
    .Y(_00524_));
 sg13g2_a21oi_1 _13189_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[6] ),
    .Y(_04454_),
    .B1(_04452_));
 sg13g2_nand2_1 _13190_ (.Y(_04455_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[7] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_nor2_1 _13191_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[7] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[7] ),
    .Y(_04456_));
 sg13g2_xor2_1 _13192_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[7] ),
    .X(_04457_));
 sg13g2_xnor2_1 _13193_ (.Y(_00525_),
    .A(_04454_),
    .B(_04457_));
 sg13g2_o21ai_1 _13194_ (.B1(_04455_),
    .Y(_04458_),
    .A1(_04454_),
    .A2(_04456_));
 sg13g2_xnor2_1 _13195_ (.Y(_04459_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[8] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_nor2b_1 _13196_ (.A(_04459_),
    .B_N(_04458_),
    .Y(_04460_));
 sg13g2_xnor2_1 _13197_ (.Y(_00526_),
    .A(_04458_),
    .B(_04459_));
 sg13g2_a21o_1 _13198_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[8] ),
    .B1(_04460_),
    .X(_04461_));
 sg13g2_xnor2_1 _13199_ (.Y(_04462_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[9] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_xnor2_1 _13200_ (.Y(_00527_),
    .A(_04461_),
    .B(_04462_));
 sg13g2_nand2_1 _13201_ (.Y(_04463_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[10] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_nor2_1 _13202_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[10] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[10] ),
    .Y(_04464_));
 sg13g2_xor2_1 _13203_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[10] ),
    .X(_04465_));
 sg13g2_a21o_1 _13204_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[9] ),
    .B1(_04461_),
    .X(_04466_));
 sg13g2_o21ai_1 _13205_ (.B1(_04466_),
    .Y(_04467_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_xnor2_1 _13206_ (.Y(_00510_),
    .A(_04465_),
    .B(_04467_));
 sg13g2_o21ai_1 _13207_ (.B1(_04463_),
    .Y(_04468_),
    .A1(_04464_),
    .A2(_04467_));
 sg13g2_xnor2_1 _13208_ (.Y(_04469_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[11] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_xnor2_1 _13209_ (.Y(_00511_),
    .A(_04468_),
    .B(_04469_));
 sg13g2_nand2_1 _13210_ (.Y(_04470_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[12] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_nor2_1 _13211_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[12] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[12] ),
    .Y(_04471_));
 sg13g2_xor2_1 _13212_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[12] ),
    .X(_04472_));
 sg13g2_a21o_1 _13213_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[11] ),
    .B1(_04468_),
    .X(_04473_));
 sg13g2_o21ai_1 _13214_ (.B1(_04473_),
    .Y(_04474_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_xnor2_1 _13215_ (.Y(_00512_),
    .A(_04472_),
    .B(_04474_));
 sg13g2_o21ai_1 _13216_ (.B1(_04470_),
    .Y(_04475_),
    .A1(_04471_),
    .A2(_04474_));
 sg13g2_xnor2_1 _13217_ (.Y(_04476_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[13] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_xnor2_1 _13218_ (.Y(_00513_),
    .A(_04475_),
    .B(_04476_));
 sg13g2_xor2_1 _13219_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[14] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[14] ),
    .X(_04477_));
 sg13g2_a21o_1 _13220_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[13] ),
    .B1(_04475_),
    .X(_04478_));
 sg13g2_o21ai_1 _13221_ (.B1(_04478_),
    .Y(_04479_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_nor2b_1 _13222_ (.A(_04479_),
    .B_N(_04477_),
    .Y(_04480_));
 sg13g2_xnor2_1 _13223_ (.Y(_00514_),
    .A(_04477_),
    .B(_04479_));
 sg13g2_a21o_1 _13224_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[14] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[14] ),
    .B1(_04480_),
    .X(_04481_));
 sg13g2_nand2_1 _13225_ (.Y(_04482_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_xnor2_1 _13226_ (.Y(_04483_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_xnor2_1 _13227_ (.Y(_00515_),
    .A(_04481_),
    .B(_04483_));
 sg13g2_nand2_1 _13228_ (.Y(_04484_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[16] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_xor2_1 _13229_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[16] ),
    .X(_04485_));
 sg13g2_o21ai_1 _13230_ (.B1(_04481_),
    .Y(_04486_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[15] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_nand2_1 _13231_ (.Y(_04487_),
    .A(_04482_),
    .B(_04486_));
 sg13g2_nand2_1 _13232_ (.Y(_04488_),
    .A(_04485_),
    .B(_04487_));
 sg13g2_xor2_1 _13233_ (.B(_04487_),
    .A(_04485_),
    .X(_00516_));
 sg13g2_xnor2_1 _13234_ (.Y(_04489_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[17] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_a21oi_1 _13235_ (.A1(_04484_),
    .A2(_04488_),
    .Y(_04490_),
    .B1(_04489_));
 sg13g2_nand3_1 _13236_ (.B(_04488_),
    .C(_04489_),
    .A(_04484_),
    .Y(_04491_));
 sg13g2_nor2b_1 _13237_ (.A(_04490_),
    .B_N(_04491_),
    .Y(_00517_));
 sg13g2_a21oi_1 _13238_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[17] ),
    .Y(_04492_),
    .B1(_04490_));
 sg13g2_xor2_1 _13239_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[18] ),
    .X(_04493_));
 sg13g2_xnor2_1 _13240_ (.Y(_00518_),
    .A(_04492_),
    .B(_04493_));
 sg13g2_nor2b_1 _13241_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][1] ),
    .Y(_04494_));
 sg13g2_xnor2_1 _13242_ (.Y(_04495_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][1] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _13243_ (.B(_04495_),
    .A(_02507_),
    .X(_00538_));
 sg13g2_a21oi_1 _13244_ (.A1(_02507_),
    .A2(_04495_),
    .Y(_04496_),
    .B1(_04494_));
 sg13g2_xnor2_1 _13245_ (.Y(_04497_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][2] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _13246_ (.A(_04496_),
    .B_N(_04497_),
    .Y(_04498_));
 sg13g2_xnor2_1 _13247_ (.Y(_00539_),
    .A(_04496_),
    .B(_04497_));
 sg13g2_a21oi_1 _13248_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][2] ),
    .A2(_02372_),
    .Y(_04499_),
    .B1(_04498_));
 sg13g2_xnor2_1 _13249_ (.Y(_04500_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][3] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _13250_ (.A(_04499_),
    .B_N(_04500_),
    .Y(_04501_));
 sg13g2_xnor2_1 _13251_ (.Y(_00540_),
    .A(_04499_),
    .B(_04500_));
 sg13g2_a21oi_1 _13252_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][3] ),
    .A2(_02373_),
    .Y(_04502_),
    .B1(_04501_));
 sg13g2_xnor2_1 _13253_ (.Y(_04503_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][4] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _13254_ (.A(_04502_),
    .B_N(_04503_),
    .Y(_04504_));
 sg13g2_xnor2_1 _13255_ (.Y(_00541_),
    .A(_04502_),
    .B(_04503_));
 sg13g2_a21oi_1 _13256_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][4] ),
    .A2(_02374_),
    .Y(_04505_),
    .B1(_04504_));
 sg13g2_xnor2_1 _13257_ (.Y(_04506_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][5] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _13258_ (.A(_04505_),
    .B_N(_04506_),
    .Y(_04507_));
 sg13g2_xnor2_1 _13259_ (.Y(_00542_),
    .A(_04505_),
    .B(_04506_));
 sg13g2_a21oi_1 _13260_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][5] ),
    .A2(_02375_),
    .Y(_04508_),
    .B1(_04507_));
 sg13g2_xnor2_1 _13261_ (.Y(_04509_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][6] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_nor2b_1 _13262_ (.A(_04508_),
    .B_N(_04509_),
    .Y(_04510_));
 sg13g2_xnor2_1 _13263_ (.Y(_00543_),
    .A(_04508_),
    .B(_04509_));
 sg13g2_a21oi_1 _13264_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][6] ),
    .A2(_02376_),
    .Y(_04511_),
    .B1(_04510_));
 sg13g2_xnor2_1 _13265_ (.Y(_04512_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][7] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _13266_ (.A(_04511_),
    .B_N(_04512_),
    .Y(_04513_));
 sg13g2_xnor2_1 _13267_ (.Y(_00544_),
    .A(_04511_),
    .B(_04512_));
 sg13g2_a21oi_1 _13268_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][7] ),
    .A2(_02377_),
    .Y(_04514_),
    .B1(_04513_));
 sg13g2_xnor2_1 _13269_ (.Y(_04515_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][8] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_nor2b_1 _13270_ (.A(_04514_),
    .B_N(_04515_),
    .Y(_04516_));
 sg13g2_xnor2_1 _13271_ (.Y(_00545_),
    .A(_04514_),
    .B(_04515_));
 sg13g2_a21oi_1 _13272_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][8] ),
    .A2(_02378_),
    .Y(_04517_),
    .B1(_04516_));
 sg13g2_nand2b_1 _13273_ (.Y(_04518_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][9] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _13274_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][9] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[9] ),
    .Y(_04519_));
 sg13g2_xnor2_1 _13275_ (.Y(_04520_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][9] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_xnor2_1 _13276_ (.Y(_00546_),
    .A(_04517_),
    .B(_04520_));
 sg13g2_nor2b_1 _13277_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][10] ),
    .Y(_04521_));
 sg13g2_nand2b_1 _13278_ (.Y(_04522_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][10] ));
 sg13g2_nand2b_1 _13279_ (.Y(_04523_),
    .B(_04522_),
    .A_N(_04521_));
 sg13g2_o21ai_1 _13280_ (.B1(_04518_),
    .Y(_04524_),
    .A1(_04517_),
    .A2(_04519_));
 sg13g2_xnor2_1 _13281_ (.Y(_00529_),
    .A(_04523_),
    .B(_04524_));
 sg13g2_a21oi_1 _13282_ (.A1(_04522_),
    .A2(_04524_),
    .Y(_04525_),
    .B1(_04521_));
 sg13g2_nand2b_1 _13283_ (.Y(_04526_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][11] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _13284_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][11] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[11] ),
    .Y(_04527_));
 sg13g2_xnor2_1 _13285_ (.Y(_04528_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][11] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_xnor2_1 _13286_ (.Y(_00530_),
    .A(_04525_),
    .B(_04528_));
 sg13g2_nor2b_1 _13287_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][12] ),
    .Y(_04529_));
 sg13g2_nand2b_1 _13288_ (.Y(_04530_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][12] ));
 sg13g2_nand2b_1 _13289_ (.Y(_04531_),
    .B(_04530_),
    .A_N(_04529_));
 sg13g2_o21ai_1 _13290_ (.B1(_04526_),
    .Y(_04532_),
    .A1(_04525_),
    .A2(_04527_));
 sg13g2_xnor2_1 _13291_ (.Y(_00531_),
    .A(_04531_),
    .B(_04532_));
 sg13g2_a21oi_1 _13292_ (.A1(_04530_),
    .A2(_04532_),
    .Y(_04533_),
    .B1(_04529_));
 sg13g2_nand2b_1 _13293_ (.Y(_04534_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][13] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _13294_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][13] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[13] ),
    .Y(_04535_));
 sg13g2_xnor2_1 _13295_ (.Y(_04536_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][13] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_xnor2_1 _13296_ (.Y(_00532_),
    .A(_04533_),
    .B(_04536_));
 sg13g2_nor2b_1 _13297_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][14] ),
    .Y(_04537_));
 sg13g2_nand2b_1 _13298_ (.Y(_04538_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][14] ));
 sg13g2_nand2b_1 _13299_ (.Y(_04539_),
    .B(_04538_),
    .A_N(_04537_));
 sg13g2_o21ai_1 _13300_ (.B1(_04534_),
    .Y(_04540_),
    .A1(_04533_),
    .A2(_04535_));
 sg13g2_xnor2_1 _13301_ (.Y(_00533_),
    .A(_04539_),
    .B(_04540_));
 sg13g2_a21oi_1 _13302_ (.A1(_04538_),
    .A2(_04540_),
    .Y(_04541_),
    .B1(_04537_));
 sg13g2_nand2b_1 _13303_ (.Y(_04542_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][15] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _13304_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][15] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[15] ),
    .Y(_04543_));
 sg13g2_xnor2_1 _13305_ (.Y(_04544_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][15] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_xnor2_1 _13306_ (.Y(_00534_),
    .A(_04541_),
    .B(_04544_));
 sg13g2_xor2_1 _13307_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][16] ),
    .X(_04545_));
 sg13g2_o21ai_1 _13308_ (.B1(_04542_),
    .Y(_04546_),
    .A1(_04541_),
    .A2(_04543_));
 sg13g2_nor2b_1 _13309_ (.A(_04545_),
    .B_N(_04546_),
    .Y(_04547_));
 sg13g2_xnor2_1 _13310_ (.Y(_00535_),
    .A(_04545_),
    .B(_04546_));
 sg13g2_a21oi_2 _13311_ (.B1(_04547_),
    .Y(_04548_),
    .A2(_02379_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][16] ));
 sg13g2_nand2b_1 _13312_ (.Y(_04549_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][17] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _13313_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][17] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[17] ),
    .Y(_04550_));
 sg13g2_xnor2_1 _13314_ (.Y(_04551_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][17] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _13315_ (.Y(_00536_),
    .A(_04548_),
    .B(_04551_));
 sg13g2_o21ai_1 _13316_ (.B1(_04549_),
    .Y(_04552_),
    .A1(_04548_),
    .A2(_04550_));
 sg13g2_xor2_1 _13317_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][18] ),
    .X(_04553_));
 sg13g2_xnor2_1 _13318_ (.Y(_00537_),
    .A(_04552_),
    .B(_04553_));
 sg13g2_nand2_1 _13319_ (.Y(_04554_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[0] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_xor2_1 _13320_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[0] ),
    .X(_00490_));
 sg13g2_nand2_1 _13321_ (.Y(_04555_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_nor2_1 _13322_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[1] ),
    .Y(_04556_));
 sg13g2_xor2_1 _13323_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[1] ),
    .X(_04557_));
 sg13g2_xnor2_1 _13324_ (.Y(_00500_),
    .A(_04554_),
    .B(_04557_));
 sg13g2_o21ai_1 _13325_ (.B1(_04555_),
    .Y(_04558_),
    .A1(_04554_),
    .A2(_04556_));
 sg13g2_xnor2_1 _13326_ (.Y(_04559_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[2] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_nor2b_1 _13327_ (.A(_04559_),
    .B_N(_04558_),
    .Y(_04560_));
 sg13g2_xnor2_1 _13328_ (.Y(_00501_),
    .A(_04558_),
    .B(_04559_));
 sg13g2_a21o_1 _13329_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[2] ),
    .B1(_04560_),
    .X(_04561_));
 sg13g2_xnor2_1 _13330_ (.Y(_04562_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[3] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_nor2b_1 _13331_ (.A(_04562_),
    .B_N(_04561_),
    .Y(_04563_));
 sg13g2_xnor2_1 _13332_ (.Y(_00502_),
    .A(_04561_),
    .B(_04562_));
 sg13g2_a21o_1 _13333_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[3] ),
    .B1(_04563_),
    .X(_04564_));
 sg13g2_xnor2_1 _13334_ (.Y(_04565_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[4] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_nor2b_1 _13335_ (.A(_04565_),
    .B_N(_04564_),
    .Y(_04566_));
 sg13g2_xnor2_1 _13336_ (.Y(_00503_),
    .A(_04564_),
    .B(_04565_));
 sg13g2_a21o_1 _13337_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[4] ),
    .B1(_04566_),
    .X(_04567_));
 sg13g2_nand2_1 _13338_ (.Y(_04568_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _13339_ (.Y(_04569_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _13340_ (.Y(_00504_),
    .A(_04567_),
    .B(_04569_));
 sg13g2_xnor2_1 _13341_ (.Y(_04570_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[6] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_o21ai_1 _13342_ (.B1(_04567_),
    .Y(_04571_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_a21oi_1 _13343_ (.A1(_04568_),
    .A2(_04571_),
    .Y(_04572_),
    .B1(_04570_));
 sg13g2_nand3_1 _13344_ (.B(_04570_),
    .C(_04571_),
    .A(_04568_),
    .Y(_04573_));
 sg13g2_nor2b_1 _13345_ (.A(_04572_),
    .B_N(_04573_),
    .Y(_00505_));
 sg13g2_a21oi_1 _13346_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[6] ),
    .Y(_04574_),
    .B1(_04572_));
 sg13g2_nand2_1 _13347_ (.Y(_04575_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_nor2_1 _13348_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[7] ),
    .Y(_04576_));
 sg13g2_xor2_1 _13349_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[7] ),
    .X(_04577_));
 sg13g2_xnor2_1 _13350_ (.Y(_00506_),
    .A(_04574_),
    .B(_04577_));
 sg13g2_o21ai_1 _13351_ (.B1(_04575_),
    .Y(_04578_),
    .A1(_04574_),
    .A2(_04576_));
 sg13g2_xnor2_1 _13352_ (.Y(_04579_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[8] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_nor2b_1 _13353_ (.A(_04579_),
    .B_N(_04578_),
    .Y(_04580_));
 sg13g2_xnor2_1 _13354_ (.Y(_00507_),
    .A(_04578_),
    .B(_04579_));
 sg13g2_a21o_1 _13355_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[8] ),
    .B1(_04580_),
    .X(_04581_));
 sg13g2_xnor2_1 _13356_ (.Y(_04582_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[9] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _13357_ (.Y(_00508_),
    .A(_04581_),
    .B(_04582_));
 sg13g2_nand2_1 _13358_ (.Y(_04583_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_nor2_1 _13359_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[10] ),
    .Y(_04584_));
 sg13g2_xor2_1 _13360_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[10] ),
    .X(_04585_));
 sg13g2_a21o_1 _13361_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[9] ),
    .B1(_04581_),
    .X(_04586_));
 sg13g2_o21ai_1 _13362_ (.B1(_04586_),
    .Y(_04587_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _13363_ (.Y(_00491_),
    .A(_04585_),
    .B(_04587_));
 sg13g2_o21ai_1 _13364_ (.B1(_04583_),
    .Y(_04588_),
    .A1(_04584_),
    .A2(_04587_));
 sg13g2_xnor2_1 _13365_ (.Y(_04589_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[11] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _13366_ (.Y(_00492_),
    .A(_04588_),
    .B(_04589_));
 sg13g2_nand2_1 _13367_ (.Y(_04590_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[12] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_nor2_1 _13368_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[12] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[12] ),
    .Y(_04591_));
 sg13g2_xor2_1 _13369_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[12] ),
    .X(_04592_));
 sg13g2_a21o_1 _13370_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[11] ),
    .B1(_04588_),
    .X(_04593_));
 sg13g2_o21ai_1 _13371_ (.B1(_04593_),
    .Y(_04594_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _13372_ (.Y(_00493_),
    .A(_04592_),
    .B(_04594_));
 sg13g2_o21ai_1 _13373_ (.B1(_04590_),
    .Y(_04595_),
    .A1(_04591_),
    .A2(_04594_));
 sg13g2_xnor2_1 _13374_ (.Y(_04596_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[13] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_xnor2_1 _13375_ (.Y(_00494_),
    .A(_04595_),
    .B(_04596_));
 sg13g2_xor2_1 _13376_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[14] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[14] ),
    .X(_04597_));
 sg13g2_a21o_1 _13377_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[13] ),
    .B1(_04595_),
    .X(_04598_));
 sg13g2_o21ai_1 _13378_ (.B1(_04598_),
    .Y(_04599_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_nor2b_1 _13379_ (.A(_04599_),
    .B_N(_04597_),
    .Y(_04600_));
 sg13g2_xnor2_1 _13380_ (.Y(_00495_),
    .A(_04597_),
    .B(_04599_));
 sg13g2_a21o_1 _13381_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[14] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[14] ),
    .B1(_04600_),
    .X(_04601_));
 sg13g2_and2_1 _13382_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[15] ),
    .X(_04602_));
 sg13g2_or2_1 _13383_ (.X(_04603_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[15] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand2b_1 _13384_ (.Y(_04604_),
    .B(_04603_),
    .A_N(_04602_));
 sg13g2_xnor2_1 _13385_ (.Y(_00496_),
    .A(_04601_),
    .B(_04604_));
 sg13g2_and2_1 _13386_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[16] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[16] ),
    .X(_04605_));
 sg13g2_xor2_1 _13387_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[16] ),
    .X(_04606_));
 sg13g2_a21o_1 _13388_ (.A2(_04603_),
    .A1(_04601_),
    .B1(_04602_),
    .X(_04607_));
 sg13g2_xor2_1 _13389_ (.B(_04607_),
    .A(_04606_),
    .X(_00497_));
 sg13g2_a21o_1 _13390_ (.A2(_04607_),
    .A1(_04606_),
    .B1(_04605_),
    .X(_04608_));
 sg13g2_xnor2_1 _13391_ (.Y(_04609_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[17] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xnor2_1 _13392_ (.Y(_00498_),
    .A(_04608_),
    .B(_04609_));
 sg13g2_a21o_1 _13393_ (.A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[17] ),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[17] ),
    .B1(_04608_),
    .X(_04610_));
 sg13g2_o21ai_1 _13394_ (.B1(_04610_),
    .Y(_04611_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xor2_1 _13395_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[18] ),
    .X(_04612_));
 sg13g2_xnor2_1 _13396_ (.Y(_00499_),
    .A(_04611_),
    .B(_04612_));
 sg13g2_nand2b_1 _13397_ (.Y(_04613_),
    .B(net4977),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_nor2b_1 _13398_ (.A(net4977),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[1] ),
    .Y(_04614_));
 sg13g2_xnor2_1 _13399_ (.Y(_04615_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[1] ),
    .B(net4976));
 sg13g2_xnor2_1 _13400_ (.Y(_00481_),
    .A(_01193_),
    .B(_04615_));
 sg13g2_xnor2_1 _13401_ (.Y(_04616_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[2] ),
    .B(net4977));
 sg13g2_o21ai_1 _13402_ (.B1(_04613_),
    .Y(_04617_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[0] ),
    .A2(_04614_));
 sg13g2_nor2b_1 _13403_ (.A(_04617_),
    .B_N(_04616_),
    .Y(_04618_));
 sg13g2_xnor2_1 _13404_ (.Y(_00482_),
    .A(_04616_),
    .B(_04617_));
 sg13g2_a21oi_1 _13405_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[2] ),
    .A2(net4946),
    .Y(_04619_),
    .B1(_04618_));
 sg13g2_nor2_1 _13406_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4946),
    .Y(_04620_));
 sg13g2_nand2_1 _13407_ (.Y(_04621_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4946));
 sg13g2_nor2b_1 _13408_ (.A(_04620_),
    .B_N(_04621_),
    .Y(_04622_));
 sg13g2_xnor2_1 _13409_ (.Y(_00483_),
    .A(_04619_),
    .B(_04622_));
 sg13g2_xnor2_1 _13410_ (.Y(_04623_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[4] ),
    .B(net4977));
 sg13g2_o21ai_1 _13411_ (.B1(_04621_),
    .Y(_04624_),
    .A1(_04619_),
    .A2(_04620_));
 sg13g2_and2_1 _13412_ (.A(_04623_),
    .B(_04624_),
    .X(_04625_));
 sg13g2_xor2_1 _13413_ (.B(_04624_),
    .A(_04623_),
    .X(_00484_));
 sg13g2_xnor2_1 _13414_ (.Y(_04626_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[5] ),
    .B(net4977));
 sg13g2_a21oi_1 _13415_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[4] ),
    .A2(net4946),
    .Y(_04627_),
    .B1(_04625_));
 sg13g2_xnor2_1 _13416_ (.Y(_00485_),
    .A(_04626_),
    .B(_04627_));
 sg13g2_o21ai_1 _13417_ (.B1(net4946),
    .Y(_04628_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[4] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_and2_1 _13418_ (.A(_04625_),
    .B(_04626_),
    .X(_04629_));
 sg13g2_nor2b_1 _13419_ (.A(_04629_),
    .B_N(_04628_),
    .Y(_04630_));
 sg13g2_nand2_1 _13420_ (.Y(_04631_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4946));
 sg13g2_nor2_1 _13421_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4946),
    .Y(_04632_));
 sg13g2_xnor2_1 _13422_ (.Y(_04633_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4976));
 sg13g2_xnor2_1 _13423_ (.Y(_00486_),
    .A(_04630_),
    .B(_04633_));
 sg13g2_nand2b_1 _13424_ (.Y(_04634_),
    .B(net4976),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_xor2_1 _13425_ (.B(net4976),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[7] ),
    .X(_04635_));
 sg13g2_o21ai_1 _13426_ (.B1(_04631_),
    .Y(_04636_),
    .A1(_04630_),
    .A2(_04632_));
 sg13g2_xnor2_1 _13427_ (.Y(_00487_),
    .A(_04635_),
    .B(_04636_));
 sg13g2_xnor2_1 _13428_ (.Y(_04637_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[8] ),
    .B(net4976));
 sg13g2_o21ai_1 _13429_ (.B1(net4946),
    .Y(_04638_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_nand3_1 _13430_ (.B(_04633_),
    .C(_04634_),
    .A(_04629_),
    .Y(_04639_));
 sg13g2_and3_1 _13431_ (.X(_04640_),
    .A(_04628_),
    .B(_04638_),
    .C(_04639_));
 sg13g2_nand2b_1 _13432_ (.Y(_04641_),
    .B(_04637_),
    .A_N(_04640_));
 sg13g2_xnor2_1 _13433_ (.Y(_00488_),
    .A(_04637_),
    .B(_04640_));
 sg13g2_xor2_1 _13434_ (.B(net4976),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[9] ),
    .X(_04642_));
 sg13g2_o21ai_1 _13435_ (.B1(_04641_),
    .Y(_04643_),
    .A1(_02380_),
    .A2(net4976));
 sg13g2_xnor2_1 _13436_ (.Y(_00489_),
    .A(_04642_),
    .B(_04643_));
 sg13g2_o21ai_1 _13437_ (.B1(net4947),
    .Y(_04644_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[8] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_or2_1 _13438_ (.X(_04645_),
    .B(_04642_),
    .A(_04641_));
 sg13g2_xnor2_1 _13439_ (.Y(_04646_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4978));
 sg13g2_inv_1 _13440_ (.Y(_04647_),
    .A(_04646_));
 sg13g2_a21oi_1 _13441_ (.A1(_04644_),
    .A2(_04645_),
    .Y(_04648_),
    .B1(_04647_));
 sg13g2_nand3_1 _13442_ (.B(_04645_),
    .C(_04647_),
    .A(_04644_),
    .Y(_04649_));
 sg13g2_nor2b_1 _13443_ (.A(_04648_),
    .B_N(_04649_),
    .Y(_00472_));
 sg13g2_xor2_1 _13444_ (.B(net4978),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[11] ),
    .X(_04650_));
 sg13g2_a21oi_1 _13445_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[10] ),
    .A2(net4947),
    .Y(_04651_),
    .B1(_04648_));
 sg13g2_xor2_1 _13446_ (.B(_04651_),
    .A(_04650_),
    .X(_00473_));
 sg13g2_xnor2_1 _13447_ (.Y(_04652_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[12] ),
    .B(net4978));
 sg13g2_xor2_1 _13448_ (.B(net4978),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[12] ),
    .X(_04653_));
 sg13g2_nor3_2 _13449_ (.A(_04645_),
    .B(_04647_),
    .C(_04650_),
    .Y(_04654_));
 sg13g2_o21ai_1 _13450_ (.B1(net4947),
    .Y(_04655_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[10] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_nand2_1 _13451_ (.Y(_04656_),
    .A(_04644_),
    .B(_04655_));
 sg13g2_inv_1 _13452_ (.Y(_04657_),
    .A(_04656_));
 sg13g2_o21ai_1 _13453_ (.B1(_04652_),
    .Y(_04658_),
    .A1(_04654_),
    .A2(_04656_));
 sg13g2_or3_1 _13454_ (.A(_04652_),
    .B(_04654_),
    .C(_04656_),
    .X(_04659_));
 sg13g2_and2_1 _13455_ (.A(_04658_),
    .B(_04659_),
    .X(_00474_));
 sg13g2_xor2_1 _13456_ (.B(net4978),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[13] ),
    .X(_04660_));
 sg13g2_o21ai_1 _13457_ (.B1(_04658_),
    .Y(_04661_),
    .A1(_02381_),
    .A2(net4978));
 sg13g2_xnor2_1 _13458_ (.Y(_00475_),
    .A(_04660_),
    .B(_04661_));
 sg13g2_nor2b_1 _13459_ (.A(net4979),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[14] ),
    .Y(_04662_));
 sg13g2_xnor2_1 _13460_ (.Y(_04663_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[14] ),
    .B(net4979));
 sg13g2_o21ai_1 _13461_ (.B1(net4947),
    .Y(_04664_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[12] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_a22oi_1 _13462_ (.Y(_04665_),
    .B1(_04658_),
    .B2(_04664_),
    .A2(net4978),
    .A1(_02382_));
 sg13g2_xor2_1 _13463_ (.B(_04665_),
    .A(_04663_),
    .X(_00476_));
 sg13g2_xnor2_1 _13464_ (.Y(_04666_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[15] ),
    .B(net4978));
 sg13g2_a21oi_1 _13465_ (.A1(_04663_),
    .A2(_04665_),
    .Y(_04667_),
    .B1(_04662_));
 sg13g2_xnor2_1 _13466_ (.Y(_00477_),
    .A(_04666_),
    .B(_04667_));
 sg13g2_nor2_1 _13467_ (.A(_04653_),
    .B(_04660_),
    .Y(_04668_));
 sg13g2_nand4_1 _13468_ (.B(_04663_),
    .C(_04666_),
    .A(_04654_),
    .Y(_04669_),
    .D(_04668_));
 sg13g2_o21ai_1 _13469_ (.B1(net4947),
    .Y(_04670_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand4_1 _13470_ (.B(_04664_),
    .C(_04669_),
    .A(_04657_),
    .Y(_04671_),
    .D(_04670_));
 sg13g2_nor2b_1 _13471_ (.A(net4979),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[16] ),
    .Y(_04672_));
 sg13g2_xnor2_1 _13472_ (.Y(_04673_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[16] ),
    .B(net4979));
 sg13g2_xor2_1 _13473_ (.B(_04673_),
    .A(_04671_),
    .X(_00478_));
 sg13g2_a21o_1 _13474_ (.A2(_04673_),
    .A1(_04671_),
    .B1(_04672_),
    .X(_04674_));
 sg13g2_xor2_1 _13475_ (.B(net4979),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[17] ),
    .X(_04675_));
 sg13g2_xnor2_1 _13476_ (.Y(_00479_),
    .A(_04674_),
    .B(_04675_));
 sg13g2_nor3_1 _13477_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[17] ),
    .B(net4979),
    .C(_04674_),
    .Y(_04676_));
 sg13g2_nand3_1 _13478_ (.B(net4979),
    .C(_04674_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[17] ),
    .Y(_04677_));
 sg13g2_nor2b_1 _13479_ (.A(_04676_),
    .B_N(_04677_),
    .Y(_04678_));
 sg13g2_xnor2_1 _13480_ (.Y(_00480_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[18] ),
    .B(_04678_));
 sg13g2_nor2b_1 _13481_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][1] ),
    .Y(_04679_));
 sg13g2_xnor2_1 _13482_ (.Y(_04680_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][1] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _13483_ (.B(_04680_),
    .A(_02508_),
    .X(_00463_));
 sg13g2_a21oi_1 _13484_ (.A1(_02508_),
    .A2(_04680_),
    .Y(_04681_),
    .B1(_04679_));
 sg13g2_xnor2_1 _13485_ (.Y(_04682_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][2] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _13486_ (.A(_04681_),
    .B_N(_04682_),
    .Y(_04683_));
 sg13g2_xnor2_1 _13487_ (.Y(_00464_),
    .A(_04681_),
    .B(_04682_));
 sg13g2_a21oi_1 _13488_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][2] ),
    .A2(_02384_),
    .Y(_04684_),
    .B1(_04683_));
 sg13g2_xnor2_1 _13489_ (.Y(_04685_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][3] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _13490_ (.A(_04684_),
    .B_N(_04685_),
    .Y(_04686_));
 sg13g2_xnor2_1 _13491_ (.Y(_00465_),
    .A(_04684_),
    .B(_04685_));
 sg13g2_a21oi_1 _13492_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][3] ),
    .A2(_02385_),
    .Y(_04687_),
    .B1(_04686_));
 sg13g2_xnor2_1 _13493_ (.Y(_04688_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][4] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _13494_ (.A(_04687_),
    .B_N(_04688_),
    .Y(_04689_));
 sg13g2_xnor2_1 _13495_ (.Y(_00466_),
    .A(_04687_),
    .B(_04688_));
 sg13g2_a21oi_1 _13496_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][4] ),
    .A2(_02386_),
    .Y(_04690_),
    .B1(_04689_));
 sg13g2_nand2b_1 _13497_ (.Y(_04691_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][5] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _13498_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][5] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[5] ),
    .Y(_04692_));
 sg13g2_xnor2_1 _13499_ (.Y(_04693_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][5] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_xnor2_1 _13500_ (.Y(_00467_),
    .A(_04690_),
    .B(_04693_));
 sg13g2_nor2b_1 _13501_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][6] ),
    .Y(_04694_));
 sg13g2_nand2b_1 _13502_ (.Y(_04695_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][6] ));
 sg13g2_nand2b_1 _13503_ (.Y(_04696_),
    .B(_04695_),
    .A_N(_04694_));
 sg13g2_o21ai_1 _13504_ (.B1(_04691_),
    .Y(_04697_),
    .A1(_04690_),
    .A2(_04692_));
 sg13g2_xnor2_1 _13505_ (.Y(_00468_),
    .A(_04696_),
    .B(_04697_));
 sg13g2_a21oi_1 _13506_ (.A1(_04695_),
    .A2(_04697_),
    .Y(_04698_),
    .B1(_04694_));
 sg13g2_xnor2_1 _13507_ (.Y(_04699_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][7] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nand2b_1 _13508_ (.Y(_04700_),
    .B(_04699_),
    .A_N(_04698_));
 sg13g2_xnor2_1 _13509_ (.Y(_00469_),
    .A(_04698_),
    .B(_04699_));
 sg13g2_o21ai_1 _13510_ (.B1(_04700_),
    .Y(_04701_),
    .A1(_02387_),
    .A2(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _13511_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][8] ),
    .Y(_04702_));
 sg13g2_nand2b_1 _13512_ (.Y(_04703_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][8] ));
 sg13g2_nand2b_1 _13513_ (.Y(_04704_),
    .B(_04703_),
    .A_N(_04702_));
 sg13g2_xnor2_1 _13514_ (.Y(_00470_),
    .A(_04701_),
    .B(_04704_));
 sg13g2_nand2b_1 _13515_ (.Y(_04705_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][9] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _13516_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][9] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[9] ),
    .Y(_04706_));
 sg13g2_xnor2_1 _13517_ (.Y(_04707_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][9] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_a21oi_1 _13518_ (.A1(_04701_),
    .A2(_04703_),
    .Y(_04708_),
    .B1(_04702_));
 sg13g2_xnor2_1 _13519_ (.Y(_00471_),
    .A(_04707_),
    .B(_04708_));
 sg13g2_nor2b_1 _13520_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][10] ),
    .Y(_04709_));
 sg13g2_nand2b_1 _13521_ (.Y(_04710_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][10] ));
 sg13g2_nand2b_1 _13522_ (.Y(_04711_),
    .B(_04710_),
    .A_N(_04709_));
 sg13g2_o21ai_1 _13523_ (.B1(_04705_),
    .Y(_04712_),
    .A1(_04706_),
    .A2(_04708_));
 sg13g2_xnor2_1 _13524_ (.Y(_00454_),
    .A(_04711_),
    .B(_04712_));
 sg13g2_a21oi_1 _13525_ (.A1(_04710_),
    .A2(_04712_),
    .Y(_04713_),
    .B1(_04709_));
 sg13g2_nand2b_1 _13526_ (.Y(_04714_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][11] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _13527_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][11] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[11] ),
    .Y(_04715_));
 sg13g2_xnor2_1 _13528_ (.Y(_04716_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][11] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_xnor2_1 _13529_ (.Y(_00455_),
    .A(_04713_),
    .B(_04716_));
 sg13g2_nor2b_1 _13530_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][12] ),
    .Y(_04717_));
 sg13g2_nand2b_1 _13531_ (.Y(_04718_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][12] ));
 sg13g2_nand2b_1 _13532_ (.Y(_04719_),
    .B(_04718_),
    .A_N(_04717_));
 sg13g2_o21ai_1 _13533_ (.B1(_04714_),
    .Y(_04720_),
    .A1(_04713_),
    .A2(_04715_));
 sg13g2_xnor2_1 _13534_ (.Y(_00456_),
    .A(_04719_),
    .B(_04720_));
 sg13g2_a21oi_1 _13535_ (.A1(_04718_),
    .A2(_04720_),
    .Y(_04721_),
    .B1(_04717_));
 sg13g2_nor2b_1 _13536_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][13] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[13] ),
    .Y(_04722_));
 sg13g2_nand2b_1 _13537_ (.Y(_04723_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][13] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _13538_ (.A(_04722_),
    .B_N(_04723_),
    .Y(_04724_));
 sg13g2_xnor2_1 _13539_ (.Y(_00457_),
    .A(_04721_),
    .B(_04724_));
 sg13g2_nor2b_1 _13540_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][14] ),
    .Y(_04725_));
 sg13g2_nand2b_1 _13541_ (.Y(_04726_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][14] ));
 sg13g2_nand2b_1 _13542_ (.Y(_04727_),
    .B(_04726_),
    .A_N(_04725_));
 sg13g2_a21oi_1 _13543_ (.A1(_04721_),
    .A2(_04723_),
    .Y(_04728_),
    .B1(_04722_));
 sg13g2_xnor2_1 _13544_ (.Y(_00458_),
    .A(_04727_),
    .B(_04728_));
 sg13g2_a21oi_1 _13545_ (.A1(_04726_),
    .A2(_04728_),
    .Y(_04729_),
    .B1(_04725_));
 sg13g2_nor2b_1 _13546_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][15] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[15] ),
    .Y(_04730_));
 sg13g2_nand2b_1 _13547_ (.Y(_04731_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][15] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _13548_ (.A(_04730_),
    .B_N(_04731_),
    .Y(_04732_));
 sg13g2_xnor2_1 _13549_ (.Y(_00459_),
    .A(_04729_),
    .B(_04732_));
 sg13g2_xor2_1 _13550_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][16] ),
    .X(_04733_));
 sg13g2_a21oi_1 _13551_ (.A1(_04729_),
    .A2(_04731_),
    .Y(_04734_),
    .B1(_04730_));
 sg13g2_nor2b_1 _13552_ (.A(_04733_),
    .B_N(_04734_),
    .Y(_04735_));
 sg13g2_xnor2_1 _13553_ (.Y(_00460_),
    .A(_04733_),
    .B(_04734_));
 sg13g2_a21oi_1 _13554_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][16] ),
    .A2(_02388_),
    .Y(_04736_),
    .B1(_04735_));
 sg13g2_nand2b_1 _13555_ (.Y(_04737_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][17] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _13556_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][17] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[17] ),
    .Y(_04738_));
 sg13g2_xnor2_1 _13557_ (.Y(_04739_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][17] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _13558_ (.Y(_00461_),
    .A(_04736_),
    .B(_04739_));
 sg13g2_o21ai_1 _13559_ (.B1(_04737_),
    .Y(_04740_),
    .A1(_04736_),
    .A2(_04738_));
 sg13g2_xor2_1 _13560_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][18] ),
    .X(_04741_));
 sg13g2_xnor2_1 _13561_ (.Y(_00462_),
    .A(_04740_),
    .B(_04741_));
 sg13g2_nand2_1 _13562_ (.Y(_04742_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[0] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_nand2_1 _13563_ (.Y(_04743_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_nor2_1 _13564_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[1] ),
    .Y(_04744_));
 sg13g2_xor2_1 _13565_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[1] ),
    .X(_04745_));
 sg13g2_xnor2_1 _13566_ (.Y(_01064_),
    .A(_04742_),
    .B(_04745_));
 sg13g2_o21ai_1 _13567_ (.B1(_04743_),
    .Y(_04746_),
    .A1(_04742_),
    .A2(_04744_));
 sg13g2_xnor2_1 _13568_ (.Y(_04747_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[2] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_nor2b_1 _13569_ (.A(_04747_),
    .B_N(_04746_),
    .Y(_04748_));
 sg13g2_xnor2_1 _13570_ (.Y(_01065_),
    .A(_04746_),
    .B(_04747_));
 sg13g2_a21o_1 _13571_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[2] ),
    .B1(_04748_),
    .X(_04749_));
 sg13g2_xnor2_1 _13572_ (.Y(_04750_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[3] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_nor2b_1 _13573_ (.A(_04750_),
    .B_N(_04749_),
    .Y(_04751_));
 sg13g2_xnor2_1 _13574_ (.Y(_01066_),
    .A(_04749_),
    .B(_04750_));
 sg13g2_a21o_1 _13575_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[3] ),
    .B1(_04751_),
    .X(_04752_));
 sg13g2_xnor2_1 _13576_ (.Y(_04753_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[4] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_nor2b_1 _13577_ (.A(_04753_),
    .B_N(_04752_),
    .Y(_04754_));
 sg13g2_xnor2_1 _13578_ (.Y(_01067_),
    .A(_04752_),
    .B(_04753_));
 sg13g2_a21o_1 _13579_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[4] ),
    .B1(_04754_),
    .X(_04755_));
 sg13g2_nand2_1 _13580_ (.Y(_04756_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _13581_ (.Y(_04757_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _13582_ (.Y(_01068_),
    .A(_04755_),
    .B(_04757_));
 sg13g2_xnor2_1 _13583_ (.Y(_04758_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[6] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_o21ai_1 _13584_ (.B1(_04755_),
    .Y(_04759_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_a21oi_1 _13585_ (.A1(_04756_),
    .A2(_04759_),
    .Y(_04760_),
    .B1(_04758_));
 sg13g2_nand3_1 _13586_ (.B(_04758_),
    .C(_04759_),
    .A(_04756_),
    .Y(_04761_));
 sg13g2_nor2b_1 _13587_ (.A(_04760_),
    .B_N(_04761_),
    .Y(_01069_));
 sg13g2_a21oi_1 _13588_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[6] ),
    .Y(_04762_),
    .B1(_04760_));
 sg13g2_nand2_1 _13589_ (.Y(_04763_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_nor2_1 _13590_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[7] ),
    .Y(_04764_));
 sg13g2_xor2_1 _13591_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[7] ),
    .X(_04765_));
 sg13g2_xnor2_1 _13592_ (.Y(_01070_),
    .A(_04762_),
    .B(_04765_));
 sg13g2_o21ai_1 _13593_ (.B1(_04763_),
    .Y(_04766_),
    .A1(_04762_),
    .A2(_04764_));
 sg13g2_xnor2_1 _13594_ (.Y(_04767_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[8] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_nor2b_1 _13595_ (.A(_04767_),
    .B_N(_04766_),
    .Y(_04768_));
 sg13g2_xnor2_1 _13596_ (.Y(_01071_),
    .A(_04766_),
    .B(_04767_));
 sg13g2_a21o_1 _13597_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[8] ),
    .B1(_04768_),
    .X(_04769_));
 sg13g2_xnor2_1 _13598_ (.Y(_04770_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[9] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _13599_ (.Y(_01072_),
    .A(_04769_),
    .B(_04770_));
 sg13g2_nand2_1 _13600_ (.Y(_04771_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_nor2_1 _13601_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[10] ),
    .Y(_04772_));
 sg13g2_xor2_1 _13602_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[10] ),
    .X(_04773_));
 sg13g2_a21o_1 _13603_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[9] ),
    .B1(_04769_),
    .X(_04774_));
 sg13g2_o21ai_1 _13604_ (.B1(_04774_),
    .Y(_04775_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _13605_ (.Y(_01055_),
    .A(_04773_),
    .B(_04775_));
 sg13g2_o21ai_1 _13606_ (.B1(_04771_),
    .Y(_04776_),
    .A1(_04772_),
    .A2(_04775_));
 sg13g2_xnor2_1 _13607_ (.Y(_04777_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[11] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _13608_ (.Y(_01056_),
    .A(_04776_),
    .B(_04777_));
 sg13g2_nand2_1 _13609_ (.Y(_04778_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[12] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_nor2_1 _13610_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[12] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[12] ),
    .Y(_04779_));
 sg13g2_xor2_1 _13611_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[12] ),
    .X(_04780_));
 sg13g2_a21o_1 _13612_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[11] ),
    .B1(_04776_),
    .X(_04781_));
 sg13g2_o21ai_1 _13613_ (.B1(_04781_),
    .Y(_04782_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _13614_ (.Y(_01057_),
    .A(_04780_),
    .B(_04782_));
 sg13g2_o21ai_1 _13615_ (.B1(_04778_),
    .Y(_04783_),
    .A1(_04779_),
    .A2(_04782_));
 sg13g2_xnor2_1 _13616_ (.Y(_04784_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[13] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_xnor2_1 _13617_ (.Y(_01058_),
    .A(_04783_),
    .B(_04784_));
 sg13g2_xnor2_1 _13618_ (.Y(_04785_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[14] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_a21o_1 _13619_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[13] ),
    .B1(_04783_),
    .X(_04786_));
 sg13g2_o21ai_1 _13620_ (.B1(_04786_),
    .Y(_04787_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_nor2_1 _13621_ (.A(_04785_),
    .B(_04787_),
    .Y(_04788_));
 sg13g2_xor2_1 _13622_ (.B(_04787_),
    .A(_04785_),
    .X(_01059_));
 sg13g2_a21oi_1 _13623_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[14] ),
    .Y(_04789_),
    .B1(_04788_));
 sg13g2_nor2_1 _13624_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[15] ),
    .Y(_04790_));
 sg13g2_nand2_1 _13625_ (.Y(_04791_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_nor2b_1 _13626_ (.A(_04790_),
    .B_N(_04791_),
    .Y(_04792_));
 sg13g2_xnor2_1 _13627_ (.Y(_01060_),
    .A(_04789_),
    .B(_04792_));
 sg13g2_and2_1 _13628_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[16] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[16] ),
    .X(_04793_));
 sg13g2_xor2_1 _13629_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[16] ),
    .X(_04794_));
 sg13g2_a21oi_1 _13630_ (.A1(_04789_),
    .A2(_04791_),
    .Y(_04795_),
    .B1(_04790_));
 sg13g2_xor2_1 _13631_ (.B(_04795_),
    .A(_04794_),
    .X(_01061_));
 sg13g2_a21o_1 _13632_ (.A2(_04795_),
    .A1(_04794_),
    .B1(_04793_),
    .X(_04796_));
 sg13g2_xnor2_1 _13633_ (.Y(_04797_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[17] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xnor2_1 _13634_ (.Y(_01062_),
    .A(_04796_),
    .B(_04797_));
 sg13g2_a21o_1 _13635_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[17] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[17] ),
    .B1(_04796_),
    .X(_04798_));
 sg13g2_o21ai_1 _13636_ (.B1(_04798_),
    .Y(_04799_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xor2_1 _13637_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[18] ),
    .X(_04800_));
 sg13g2_xnor2_1 _13638_ (.Y(_01063_),
    .A(_04799_),
    .B(_04800_));
 sg13g2_xor2_1 _13639_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[0] ),
    .X(_01054_));
 sg13g2_nand2_1 _13640_ (.Y(_04801_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[0] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_xor2_1 _13641_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[0] ),
    .X(_00603_));
 sg13g2_nand2_1 _13642_ (.Y(_04802_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_nor2_1 _13643_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[1] ),
    .Y(_04803_));
 sg13g2_xor2_1 _13644_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[1] ),
    .X(_04804_));
 sg13g2_xnor2_1 _13645_ (.Y(_00613_),
    .A(_04801_),
    .B(_04804_));
 sg13g2_o21ai_1 _13646_ (.B1(_04802_),
    .Y(_04805_),
    .A1(_04801_),
    .A2(_04803_));
 sg13g2_xnor2_1 _13647_ (.Y(_04806_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[2] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_nor2b_1 _13648_ (.A(_04806_),
    .B_N(_04805_),
    .Y(_04807_));
 sg13g2_xnor2_1 _13649_ (.Y(_00614_),
    .A(_04805_),
    .B(_04806_));
 sg13g2_a21o_1 _13650_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[2] ),
    .B1(_04807_),
    .X(_04808_));
 sg13g2_xnor2_1 _13651_ (.Y(_04809_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[3] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_nor2b_1 _13652_ (.A(_04809_),
    .B_N(_04808_),
    .Y(_04810_));
 sg13g2_xnor2_1 _13653_ (.Y(_00615_),
    .A(_04808_),
    .B(_04809_));
 sg13g2_a21o_1 _13654_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[3] ),
    .B1(_04810_),
    .X(_04811_));
 sg13g2_xnor2_1 _13655_ (.Y(_04812_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[4] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_nor2b_1 _13656_ (.A(_04812_),
    .B_N(_04811_),
    .Y(_04813_));
 sg13g2_xnor2_1 _13657_ (.Y(_00616_),
    .A(_04811_),
    .B(_04812_));
 sg13g2_a21o_1 _13658_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[4] ),
    .B1(_04813_),
    .X(_04814_));
 sg13g2_nand2_1 _13659_ (.Y(_04815_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[5] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_xnor2_1 _13660_ (.Y(_04816_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[5] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_xnor2_1 _13661_ (.Y(_00617_),
    .A(_04814_),
    .B(_04816_));
 sg13g2_xnor2_1 _13662_ (.Y(_04817_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[6] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_o21ai_1 _13663_ (.B1(_04814_),
    .Y(_04818_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_a21oi_1 _13664_ (.A1(_04815_),
    .A2(_04818_),
    .Y(_04819_),
    .B1(_04817_));
 sg13g2_nand3_1 _13665_ (.B(_04817_),
    .C(_04818_),
    .A(_04815_),
    .Y(_04820_));
 sg13g2_nor2b_1 _13666_ (.A(_04819_),
    .B_N(_04820_),
    .Y(_00618_));
 sg13g2_a21oi_1 _13667_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[6] ),
    .Y(_04821_),
    .B1(_04819_));
 sg13g2_nand2_1 _13668_ (.Y(_04822_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[7] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_nor2_1 _13669_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[7] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[7] ),
    .Y(_04823_));
 sg13g2_xor2_1 _13670_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[7] ),
    .X(_04824_));
 sg13g2_xnor2_1 _13671_ (.Y(_00619_),
    .A(_04821_),
    .B(_04824_));
 sg13g2_o21ai_1 _13672_ (.B1(_04822_),
    .Y(_04825_),
    .A1(_04821_),
    .A2(_04823_));
 sg13g2_xnor2_1 _13673_ (.Y(_04826_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[8] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_nor2b_1 _13674_ (.A(_04826_),
    .B_N(_04825_),
    .Y(_04827_));
 sg13g2_xnor2_1 _13675_ (.Y(_00620_),
    .A(_04825_),
    .B(_04826_));
 sg13g2_xnor2_1 _13676_ (.Y(_04828_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[9] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_a21o_1 _13677_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[8] ),
    .B1(_04827_),
    .X(_04829_));
 sg13g2_xnor2_1 _13678_ (.Y(_00621_),
    .A(_04828_),
    .B(_04829_));
 sg13g2_nand2_1 _13679_ (.Y(_04830_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[10] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_nor2_1 _13680_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[10] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[10] ),
    .Y(_04831_));
 sg13g2_xor2_1 _13681_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[10] ),
    .X(_04832_));
 sg13g2_a21o_1 _13682_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[9] ),
    .B1(_04829_),
    .X(_04833_));
 sg13g2_o21ai_1 _13683_ (.B1(_04833_),
    .Y(_04834_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_xnor2_1 _13684_ (.Y(_00604_),
    .A(_04832_),
    .B(_04834_));
 sg13g2_xnor2_1 _13685_ (.Y(_04835_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[11] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_o21ai_1 _13686_ (.B1(_04830_),
    .Y(_04836_),
    .A1(_04831_),
    .A2(_04834_));
 sg13g2_xnor2_1 _13687_ (.Y(_00605_),
    .A(_04835_),
    .B(_04836_));
 sg13g2_nand2_1 _13688_ (.Y(_04837_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[12] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_nor2_1 _13689_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[12] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[12] ),
    .Y(_04838_));
 sg13g2_xor2_1 _13690_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[12] ),
    .X(_04839_));
 sg13g2_a21o_1 _13691_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[11] ),
    .B1(_04836_),
    .X(_04840_));
 sg13g2_o21ai_1 _13692_ (.B1(_04840_),
    .Y(_04841_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_xnor2_1 _13693_ (.Y(_00606_),
    .A(_04839_),
    .B(_04841_));
 sg13g2_xnor2_1 _13694_ (.Y(_04842_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[13] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_o21ai_1 _13695_ (.B1(_04837_),
    .Y(_04843_),
    .A1(_04838_),
    .A2(_04841_));
 sg13g2_xnor2_1 _13696_ (.Y(_00607_),
    .A(_04842_),
    .B(_04843_));
 sg13g2_xnor2_1 _13697_ (.Y(_04844_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[14] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_a21o_1 _13698_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[13] ),
    .B1(_04843_),
    .X(_04845_));
 sg13g2_o21ai_1 _13699_ (.B1(_04845_),
    .Y(_04846_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_nor2_1 _13700_ (.A(_04844_),
    .B(_04846_),
    .Y(_04847_));
 sg13g2_xor2_1 _13701_ (.B(_04846_),
    .A(_04844_),
    .X(_00608_));
 sg13g2_nor2_1 _13702_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[15] ),
    .Y(_04848_));
 sg13g2_nand2_1 _13703_ (.Y(_04849_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_nor2b_1 _13704_ (.A(_04848_),
    .B_N(_04849_),
    .Y(_04850_));
 sg13g2_a21oi_1 _13705_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[14] ),
    .Y(_04851_),
    .B1(_04847_));
 sg13g2_xnor2_1 _13706_ (.Y(_00609_),
    .A(_04850_),
    .B(_04851_));
 sg13g2_nand2_1 _13707_ (.Y(_04852_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[16] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_xor2_1 _13708_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[16] ),
    .X(_04853_));
 sg13g2_o21ai_1 _13709_ (.B1(_04849_),
    .Y(_04854_),
    .A1(_04848_),
    .A2(_04851_));
 sg13g2_nand2_1 _13710_ (.Y(_04855_),
    .A(_04853_),
    .B(_04854_));
 sg13g2_xor2_1 _13711_ (.B(_04854_),
    .A(_04853_),
    .X(_00610_));
 sg13g2_xnor2_1 _13712_ (.Y(_04856_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[17] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_a21oi_1 _13713_ (.A1(_04852_),
    .A2(_04855_),
    .Y(_04857_),
    .B1(_04856_));
 sg13g2_nand3_1 _13714_ (.B(_04855_),
    .C(_04856_),
    .A(_04852_),
    .Y(_04858_));
 sg13g2_nor2b_1 _13715_ (.A(_04857_),
    .B_N(_04858_),
    .Y(_00611_));
 sg13g2_a21oi_1 _13716_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[17] ),
    .Y(_04859_),
    .B1(_04857_));
 sg13g2_xor2_1 _13717_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[18] ),
    .X(_04860_));
 sg13g2_xnor2_1 _13718_ (.Y(_00612_),
    .A(_04859_),
    .B(_04860_));
 sg13g2_nor2b_1 _13719_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][1] ),
    .Y(_04861_));
 sg13g2_xnor2_1 _13720_ (.Y(_04862_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][1] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _13721_ (.B(_04862_),
    .A(_02509_),
    .X(_00632_));
 sg13g2_a21oi_1 _13722_ (.A1(_02509_),
    .A2(_04862_),
    .Y(_04863_),
    .B1(_04861_));
 sg13g2_xnor2_1 _13723_ (.Y(_04864_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][2] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _13724_ (.A(_04863_),
    .B_N(_04864_),
    .Y(_04865_));
 sg13g2_xnor2_1 _13725_ (.Y(_00633_),
    .A(_04863_),
    .B(_04864_));
 sg13g2_a21oi_1 _13726_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][2] ),
    .A2(_02392_),
    .Y(_04866_),
    .B1(_04865_));
 sg13g2_xnor2_1 _13727_ (.Y(_04867_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][3] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _13728_ (.A(_04866_),
    .B_N(_04867_),
    .Y(_04868_));
 sg13g2_xnor2_1 _13729_ (.Y(_00634_),
    .A(_04866_),
    .B(_04867_));
 sg13g2_a21oi_1 _13730_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][3] ),
    .A2(_02393_),
    .Y(_04869_),
    .B1(_04868_));
 sg13g2_xnor2_1 _13731_ (.Y(_04870_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][4] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _13732_ (.A(_04869_),
    .B_N(_04870_),
    .Y(_04871_));
 sg13g2_xnor2_1 _13733_ (.Y(_00635_),
    .A(_04869_),
    .B(_04870_));
 sg13g2_a21oi_1 _13734_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][4] ),
    .A2(_02394_),
    .Y(_04872_),
    .B1(_04871_));
 sg13g2_xnor2_1 _13735_ (.Y(_04873_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][5] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _13736_ (.A(_04872_),
    .B_N(_04873_),
    .Y(_04874_));
 sg13g2_xnor2_1 _13737_ (.Y(_00636_),
    .A(_04872_),
    .B(_04873_));
 sg13g2_a21oi_1 _13738_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][5] ),
    .A2(_02395_),
    .Y(_04875_),
    .B1(_04874_));
 sg13g2_xnor2_1 _13739_ (.Y(_04876_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][6] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_nor2b_1 _13740_ (.A(_04875_),
    .B_N(_04876_),
    .Y(_04877_));
 sg13g2_xnor2_1 _13741_ (.Y(_00637_),
    .A(_04875_),
    .B(_04876_));
 sg13g2_a21oi_2 _13742_ (.B1(_04877_),
    .Y(_04878_),
    .A2(_02396_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][6] ));
 sg13g2_xnor2_1 _13743_ (.Y(_04879_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][7] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _13744_ (.A(_04878_),
    .B_N(_04879_),
    .Y(_04880_));
 sg13g2_xnor2_1 _13745_ (.Y(_00638_),
    .A(_04878_),
    .B(_04879_));
 sg13g2_a21oi_2 _13746_ (.B1(_04880_),
    .Y(_04881_),
    .A2(_02397_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][7] ));
 sg13g2_xnor2_1 _13747_ (.Y(_04882_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][8] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_nor2b_1 _13748_ (.A(_04881_),
    .B_N(_04882_),
    .Y(_04883_));
 sg13g2_xnor2_1 _13749_ (.Y(_00639_),
    .A(_04881_),
    .B(_04882_));
 sg13g2_a21oi_2 _13750_ (.B1(_04883_),
    .Y(_04884_),
    .A2(_02398_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][8] ));
 sg13g2_nand2b_1 _13751_ (.Y(_04885_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][9] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _13752_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][9] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[9] ),
    .Y(_04886_));
 sg13g2_xnor2_1 _13753_ (.Y(_04887_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][9] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_xnor2_1 _13754_ (.Y(_00640_),
    .A(_04884_),
    .B(_04887_));
 sg13g2_nor2b_1 _13755_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][10] ),
    .Y(_04888_));
 sg13g2_nand2b_1 _13756_ (.Y(_04889_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][10] ));
 sg13g2_nand2b_1 _13757_ (.Y(_04890_),
    .B(_04889_),
    .A_N(_04888_));
 sg13g2_o21ai_1 _13758_ (.B1(_04885_),
    .Y(_04891_),
    .A1(_04884_),
    .A2(_04886_));
 sg13g2_xnor2_1 _13759_ (.Y(_00623_),
    .A(_04890_),
    .B(_04891_));
 sg13g2_a21oi_1 _13760_ (.A1(_04889_),
    .A2(_04891_),
    .Y(_04892_),
    .B1(_04888_));
 sg13g2_nand2b_1 _13761_ (.Y(_04893_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][11] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _13762_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][11] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[11] ),
    .Y(_04894_));
 sg13g2_xnor2_1 _13763_ (.Y(_04895_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][11] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_xnor2_1 _13764_ (.Y(_00624_),
    .A(_04892_),
    .B(_04895_));
 sg13g2_nor2b_1 _13765_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][12] ),
    .Y(_04896_));
 sg13g2_nand2b_1 _13766_ (.Y(_04897_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][12] ));
 sg13g2_nand2b_1 _13767_ (.Y(_04898_),
    .B(_04897_),
    .A_N(_04896_));
 sg13g2_o21ai_1 _13768_ (.B1(_04893_),
    .Y(_04899_),
    .A1(_04892_),
    .A2(_04894_));
 sg13g2_xnor2_1 _13769_ (.Y(_00625_),
    .A(_04898_),
    .B(_04899_));
 sg13g2_a21oi_2 _13770_ (.B1(_04896_),
    .Y(_04900_),
    .A2(_04899_),
    .A1(_04897_));
 sg13g2_nand2b_1 _13771_ (.Y(_04901_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][13] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _13772_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][13] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[13] ),
    .Y(_04902_));
 sg13g2_xnor2_1 _13773_ (.Y(_04903_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][13] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_xnor2_1 _13774_ (.Y(_00626_),
    .A(_04900_),
    .B(_04903_));
 sg13g2_nor2b_1 _13775_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][14] ),
    .Y(_04904_));
 sg13g2_nand2b_1 _13776_ (.Y(_04905_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][14] ));
 sg13g2_nand2b_1 _13777_ (.Y(_04906_),
    .B(_04905_),
    .A_N(_04904_));
 sg13g2_o21ai_1 _13778_ (.B1(_04901_),
    .Y(_04907_),
    .A1(_04900_),
    .A2(_04902_));
 sg13g2_xnor2_1 _13779_ (.Y(_00627_),
    .A(_04906_),
    .B(_04907_));
 sg13g2_a21oi_2 _13780_ (.B1(_04904_),
    .Y(_04908_),
    .A2(_04907_),
    .A1(_04905_));
 sg13g2_nand2b_1 _13781_ (.Y(_04909_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][15] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _13782_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][15] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[15] ),
    .Y(_04910_));
 sg13g2_xnor2_1 _13783_ (.Y(_04911_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][15] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_xnor2_1 _13784_ (.Y(_00628_),
    .A(_04908_),
    .B(_04911_));
 sg13g2_xor2_1 _13785_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][16] ),
    .X(_04912_));
 sg13g2_o21ai_1 _13786_ (.B1(_04909_),
    .Y(_04913_),
    .A1(_04908_),
    .A2(_04910_));
 sg13g2_nor2b_1 _13787_ (.A(_04912_),
    .B_N(_04913_),
    .Y(_04914_));
 sg13g2_xnor2_1 _13788_ (.Y(_00629_),
    .A(_04912_),
    .B(_04913_));
 sg13g2_a21oi_1 _13789_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][16] ),
    .A2(_02399_),
    .Y(_04915_),
    .B1(_04914_));
 sg13g2_nand2b_1 _13790_ (.Y(_04916_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][17] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _13791_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][17] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[17] ),
    .Y(_04917_));
 sg13g2_xnor2_1 _13792_ (.Y(_04918_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][17] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _13793_ (.Y(_00630_),
    .A(_04915_),
    .B(_04918_));
 sg13g2_o21ai_1 _13794_ (.B1(_04916_),
    .Y(_04919_),
    .A1(_04915_),
    .A2(_04917_));
 sg13g2_xor2_1 _13795_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][18] ),
    .X(_04920_));
 sg13g2_xnor2_1 _13796_ (.Y(_00631_),
    .A(_04919_),
    .B(_04920_));
 sg13g2_nand2_1 _13797_ (.Y(_04921_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[0] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_xor2_1 _13798_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[0] ),
    .X(_00584_));
 sg13g2_nand2_1 _13799_ (.Y(_04922_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_nor2_1 _13800_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[1] ),
    .Y(_04923_));
 sg13g2_xor2_1 _13801_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[1] ),
    .X(_04924_));
 sg13g2_xnor2_1 _13802_ (.Y(_00594_),
    .A(_04921_),
    .B(_04924_));
 sg13g2_o21ai_1 _13803_ (.B1(_04922_),
    .Y(_04925_),
    .A1(_04921_),
    .A2(_04923_));
 sg13g2_xnor2_1 _13804_ (.Y(_04926_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[2] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_nor2b_1 _13805_ (.A(_04926_),
    .B_N(_04925_),
    .Y(_04927_));
 sg13g2_xnor2_1 _13806_ (.Y(_00595_),
    .A(_04925_),
    .B(_04926_));
 sg13g2_a21o_1 _13807_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[2] ),
    .B1(_04927_),
    .X(_04928_));
 sg13g2_xnor2_1 _13808_ (.Y(_04929_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[3] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_nor2b_1 _13809_ (.A(_04929_),
    .B_N(_04928_),
    .Y(_04930_));
 sg13g2_xnor2_1 _13810_ (.Y(_00596_),
    .A(_04928_),
    .B(_04929_));
 sg13g2_a21o_1 _13811_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[3] ),
    .B1(_04930_),
    .X(_04931_));
 sg13g2_xnor2_1 _13812_ (.Y(_04932_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[4] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_nor2b_1 _13813_ (.A(_04932_),
    .B_N(_04931_),
    .Y(_04933_));
 sg13g2_xnor2_1 _13814_ (.Y(_00597_),
    .A(_04931_),
    .B(_04932_));
 sg13g2_a21o_1 _13815_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[4] ),
    .B1(_04933_),
    .X(_04934_));
 sg13g2_nand2_1 _13816_ (.Y(_04935_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _13817_ (.Y(_04936_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _13818_ (.Y(_00598_),
    .A(_04934_),
    .B(_04936_));
 sg13g2_xnor2_1 _13819_ (.Y(_04937_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[6] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_o21ai_1 _13820_ (.B1(_04934_),
    .Y(_04938_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_a21oi_1 _13821_ (.A1(_04935_),
    .A2(_04938_),
    .Y(_04939_),
    .B1(_04937_));
 sg13g2_nand3_1 _13822_ (.B(_04937_),
    .C(_04938_),
    .A(_04935_),
    .Y(_04940_));
 sg13g2_nor2b_1 _13823_ (.A(_04939_),
    .B_N(_04940_),
    .Y(_00599_));
 sg13g2_a21oi_1 _13824_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[6] ),
    .Y(_04941_),
    .B1(_04939_));
 sg13g2_nand2_1 _13825_ (.Y(_04942_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_nor2_1 _13826_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[7] ),
    .Y(_04943_));
 sg13g2_xor2_1 _13827_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[7] ),
    .X(_04944_));
 sg13g2_xnor2_1 _13828_ (.Y(_00600_),
    .A(_04941_),
    .B(_04944_));
 sg13g2_o21ai_1 _13829_ (.B1(_04942_),
    .Y(_04945_),
    .A1(_04941_),
    .A2(_04943_));
 sg13g2_xnor2_1 _13830_ (.Y(_04946_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[8] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_nor2b_1 _13831_ (.A(_04946_),
    .B_N(_04945_),
    .Y(_04947_));
 sg13g2_xnor2_1 _13832_ (.Y(_00601_),
    .A(_04945_),
    .B(_04946_));
 sg13g2_a21o_1 _13833_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[8] ),
    .B1(_04947_),
    .X(_04948_));
 sg13g2_xnor2_1 _13834_ (.Y(_04949_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[9] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _13835_ (.Y(_00602_),
    .A(_04948_),
    .B(_04949_));
 sg13g2_nand2_1 _13836_ (.Y(_04950_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_nor2_1 _13837_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[10] ),
    .Y(_04951_));
 sg13g2_xor2_1 _13838_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[10] ),
    .X(_04952_));
 sg13g2_a21o_1 _13839_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[9] ),
    .B1(_04948_),
    .X(_04953_));
 sg13g2_o21ai_1 _13840_ (.B1(_04953_),
    .Y(_04954_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _13841_ (.Y(_00585_),
    .A(_04952_),
    .B(_04954_));
 sg13g2_o21ai_1 _13842_ (.B1(_04950_),
    .Y(_04955_),
    .A1(_04951_),
    .A2(_04954_));
 sg13g2_xnor2_1 _13843_ (.Y(_04956_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[11] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _13844_ (.Y(_00586_),
    .A(_04955_),
    .B(_04956_));
 sg13g2_xor2_1 _13845_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[12] ),
    .X(_04957_));
 sg13g2_a21o_1 _13846_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[11] ),
    .B1(_04955_),
    .X(_04958_));
 sg13g2_o21ai_1 _13847_ (.B1(_04958_),
    .Y(_04959_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_nand2b_1 _13848_ (.Y(_04960_),
    .B(_04957_),
    .A_N(_04959_));
 sg13g2_xnor2_1 _13849_ (.Y(_00587_),
    .A(_04957_),
    .B(_04959_));
 sg13g2_o21ai_1 _13850_ (.B1(_04960_),
    .Y(_04961_),
    .A1(_02401_),
    .A2(_02402_));
 sg13g2_xnor2_1 _13851_ (.Y(_04962_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[13] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_xnor2_1 _13852_ (.Y(_00588_),
    .A(_04961_),
    .B(_04962_));
 sg13g2_xnor2_1 _13853_ (.Y(_04963_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[14] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_a21o_1 _13854_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[13] ),
    .B1(_04961_),
    .X(_04964_));
 sg13g2_o21ai_1 _13855_ (.B1(_04964_),
    .Y(_04965_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_nor2_1 _13856_ (.A(_04963_),
    .B(_04965_),
    .Y(_04966_));
 sg13g2_xor2_1 _13857_ (.B(_04965_),
    .A(_04963_),
    .X(_00589_));
 sg13g2_a21oi_1 _13858_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[14] ),
    .Y(_04967_),
    .B1(_04966_));
 sg13g2_nand2_1 _13859_ (.Y(_04968_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_nor2_1 _13860_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[15] ),
    .Y(_04969_));
 sg13g2_xor2_1 _13861_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[15] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[15] ),
    .X(_04970_));
 sg13g2_xnor2_1 _13862_ (.Y(_00590_),
    .A(_04967_),
    .B(_04970_));
 sg13g2_and2_1 _13863_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[16] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[16] ),
    .X(_04971_));
 sg13g2_xor2_1 _13864_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[16] ),
    .X(_04972_));
 sg13g2_o21ai_1 _13865_ (.B1(_04968_),
    .Y(_04973_),
    .A1(_04967_),
    .A2(_04969_));
 sg13g2_xor2_1 _13866_ (.B(_04973_),
    .A(_04972_),
    .X(_00591_));
 sg13g2_a21o_1 _13867_ (.A2(_04973_),
    .A1(_04972_),
    .B1(_04971_),
    .X(_04974_));
 sg13g2_xnor2_1 _13868_ (.Y(_04975_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[17] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xnor2_1 _13869_ (.Y(_00592_),
    .A(_04974_),
    .B(_04975_));
 sg13g2_a21o_1 _13870_ (.A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[17] ),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[17] ),
    .B1(_04974_),
    .X(_04976_));
 sg13g2_o21ai_1 _13871_ (.B1(_04976_),
    .Y(_04977_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xor2_1 _13872_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[18] ),
    .X(_04978_));
 sg13g2_xnor2_1 _13873_ (.Y(_00593_),
    .A(_04977_),
    .B(_04978_));
 sg13g2_nand2b_1 _13874_ (.Y(_04979_),
    .B(net4970),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_nor2b_1 _13875_ (.A(net4970),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[1] ),
    .Y(_04980_));
 sg13g2_xnor2_1 _13876_ (.Y(_04981_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[1] ),
    .B(net4970));
 sg13g2_xnor2_1 _13877_ (.Y(_00575_),
    .A(_01192_),
    .B(_04981_));
 sg13g2_xnor2_1 _13878_ (.Y(_04982_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[2] ),
    .B(net4970));
 sg13g2_o21ai_1 _13879_ (.B1(_04979_),
    .Y(_04983_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[0] ),
    .A2(_04980_));
 sg13g2_nor2b_1 _13880_ (.A(_04983_),
    .B_N(_04982_),
    .Y(_04984_));
 sg13g2_xnor2_1 _13881_ (.Y(_00576_),
    .A(_04982_),
    .B(_04983_));
 sg13g2_a21oi_1 _13882_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[2] ),
    .A2(net4945),
    .Y(_04985_),
    .B1(_04984_));
 sg13g2_nor2_1 _13883_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4945),
    .Y(_04986_));
 sg13g2_nand2_1 _13884_ (.Y(_04987_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4945));
 sg13g2_nor2b_1 _13885_ (.A(_04986_),
    .B_N(_04987_),
    .Y(_04988_));
 sg13g2_xnor2_1 _13886_ (.Y(_00577_),
    .A(_04985_),
    .B(_04988_));
 sg13g2_xnor2_1 _13887_ (.Y(_04989_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[4] ),
    .B(net4971));
 sg13g2_o21ai_1 _13888_ (.B1(_04987_),
    .Y(_04990_),
    .A1(_04985_),
    .A2(_04986_));
 sg13g2_and2_1 _13889_ (.A(_04989_),
    .B(_04990_),
    .X(_04991_));
 sg13g2_xor2_1 _13890_ (.B(_04990_),
    .A(_04989_),
    .X(_00578_));
 sg13g2_xnor2_1 _13891_ (.Y(_04992_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[5] ),
    .B(net4971));
 sg13g2_a21oi_1 _13892_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[4] ),
    .A2(net4945),
    .Y(_04993_),
    .B1(_04991_));
 sg13g2_xnor2_1 _13893_ (.Y(_00579_),
    .A(_04992_),
    .B(_04993_));
 sg13g2_o21ai_1 _13894_ (.B1(net4945),
    .Y(_04994_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[4] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_and2_1 _13895_ (.A(_04991_),
    .B(_04992_),
    .X(_04995_));
 sg13g2_nor2b_1 _13896_ (.A(_04995_),
    .B_N(_04994_),
    .Y(_04996_));
 sg13g2_nand2_1 _13897_ (.Y(_04997_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4944));
 sg13g2_nor2_1 _13898_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4944),
    .Y(_04998_));
 sg13g2_xnor2_1 _13899_ (.Y(_04999_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4970));
 sg13g2_xnor2_1 _13900_ (.Y(_00580_),
    .A(_04996_),
    .B(_04999_));
 sg13g2_nand2b_1 _13901_ (.Y(_05000_),
    .B(net4970),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_xor2_1 _13902_ (.B(net4971),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[7] ),
    .X(_05001_));
 sg13g2_o21ai_1 _13903_ (.B1(_04997_),
    .Y(_05002_),
    .A1(_04996_),
    .A2(_04998_));
 sg13g2_xnor2_1 _13904_ (.Y(_00581_),
    .A(_05001_),
    .B(_05002_));
 sg13g2_xnor2_1 _13905_ (.Y(_05003_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[8] ),
    .B(net4970));
 sg13g2_o21ai_1 _13906_ (.B1(net4944),
    .Y(_05004_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_nand3_1 _13907_ (.B(_04999_),
    .C(_05000_),
    .A(_04995_),
    .Y(_05005_));
 sg13g2_and3_1 _13908_ (.X(_05006_),
    .A(_04994_),
    .B(_05004_),
    .C(_05005_));
 sg13g2_nand2b_1 _13909_ (.Y(_05007_),
    .B(_05003_),
    .A_N(_05006_));
 sg13g2_xnor2_1 _13910_ (.Y(_00582_),
    .A(_05003_),
    .B(_05006_));
 sg13g2_xor2_1 _13911_ (.B(net4969),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[9] ),
    .X(_05008_));
 sg13g2_o21ai_1 _13912_ (.B1(_05007_),
    .Y(_05009_),
    .A1(_02400_),
    .A2(net4969));
 sg13g2_xnor2_1 _13913_ (.Y(_00583_),
    .A(_05008_),
    .B(_05009_));
 sg13g2_o21ai_1 _13914_ (.B1(net4944),
    .Y(_05010_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[8] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_or2_1 _13915_ (.X(_05011_),
    .B(_05008_),
    .A(_05007_));
 sg13g2_xnor2_1 _13916_ (.Y(_05012_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4969));
 sg13g2_inv_1 _13917_ (.Y(_05013_),
    .A(_05012_));
 sg13g2_a21oi_1 _13918_ (.A1(_05010_),
    .A2(_05011_),
    .Y(_05014_),
    .B1(_05013_));
 sg13g2_nand3_1 _13919_ (.B(_05011_),
    .C(_05013_),
    .A(_05010_),
    .Y(_05015_));
 sg13g2_nor2b_1 _13920_ (.A(_05014_),
    .B_N(_05015_),
    .Y(_00566_));
 sg13g2_xor2_1 _13921_ (.B(net4969),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[11] ),
    .X(_05016_));
 sg13g2_a21oi_1 _13922_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[10] ),
    .A2(net4944),
    .Y(_05017_),
    .B1(_05014_));
 sg13g2_xor2_1 _13923_ (.B(_05017_),
    .A(_05016_),
    .X(_00567_));
 sg13g2_xnor2_1 _13924_ (.Y(_05018_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[12] ),
    .B(net4967));
 sg13g2_xor2_1 _13925_ (.B(net4967),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[12] ),
    .X(_05019_));
 sg13g2_nor3_2 _13926_ (.A(_05011_),
    .B(_05013_),
    .C(_05016_),
    .Y(_05020_));
 sg13g2_o21ai_1 _13927_ (.B1(net4944),
    .Y(_05021_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[10] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_nand2_1 _13928_ (.Y(_05022_),
    .A(_05010_),
    .B(_05021_));
 sg13g2_inv_1 _13929_ (.Y(_05023_),
    .A(_05022_));
 sg13g2_o21ai_1 _13930_ (.B1(_05018_),
    .Y(_05024_),
    .A1(_05020_),
    .A2(_05022_));
 sg13g2_or3_1 _13931_ (.A(_05018_),
    .B(_05020_),
    .C(_05022_),
    .X(_05025_));
 sg13g2_and2_1 _13932_ (.A(_05024_),
    .B(_05025_),
    .X(_00568_));
 sg13g2_xor2_1 _13933_ (.B(net4968),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[13] ),
    .X(_05026_));
 sg13g2_o21ai_1 _13934_ (.B1(_05024_),
    .Y(_05027_),
    .A1(_02401_),
    .A2(net4968));
 sg13g2_xnor2_1 _13935_ (.Y(_00569_),
    .A(_05026_),
    .B(_05027_));
 sg13g2_nor2b_1 _13936_ (.A(net4968),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[14] ),
    .Y(_05028_));
 sg13g2_xnor2_1 _13937_ (.Y(_05029_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[14] ),
    .B(net4967));
 sg13g2_o21ai_1 _13938_ (.B1(net4944),
    .Y(_05030_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[12] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_a22oi_1 _13939_ (.Y(_05031_),
    .B1(_05024_),
    .B2(_05030_),
    .A2(net4968),
    .A1(_02403_));
 sg13g2_xor2_1 _13940_ (.B(_05031_),
    .A(_05029_),
    .X(_00570_));
 sg13g2_xnor2_1 _13941_ (.Y(_05032_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[15] ),
    .B(net4968));
 sg13g2_a21oi_1 _13942_ (.A1(_05029_),
    .A2(_05031_),
    .Y(_05033_),
    .B1(_05028_));
 sg13g2_xnor2_1 _13943_ (.Y(_00571_),
    .A(_05032_),
    .B(_05033_));
 sg13g2_nor2_1 _13944_ (.A(_05019_),
    .B(_05026_),
    .Y(_05034_));
 sg13g2_nand4_1 _13945_ (.B(_05029_),
    .C(_05032_),
    .A(_05020_),
    .Y(_05035_),
    .D(_05034_));
 sg13g2_o21ai_1 _13946_ (.B1(net4944),
    .Y(_05036_),
    .A1(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand4_1 _13947_ (.B(_05030_),
    .C(_05035_),
    .A(_05023_),
    .Y(_05037_),
    .D(_05036_));
 sg13g2_nor2b_1 _13948_ (.A(net4967),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[16] ),
    .Y(_05038_));
 sg13g2_xnor2_1 _13949_ (.Y(_05039_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[16] ),
    .B(net4967));
 sg13g2_xor2_1 _13950_ (.B(_05039_),
    .A(_05037_),
    .X(_00572_));
 sg13g2_a21o_1 _13951_ (.A2(_05039_),
    .A1(_05037_),
    .B1(_05038_),
    .X(_05040_));
 sg13g2_xor2_1 _13952_ (.B(net4967),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[17] ),
    .X(_05041_));
 sg13g2_xnor2_1 _13953_ (.Y(_00573_),
    .A(_05040_),
    .B(_05041_));
 sg13g2_nor3_1 _13954_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[17] ),
    .B(net4967),
    .C(_05040_),
    .Y(_05042_));
 sg13g2_nand3_1 _13955_ (.B(net4967),
    .C(_05040_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[17] ),
    .Y(_05043_));
 sg13g2_nor2b_1 _13956_ (.A(_05042_),
    .B_N(_05043_),
    .Y(_05044_));
 sg13g2_xnor2_1 _13957_ (.Y(_00574_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[18] ),
    .B(_05044_));
 sg13g2_nor2b_1 _13958_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][1] ),
    .Y(_05045_));
 sg13g2_xnor2_1 _13959_ (.Y(_05046_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][1] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _13960_ (.B(_05046_),
    .A(_02510_),
    .X(_00557_));
 sg13g2_a21oi_1 _13961_ (.A1(_02510_),
    .A2(_05046_),
    .Y(_05047_),
    .B1(_05045_));
 sg13g2_xnor2_1 _13962_ (.Y(_05048_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][2] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _13963_ (.A(_05047_),
    .B_N(_05048_),
    .Y(_05049_));
 sg13g2_xnor2_1 _13964_ (.Y(_00558_),
    .A(_05047_),
    .B(_05048_));
 sg13g2_a21oi_1 _13965_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][2] ),
    .A2(_02405_),
    .Y(_05050_),
    .B1(_05049_));
 sg13g2_xnor2_1 _13966_ (.Y(_05051_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][3] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _13967_ (.A(_05050_),
    .B_N(_05051_),
    .Y(_05052_));
 sg13g2_xnor2_1 _13968_ (.Y(_00559_),
    .A(_05050_),
    .B(_05051_));
 sg13g2_a21oi_1 _13969_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][3] ),
    .A2(_02406_),
    .Y(_05053_),
    .B1(_05052_));
 sg13g2_xnor2_1 _13970_ (.Y(_05054_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][4] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _13971_ (.A(_05053_),
    .B_N(_05054_),
    .Y(_05055_));
 sg13g2_xnor2_1 _13972_ (.Y(_00560_),
    .A(_05053_),
    .B(_05054_));
 sg13g2_a21oi_1 _13973_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][4] ),
    .A2(_02407_),
    .Y(_05056_),
    .B1(_05055_));
 sg13g2_xnor2_1 _13974_ (.Y(_05057_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][5] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _13975_ (.A(_05056_),
    .B_N(_05057_),
    .Y(_05058_));
 sg13g2_xnor2_1 _13976_ (.Y(_00561_),
    .A(_05056_),
    .B(_05057_));
 sg13g2_a21oi_1 _13977_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][5] ),
    .A2(_02408_),
    .Y(_05059_),
    .B1(_05058_));
 sg13g2_xnor2_1 _13978_ (.Y(_05060_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][6] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_nor2b_1 _13979_ (.A(_05059_),
    .B_N(_05060_),
    .Y(_05061_));
 sg13g2_xnor2_1 _13980_ (.Y(_00562_),
    .A(_05059_),
    .B(_05060_));
 sg13g2_a21oi_1 _13981_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][6] ),
    .A2(_02409_),
    .Y(_05062_),
    .B1(_05061_));
 sg13g2_xnor2_1 _13982_ (.Y(_05063_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][7] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _13983_ (.A(_05062_),
    .B_N(_05063_),
    .Y(_05064_));
 sg13g2_xnor2_1 _13984_ (.Y(_00563_),
    .A(_05062_),
    .B(_05063_));
 sg13g2_a21oi_1 _13985_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][7] ),
    .A2(_02410_),
    .Y(_05065_),
    .B1(_05064_));
 sg13g2_xnor2_1 _13986_ (.Y(_05066_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][8] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_nor2b_1 _13987_ (.A(_05065_),
    .B_N(_05066_),
    .Y(_05067_));
 sg13g2_xnor2_1 _13988_ (.Y(_00564_),
    .A(_05065_),
    .B(_05066_));
 sg13g2_nor2b_1 _13989_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][9] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[9] ),
    .Y(_05068_));
 sg13g2_nand2b_1 _13990_ (.Y(_05069_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][9] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _13991_ (.A(_05068_),
    .B_N(_05069_),
    .Y(_05070_));
 sg13g2_a21oi_1 _13992_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][8] ),
    .A2(_02411_),
    .Y(_05071_),
    .B1(_05067_));
 sg13g2_xnor2_1 _13993_ (.Y(_00565_),
    .A(_05070_),
    .B(_05071_));
 sg13g2_nor2b_1 _13994_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][10] ),
    .Y(_05072_));
 sg13g2_nand2b_1 _13995_ (.Y(_05073_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][10] ));
 sg13g2_nand2b_1 _13996_ (.Y(_05074_),
    .B(_05073_),
    .A_N(_05072_));
 sg13g2_o21ai_1 _13997_ (.B1(_05069_),
    .Y(_05075_),
    .A1(_05068_),
    .A2(_05071_));
 sg13g2_xnor2_1 _13998_ (.Y(_00548_),
    .A(_05074_),
    .B(_05075_));
 sg13g2_a21oi_1 _13999_ (.A1(_05073_),
    .A2(_05075_),
    .Y(_05076_),
    .B1(_05072_));
 sg13g2_nand2b_1 _14000_ (.Y(_05077_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][11] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _14001_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][11] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[11] ),
    .Y(_05078_));
 sg13g2_xnor2_1 _14002_ (.Y(_05079_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][11] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_xnor2_1 _14003_ (.Y(_00549_),
    .A(_05076_),
    .B(_05079_));
 sg13g2_nor2b_1 _14004_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][12] ),
    .Y(_05080_));
 sg13g2_nand2b_1 _14005_ (.Y(_05081_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][12] ));
 sg13g2_nand2b_1 _14006_ (.Y(_05082_),
    .B(_05081_),
    .A_N(_05080_));
 sg13g2_o21ai_1 _14007_ (.B1(_05077_),
    .Y(_05083_),
    .A1(_05076_),
    .A2(_05078_));
 sg13g2_xnor2_1 _14008_ (.Y(_00550_),
    .A(_05082_),
    .B(_05083_));
 sg13g2_a21oi_1 _14009_ (.A1(_05081_),
    .A2(_05083_),
    .Y(_05084_),
    .B1(_05080_));
 sg13g2_nand2b_1 _14010_ (.Y(_05085_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][13] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _14011_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][13] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[13] ),
    .Y(_05086_));
 sg13g2_xnor2_1 _14012_ (.Y(_05087_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][13] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_xnor2_1 _14013_ (.Y(_00551_),
    .A(_05084_),
    .B(_05087_));
 sg13g2_nor2b_1 _14014_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][14] ),
    .Y(_05088_));
 sg13g2_nand2b_1 _14015_ (.Y(_05089_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][14] ));
 sg13g2_nand2b_1 _14016_ (.Y(_05090_),
    .B(_05089_),
    .A_N(_05088_));
 sg13g2_o21ai_1 _14017_ (.B1(_05085_),
    .Y(_05091_),
    .A1(_05084_),
    .A2(_05086_));
 sg13g2_xnor2_1 _14018_ (.Y(_00552_),
    .A(_05090_),
    .B(_05091_));
 sg13g2_a21oi_1 _14019_ (.A1(_05089_),
    .A2(_05091_),
    .Y(_05092_),
    .B1(_05088_));
 sg13g2_nor2b_1 _14020_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][15] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[15] ),
    .Y(_05093_));
 sg13g2_nand2b_1 _14021_ (.Y(_05094_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][15] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _14022_ (.A(_05093_),
    .B_N(_05094_),
    .Y(_05095_));
 sg13g2_xnor2_1 _14023_ (.Y(_00553_),
    .A(_05092_),
    .B(_05095_));
 sg13g2_xor2_1 _14024_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][16] ),
    .X(_05096_));
 sg13g2_a21oi_1 _14025_ (.A1(_05092_),
    .A2(_05094_),
    .Y(_05097_),
    .B1(_05093_));
 sg13g2_nor2b_1 _14026_ (.A(_05096_),
    .B_N(_05097_),
    .Y(_05098_));
 sg13g2_xnor2_1 _14027_ (.Y(_00554_),
    .A(_05096_),
    .B(_05097_));
 sg13g2_a21oi_1 _14028_ (.A1(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][16] ),
    .A2(_02412_),
    .Y(_05099_),
    .B1(_05098_));
 sg13g2_nand2b_1 _14029_ (.Y(_05100_),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][17] ),
    .A_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _14030_ (.A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][17] ),
    .B_N(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[17] ),
    .Y(_05101_));
 sg13g2_xnor2_1 _14031_ (.Y(_05102_),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][17] ),
    .B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _14032_ (.Y(_00555_),
    .A(_05099_),
    .B(_05102_));
 sg13g2_o21ai_1 _14033_ (.B1(_05100_),
    .Y(_05103_),
    .A1(_05099_),
    .A2(_05101_));
 sg13g2_xor2_1 _14034_ (.B(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][18] ),
    .X(_05104_));
 sg13g2_xnor2_1 _14035_ (.Y(_00556_),
    .A(_05103_),
    .B(_05104_));
 sg13g2_nand2_1 _14036_ (.Y(_05105_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[0] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_xor2_1 _14037_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[0] ),
    .X(_00697_));
 sg13g2_nand2_1 _14038_ (.Y(_05106_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_nor2_1 _14039_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[1] ),
    .Y(_05107_));
 sg13g2_xor2_1 _14040_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[1] ),
    .X(_05108_));
 sg13g2_xnor2_1 _14041_ (.Y(_00707_),
    .A(_05105_),
    .B(_05108_));
 sg13g2_o21ai_1 _14042_ (.B1(_05106_),
    .Y(_05109_),
    .A1(_05105_),
    .A2(_05107_));
 sg13g2_xnor2_1 _14043_ (.Y(_05110_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[2] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_nor2b_1 _14044_ (.A(_05110_),
    .B_N(_05109_),
    .Y(_05111_));
 sg13g2_xnor2_1 _14045_ (.Y(_00708_),
    .A(_05109_),
    .B(_05110_));
 sg13g2_a21o_1 _14046_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[2] ),
    .B1(_05111_),
    .X(_05112_));
 sg13g2_xnor2_1 _14047_ (.Y(_05113_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[3] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_nor2b_1 _14048_ (.A(_05113_),
    .B_N(_05112_),
    .Y(_05114_));
 sg13g2_xnor2_1 _14049_ (.Y(_00709_),
    .A(_05112_),
    .B(_05113_));
 sg13g2_a21o_1 _14050_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[3] ),
    .B1(_05114_),
    .X(_05115_));
 sg13g2_xnor2_1 _14051_ (.Y(_05116_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[4] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_nor2b_1 _14052_ (.A(_05116_),
    .B_N(_05115_),
    .Y(_05117_));
 sg13g2_xnor2_1 _14053_ (.Y(_00710_),
    .A(_05115_),
    .B(_05116_));
 sg13g2_a21o_1 _14054_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[4] ),
    .B1(_05117_),
    .X(_05118_));
 sg13g2_xnor2_1 _14055_ (.Y(_05119_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[5] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_nor2b_1 _14056_ (.A(_05119_),
    .B_N(_05118_),
    .Y(_05120_));
 sg13g2_xnor2_1 _14057_ (.Y(_00711_),
    .A(_05118_),
    .B(_05119_));
 sg13g2_a21o_1 _14058_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[5] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[5] ),
    .B1(_05120_),
    .X(_05121_));
 sg13g2_xnor2_1 _14059_ (.Y(_05122_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[6] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_nor2b_1 _14060_ (.A(_05122_),
    .B_N(_05121_),
    .Y(_05123_));
 sg13g2_xnor2_1 _14061_ (.Y(_00712_),
    .A(_05121_),
    .B(_05122_));
 sg13g2_a21o_1 _14062_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[6] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[6] ),
    .B1(_05123_),
    .X(_05124_));
 sg13g2_xnor2_1 _14063_ (.Y(_05125_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[7] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_nor2b_1 _14064_ (.A(_05125_),
    .B_N(_05124_),
    .Y(_05126_));
 sg13g2_xnor2_1 _14065_ (.Y(_00713_),
    .A(_05124_),
    .B(_05125_));
 sg13g2_a21o_1 _14066_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[7] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[7] ),
    .B1(_05126_),
    .X(_05127_));
 sg13g2_xnor2_1 _14067_ (.Y(_05128_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[8] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_nor2b_1 _14068_ (.A(_05128_),
    .B_N(_05127_),
    .Y(_05129_));
 sg13g2_xnor2_1 _14069_ (.Y(_00714_),
    .A(_05127_),
    .B(_05128_));
 sg13g2_a21o_1 _14070_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[8] ),
    .B1(_05129_),
    .X(_05130_));
 sg13g2_nand2_1 _14071_ (.Y(_05131_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[9] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_xnor2_1 _14072_ (.Y(_05132_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[9] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_xnor2_1 _14073_ (.Y(_00715_),
    .A(_05130_),
    .B(_05132_));
 sg13g2_xnor2_1 _14074_ (.Y(_05133_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[10] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_o21ai_1 _14075_ (.B1(_05130_),
    .Y(_05134_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_a21oi_1 _14076_ (.A1(_05131_),
    .A2(_05134_),
    .Y(_05135_),
    .B1(_05133_));
 sg13g2_nand3_1 _14077_ (.B(_05133_),
    .C(_05134_),
    .A(_05131_),
    .Y(_05136_));
 sg13g2_nor2b_1 _14078_ (.A(_05135_),
    .B_N(_05136_),
    .Y(_00698_));
 sg13g2_a21oi_2 _14079_ (.B1(_05135_),
    .Y(_05137_),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[10] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_nand2_1 _14080_ (.Y(_05138_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[11] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_nor2_1 _14081_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[11] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[11] ),
    .Y(_05139_));
 sg13g2_xor2_1 _14082_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[11] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[11] ),
    .X(_05140_));
 sg13g2_xnor2_1 _14083_ (.Y(_00699_),
    .A(_05137_),
    .B(_05140_));
 sg13g2_xnor2_1 _14084_ (.Y(_05141_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[12] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_o21ai_1 _14085_ (.B1(_05138_),
    .Y(_05142_),
    .A1(_05137_),
    .A2(_05139_));
 sg13g2_nor2b_1 _14086_ (.A(_05141_),
    .B_N(_05142_),
    .Y(_05143_));
 sg13g2_xnor2_1 _14087_ (.Y(_00700_),
    .A(_05141_),
    .B(_05142_));
 sg13g2_a21o_1 _14088_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[12] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[12] ),
    .B1(_05143_),
    .X(_05144_));
 sg13g2_xnor2_1 _14089_ (.Y(_05145_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[13] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_xnor2_1 _14090_ (.Y(_00701_),
    .A(_05144_),
    .B(_05145_));
 sg13g2_xor2_1 _14091_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[14] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[14] ),
    .X(_05146_));
 sg13g2_a21o_1 _14092_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[13] ),
    .B1(_05144_),
    .X(_05147_));
 sg13g2_o21ai_1 _14093_ (.B1(_05147_),
    .Y(_05148_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_nor2b_1 _14094_ (.A(_05148_),
    .B_N(_05146_),
    .Y(_05149_));
 sg13g2_xnor2_1 _14095_ (.Y(_00702_),
    .A(_05146_),
    .B(_05148_));
 sg13g2_a21o_1 _14096_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[14] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[14] ),
    .B1(_05149_),
    .X(_05150_));
 sg13g2_nand2_1 _14097_ (.Y(_05151_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_xnor2_1 _14098_ (.Y(_05152_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_xnor2_1 _14099_ (.Y(_00703_),
    .A(_05150_),
    .B(_05152_));
 sg13g2_nand2_1 _14100_ (.Y(_05153_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[16] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_xor2_1 _14101_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[16] ),
    .X(_05154_));
 sg13g2_o21ai_1 _14102_ (.B1(_05150_),
    .Y(_05155_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[15] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_nand2_1 _14103_ (.Y(_05156_),
    .A(_05151_),
    .B(_05155_));
 sg13g2_nand2_1 _14104_ (.Y(_05157_),
    .A(_05154_),
    .B(_05156_));
 sg13g2_xor2_1 _14105_ (.B(_05156_),
    .A(_05154_),
    .X(_00704_));
 sg13g2_xnor2_1 _14106_ (.Y(_05158_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[17] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_a21oi_1 _14107_ (.A1(_05153_),
    .A2(_05157_),
    .Y(_05159_),
    .B1(_05158_));
 sg13g2_nand3_1 _14108_ (.B(_05157_),
    .C(_05158_),
    .A(_05153_),
    .Y(_05160_));
 sg13g2_nor2b_1 _14109_ (.A(_05159_),
    .B_N(_05160_),
    .Y(_00705_));
 sg13g2_a21oi_1 _14110_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[17] ),
    .Y(_05161_),
    .B1(_05159_));
 sg13g2_xor2_1 _14111_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[18] ),
    .X(_05162_));
 sg13g2_xnor2_1 _14112_ (.Y(_00706_),
    .A(_05161_),
    .B(_05162_));
 sg13g2_nor2b_1 _14113_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][1] ),
    .Y(_05163_));
 sg13g2_xnor2_1 _14114_ (.Y(_05164_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][1] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _14115_ (.B(_05164_),
    .A(_02511_),
    .X(_00726_));
 sg13g2_a21oi_2 _14116_ (.B1(_05163_),
    .Y(_05165_),
    .A2(_05164_),
    .A1(_02511_));
 sg13g2_xnor2_1 _14117_ (.Y(_05166_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][2] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _14118_ (.A(_05165_),
    .B_N(_05166_),
    .Y(_05167_));
 sg13g2_xnor2_1 _14119_ (.Y(_00727_),
    .A(_05165_),
    .B(_05166_));
 sg13g2_a21oi_2 _14120_ (.B1(_05167_),
    .Y(_05168_),
    .A2(_02413_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][2] ));
 sg13g2_xnor2_1 _14121_ (.Y(_05169_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][3] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _14122_ (.A(_05168_),
    .B_N(_05169_),
    .Y(_05170_));
 sg13g2_xnor2_1 _14123_ (.Y(_00728_),
    .A(_05168_),
    .B(_05169_));
 sg13g2_a21oi_2 _14124_ (.B1(_05170_),
    .Y(_05171_),
    .A2(_02414_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][3] ));
 sg13g2_xnor2_1 _14125_ (.Y(_05172_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][4] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _14126_ (.A(_05171_),
    .B_N(_05172_),
    .Y(_05173_));
 sg13g2_xnor2_1 _14127_ (.Y(_00729_),
    .A(_05171_),
    .B(_05172_));
 sg13g2_a21oi_2 _14128_ (.B1(_05173_),
    .Y(_05174_),
    .A2(_02415_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][4] ));
 sg13g2_nand2b_1 _14129_ (.Y(_05175_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][5] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _14130_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][5] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[5] ),
    .Y(_05176_));
 sg13g2_xnor2_1 _14131_ (.Y(_05177_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][5] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_xnor2_1 _14132_ (.Y(_00730_),
    .A(_05174_),
    .B(_05177_));
 sg13g2_nor2b_1 _14133_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[6] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][6] ),
    .Y(_05178_));
 sg13g2_nand2b_1 _14134_ (.Y(_05179_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[6] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][6] ));
 sg13g2_nand2b_1 _14135_ (.Y(_05180_),
    .B(_05179_),
    .A_N(_05178_));
 sg13g2_o21ai_1 _14136_ (.B1(_05175_),
    .Y(_05181_),
    .A1(_05174_),
    .A2(_05176_));
 sg13g2_xnor2_1 _14137_ (.Y(_00731_),
    .A(_05180_),
    .B(_05181_));
 sg13g2_a21oi_1 _14138_ (.A1(_05179_),
    .A2(_05181_),
    .Y(_05182_),
    .B1(_05178_));
 sg13g2_xnor2_1 _14139_ (.Y(_05183_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][7] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nand2b_1 _14140_ (.Y(_05184_),
    .B(_05183_),
    .A_N(_05182_));
 sg13g2_xnor2_1 _14141_ (.Y(_00732_),
    .A(_05182_),
    .B(_05183_));
 sg13g2_o21ai_1 _14142_ (.B1(_05184_),
    .Y(_05185_),
    .A1(_02416_),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _14143_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[8] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][8] ),
    .Y(_05186_));
 sg13g2_nand2b_1 _14144_ (.Y(_05187_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[8] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][8] ));
 sg13g2_nand2b_1 _14145_ (.Y(_05188_),
    .B(_05187_),
    .A_N(_05186_));
 sg13g2_xnor2_1 _14146_ (.Y(_00733_),
    .A(_05185_),
    .B(_05188_));
 sg13g2_a21oi_2 _14147_ (.B1(_05186_),
    .Y(_05189_),
    .A2(_05187_),
    .A1(_05185_));
 sg13g2_nand2b_1 _14148_ (.Y(_05190_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][9] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _14149_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][9] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[9] ),
    .Y(_05191_));
 sg13g2_xnor2_1 _14150_ (.Y(_05192_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][9] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_xnor2_1 _14151_ (.Y(_00734_),
    .A(_05189_),
    .B(_05192_));
 sg13g2_nor2b_1 _14152_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][10] ),
    .Y(_05193_));
 sg13g2_nand2b_1 _14153_ (.Y(_05194_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][10] ));
 sg13g2_nand2b_1 _14154_ (.Y(_05195_),
    .B(_05194_),
    .A_N(_05193_));
 sg13g2_a21oi_2 _14155_ (.B1(_05191_),
    .Y(_05196_),
    .A2(_05190_),
    .A1(_05189_));
 sg13g2_xnor2_1 _14156_ (.Y(_00717_),
    .A(_05195_),
    .B(_05196_));
 sg13g2_a21oi_2 _14157_ (.B1(_05193_),
    .Y(_05197_),
    .A2(_05196_),
    .A1(_05194_));
 sg13g2_nor2b_1 _14158_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][11] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[11] ),
    .Y(_05198_));
 sg13g2_nand2b_1 _14159_ (.Y(_05199_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][11] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _14160_ (.A(_05198_),
    .B_N(_05199_),
    .Y(_05200_));
 sg13g2_xnor2_1 _14161_ (.Y(_00718_),
    .A(_05197_),
    .B(_05200_));
 sg13g2_nor2b_1 _14162_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][12] ),
    .Y(_05201_));
 sg13g2_nand2b_1 _14163_ (.Y(_05202_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][12] ));
 sg13g2_nand2b_1 _14164_ (.Y(_05203_),
    .B(_05202_),
    .A_N(_05201_));
 sg13g2_a21oi_2 _14165_ (.B1(_05198_),
    .Y(_05204_),
    .A2(_05199_),
    .A1(_05197_));
 sg13g2_xnor2_1 _14166_ (.Y(_00719_),
    .A(_05203_),
    .B(_05204_));
 sg13g2_a21oi_2 _14167_ (.B1(_05201_),
    .Y(_05205_),
    .A2(_05204_),
    .A1(_05202_));
 sg13g2_nor2b_1 _14168_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][13] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[13] ),
    .Y(_05206_));
 sg13g2_nand2b_1 _14169_ (.Y(_05207_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][13] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _14170_ (.A(_05206_),
    .B_N(_05207_),
    .Y(_05208_));
 sg13g2_xnor2_1 _14171_ (.Y(_00720_),
    .A(_05205_),
    .B(_05208_));
 sg13g2_nor2b_1 _14172_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][14] ),
    .Y(_05209_));
 sg13g2_nand2b_1 _14173_ (.Y(_05210_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][14] ));
 sg13g2_nand2b_1 _14174_ (.Y(_05211_),
    .B(_05210_),
    .A_N(_05209_));
 sg13g2_a21oi_2 _14175_ (.B1(_05206_),
    .Y(_05212_),
    .A2(_05207_),
    .A1(_05205_));
 sg13g2_xnor2_1 _14176_ (.Y(_00721_),
    .A(_05211_),
    .B(_05212_));
 sg13g2_a21oi_2 _14177_ (.B1(_05209_),
    .Y(_05213_),
    .A2(_05212_),
    .A1(_05210_));
 sg13g2_nor2b_1 _14178_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][15] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[15] ),
    .Y(_05214_));
 sg13g2_nand2b_1 _14179_ (.Y(_05215_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][15] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _14180_ (.A(_05214_),
    .B_N(_05215_),
    .Y(_05216_));
 sg13g2_xnor2_1 _14181_ (.Y(_00722_),
    .A(_05213_),
    .B(_05216_));
 sg13g2_nor2b_1 _14182_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[16] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][16] ),
    .Y(_05217_));
 sg13g2_nand2b_1 _14183_ (.Y(_05218_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[16] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][16] ));
 sg13g2_nand2b_1 _14184_ (.Y(_05219_),
    .B(_05218_),
    .A_N(_05217_));
 sg13g2_a21oi_2 _14185_ (.B1(_05214_),
    .Y(_05220_),
    .A2(_05215_),
    .A1(_05213_));
 sg13g2_xnor2_1 _14186_ (.Y(_00723_),
    .A(_05219_),
    .B(_05220_));
 sg13g2_a21oi_2 _14187_ (.B1(_05217_),
    .Y(_05221_),
    .A2(_05220_),
    .A1(_05218_));
 sg13g2_nand2b_1 _14188_ (.Y(_05222_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][17] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _14189_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][17] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[17] ),
    .Y(_05223_));
 sg13g2_xnor2_1 _14190_ (.Y(_05224_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][17] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _14191_ (.Y(_00724_),
    .A(_05221_),
    .B(_05224_));
 sg13g2_o21ai_1 _14192_ (.B1(_05222_),
    .Y(_05225_),
    .A1(_05221_),
    .A2(_05223_));
 sg13g2_xor2_1 _14193_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][18] ),
    .X(_05226_));
 sg13g2_xnor2_1 _14194_ (.Y(_00725_),
    .A(_05225_),
    .B(_05226_));
 sg13g2_nand2_1 _14195_ (.Y(_05227_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[0] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_xor2_1 _14196_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[0] ),
    .X(_00678_));
 sg13g2_nand2_1 _14197_ (.Y(_05228_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_nor2_1 _14198_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[1] ),
    .Y(_05229_));
 sg13g2_xor2_1 _14199_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[1] ),
    .X(_05230_));
 sg13g2_xnor2_1 _14200_ (.Y(_00688_),
    .A(_05227_),
    .B(_05230_));
 sg13g2_o21ai_1 _14201_ (.B1(_05228_),
    .Y(_05231_),
    .A1(_05227_),
    .A2(_05229_));
 sg13g2_xnor2_1 _14202_ (.Y(_05232_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[2] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_nor2b_1 _14203_ (.A(_05232_),
    .B_N(_05231_),
    .Y(_05233_));
 sg13g2_xnor2_1 _14204_ (.Y(_00689_),
    .A(_05231_),
    .B(_05232_));
 sg13g2_a21o_1 _14205_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[2] ),
    .B1(_05233_),
    .X(_05234_));
 sg13g2_xnor2_1 _14206_ (.Y(_05235_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[3] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_nor2b_1 _14207_ (.A(_05235_),
    .B_N(_05234_),
    .Y(_05236_));
 sg13g2_xnor2_1 _14208_ (.Y(_00690_),
    .A(_05234_),
    .B(_05235_));
 sg13g2_a21o_1 _14209_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[3] ),
    .B1(_05236_),
    .X(_05237_));
 sg13g2_xnor2_1 _14210_ (.Y(_05238_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[4] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_nor2b_1 _14211_ (.A(_05238_),
    .B_N(_05237_),
    .Y(_05239_));
 sg13g2_xnor2_1 _14212_ (.Y(_00691_),
    .A(_05237_),
    .B(_05238_));
 sg13g2_a21o_1 _14213_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[4] ),
    .B1(_05239_),
    .X(_05240_));
 sg13g2_nand2_1 _14214_ (.Y(_05241_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _14215_ (.Y(_05242_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _14216_ (.Y(_00692_),
    .A(_05240_),
    .B(_05242_));
 sg13g2_xnor2_1 _14217_ (.Y(_05243_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[6] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_o21ai_1 _14218_ (.B1(_05240_),
    .Y(_05244_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_a21oi_1 _14219_ (.A1(_05241_),
    .A2(_05244_),
    .Y(_05245_),
    .B1(_05243_));
 sg13g2_nand3_1 _14220_ (.B(_05243_),
    .C(_05244_),
    .A(_05241_),
    .Y(_05246_));
 sg13g2_nor2b_1 _14221_ (.A(_05245_),
    .B_N(_05246_),
    .Y(_00693_));
 sg13g2_a21oi_2 _14222_ (.B1(_05245_),
    .Y(_05247_),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[6] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_nand2_1 _14223_ (.Y(_05248_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_nor2_1 _14224_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[7] ),
    .Y(_05249_));
 sg13g2_xor2_1 _14225_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[7] ),
    .X(_05250_));
 sg13g2_xnor2_1 _14226_ (.Y(_00694_),
    .A(_05247_),
    .B(_05250_));
 sg13g2_o21ai_1 _14227_ (.B1(_05248_),
    .Y(_05251_),
    .A1(_05247_),
    .A2(_05249_));
 sg13g2_xnor2_1 _14228_ (.Y(_05252_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[8] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_nor2b_1 _14229_ (.A(_05252_),
    .B_N(_05251_),
    .Y(_05253_));
 sg13g2_xnor2_1 _14230_ (.Y(_00695_),
    .A(_05251_),
    .B(_05252_));
 sg13g2_a21o_1 _14231_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[8] ),
    .B1(_05253_),
    .X(_05254_));
 sg13g2_xnor2_1 _14232_ (.Y(_05255_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[9] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _14233_ (.Y(_00696_),
    .A(_05254_),
    .B(_05255_));
 sg13g2_nand2_1 _14234_ (.Y(_05256_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_nor2_1 _14235_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[10] ),
    .Y(_05257_));
 sg13g2_xor2_1 _14236_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[10] ),
    .X(_05258_));
 sg13g2_a21o_1 _14237_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[9] ),
    .B1(_05254_),
    .X(_05259_));
 sg13g2_o21ai_1 _14238_ (.B1(_05259_),
    .Y(_05260_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _14239_ (.Y(_00679_),
    .A(_05258_),
    .B(_05260_));
 sg13g2_o21ai_1 _14240_ (.B1(_05256_),
    .Y(_05261_),
    .A1(_05257_),
    .A2(_05260_));
 sg13g2_xnor2_1 _14241_ (.Y(_05262_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[11] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _14242_ (.Y(_00680_),
    .A(_05261_),
    .B(_05262_));
 sg13g2_nand2_1 _14243_ (.Y(_05263_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[12] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_nor2_1 _14244_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[12] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[12] ),
    .Y(_05264_));
 sg13g2_xor2_1 _14245_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[12] ),
    .X(_05265_));
 sg13g2_a21o_1 _14246_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[11] ),
    .B1(_05261_),
    .X(_05266_));
 sg13g2_o21ai_1 _14247_ (.B1(_05266_),
    .Y(_05267_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _14248_ (.Y(_00681_),
    .A(_05265_),
    .B(_05267_));
 sg13g2_o21ai_1 _14249_ (.B1(_05263_),
    .Y(_05268_),
    .A1(_05264_),
    .A2(_05267_));
 sg13g2_xnor2_1 _14250_ (.Y(_05269_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[13] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_xnor2_1 _14251_ (.Y(_00682_),
    .A(_05268_),
    .B(_05269_));
 sg13g2_xor2_1 _14252_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[14] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[14] ),
    .X(_05270_));
 sg13g2_a21o_1 _14253_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[13] ),
    .B1(_05268_),
    .X(_05271_));
 sg13g2_o21ai_1 _14254_ (.B1(_05271_),
    .Y(_05272_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_nor2b_1 _14255_ (.A(_05272_),
    .B_N(_05270_),
    .Y(_05273_));
 sg13g2_xnor2_1 _14256_ (.Y(_00683_),
    .A(_05270_),
    .B(_05272_));
 sg13g2_a21o_1 _14257_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[14] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[14] ),
    .B1(_05273_),
    .X(_05274_));
 sg13g2_and2_1 _14258_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[15] ),
    .X(_05275_));
 sg13g2_or2_1 _14259_ (.X(_05276_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[15] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand2b_1 _14260_ (.Y(_05277_),
    .B(_05276_),
    .A_N(_05275_));
 sg13g2_xnor2_1 _14261_ (.Y(_00684_),
    .A(_05274_),
    .B(_05277_));
 sg13g2_and2_1 _14262_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[16] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[16] ),
    .X(_05278_));
 sg13g2_xor2_1 _14263_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[16] ),
    .X(_05279_));
 sg13g2_a21o_1 _14264_ (.A2(_05276_),
    .A1(_05274_),
    .B1(_05275_),
    .X(_05280_));
 sg13g2_xor2_1 _14265_ (.B(_05280_),
    .A(_05279_),
    .X(_00685_));
 sg13g2_a21o_1 _14266_ (.A2(_05280_),
    .A1(_05279_),
    .B1(_05278_),
    .X(_05281_));
 sg13g2_xnor2_1 _14267_ (.Y(_05282_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[17] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xnor2_1 _14268_ (.Y(_00686_),
    .A(_05281_),
    .B(_05282_));
 sg13g2_a21o_1 _14269_ (.A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[17] ),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[17] ),
    .B1(_05281_),
    .X(_05283_));
 sg13g2_o21ai_1 _14270_ (.B1(_05283_),
    .Y(_05284_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xor2_1 _14271_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[18] ),
    .X(_05285_));
 sg13g2_xnor2_1 _14272_ (.Y(_00687_),
    .A(_05284_),
    .B(_05285_));
 sg13g2_nand2b_1 _14273_ (.Y(_05286_),
    .B(net4962),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_nor2b_1 _14274_ (.A(net4961),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[1] ),
    .Y(_05287_));
 sg13g2_xnor2_1 _14275_ (.Y(_05288_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[1] ),
    .B(net4961));
 sg13g2_xnor2_1 _14276_ (.Y(_00669_),
    .A(_01191_),
    .B(_05288_));
 sg13g2_xnor2_1 _14277_ (.Y(_05289_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[2] ),
    .B(net4961));
 sg13g2_o21ai_1 _14278_ (.B1(_05286_),
    .Y(_05290_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[0] ),
    .A2(_05287_));
 sg13g2_nor2b_1 _14279_ (.A(_05290_),
    .B_N(_05289_),
    .Y(_05291_));
 sg13g2_xnor2_1 _14280_ (.Y(_00670_),
    .A(_05289_),
    .B(_05290_));
 sg13g2_a21oi_1 _14281_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[2] ),
    .A2(net4943),
    .Y(_05292_),
    .B1(_05291_));
 sg13g2_nor2_1 _14282_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4943),
    .Y(_05293_));
 sg13g2_nand2_1 _14283_ (.Y(_05294_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4943));
 sg13g2_nor2b_1 _14284_ (.A(_05293_),
    .B_N(_05294_),
    .Y(_05295_));
 sg13g2_xnor2_1 _14285_ (.Y(_00671_),
    .A(_05292_),
    .B(_05295_));
 sg13g2_xnor2_1 _14286_ (.Y(_05296_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[4] ),
    .B(net4961));
 sg13g2_o21ai_1 _14287_ (.B1(_05294_),
    .Y(_05297_),
    .A1(_05292_),
    .A2(_05293_));
 sg13g2_and2_1 _14288_ (.A(_05296_),
    .B(_05297_),
    .X(_05298_));
 sg13g2_xor2_1 _14289_ (.B(_05297_),
    .A(_05296_),
    .X(_00672_));
 sg13g2_xnor2_1 _14290_ (.Y(_05299_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[5] ),
    .B(net4961));
 sg13g2_a21oi_1 _14291_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[4] ),
    .A2(net4943),
    .Y(_05300_),
    .B1(_05298_));
 sg13g2_xnor2_1 _14292_ (.Y(_00673_),
    .A(_05299_),
    .B(_05300_));
 sg13g2_o21ai_1 _14293_ (.B1(net4943),
    .Y(_05301_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[4] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_and2_1 _14294_ (.A(_05298_),
    .B(_05299_),
    .X(_05302_));
 sg13g2_nor2b_1 _14295_ (.A(_05302_),
    .B_N(_05301_),
    .Y(_05303_));
 sg13g2_nand2_1 _14296_ (.Y(_05304_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4943));
 sg13g2_nor2_1 _14297_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4942),
    .Y(_05305_));
 sg13g2_xnor2_1 _14298_ (.Y(_05306_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4961));
 sg13g2_xnor2_1 _14299_ (.Y(_00674_),
    .A(_05303_),
    .B(_05306_));
 sg13g2_nand2b_1 _14300_ (.Y(_05307_),
    .B(net4961),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_xor2_1 _14301_ (.B(net4961),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[7] ),
    .X(_05308_));
 sg13g2_o21ai_1 _14302_ (.B1(_05304_),
    .Y(_05309_),
    .A1(_05303_),
    .A2(_05305_));
 sg13g2_xnor2_1 _14303_ (.Y(_00675_),
    .A(_05308_),
    .B(_05309_));
 sg13g2_xnor2_1 _14304_ (.Y(_05310_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[8] ),
    .B(net4962));
 sg13g2_o21ai_1 _14305_ (.B1(net4943),
    .Y(_05311_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_nand3_1 _14306_ (.B(_05306_),
    .C(_05307_),
    .A(_05302_),
    .Y(_05312_));
 sg13g2_and3_1 _14307_ (.X(_05313_),
    .A(_05301_),
    .B(_05311_),
    .C(_05312_));
 sg13g2_nand2b_1 _14308_ (.Y(_05314_),
    .B(_05310_),
    .A_N(_05313_));
 sg13g2_xnor2_1 _14309_ (.Y(_00676_),
    .A(_05310_),
    .B(_05313_));
 sg13g2_xor2_1 _14310_ (.B(net4962),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[9] ),
    .X(_05315_));
 sg13g2_o21ai_1 _14311_ (.B1(_05314_),
    .Y(_05316_),
    .A1(_02417_),
    .A2(net4962));
 sg13g2_xnor2_1 _14312_ (.Y(_00677_),
    .A(_05315_),
    .B(_05316_));
 sg13g2_o21ai_1 _14313_ (.B1(net4942),
    .Y(_05317_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[8] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_nor2_1 _14314_ (.A(_05314_),
    .B(_05315_),
    .Y(_05318_));
 sg13g2_nor2b_1 _14315_ (.A(_05318_),
    .B_N(_05317_),
    .Y(_05319_));
 sg13g2_nand2_1 _14316_ (.Y(_05320_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4942));
 sg13g2_nor2_1 _14317_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4942),
    .Y(_05321_));
 sg13g2_xnor2_1 _14318_ (.Y(_05322_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4960));
 sg13g2_xnor2_1 _14319_ (.Y(_00660_),
    .A(_05319_),
    .B(_05322_));
 sg13g2_xor2_1 _14320_ (.B(net4960),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[11] ),
    .X(_05323_));
 sg13g2_o21ai_1 _14321_ (.B1(_05320_),
    .Y(_05324_),
    .A1(_05319_),
    .A2(_05321_));
 sg13g2_xnor2_1 _14322_ (.Y(_00661_),
    .A(_05323_),
    .B(_05324_));
 sg13g2_xnor2_1 _14323_ (.Y(_05325_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[12] ),
    .B(net4960));
 sg13g2_nand2_1 _14324_ (.Y(_05326_),
    .A(_05318_),
    .B(_05322_));
 sg13g2_nor2_1 _14325_ (.A(_05323_),
    .B(_05326_),
    .Y(_05327_));
 sg13g2_o21ai_1 _14326_ (.B1(net4942),
    .Y(_05328_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[10] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_nand2_1 _14327_ (.Y(_05329_),
    .A(_05317_),
    .B(_05328_));
 sg13g2_inv_1 _14328_ (.Y(_05330_),
    .A(_05329_));
 sg13g2_o21ai_1 _14329_ (.B1(_05325_),
    .Y(_05331_),
    .A1(_05327_),
    .A2(_05329_));
 sg13g2_or3_1 _14330_ (.A(_05325_),
    .B(_05327_),
    .C(_05329_),
    .X(_05332_));
 sg13g2_and2_1 _14331_ (.A(_05331_),
    .B(_05332_),
    .X(_00662_));
 sg13g2_nand2_1 _14332_ (.Y(_05333_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[13] ),
    .B(net4942));
 sg13g2_nand2_1 _14333_ (.Y(_05334_),
    .A(_02419_),
    .B(net4960));
 sg13g2_nand2_1 _14334_ (.Y(_05335_),
    .A(_05333_),
    .B(_05334_));
 sg13g2_o21ai_1 _14335_ (.B1(_05331_),
    .Y(_05336_),
    .A1(_02418_),
    .A2(net4960));
 sg13g2_xnor2_1 _14336_ (.Y(_00663_),
    .A(_05335_),
    .B(_05336_));
 sg13g2_nor2b_1 _14337_ (.A(net4959),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[14] ),
    .Y(_05337_));
 sg13g2_xnor2_1 _14338_ (.Y(_05338_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[14] ),
    .B(net4959));
 sg13g2_o21ai_1 _14339_ (.B1(net4942),
    .Y(_05339_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[12] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_a22oi_1 _14340_ (.Y(_05340_),
    .B1(_05331_),
    .B2(_05339_),
    .A2(net4960),
    .A1(_02419_));
 sg13g2_xor2_1 _14341_ (.B(_05340_),
    .A(_05338_),
    .X(_00664_));
 sg13g2_xnor2_1 _14342_ (.Y(_05341_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[15] ),
    .B(net4959));
 sg13g2_a21oi_1 _14343_ (.A1(_05338_),
    .A2(_05340_),
    .Y(_05342_),
    .B1(_05337_));
 sg13g2_xnor2_1 _14344_ (.Y(_00665_),
    .A(_05341_),
    .B(_05342_));
 sg13g2_and4_1 _14345_ (.A(_05325_),
    .B(_05333_),
    .C(_05334_),
    .D(_05341_),
    .X(_05343_));
 sg13g2_nand3_1 _14346_ (.B(_05338_),
    .C(_05343_),
    .A(_05327_),
    .Y(_05344_));
 sg13g2_o21ai_1 _14347_ (.B1(net4942),
    .Y(_05345_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand4_1 _14348_ (.B(_05339_),
    .C(_05344_),
    .A(_05330_),
    .Y(_05346_),
    .D(_05345_));
 sg13g2_nor2b_1 _14349_ (.A(net4959),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[16] ),
    .Y(_05347_));
 sg13g2_xnor2_1 _14350_ (.Y(_05348_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[16] ),
    .B(net4959));
 sg13g2_xor2_1 _14351_ (.B(_05348_),
    .A(_05346_),
    .X(_00666_));
 sg13g2_a21o_1 _14352_ (.A2(_05348_),
    .A1(_05346_),
    .B1(_05347_),
    .X(_05349_));
 sg13g2_xor2_1 _14353_ (.B(net4959),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[17] ),
    .X(_05350_));
 sg13g2_xnor2_1 _14354_ (.Y(_00667_),
    .A(_05349_),
    .B(_05350_));
 sg13g2_nor3_1 _14355_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[17] ),
    .B(net4959),
    .C(_05349_),
    .Y(_05351_));
 sg13g2_nand3_1 _14356_ (.B(net4959),
    .C(_05349_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[17] ),
    .Y(_05352_));
 sg13g2_nor2b_1 _14357_ (.A(_05351_),
    .B_N(_05352_),
    .Y(_05353_));
 sg13g2_xnor2_1 _14358_ (.Y(_00668_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[18] ),
    .B(_05353_));
 sg13g2_nor2b_1 _14359_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][1] ),
    .Y(_05354_));
 sg13g2_xnor2_1 _14360_ (.Y(_05355_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][1] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _14361_ (.B(_05355_),
    .A(_02512_),
    .X(_00651_));
 sg13g2_a21oi_1 _14362_ (.A1(_02512_),
    .A2(_05355_),
    .Y(_05356_),
    .B1(_05354_));
 sg13g2_xnor2_1 _14363_ (.Y(_05357_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][2] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _14364_ (.A(_05356_),
    .B_N(_05357_),
    .Y(_05358_));
 sg13g2_xnor2_1 _14365_ (.Y(_00652_),
    .A(_05356_),
    .B(_05357_));
 sg13g2_a21oi_1 _14366_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][2] ),
    .A2(_02421_),
    .Y(_05359_),
    .B1(_05358_));
 sg13g2_xnor2_1 _14367_ (.Y(_05360_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][3] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _14368_ (.A(_05359_),
    .B_N(_05360_),
    .Y(_05361_));
 sg13g2_xnor2_1 _14369_ (.Y(_00653_),
    .A(_05359_),
    .B(_05360_));
 sg13g2_a21oi_1 _14370_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][3] ),
    .A2(_02422_),
    .Y(_05362_),
    .B1(_05361_));
 sg13g2_xnor2_1 _14371_ (.Y(_05363_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][4] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _14372_ (.A(_05362_),
    .B_N(_05363_),
    .Y(_05364_));
 sg13g2_xnor2_1 _14373_ (.Y(_00654_),
    .A(_05362_),
    .B(_05363_));
 sg13g2_a21oi_1 _14374_ (.A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][4] ),
    .A2(_02423_),
    .Y(_05365_),
    .B1(_05364_));
 sg13g2_nand2b_1 _14375_ (.Y(_05366_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][5] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _14376_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][5] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[5] ),
    .Y(_05367_));
 sg13g2_xnor2_1 _14377_ (.Y(_05368_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][5] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_xnor2_1 _14378_ (.Y(_00655_),
    .A(_05365_),
    .B(_05368_));
 sg13g2_nor2b_1 _14379_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][6] ),
    .Y(_05369_));
 sg13g2_nand2b_1 _14380_ (.Y(_05370_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][6] ));
 sg13g2_nand2b_1 _14381_ (.Y(_05371_),
    .B(_05370_),
    .A_N(_05369_));
 sg13g2_o21ai_1 _14382_ (.B1(_05366_),
    .Y(_05372_),
    .A1(_05365_),
    .A2(_05367_));
 sg13g2_xnor2_1 _14383_ (.Y(_00656_),
    .A(_05371_),
    .B(_05372_));
 sg13g2_a21oi_1 _14384_ (.A1(_05370_),
    .A2(_05372_),
    .Y(_05373_),
    .B1(_05369_));
 sg13g2_xnor2_1 _14385_ (.Y(_05374_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][7] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nand2b_1 _14386_ (.Y(_05375_),
    .B(_05374_),
    .A_N(_05373_));
 sg13g2_xnor2_1 _14387_ (.Y(_00657_),
    .A(_05373_),
    .B(_05374_));
 sg13g2_o21ai_1 _14388_ (.B1(_05375_),
    .Y(_05376_),
    .A1(_02424_),
    .A2(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _14389_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][8] ),
    .Y(_05377_));
 sg13g2_nand2b_1 _14390_ (.Y(_05378_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][8] ));
 sg13g2_nand2b_1 _14391_ (.Y(_05379_),
    .B(_05378_),
    .A_N(_05377_));
 sg13g2_xnor2_1 _14392_ (.Y(_00658_),
    .A(_05376_),
    .B(_05379_));
 sg13g2_a21oi_2 _14393_ (.B1(_05377_),
    .Y(_05380_),
    .A2(_05378_),
    .A1(_05376_));
 sg13g2_nor2b_1 _14394_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][9] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[9] ),
    .Y(_05381_));
 sg13g2_nand2b_1 _14395_ (.Y(_05382_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][9] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _14396_ (.A(_05381_),
    .B_N(_05382_),
    .Y(_05383_));
 sg13g2_xnor2_1 _14397_ (.Y(_00659_),
    .A(_05380_),
    .B(_05383_));
 sg13g2_nor2b_1 _14398_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][10] ),
    .Y(_05384_));
 sg13g2_nand2b_1 _14399_ (.Y(_05385_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][10] ));
 sg13g2_nand2b_1 _14400_ (.Y(_05386_),
    .B(_05385_),
    .A_N(_05384_));
 sg13g2_a21oi_2 _14401_ (.B1(_05381_),
    .Y(_05387_),
    .A2(_05382_),
    .A1(_05380_));
 sg13g2_xnor2_1 _14402_ (.Y(_00642_),
    .A(_05386_),
    .B(_05387_));
 sg13g2_a21oi_2 _14403_ (.B1(_05384_),
    .Y(_05388_),
    .A2(_05387_),
    .A1(_05385_));
 sg13g2_nand2b_1 _14404_ (.Y(_05389_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][11] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _14405_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][11] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[11] ),
    .Y(_05390_));
 sg13g2_xnor2_1 _14406_ (.Y(_05391_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][11] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_xnor2_1 _14407_ (.Y(_00643_),
    .A(_05388_),
    .B(_05391_));
 sg13g2_nor2b_1 _14408_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][12] ),
    .Y(_05392_));
 sg13g2_nand2b_1 _14409_ (.Y(_05393_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][12] ));
 sg13g2_nand2b_1 _14410_ (.Y(_05394_),
    .B(_05393_),
    .A_N(_05392_));
 sg13g2_a21oi_2 _14411_ (.B1(_05390_),
    .Y(_05395_),
    .A2(_05389_),
    .A1(_05388_));
 sg13g2_xnor2_1 _14412_ (.Y(_00644_),
    .A(_05394_),
    .B(_05395_));
 sg13g2_a21oi_2 _14413_ (.B1(_05392_),
    .Y(_05396_),
    .A2(_05395_),
    .A1(_05393_));
 sg13g2_nand2b_1 _14414_ (.Y(_05397_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][13] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _14415_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][13] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[13] ),
    .Y(_05398_));
 sg13g2_xnor2_1 _14416_ (.Y(_05399_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][13] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_xnor2_1 _14417_ (.Y(_00645_),
    .A(_05396_),
    .B(_05399_));
 sg13g2_nor2b_1 _14418_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][14] ),
    .Y(_05400_));
 sg13g2_nand2b_1 _14419_ (.Y(_05401_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][14] ));
 sg13g2_nand2b_1 _14420_ (.Y(_05402_),
    .B(_05401_),
    .A_N(_05400_));
 sg13g2_a21oi_1 _14421_ (.A1(_05396_),
    .A2(_05397_),
    .Y(_05403_),
    .B1(_05398_));
 sg13g2_xnor2_1 _14422_ (.Y(_00646_),
    .A(_05402_),
    .B(_05403_));
 sg13g2_a21oi_1 _14423_ (.A1(_05401_),
    .A2(_05403_),
    .Y(_05404_),
    .B1(_05400_));
 sg13g2_nor2b_1 _14424_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][15] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[15] ),
    .Y(_05405_));
 sg13g2_nand2b_1 _14425_ (.Y(_05406_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][15] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _14426_ (.A(_05405_),
    .B_N(_05406_),
    .Y(_05407_));
 sg13g2_xnor2_1 _14427_ (.Y(_00647_),
    .A(_05404_),
    .B(_05407_));
 sg13g2_xor2_1 _14428_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][16] ),
    .X(_05408_));
 sg13g2_a21oi_1 _14429_ (.A1(_05404_),
    .A2(_05406_),
    .Y(_05409_),
    .B1(_05405_));
 sg13g2_nor2b_1 _14430_ (.A(_05408_),
    .B_N(_05409_),
    .Y(_05410_));
 sg13g2_xnor2_1 _14431_ (.Y(_00648_),
    .A(_05408_),
    .B(_05409_));
 sg13g2_a21oi_2 _14432_ (.B1(_05410_),
    .Y(_05411_),
    .A2(_02425_),
    .A1(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][16] ));
 sg13g2_nand2b_1 _14433_ (.Y(_05412_),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][17] ),
    .A_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _14434_ (.A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][17] ),
    .B_N(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[17] ),
    .Y(_05413_));
 sg13g2_xnor2_1 _14435_ (.Y(_05414_),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][17] ),
    .B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _14436_ (.Y(_00649_),
    .A(_05411_),
    .B(_05414_));
 sg13g2_o21ai_1 _14437_ (.B1(_05412_),
    .Y(_05415_),
    .A1(_05411_),
    .A2(_05413_));
 sg13g2_xor2_1 _14438_ (.B(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][18] ),
    .X(_05416_));
 sg13g2_xnor2_1 _14439_ (.Y(_00650_),
    .A(_05415_),
    .B(_05416_));
 sg13g2_and2_1 _14440_ (.A(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.u_mux_shift.sum_res ),
    .B(net4932),
    .X(_00255_));
 sg13g2_nand2_1 _14441_ (.Y(_05417_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[0] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_xor2_1 _14442_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[0] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[0] ),
    .X(_00791_));
 sg13g2_nand2_1 _14443_ (.Y(_05418_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[1] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_nor2_1 _14444_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[1] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[1] ),
    .Y(_05419_));
 sg13g2_xor2_1 _14445_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[1] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[1] ),
    .X(_05420_));
 sg13g2_xnor2_1 _14446_ (.Y(_00801_),
    .A(_05417_),
    .B(_05420_));
 sg13g2_o21ai_1 _14447_ (.B1(_05418_),
    .Y(_05421_),
    .A1(_05417_),
    .A2(_05419_));
 sg13g2_xnor2_1 _14448_ (.Y(_05422_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[2] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_nor2b_1 _14449_ (.A(_05422_),
    .B_N(_05421_),
    .Y(_05423_));
 sg13g2_xnor2_1 _14450_ (.Y(_00802_),
    .A(_05421_),
    .B(_05422_));
 sg13g2_a21o_1 _14451_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[2] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[2] ),
    .B1(_05423_),
    .X(_05424_));
 sg13g2_xnor2_1 _14452_ (.Y(_05425_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[3] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_nor2b_1 _14453_ (.A(_05425_),
    .B_N(_05424_),
    .Y(_05426_));
 sg13g2_xnor2_1 _14454_ (.Y(_00803_),
    .A(_05424_),
    .B(_05425_));
 sg13g2_a21o_1 _14455_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[3] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[3] ),
    .B1(_05426_),
    .X(_05427_));
 sg13g2_xnor2_1 _14456_ (.Y(_05428_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[4] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_nor2b_1 _14457_ (.A(_05428_),
    .B_N(_05427_),
    .Y(_05429_));
 sg13g2_xnor2_1 _14458_ (.Y(_00804_),
    .A(_05427_),
    .B(_05428_));
 sg13g2_a21o_1 _14459_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[4] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[4] ),
    .B1(_05429_),
    .X(_05430_));
 sg13g2_nand2_1 _14460_ (.Y(_05431_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[5] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_xnor2_1 _14461_ (.Y(_05432_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[5] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_xnor2_1 _14462_ (.Y(_00805_),
    .A(_05430_),
    .B(_05432_));
 sg13g2_xnor2_1 _14463_ (.Y(_05433_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[6] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_o21ai_1 _14464_ (.B1(_05430_),
    .Y(_05434_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[5] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_a21oi_1 _14465_ (.A1(_05431_),
    .A2(_05434_),
    .Y(_05435_),
    .B1(_05433_));
 sg13g2_nand3_1 _14466_ (.B(_05433_),
    .C(_05434_),
    .A(_05431_),
    .Y(_05436_));
 sg13g2_nor2b_1 _14467_ (.A(_05435_),
    .B_N(_05436_),
    .Y(_00806_));
 sg13g2_a21oi_1 _14468_ (.A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[6] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[6] ),
    .Y(_05437_),
    .B1(_05435_));
 sg13g2_nand2_1 _14469_ (.Y(_05438_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[7] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_nor2_1 _14470_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[7] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[7] ),
    .Y(_05439_));
 sg13g2_xor2_1 _14471_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[7] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[7] ),
    .X(_05440_));
 sg13g2_xnor2_1 _14472_ (.Y(_00807_),
    .A(_05437_),
    .B(_05440_));
 sg13g2_o21ai_1 _14473_ (.B1(_05438_),
    .Y(_05441_),
    .A1(_05437_),
    .A2(_05439_));
 sg13g2_xnor2_1 _14474_ (.Y(_05442_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[8] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_nor2b_1 _14475_ (.A(_05442_),
    .B_N(_05441_),
    .Y(_05443_));
 sg13g2_xnor2_1 _14476_ (.Y(_00808_),
    .A(_05441_),
    .B(_05442_));
 sg13g2_a21o_1 _14477_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[8] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[8] ),
    .B1(_05443_),
    .X(_05444_));
 sg13g2_xnor2_1 _14478_ (.Y(_05445_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[9] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_xnor2_1 _14479_ (.Y(_00809_),
    .A(_05444_),
    .B(_05445_));
 sg13g2_nand2_1 _14480_ (.Y(_05446_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[10] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_nor2_1 _14481_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[10] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[10] ),
    .Y(_05447_));
 sg13g2_xor2_1 _14482_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[10] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[10] ),
    .X(_05448_));
 sg13g2_a21o_1 _14483_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[9] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[9] ),
    .B1(_05444_),
    .X(_05449_));
 sg13g2_o21ai_1 _14484_ (.B1(_05449_),
    .Y(_05450_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[9] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_xnor2_1 _14485_ (.Y(_00792_),
    .A(_05448_),
    .B(_05450_));
 sg13g2_o21ai_1 _14486_ (.B1(_05446_),
    .Y(_05451_),
    .A1(_05447_),
    .A2(_05450_));
 sg13g2_xnor2_1 _14487_ (.Y(_05452_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[11] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_xnor2_1 _14488_ (.Y(_00793_),
    .A(_05451_),
    .B(_05452_));
 sg13g2_nand2_1 _14489_ (.Y(_05453_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[12] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_nor2_1 _14490_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[12] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[12] ),
    .Y(_05454_));
 sg13g2_xor2_1 _14491_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[12] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[12] ),
    .X(_05455_));
 sg13g2_a21o_1 _14492_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[11] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[11] ),
    .B1(_05451_),
    .X(_05456_));
 sg13g2_o21ai_1 _14493_ (.B1(_05456_),
    .Y(_05457_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[11] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_xnor2_1 _14494_ (.Y(_00794_),
    .A(_05455_),
    .B(_05457_));
 sg13g2_o21ai_1 _14495_ (.B1(_05453_),
    .Y(_05458_),
    .A1(_05454_),
    .A2(_05457_));
 sg13g2_xnor2_1 _14496_ (.Y(_05459_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[13] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_xnor2_1 _14497_ (.Y(_00795_),
    .A(_05458_),
    .B(_05459_));
 sg13g2_xor2_1 _14498_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[14] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[14] ),
    .X(_05460_));
 sg13g2_a21o_1 _14499_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[13] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[13] ),
    .B1(_05458_),
    .X(_05461_));
 sg13g2_o21ai_1 _14500_ (.B1(_05461_),
    .Y(_05462_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[13] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_nor2b_1 _14501_ (.A(_05462_),
    .B_N(_05460_),
    .Y(_05463_));
 sg13g2_xnor2_1 _14502_ (.Y(_00796_),
    .A(_05460_),
    .B(_05462_));
 sg13g2_a21o_1 _14503_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[14] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[14] ),
    .B1(_05463_),
    .X(_05464_));
 sg13g2_nand2_1 _14504_ (.Y(_05465_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[15] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_xnor2_1 _14505_ (.Y(_05466_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[15] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_xnor2_1 _14506_ (.Y(_00797_),
    .A(_05464_),
    .B(_05466_));
 sg13g2_nand2_1 _14507_ (.Y(_05467_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[16] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_xor2_1 _14508_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[16] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[16] ),
    .X(_05468_));
 sg13g2_o21ai_1 _14509_ (.B1(_05464_),
    .Y(_05469_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[15] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_nand2_1 _14510_ (.Y(_05470_),
    .A(_05465_),
    .B(_05469_));
 sg13g2_nand2_1 _14511_ (.Y(_05471_),
    .A(_05468_),
    .B(_05470_));
 sg13g2_xor2_1 _14512_ (.B(_05470_),
    .A(_05468_),
    .X(_00798_));
 sg13g2_xnor2_1 _14513_ (.Y(_05472_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[17] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_a21oi_1 _14514_ (.A1(_05467_),
    .A2(_05471_),
    .Y(_05473_),
    .B1(_05472_));
 sg13g2_nand3_1 _14515_ (.B(_05471_),
    .C(_05472_),
    .A(_05467_),
    .Y(_05474_));
 sg13g2_nor2b_1 _14516_ (.A(_05473_),
    .B_N(_05474_),
    .Y(_00799_));
 sg13g2_a21oi_1 _14517_ (.A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[17] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[17] ),
    .Y(_05475_),
    .B1(_05473_));
 sg13g2_xor2_1 _14518_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[18] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[18] ),
    .X(_05476_));
 sg13g2_xnor2_1 _14519_ (.Y(_00800_),
    .A(_05475_),
    .B(_05476_));
 sg13g2_nor2b_1 _14520_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][1] ),
    .Y(_05477_));
 sg13g2_xnor2_1 _14521_ (.Y(_05478_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][1] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _14522_ (.B(_05478_),
    .A(_02513_),
    .X(_00820_));
 sg13g2_a21oi_1 _14523_ (.A1(_02513_),
    .A2(_05478_),
    .Y(_05479_),
    .B1(_05477_));
 sg13g2_xnor2_1 _14524_ (.Y(_05480_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][2] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _14525_ (.A(_05479_),
    .B_N(_05480_),
    .Y(_05481_));
 sg13g2_xnor2_1 _14526_ (.Y(_00821_),
    .A(_05479_),
    .B(_05480_));
 sg13g2_a21oi_1 _14527_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][2] ),
    .A2(_02426_),
    .Y(_05482_),
    .B1(_05481_));
 sg13g2_xnor2_1 _14528_ (.Y(_05483_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][3] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _14529_ (.A(_05482_),
    .B_N(_05483_),
    .Y(_05484_));
 sg13g2_xnor2_1 _14530_ (.Y(_00822_),
    .A(_05482_),
    .B(_05483_));
 sg13g2_a21oi_1 _14531_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][3] ),
    .A2(_02427_),
    .Y(_05485_),
    .B1(_05484_));
 sg13g2_xnor2_1 _14532_ (.Y(_05486_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][4] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _14533_ (.A(_05485_),
    .B_N(_05486_),
    .Y(_05487_));
 sg13g2_xnor2_1 _14534_ (.Y(_00823_),
    .A(_05485_),
    .B(_05486_));
 sg13g2_a21oi_1 _14535_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][4] ),
    .A2(_02428_),
    .Y(_05488_),
    .B1(_05487_));
 sg13g2_xnor2_1 _14536_ (.Y(_05489_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][5] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _14537_ (.A(_05488_),
    .B_N(_05489_),
    .Y(_05490_));
 sg13g2_xnor2_1 _14538_ (.Y(_00824_),
    .A(_05488_),
    .B(_05489_));
 sg13g2_a21oi_1 _14539_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][5] ),
    .A2(_02429_),
    .Y(_05491_),
    .B1(_05490_));
 sg13g2_xnor2_1 _14540_ (.Y(_05492_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][6] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_nor2b_1 _14541_ (.A(_05491_),
    .B_N(_05492_),
    .Y(_05493_));
 sg13g2_xnor2_1 _14542_ (.Y(_00825_),
    .A(_05491_),
    .B(_05492_));
 sg13g2_a21oi_1 _14543_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][6] ),
    .A2(_02430_),
    .Y(_05494_),
    .B1(_05493_));
 sg13g2_xnor2_1 _14544_ (.Y(_05495_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][7] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _14545_ (.A(_05494_),
    .B_N(_05495_),
    .Y(_05496_));
 sg13g2_xnor2_1 _14546_ (.Y(_00826_),
    .A(_05494_),
    .B(_05495_));
 sg13g2_a21oi_1 _14547_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][7] ),
    .A2(_02431_),
    .Y(_05497_),
    .B1(_05496_));
 sg13g2_xnor2_1 _14548_ (.Y(_05498_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][8] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_nor2b_1 _14549_ (.A(_05497_),
    .B_N(_05498_),
    .Y(_05499_));
 sg13g2_xnor2_1 _14550_ (.Y(_00827_),
    .A(_05497_),
    .B(_05498_));
 sg13g2_a21oi_1 _14551_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][8] ),
    .A2(_02432_),
    .Y(_05500_),
    .B1(_05499_));
 sg13g2_nor2b_1 _14552_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][9] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[9] ),
    .Y(_05501_));
 sg13g2_nand2b_1 _14553_ (.Y(_05502_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][9] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _14554_ (.A(_05501_),
    .B_N(_05502_),
    .Y(_05503_));
 sg13g2_xnor2_1 _14555_ (.Y(_00828_),
    .A(_05500_),
    .B(_05503_));
 sg13g2_nor2b_1 _14556_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][10] ),
    .Y(_05504_));
 sg13g2_nand2b_1 _14557_ (.Y(_05505_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][10] ));
 sg13g2_nand2b_1 _14558_ (.Y(_05506_),
    .B(_05505_),
    .A_N(_05504_));
 sg13g2_a21oi_1 _14559_ (.A1(_05500_),
    .A2(_05502_),
    .Y(_05507_),
    .B1(_05501_));
 sg13g2_xnor2_1 _14560_ (.Y(_00811_),
    .A(_05506_),
    .B(_05507_));
 sg13g2_a21oi_1 _14561_ (.A1(_05505_),
    .A2(_05507_),
    .Y(_05508_),
    .B1(_05504_));
 sg13g2_nor2b_1 _14562_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][11] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[11] ),
    .Y(_05509_));
 sg13g2_nand2b_1 _14563_ (.Y(_05510_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][11] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _14564_ (.A(_05509_),
    .B_N(_05510_),
    .Y(_05511_));
 sg13g2_xnor2_1 _14565_ (.Y(_00812_),
    .A(_05508_),
    .B(_05511_));
 sg13g2_nor2b_1 _14566_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][12] ),
    .Y(_05512_));
 sg13g2_nand2b_1 _14567_ (.Y(_05513_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][12] ));
 sg13g2_nand2b_1 _14568_ (.Y(_05514_),
    .B(_05513_),
    .A_N(_05512_));
 sg13g2_a21oi_1 _14569_ (.A1(_05508_),
    .A2(_05510_),
    .Y(_05515_),
    .B1(_05509_));
 sg13g2_xnor2_1 _14570_ (.Y(_00813_),
    .A(_05514_),
    .B(_05515_));
 sg13g2_a21oi_1 _14571_ (.A1(_05513_),
    .A2(_05515_),
    .Y(_05516_),
    .B1(_05512_));
 sg13g2_nand2b_1 _14572_ (.Y(_05517_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][13] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _14573_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][13] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[13] ),
    .Y(_05518_));
 sg13g2_xnor2_1 _14574_ (.Y(_05519_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][13] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_xnor2_1 _14575_ (.Y(_00814_),
    .A(_05516_),
    .B(_05519_));
 sg13g2_nor2b_1 _14576_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][14] ),
    .Y(_05520_));
 sg13g2_nand2b_1 _14577_ (.Y(_05521_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][14] ));
 sg13g2_nand2b_1 _14578_ (.Y(_05522_),
    .B(_05521_),
    .A_N(_05520_));
 sg13g2_a21oi_1 _14579_ (.A1(_05516_),
    .A2(_05517_),
    .Y(_05523_),
    .B1(_05518_));
 sg13g2_xnor2_1 _14580_ (.Y(_00815_),
    .A(_05522_),
    .B(_05523_));
 sg13g2_a21oi_1 _14581_ (.A1(_05521_),
    .A2(_05523_),
    .Y(_05524_),
    .B1(_05520_));
 sg13g2_nor2b_1 _14582_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][15] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[15] ),
    .Y(_05525_));
 sg13g2_nand2b_1 _14583_ (.Y(_05526_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][15] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _14584_ (.A(_05525_),
    .B_N(_05526_),
    .Y(_05527_));
 sg13g2_xnor2_1 _14585_ (.Y(_00816_),
    .A(_05524_),
    .B(_05527_));
 sg13g2_xor2_1 _14586_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][16] ),
    .X(_05528_));
 sg13g2_a21oi_1 _14587_ (.A1(_05524_),
    .A2(_05526_),
    .Y(_05529_),
    .B1(_05525_));
 sg13g2_nor2b_1 _14588_ (.A(_05528_),
    .B_N(_05529_),
    .Y(_05530_));
 sg13g2_xnor2_1 _14589_ (.Y(_00817_),
    .A(_05528_),
    .B(_05529_));
 sg13g2_a21oi_1 _14590_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][16] ),
    .A2(_02433_),
    .Y(_05531_),
    .B1(_05530_));
 sg13g2_nand2b_1 _14591_ (.Y(_05532_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][17] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _14592_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][17] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[17] ),
    .Y(_05533_));
 sg13g2_xnor2_1 _14593_ (.Y(_05534_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][17] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _14594_ (.Y(_00818_),
    .A(_05531_),
    .B(_05534_));
 sg13g2_o21ai_1 _14595_ (.B1(_05532_),
    .Y(_05535_),
    .A1(_05531_),
    .A2(_05533_));
 sg13g2_xor2_1 _14596_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][18] ),
    .X(_05536_));
 sg13g2_xnor2_1 _14597_ (.Y(_00819_),
    .A(_05535_),
    .B(_05536_));
 sg13g2_nand2_1 _14598_ (.Y(_05537_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[0] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_xor2_1 _14599_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[0] ),
    .X(_00885_));
 sg13g2_nand2_1 _14600_ (.Y(_05538_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_nor2_1 _14601_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[1] ),
    .Y(_05539_));
 sg13g2_xor2_1 _14602_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[1] ),
    .X(_05540_));
 sg13g2_xnor2_1 _14603_ (.Y(_00895_),
    .A(_05537_),
    .B(_05540_));
 sg13g2_o21ai_1 _14604_ (.B1(_05538_),
    .Y(_05541_),
    .A1(_05537_),
    .A2(_05539_));
 sg13g2_xnor2_1 _14605_ (.Y(_05542_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[2] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_nor2b_1 _14606_ (.A(_05542_),
    .B_N(_05541_),
    .Y(_05543_));
 sg13g2_xnor2_1 _14607_ (.Y(_00896_),
    .A(_05541_),
    .B(_05542_));
 sg13g2_a21o_1 _14608_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[2] ),
    .B1(_05543_),
    .X(_05544_));
 sg13g2_xnor2_1 _14609_ (.Y(_05545_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[3] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_nor2b_1 _14610_ (.A(_05545_),
    .B_N(_05544_),
    .Y(_05546_));
 sg13g2_xnor2_1 _14611_ (.Y(_00897_),
    .A(_05544_),
    .B(_05545_));
 sg13g2_a21o_1 _14612_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[3] ),
    .B1(_05546_),
    .X(_05547_));
 sg13g2_xnor2_1 _14613_ (.Y(_05548_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[4] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_nor2b_1 _14614_ (.A(_05548_),
    .B_N(_05547_),
    .Y(_05549_));
 sg13g2_xnor2_1 _14615_ (.Y(_00898_),
    .A(_05547_),
    .B(_05548_));
 sg13g2_a21o_1 _14616_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[4] ),
    .B1(_05549_),
    .X(_05550_));
 sg13g2_nand2_1 _14617_ (.Y(_05551_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[5] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_xnor2_1 _14618_ (.Y(_05552_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[5] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_xnor2_1 _14619_ (.Y(_00899_),
    .A(_05550_),
    .B(_05552_));
 sg13g2_xnor2_1 _14620_ (.Y(_05553_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[6] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_o21ai_1 _14621_ (.B1(_05550_),
    .Y(_05554_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_a21oi_1 _14622_ (.A1(_05551_),
    .A2(_05554_),
    .Y(_05555_),
    .B1(_05553_));
 sg13g2_nand3_1 _14623_ (.B(_05553_),
    .C(_05554_),
    .A(_05551_),
    .Y(_05556_));
 sg13g2_nor2b_1 _14624_ (.A(_05555_),
    .B_N(_05556_),
    .Y(_00900_));
 sg13g2_a21oi_1 _14625_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[6] ),
    .Y(_05557_),
    .B1(_05555_));
 sg13g2_nand2_1 _14626_ (.Y(_05558_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[7] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_nor2_1 _14627_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[7] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[7] ),
    .Y(_05559_));
 sg13g2_xor2_1 _14628_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[7] ),
    .X(_05560_));
 sg13g2_xnor2_1 _14629_ (.Y(_00901_),
    .A(_05557_),
    .B(_05560_));
 sg13g2_o21ai_1 _14630_ (.B1(_05558_),
    .Y(_05561_),
    .A1(_05557_),
    .A2(_05559_));
 sg13g2_xnor2_1 _14631_ (.Y(_05562_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[8] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_nor2b_1 _14632_ (.A(_05562_),
    .B_N(_05561_),
    .Y(_05563_));
 sg13g2_xnor2_1 _14633_ (.Y(_00902_),
    .A(_05561_),
    .B(_05562_));
 sg13g2_a21o_1 _14634_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[8] ),
    .B1(_05563_),
    .X(_05564_));
 sg13g2_xnor2_1 _14635_ (.Y(_05565_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[9] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_xnor2_1 _14636_ (.Y(_00903_),
    .A(_05564_),
    .B(_05565_));
 sg13g2_nand2_1 _14637_ (.Y(_05566_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[10] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_nor2_1 _14638_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[10] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[10] ),
    .Y(_05567_));
 sg13g2_xor2_1 _14639_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[10] ),
    .X(_05568_));
 sg13g2_a21o_1 _14640_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[9] ),
    .B1(_05564_),
    .X(_05569_));
 sg13g2_o21ai_1 _14641_ (.B1(_05569_),
    .Y(_05570_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_xnor2_1 _14642_ (.Y(_00886_),
    .A(_05568_),
    .B(_05570_));
 sg13g2_o21ai_1 _14643_ (.B1(_05566_),
    .Y(_05571_),
    .A1(_05567_),
    .A2(_05570_));
 sg13g2_xnor2_1 _14644_ (.Y(_05572_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[11] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_xnor2_1 _14645_ (.Y(_00887_),
    .A(_05571_),
    .B(_05572_));
 sg13g2_nand2_1 _14646_ (.Y(_05573_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[12] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_nor2_1 _14647_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[12] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[12] ),
    .Y(_05574_));
 sg13g2_xor2_1 _14648_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[12] ),
    .X(_05575_));
 sg13g2_a21o_1 _14649_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[11] ),
    .B1(_05571_),
    .X(_05576_));
 sg13g2_o21ai_1 _14650_ (.B1(_05576_),
    .Y(_05577_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_xnor2_1 _14651_ (.Y(_00888_),
    .A(_05575_),
    .B(_05577_));
 sg13g2_o21ai_1 _14652_ (.B1(_05573_),
    .Y(_05578_),
    .A1(_05574_),
    .A2(_05577_));
 sg13g2_xnor2_1 _14653_ (.Y(_05579_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[13] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_xnor2_1 _14654_ (.Y(_00889_),
    .A(_05578_),
    .B(_05579_));
 sg13g2_xor2_1 _14655_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[14] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[14] ),
    .X(_05580_));
 sg13g2_a21o_1 _14656_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[13] ),
    .B1(_05578_),
    .X(_05581_));
 sg13g2_o21ai_1 _14657_ (.B1(_05581_),
    .Y(_05582_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_nor2b_1 _14658_ (.A(_05582_),
    .B_N(_05580_),
    .Y(_05583_));
 sg13g2_xnor2_1 _14659_ (.Y(_00890_),
    .A(_05580_),
    .B(_05582_));
 sg13g2_a21o_1 _14660_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[14] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[14] ),
    .B1(_05583_),
    .X(_05584_));
 sg13g2_nand2_1 _14661_ (.Y(_05585_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_xnor2_1 _14662_ (.Y(_05586_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_xnor2_1 _14663_ (.Y(_00891_),
    .A(_05584_),
    .B(_05586_));
 sg13g2_nand2_1 _14664_ (.Y(_05587_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[16] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_xor2_1 _14665_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[16] ),
    .X(_05588_));
 sg13g2_o21ai_1 _14666_ (.B1(_05584_),
    .Y(_05589_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[15] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_nand2_1 _14667_ (.Y(_05590_),
    .A(_05585_),
    .B(_05589_));
 sg13g2_nand2_1 _14668_ (.Y(_05591_),
    .A(_05588_),
    .B(_05590_));
 sg13g2_xor2_1 _14669_ (.B(_05590_),
    .A(_05588_),
    .X(_00892_));
 sg13g2_xnor2_1 _14670_ (.Y(_05592_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[17] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_a21oi_1 _14671_ (.A1(_05587_),
    .A2(_05591_),
    .Y(_05593_),
    .B1(_05592_));
 sg13g2_nand3_1 _14672_ (.B(_05591_),
    .C(_05592_),
    .A(_05587_),
    .Y(_05594_));
 sg13g2_nor2b_1 _14673_ (.A(_05593_),
    .B_N(_05594_),
    .Y(_00893_));
 sg13g2_a21oi_1 _14674_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[17] ),
    .Y(_05595_),
    .B1(_05593_));
 sg13g2_xor2_1 _14675_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[18] ),
    .X(_05596_));
 sg13g2_xnor2_1 _14676_ (.Y(_00894_),
    .A(_05595_),
    .B(_05596_));
 sg13g2_nand2b_1 _14677_ (.Y(_05597_),
    .B(net4974),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_nor2b_1 _14678_ (.A(net4974),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[1] ),
    .Y(_05598_));
 sg13g2_xnor2_1 _14679_ (.Y(_05599_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[1] ),
    .B(net4974));
 sg13g2_xnor2_1 _14680_ (.Y(_00951_),
    .A(_01188_),
    .B(_05599_));
 sg13g2_xnor2_1 _14681_ (.Y(_05600_),
    .A(net4974),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_o21ai_1 _14682_ (.B1(_05597_),
    .Y(_05601_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[0] ),
    .A2(_05598_));
 sg13g2_nor2b_1 _14683_ (.A(_05601_),
    .B_N(_05600_),
    .Y(_05602_));
 sg13g2_xnor2_1 _14684_ (.Y(_00952_),
    .A(_05600_),
    .B(_05601_));
 sg13g2_a21oi_1 _14685_ (.A1(net4941),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[2] ),
    .Y(_05603_),
    .B1(_05602_));
 sg13g2_nor2_1 _14686_ (.A(net4941),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[3] ),
    .Y(_05604_));
 sg13g2_nand2_1 _14687_ (.Y(_05605_),
    .A(net4941),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_nor2b_1 _14688_ (.A(_05604_),
    .B_N(_05605_),
    .Y(_05606_));
 sg13g2_xnor2_1 _14689_ (.Y(_00953_),
    .A(_05603_),
    .B(_05606_));
 sg13g2_xor2_1 _14690_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[4] ),
    .A(net4975),
    .X(_05607_));
 sg13g2_a21oi_1 _14691_ (.A1(_05603_),
    .A2(_05605_),
    .Y(_05608_),
    .B1(_05604_));
 sg13g2_nor2b_1 _14692_ (.A(_05607_),
    .B_N(_05608_),
    .Y(_05609_));
 sg13g2_xnor2_1 _14693_ (.Y(_00954_),
    .A(_05607_),
    .B(_05608_));
 sg13g2_xnor2_1 _14694_ (.Y(_05610_),
    .A(net4974),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_a21oi_1 _14695_ (.A1(net4940),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[4] ),
    .Y(_05611_),
    .B1(_05609_));
 sg13g2_xnor2_1 _14696_ (.Y(_00955_),
    .A(_05610_),
    .B(_05611_));
 sg13g2_o21ai_1 _14697_ (.B1(net4940),
    .Y(_05612_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[4] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_and2_1 _14698_ (.A(_05609_),
    .B(_05610_),
    .X(_05613_));
 sg13g2_nor2b_1 _14699_ (.A(_05613_),
    .B_N(_05612_),
    .Y(_05614_));
 sg13g2_nand2_1 _14700_ (.Y(_05615_),
    .A(net4941),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_nor2_1 _14701_ (.A(net4941),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[6] ),
    .Y(_05616_));
 sg13g2_xnor2_1 _14702_ (.Y(_05617_),
    .A(net4974),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_xnor2_1 _14703_ (.Y(_00956_),
    .A(_05614_),
    .B(_05617_));
 sg13g2_nand2b_1 _14704_ (.Y(_05618_),
    .B(net4974),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_xor2_1 _14705_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[7] ),
    .A(net4974),
    .X(_05619_));
 sg13g2_o21ai_1 _14706_ (.B1(_05615_),
    .Y(_05620_),
    .A1(_05614_),
    .A2(_05616_));
 sg13g2_xnor2_1 _14707_ (.Y(_00957_),
    .A(_05619_),
    .B(_05620_));
 sg13g2_xnor2_1 _14708_ (.Y(_05621_),
    .A(net4975),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_o21ai_1 _14709_ (.B1(net4940),
    .Y(_05622_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_nand3_1 _14710_ (.B(_05617_),
    .C(_05618_),
    .A(_05613_),
    .Y(_05623_));
 sg13g2_and3_1 _14711_ (.X(_05624_),
    .A(_05612_),
    .B(_05622_),
    .C(_05623_));
 sg13g2_nand2b_1 _14712_ (.Y(_05625_),
    .B(_05621_),
    .A_N(_05624_));
 sg13g2_xnor2_1 _14713_ (.Y(_00958_),
    .A(_05621_),
    .B(_05624_));
 sg13g2_xor2_1 _14714_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[9] ),
    .A(net4975),
    .X(_05626_));
 sg13g2_o21ai_1 _14715_ (.B1(_05625_),
    .Y(_05627_),
    .A1(net4975),
    .A2(_02435_));
 sg13g2_xnor2_1 _14716_ (.Y(_00959_),
    .A(_05626_),
    .B(_05627_));
 sg13g2_o21ai_1 _14717_ (.B1(net4940),
    .Y(_05628_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[8] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_or2_1 _14718_ (.X(_05629_),
    .B(_05626_),
    .A(_05625_));
 sg13g2_nand2_1 _14719_ (.Y(_05630_),
    .A(_05628_),
    .B(_05629_));
 sg13g2_nor2b_1 _14720_ (.A(net4973),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[10] ),
    .Y(_05631_));
 sg13g2_xnor2_1 _14721_ (.Y(_05632_),
    .A(net4973),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_xor2_1 _14722_ (.B(_05632_),
    .A(_05630_),
    .X(_00942_));
 sg13g2_xnor2_1 _14723_ (.Y(_05633_),
    .A(net4973),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_a21oi_1 _14724_ (.A1(_05630_),
    .A2(_05632_),
    .Y(_05634_),
    .B1(_05631_));
 sg13g2_xnor2_1 _14725_ (.Y(_00943_),
    .A(_05633_),
    .B(_05634_));
 sg13g2_xnor2_1 _14726_ (.Y(_05635_),
    .A(net4973),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_nor2b_1 _14727_ (.A(_05629_),
    .B_N(_05633_),
    .Y(_05636_));
 sg13g2_o21ai_1 _14728_ (.B1(net4940),
    .Y(_05637_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[10] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_nand2_1 _14729_ (.Y(_05638_),
    .A(_05628_),
    .B(_05637_));
 sg13g2_a21oi_1 _14730_ (.A1(_05632_),
    .A2(_05636_),
    .Y(_05639_),
    .B1(_05638_));
 sg13g2_nand2b_1 _14731_ (.Y(_05640_),
    .B(_05635_),
    .A_N(_05639_));
 sg13g2_xnor2_1 _14732_ (.Y(_00944_),
    .A(_05635_),
    .B(_05639_));
 sg13g2_xor2_1 _14733_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[13] ),
    .A(net4973),
    .X(_05641_));
 sg13g2_o21ai_1 _14734_ (.B1(_05640_),
    .Y(_05642_),
    .A1(net4973),
    .A2(_02436_));
 sg13g2_xnor2_1 _14735_ (.Y(_00945_),
    .A(_05641_),
    .B(_05642_));
 sg13g2_o21ai_1 _14736_ (.B1(net4940),
    .Y(_05643_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[12] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_o21ai_1 _14737_ (.B1(_05643_),
    .Y(_05644_),
    .A1(_05640_),
    .A2(_05641_));
 sg13g2_nor2b_1 _14738_ (.A(net4972),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[14] ),
    .Y(_05645_));
 sg13g2_nand2b_1 _14739_ (.Y(_05646_),
    .B(net4972),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_nand2b_1 _14740_ (.Y(_05647_),
    .B(_05646_),
    .A_N(_05645_));
 sg13g2_xnor2_1 _14741_ (.Y(_00946_),
    .A(_05644_),
    .B(_05647_));
 sg13g2_xnor2_1 _14742_ (.Y(_05648_),
    .A(net4972),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_a21oi_1 _14743_ (.A1(_05644_),
    .A2(_05646_),
    .Y(_05649_),
    .B1(_05645_));
 sg13g2_xnor2_1 _14744_ (.Y(_00947_),
    .A(_05648_),
    .B(_05649_));
 sg13g2_xnor2_1 _14745_ (.Y(_05650_),
    .A(net4972),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_nand2b_1 _14746_ (.Y(_05651_),
    .B(_05648_),
    .A_N(_05647_));
 sg13g2_nor2_1 _14747_ (.A(_05641_),
    .B(_05651_),
    .Y(_05652_));
 sg13g2_and4_1 _14748_ (.A(_05632_),
    .B(_05635_),
    .C(_05636_),
    .D(_05652_),
    .X(_05653_));
 sg13g2_o21ai_1 _14749_ (.B1(net4940),
    .Y(_05654_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand2_1 _14750_ (.Y(_05655_),
    .A(_05643_),
    .B(_05654_));
 sg13g2_nor3_2 _14751_ (.A(_05638_),
    .B(_05653_),
    .C(_05655_),
    .Y(_05656_));
 sg13g2_nand2b_1 _14752_ (.Y(_05657_),
    .B(_05650_),
    .A_N(_05656_));
 sg13g2_xnor2_1 _14753_ (.Y(_00948_),
    .A(_05650_),
    .B(_05656_));
 sg13g2_xor2_1 _14754_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[17] ),
    .A(net4972),
    .X(_05658_));
 sg13g2_o21ai_1 _14755_ (.B1(_05657_),
    .Y(_05659_),
    .A1(net4972),
    .A2(_02437_));
 sg13g2_xnor2_1 _14756_ (.Y(_00949_),
    .A(_05658_),
    .B(_05659_));
 sg13g2_o21ai_1 _14757_ (.B1(net4940),
    .Y(_05660_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[16] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_o21ai_1 _14758_ (.B1(_05660_),
    .Y(_05661_),
    .A1(_05657_),
    .A2(_05658_));
 sg13g2_xor2_1 _14759_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[18] ),
    .A(net4972),
    .X(_05662_));
 sg13g2_xnor2_1 _14760_ (.Y(_00950_),
    .A(_05661_),
    .B(_05662_));
 sg13g2_nor2b_1 _14761_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][1] ),
    .Y(_05663_));
 sg13g2_xnor2_1 _14762_ (.Y(_05664_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][1] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _14763_ (.B(_05664_),
    .A(_02520_),
    .X(_00839_));
 sg13g2_a21oi_1 _14764_ (.A1(_02520_),
    .A2(_05664_),
    .Y(_05665_),
    .B1(_05663_));
 sg13g2_xnor2_1 _14765_ (.Y(_05666_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][2] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _14766_ (.A(_05665_),
    .B_N(_05666_),
    .Y(_05667_));
 sg13g2_xnor2_1 _14767_ (.Y(_00840_),
    .A(_05665_),
    .B(_05666_));
 sg13g2_a21oi_1 _14768_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][2] ),
    .A2(_02438_),
    .Y(_05668_),
    .B1(_05667_));
 sg13g2_xnor2_1 _14769_ (.Y(_05669_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][3] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _14770_ (.A(_05668_),
    .B_N(_05669_),
    .Y(_05670_));
 sg13g2_xnor2_1 _14771_ (.Y(_00841_),
    .A(_05668_),
    .B(_05669_));
 sg13g2_a21oi_1 _14772_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][3] ),
    .A2(_02439_),
    .Y(_05671_),
    .B1(_05670_));
 sg13g2_xnor2_1 _14773_ (.Y(_05672_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][4] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _14774_ (.A(_05671_),
    .B_N(_05672_),
    .Y(_05673_));
 sg13g2_xnor2_1 _14775_ (.Y(_00842_),
    .A(_05671_),
    .B(_05672_));
 sg13g2_a21oi_1 _14776_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][4] ),
    .A2(_02440_),
    .Y(_05674_),
    .B1(_05673_));
 sg13g2_xnor2_1 _14777_ (.Y(_05675_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][5] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _14778_ (.A(_05674_),
    .B_N(_05675_),
    .Y(_05676_));
 sg13g2_xnor2_1 _14779_ (.Y(_00843_),
    .A(_05674_),
    .B(_05675_));
 sg13g2_a21oi_1 _14780_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][5] ),
    .A2(_02441_),
    .Y(_05677_),
    .B1(_05676_));
 sg13g2_xnor2_1 _14781_ (.Y(_05678_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][6] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_nor2b_1 _14782_ (.A(_05677_),
    .B_N(_05678_),
    .Y(_05679_));
 sg13g2_xnor2_1 _14783_ (.Y(_00844_),
    .A(_05677_),
    .B(_05678_));
 sg13g2_a21oi_1 _14784_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][6] ),
    .A2(_02442_),
    .Y(_05680_),
    .B1(_05679_));
 sg13g2_xnor2_1 _14785_ (.Y(_05681_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][7] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _14786_ (.A(_05680_),
    .B_N(_05681_),
    .Y(_05682_));
 sg13g2_xnor2_1 _14787_ (.Y(_00845_),
    .A(_05680_),
    .B(_05681_));
 sg13g2_a21oi_1 _14788_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][7] ),
    .A2(_02443_),
    .Y(_05683_),
    .B1(_05682_));
 sg13g2_xnor2_1 _14789_ (.Y(_05684_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][8] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_nor2b_1 _14790_ (.A(_05683_),
    .B_N(_05684_),
    .Y(_05685_));
 sg13g2_xnor2_1 _14791_ (.Y(_00846_),
    .A(_05683_),
    .B(_05684_));
 sg13g2_a21oi_1 _14792_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][8] ),
    .A2(_02444_),
    .Y(_05686_),
    .B1(_05685_));
 sg13g2_nand2b_1 _14793_ (.Y(_05687_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][9] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _14794_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][9] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[9] ),
    .Y(_05688_));
 sg13g2_xnor2_1 _14795_ (.Y(_05689_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][9] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_xnor2_1 _14796_ (.Y(_00847_),
    .A(_05686_),
    .B(_05689_));
 sg13g2_nor2b_1 _14797_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][10] ),
    .Y(_05690_));
 sg13g2_nand2b_1 _14798_ (.Y(_05691_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][10] ));
 sg13g2_nand2b_1 _14799_ (.Y(_05692_),
    .B(_05691_),
    .A_N(_05690_));
 sg13g2_o21ai_1 _14800_ (.B1(_05687_),
    .Y(_05693_),
    .A1(_05686_),
    .A2(_05688_));
 sg13g2_xnor2_1 _14801_ (.Y(_00830_),
    .A(_05692_),
    .B(_05693_));
 sg13g2_a21oi_1 _14802_ (.A1(_05691_),
    .A2(_05693_),
    .Y(_05694_),
    .B1(_05690_));
 sg13g2_nand2b_1 _14803_ (.Y(_05695_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][11] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _14804_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][11] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[11] ),
    .Y(_05696_));
 sg13g2_xnor2_1 _14805_ (.Y(_05697_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][11] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_xnor2_1 _14806_ (.Y(_00831_),
    .A(_05694_),
    .B(_05697_));
 sg13g2_nor2b_1 _14807_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][12] ),
    .Y(_05698_));
 sg13g2_nand2b_1 _14808_ (.Y(_05699_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][12] ));
 sg13g2_nand2b_1 _14809_ (.Y(_05700_),
    .B(_05699_),
    .A_N(_05698_));
 sg13g2_o21ai_1 _14810_ (.B1(_05695_),
    .Y(_05701_),
    .A1(_05694_),
    .A2(_05696_));
 sg13g2_xnor2_1 _14811_ (.Y(_00832_),
    .A(_05700_),
    .B(_05701_));
 sg13g2_a21oi_1 _14812_ (.A1(_05699_),
    .A2(_05701_),
    .Y(_05702_),
    .B1(_05698_));
 sg13g2_nand2b_1 _14813_ (.Y(_05703_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][13] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _14814_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][13] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[13] ),
    .Y(_05704_));
 sg13g2_xnor2_1 _14815_ (.Y(_05705_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][13] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_xnor2_1 _14816_ (.Y(_00833_),
    .A(_05702_),
    .B(_05705_));
 sg13g2_nor2b_1 _14817_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][14] ),
    .Y(_05706_));
 sg13g2_nand2b_1 _14818_ (.Y(_05707_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][14] ));
 sg13g2_nand2b_1 _14819_ (.Y(_05708_),
    .B(_05707_),
    .A_N(_05706_));
 sg13g2_a21oi_1 _14820_ (.A1(_05702_),
    .A2(_05703_),
    .Y(_05709_),
    .B1(_05704_));
 sg13g2_xnor2_1 _14821_ (.Y(_00834_),
    .A(_05708_),
    .B(_05709_));
 sg13g2_a21oi_1 _14822_ (.A1(_05707_),
    .A2(_05709_),
    .Y(_05710_),
    .B1(_05706_));
 sg13g2_nor2b_1 _14823_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][15] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[15] ),
    .Y(_05711_));
 sg13g2_nand2b_1 _14824_ (.Y(_05712_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][15] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _14825_ (.A(_05711_),
    .B_N(_05712_),
    .Y(_05713_));
 sg13g2_xnor2_1 _14826_ (.Y(_00835_),
    .A(_05710_),
    .B(_05713_));
 sg13g2_xor2_1 _14827_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][16] ),
    .X(_05714_));
 sg13g2_a21oi_1 _14828_ (.A1(_05710_),
    .A2(_05712_),
    .Y(_05715_),
    .B1(_05711_));
 sg13g2_nor2b_1 _14829_ (.A(_05714_),
    .B_N(_05715_),
    .Y(_05716_));
 sg13g2_xnor2_1 _14830_ (.Y(_00836_),
    .A(_05714_),
    .B(_05715_));
 sg13g2_a21oi_1 _14831_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][16] ),
    .A2(_02445_),
    .Y(_05717_),
    .B1(_05716_));
 sg13g2_nand2b_1 _14832_ (.Y(_05718_),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][17] ),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _14833_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][17] ),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[17] ),
    .Y(_05719_));
 sg13g2_xnor2_1 _14834_ (.Y(_05720_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][17] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _14835_ (.Y(_00837_),
    .A(_05717_),
    .B(_05720_));
 sg13g2_o21ai_1 _14836_ (.B1(_05718_),
    .Y(_05721_),
    .A1(_05717_),
    .A2(_05719_));
 sg13g2_xor2_1 _14837_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][18] ),
    .X(_05722_));
 sg13g2_xnor2_1 _14838_ (.Y(_00838_),
    .A(_05721_),
    .B(_05722_));
 sg13g2_nand2b_1 _14839_ (.Y(_05723_),
    .B(net4983),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_nor2b_1 _14840_ (.A(net4983),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[1] ),
    .Y(_05724_));
 sg13g2_xnor2_1 _14841_ (.Y(_05725_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[1] ),
    .B(net4982));
 sg13g2_xnor2_1 _14842_ (.Y(_00857_),
    .A(_01189_),
    .B(_05725_));
 sg13g2_xnor2_1 _14843_ (.Y(_05726_),
    .A(net4982),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_o21ai_1 _14844_ (.B1(_05723_),
    .Y(_05727_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[0] ),
    .A2(_05724_));
 sg13g2_nor2b_1 _14845_ (.A(_05727_),
    .B_N(_05726_),
    .Y(_05728_));
 sg13g2_xnor2_1 _14846_ (.Y(_00858_),
    .A(_05726_),
    .B(_05727_));
 sg13g2_a21oi_1 _14847_ (.A1(net4939),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[2] ),
    .Y(_05729_),
    .B1(_05728_));
 sg13g2_nor2_1 _14848_ (.A(net4939),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[3] ),
    .Y(_05730_));
 sg13g2_nand2_1 _14849_ (.Y(_05731_),
    .A(net4939),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_nor2b_1 _14850_ (.A(_05730_),
    .B_N(_05731_),
    .Y(_05732_));
 sg13g2_xnor2_1 _14851_ (.Y(_00859_),
    .A(_05729_),
    .B(_05732_));
 sg13g2_xor2_1 _14852_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[4] ),
    .A(net4983),
    .X(_05733_));
 sg13g2_a21oi_1 _14853_ (.A1(_05729_),
    .A2(_05731_),
    .Y(_05734_),
    .B1(_05730_));
 sg13g2_nor2b_1 _14854_ (.A(_05733_),
    .B_N(_05734_),
    .Y(_05735_));
 sg13g2_xnor2_1 _14855_ (.Y(_00860_),
    .A(_05733_),
    .B(_05734_));
 sg13g2_xnor2_1 _14856_ (.Y(_05736_),
    .A(net4982),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_a21oi_1 _14857_ (.A1(net4939),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[4] ),
    .Y(_05737_),
    .B1(_05735_));
 sg13g2_xnor2_1 _14858_ (.Y(_00861_),
    .A(_05736_),
    .B(_05737_));
 sg13g2_o21ai_1 _14859_ (.B1(net4939),
    .Y(_05738_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[4] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_and2_1 _14860_ (.A(_05735_),
    .B(_05736_),
    .X(_05739_));
 sg13g2_nor2b_1 _14861_ (.A(_05739_),
    .B_N(_05738_),
    .Y(_05740_));
 sg13g2_nand2_1 _14862_ (.Y(_05741_),
    .A(net4938),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_nor2_1 _14863_ (.A(net4938),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[6] ),
    .Y(_05742_));
 sg13g2_xnor2_1 _14864_ (.Y(_05743_),
    .A(net4982),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_xnor2_1 _14865_ (.Y(_00862_),
    .A(_05740_),
    .B(_05743_));
 sg13g2_nand2b_1 _14866_ (.Y(_05744_),
    .B(net4982),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_xor2_1 _14867_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[7] ),
    .A(net4982),
    .X(_05745_));
 sg13g2_o21ai_1 _14868_ (.B1(_05741_),
    .Y(_05746_),
    .A1(_05740_),
    .A2(_05742_));
 sg13g2_xnor2_1 _14869_ (.Y(_00863_),
    .A(_05745_),
    .B(_05746_));
 sg13g2_xnor2_1 _14870_ (.Y(_05747_),
    .A(net4982),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_o21ai_1 _14871_ (.B1(net4938),
    .Y(_05748_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_nand3_1 _14872_ (.B(_05743_),
    .C(_05744_),
    .A(_05739_),
    .Y(_05749_));
 sg13g2_and3_1 _14873_ (.X(_05750_),
    .A(_05738_),
    .B(_05748_),
    .C(_05749_));
 sg13g2_nand2b_1 _14874_ (.Y(_05751_),
    .B(_05747_),
    .A_N(_05750_));
 sg13g2_xnor2_1 _14875_ (.Y(_00864_),
    .A(_05747_),
    .B(_05750_));
 sg13g2_xor2_1 _14876_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[9] ),
    .A(net4981),
    .X(_05752_));
 sg13g2_o21ai_1 _14877_ (.B1(_05751_),
    .Y(_05753_),
    .A1(net4981),
    .A2(_02447_));
 sg13g2_xnor2_1 _14878_ (.Y(_00865_),
    .A(_05752_),
    .B(_05753_));
 sg13g2_o21ai_1 _14879_ (.B1(net4938),
    .Y(_05754_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[8] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_or2_1 _14880_ (.X(_05755_),
    .B(_05752_),
    .A(_05751_));
 sg13g2_nand2_1 _14881_ (.Y(_05756_),
    .A(_05754_),
    .B(_05755_));
 sg13g2_nor2b_1 _14882_ (.A(net4981),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[10] ),
    .Y(_05757_));
 sg13g2_xnor2_1 _14883_ (.Y(_05758_),
    .A(net4981),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_xor2_1 _14884_ (.B(_05758_),
    .A(_05756_),
    .X(_00848_));
 sg13g2_xnor2_1 _14885_ (.Y(_05759_),
    .A(net4981),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_a21oi_1 _14886_ (.A1(_05756_),
    .A2(_05758_),
    .Y(_05760_),
    .B1(_05757_));
 sg13g2_xnor2_1 _14887_ (.Y(_00849_),
    .A(_05759_),
    .B(_05760_));
 sg13g2_xnor2_1 _14888_ (.Y(_05761_),
    .A(net4981),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_nor2b_1 _14889_ (.A(_05755_),
    .B_N(_05759_),
    .Y(_05762_));
 sg13g2_o21ai_1 _14890_ (.B1(net4938),
    .Y(_05763_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[10] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_nand2_1 _14891_ (.Y(_05764_),
    .A(_05754_),
    .B(_05763_));
 sg13g2_a21oi_1 _14892_ (.A1(_05758_),
    .A2(_05762_),
    .Y(_05765_),
    .B1(_05764_));
 sg13g2_nand2b_1 _14893_ (.Y(_05766_),
    .B(_05761_),
    .A_N(_05765_));
 sg13g2_xnor2_1 _14894_ (.Y(_00850_),
    .A(_05761_),
    .B(_05765_));
 sg13g2_xor2_1 _14895_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[13] ),
    .A(net4980),
    .X(_05767_));
 sg13g2_o21ai_1 _14896_ (.B1(_05766_),
    .Y(_05768_),
    .A1(net4980),
    .A2(_02448_));
 sg13g2_xnor2_1 _14897_ (.Y(_00851_),
    .A(_05767_),
    .B(_05768_));
 sg13g2_o21ai_1 _14898_ (.B1(net4938),
    .Y(_05769_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[12] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_o21ai_1 _14899_ (.B1(_05769_),
    .Y(_05770_),
    .A1(_05766_),
    .A2(_05767_));
 sg13g2_nor2b_1 _14900_ (.A(net4980),
    .B_N(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[14] ),
    .Y(_05771_));
 sg13g2_nand2b_1 _14901_ (.Y(_05772_),
    .B(net4980),
    .A_N(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_nand2b_1 _14902_ (.Y(_05773_),
    .B(_05772_),
    .A_N(_05771_));
 sg13g2_xnor2_1 _14903_ (.Y(_00852_),
    .A(_05770_),
    .B(_05773_));
 sg13g2_xnor2_1 _14904_ (.Y(_05774_),
    .A(net4981),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_a21oi_1 _14905_ (.A1(_05770_),
    .A2(_05772_),
    .Y(_05775_),
    .B1(_05771_));
 sg13g2_xnor2_1 _14906_ (.Y(_00853_),
    .A(_05774_),
    .B(_05775_));
 sg13g2_xnor2_1 _14907_ (.Y(_05776_),
    .A(net4980),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_nand2b_1 _14908_ (.Y(_05777_),
    .B(_05774_),
    .A_N(_05773_));
 sg13g2_nor2_1 _14909_ (.A(_05767_),
    .B(_05777_),
    .Y(_05778_));
 sg13g2_and4_1 _14910_ (.A(_05758_),
    .B(_05761_),
    .C(_05762_),
    .D(_05778_),
    .X(_05779_));
 sg13g2_o21ai_1 _14911_ (.B1(net4938),
    .Y(_05780_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand2_1 _14912_ (.Y(_05781_),
    .A(_05769_),
    .B(_05780_));
 sg13g2_nor3_2 _14913_ (.A(_05764_),
    .B(_05779_),
    .C(_05781_),
    .Y(_05782_));
 sg13g2_nand2b_1 _14914_ (.Y(_05783_),
    .B(_05776_),
    .A_N(_05782_));
 sg13g2_xnor2_1 _14915_ (.Y(_00854_),
    .A(_05776_),
    .B(_05782_));
 sg13g2_xor2_1 _14916_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[17] ),
    .A(net4980),
    .X(_05784_));
 sg13g2_o21ai_1 _14917_ (.B1(_05783_),
    .Y(_05785_),
    .A1(net4980),
    .A2(_02449_));
 sg13g2_xnor2_1 _14918_ (.Y(_00855_),
    .A(_05784_),
    .B(_05785_));
 sg13g2_o21ai_1 _14919_ (.B1(net4938),
    .Y(_05786_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[16] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_o21ai_1 _14920_ (.B1(_05786_),
    .Y(_05787_),
    .A1(_05783_),
    .A2(_05784_));
 sg13g2_xor2_1 _14921_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[18] ),
    .A(net4980),
    .X(_05788_));
 sg13g2_xnor2_1 _14922_ (.Y(_00856_),
    .A(_05787_),
    .B(_05788_));
 sg13g2_nand2_1 _14923_ (.Y(_05789_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[0] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_xor2_1 _14924_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[0] ),
    .X(_00960_));
 sg13g2_nand2_1 _14925_ (.Y(_05790_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_nor2_1 _14926_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[1] ),
    .Y(_05791_));
 sg13g2_xor2_1 _14927_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[1] ),
    .X(_05792_));
 sg13g2_xnor2_1 _14928_ (.Y(_00970_),
    .A(_05789_),
    .B(_05792_));
 sg13g2_o21ai_1 _14929_ (.B1(_05790_),
    .Y(_05793_),
    .A1(_05789_),
    .A2(_05791_));
 sg13g2_xnor2_1 _14930_ (.Y(_05794_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[2] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_nor2b_1 _14931_ (.A(_05794_),
    .B_N(_05793_),
    .Y(_05795_));
 sg13g2_xnor2_1 _14932_ (.Y(_00971_),
    .A(_05793_),
    .B(_05794_));
 sg13g2_a21o_1 _14933_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[2] ),
    .B1(_05795_),
    .X(_05796_));
 sg13g2_xnor2_1 _14934_ (.Y(_05797_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[3] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_nor2b_1 _14935_ (.A(_05797_),
    .B_N(_05796_),
    .Y(_05798_));
 sg13g2_xnor2_1 _14936_ (.Y(_00972_),
    .A(_05796_),
    .B(_05797_));
 sg13g2_a21o_1 _14937_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[3] ),
    .B1(_05798_),
    .X(_05799_));
 sg13g2_xnor2_1 _14938_ (.Y(_05800_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[4] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_nor2b_1 _14939_ (.A(_05800_),
    .B_N(_05799_),
    .Y(_05801_));
 sg13g2_xnor2_1 _14940_ (.Y(_00973_),
    .A(_05799_),
    .B(_05800_));
 sg13g2_a21o_1 _14941_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[4] ),
    .B1(_05801_),
    .X(_05802_));
 sg13g2_nand2_1 _14942_ (.Y(_05803_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _14943_ (.Y(_05804_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _14944_ (.Y(_00974_),
    .A(_05802_),
    .B(_05804_));
 sg13g2_xnor2_1 _14945_ (.Y(_05805_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[6] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_o21ai_1 _14946_ (.B1(_05802_),
    .Y(_05806_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_a21oi_1 _14947_ (.A1(_05803_),
    .A2(_05806_),
    .Y(_05807_),
    .B1(_05805_));
 sg13g2_nand3_1 _14948_ (.B(_05805_),
    .C(_05806_),
    .A(_05803_),
    .Y(_05808_));
 sg13g2_nor2b_1 _14949_ (.A(_05807_),
    .B_N(_05808_),
    .Y(_00975_));
 sg13g2_a21oi_2 _14950_ (.B1(_05807_),
    .Y(_05809_),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[6] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_nand2_1 _14951_ (.Y(_05810_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_nor2_1 _14952_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[7] ),
    .Y(_05811_));
 sg13g2_xor2_1 _14953_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[7] ),
    .X(_05812_));
 sg13g2_xnor2_1 _14954_ (.Y(_00976_),
    .A(_05809_),
    .B(_05812_));
 sg13g2_o21ai_1 _14955_ (.B1(_05810_),
    .Y(_05813_),
    .A1(_05809_),
    .A2(_05811_));
 sg13g2_xnor2_1 _14956_ (.Y(_05814_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[8] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_nor2b_1 _14957_ (.A(_05814_),
    .B_N(_05813_),
    .Y(_05815_));
 sg13g2_xnor2_1 _14958_ (.Y(_00977_),
    .A(_05813_),
    .B(_05814_));
 sg13g2_a21o_1 _14959_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[8] ),
    .B1(_05815_),
    .X(_05816_));
 sg13g2_xnor2_1 _14960_ (.Y(_05817_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[9] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _14961_ (.Y(_00978_),
    .A(_05816_),
    .B(_05817_));
 sg13g2_nand2_1 _14962_ (.Y(_05818_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_nor2_1 _14963_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[10] ),
    .Y(_05819_));
 sg13g2_xor2_1 _14964_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[10] ),
    .X(_05820_));
 sg13g2_a21o_1 _14965_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[9] ),
    .B1(_05816_),
    .X(_05821_));
 sg13g2_o21ai_1 _14966_ (.B1(_05821_),
    .Y(_05822_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _14967_ (.Y(_00961_),
    .A(_05820_),
    .B(_05822_));
 sg13g2_o21ai_1 _14968_ (.B1(_05818_),
    .Y(_05823_),
    .A1(_05819_),
    .A2(_05822_));
 sg13g2_xnor2_1 _14969_ (.Y(_05824_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[11] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _14970_ (.Y(_00962_),
    .A(_05823_),
    .B(_05824_));
 sg13g2_xor2_1 _14971_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[12] ),
    .X(_05825_));
 sg13g2_a21o_1 _14972_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[11] ),
    .B1(_05823_),
    .X(_05826_));
 sg13g2_o21ai_1 _14973_ (.B1(_05826_),
    .Y(_05827_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_nand2b_1 _14974_ (.Y(_05828_),
    .B(_05825_),
    .A_N(_05827_));
 sg13g2_xnor2_1 _14975_ (.Y(_00963_),
    .A(_05825_),
    .B(_05827_));
 sg13g2_o21ai_1 _14976_ (.B1(_05828_),
    .Y(_05829_),
    .A1(_02436_),
    .A2(_02450_));
 sg13g2_xnor2_1 _14977_ (.Y(_05830_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[13] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_xnor2_1 _14978_ (.Y(_00964_),
    .A(_05829_),
    .B(_05830_));
 sg13g2_xnor2_1 _14979_ (.Y(_05831_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[14] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_a21o_1 _14980_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[13] ),
    .B1(_05829_),
    .X(_05832_));
 sg13g2_o21ai_1 _14981_ (.B1(_05832_),
    .Y(_05833_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_nor2_1 _14982_ (.A(_05831_),
    .B(_05833_),
    .Y(_05834_));
 sg13g2_xor2_1 _14983_ (.B(_05833_),
    .A(_05831_),
    .X(_00965_));
 sg13g2_a21oi_1 _14984_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[14] ),
    .Y(_05835_),
    .B1(_05834_));
 sg13g2_nand2_1 _14985_ (.Y(_05836_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_nor2_1 _14986_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[15] ),
    .Y(_05837_));
 sg13g2_xor2_1 _14987_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[15] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[15] ),
    .X(_05838_));
 sg13g2_xnor2_1 _14988_ (.Y(_00966_),
    .A(_05835_),
    .B(_05838_));
 sg13g2_and2_1 _14989_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[16] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[16] ),
    .X(_05839_));
 sg13g2_xor2_1 _14990_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[16] ),
    .X(_05840_));
 sg13g2_o21ai_1 _14991_ (.B1(_05836_),
    .Y(_05841_),
    .A1(_05835_),
    .A2(_05837_));
 sg13g2_xor2_1 _14992_ (.B(_05841_),
    .A(_05840_),
    .X(_00967_));
 sg13g2_a21o_1 _14993_ (.A2(_05841_),
    .A1(_05840_),
    .B1(_05839_),
    .X(_05842_));
 sg13g2_xnor2_1 _14994_ (.Y(_05843_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[17] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xnor2_1 _14995_ (.Y(_00968_),
    .A(_05842_),
    .B(_05843_));
 sg13g2_a21o_1 _14996_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[17] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[17] ),
    .B1(_05842_),
    .X(_05844_));
 sg13g2_o21ai_1 _14997_ (.B1(_05844_),
    .Y(_05845_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xor2_1 _14998_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[18] ),
    .X(_05846_));
 sg13g2_xnor2_1 _14999_ (.Y(_00969_),
    .A(_05845_),
    .B(_05846_));
 sg13g2_nor2b_1 _15000_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][1] ),
    .Y(_05847_));
 sg13g2_xnor2_1 _15001_ (.Y(_05848_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][1] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _15002_ (.B(_05848_),
    .A(_02514_),
    .X(_00745_));
 sg13g2_a21oi_2 _15003_ (.B1(_05847_),
    .Y(_05849_),
    .A2(_05848_),
    .A1(_02514_));
 sg13g2_xnor2_1 _15004_ (.Y(_05850_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][2] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _15005_ (.A(_05849_),
    .B_N(_05850_),
    .Y(_05851_));
 sg13g2_xnor2_1 _15006_ (.Y(_00746_),
    .A(_05849_),
    .B(_05850_));
 sg13g2_a21oi_2 _15007_ (.B1(_05851_),
    .Y(_05852_),
    .A2(_02451_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][2] ));
 sg13g2_xnor2_1 _15008_ (.Y(_05853_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][3] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _15009_ (.A(_05852_),
    .B_N(_05853_),
    .Y(_05854_));
 sg13g2_xnor2_1 _15010_ (.Y(_00747_),
    .A(_05852_),
    .B(_05853_));
 sg13g2_a21oi_2 _15011_ (.B1(_05854_),
    .Y(_05855_),
    .A2(_02452_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][3] ));
 sg13g2_xnor2_1 _15012_ (.Y(_05856_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][4] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _15013_ (.A(_05855_),
    .B_N(_05856_),
    .Y(_05857_));
 sg13g2_xnor2_1 _15014_ (.Y(_00748_),
    .A(_05855_),
    .B(_05856_));
 sg13g2_a21oi_2 _15015_ (.B1(_05857_),
    .Y(_05858_),
    .A2(_02453_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][4] ));
 sg13g2_nand2b_1 _15016_ (.Y(_05859_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][5] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _15017_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][5] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[5] ),
    .Y(_05860_));
 sg13g2_xnor2_1 _15018_ (.Y(_05861_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][5] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_xnor2_1 _15019_ (.Y(_00749_),
    .A(_05858_),
    .B(_05861_));
 sg13g2_nor2b_1 _15020_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][6] ),
    .Y(_05862_));
 sg13g2_nand2b_1 _15021_ (.Y(_05863_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][6] ));
 sg13g2_nand2b_1 _15022_ (.Y(_05864_),
    .B(_05863_),
    .A_N(_05862_));
 sg13g2_o21ai_1 _15023_ (.B1(_05859_),
    .Y(_05865_),
    .A1(_05858_),
    .A2(_05860_));
 sg13g2_xnor2_1 _15024_ (.Y(_00750_),
    .A(_05864_),
    .B(_05865_));
 sg13g2_a21oi_1 _15025_ (.A1(_05863_),
    .A2(_05865_),
    .Y(_05866_),
    .B1(_05862_));
 sg13g2_xnor2_1 _15026_ (.Y(_05867_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][7] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nand2b_1 _15027_ (.Y(_05868_),
    .B(_05867_),
    .A_N(_05866_));
 sg13g2_xnor2_1 _15028_ (.Y(_00751_),
    .A(_05866_),
    .B(_05867_));
 sg13g2_o21ai_1 _15029_ (.B1(_05868_),
    .Y(_05869_),
    .A1(_02454_),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _15030_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][8] ),
    .Y(_05870_));
 sg13g2_nand2b_1 _15031_ (.Y(_05871_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][8] ));
 sg13g2_nand2b_1 _15032_ (.Y(_05872_),
    .B(_05871_),
    .A_N(_05870_));
 sg13g2_xnor2_1 _15033_ (.Y(_00752_),
    .A(_05869_),
    .B(_05872_));
 sg13g2_a21oi_2 _15034_ (.B1(_05870_),
    .Y(_05873_),
    .A2(_05871_),
    .A1(_05869_));
 sg13g2_nand2b_1 _15035_ (.Y(_05874_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][9] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _15036_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][9] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[9] ),
    .Y(_05875_));
 sg13g2_xnor2_1 _15037_ (.Y(_05876_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][9] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_xnor2_1 _15038_ (.Y(_00753_),
    .A(_05873_),
    .B(_05876_));
 sg13g2_nor2b_1 _15039_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][10] ),
    .Y(_05877_));
 sg13g2_nand2b_1 _15040_ (.Y(_05878_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][10] ));
 sg13g2_nand2b_1 _15041_ (.Y(_05879_),
    .B(_05878_),
    .A_N(_05877_));
 sg13g2_o21ai_1 _15042_ (.B1(_05874_),
    .Y(_05880_),
    .A1(_05873_),
    .A2(_05875_));
 sg13g2_xnor2_1 _15043_ (.Y(_00736_),
    .A(_05879_),
    .B(_05880_));
 sg13g2_a21oi_2 _15044_ (.B1(_05877_),
    .Y(_05881_),
    .A2(_05880_),
    .A1(_05878_));
 sg13g2_nand2b_1 _15045_ (.Y(_05882_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][11] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _15046_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][11] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[11] ),
    .Y(_05883_));
 sg13g2_xnor2_1 _15047_ (.Y(_05884_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][11] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_xnor2_1 _15048_ (.Y(_00737_),
    .A(_05881_),
    .B(_05884_));
 sg13g2_nor2b_1 _15049_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][12] ),
    .Y(_05885_));
 sg13g2_nand2b_1 _15050_ (.Y(_05886_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][12] ));
 sg13g2_nand2b_1 _15051_ (.Y(_05887_),
    .B(_05886_),
    .A_N(_05885_));
 sg13g2_o21ai_1 _15052_ (.B1(_05882_),
    .Y(_05888_),
    .A1(_05881_),
    .A2(_05883_));
 sg13g2_xnor2_1 _15053_ (.Y(_00738_),
    .A(_05887_),
    .B(_05888_));
 sg13g2_a21oi_2 _15054_ (.B1(_05885_),
    .Y(_05889_),
    .A2(_05888_),
    .A1(_05886_));
 sg13g2_nand2b_1 _15055_ (.Y(_05890_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][13] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _15056_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][13] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[13] ),
    .Y(_05891_));
 sg13g2_xnor2_1 _15057_ (.Y(_05892_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][13] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_xnor2_1 _15058_ (.Y(_00739_),
    .A(_05889_),
    .B(_05892_));
 sg13g2_nor2b_1 _15059_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][14] ),
    .Y(_05893_));
 sg13g2_nand2b_1 _15060_ (.Y(_05894_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][14] ));
 sg13g2_nand2b_1 _15061_ (.Y(_05895_),
    .B(_05894_),
    .A_N(_05893_));
 sg13g2_o21ai_1 _15062_ (.B1(_05890_),
    .Y(_05896_),
    .A1(_05889_),
    .A2(_05891_));
 sg13g2_xnor2_1 _15063_ (.Y(_00740_),
    .A(_05895_),
    .B(_05896_));
 sg13g2_a21oi_2 _15064_ (.B1(_05893_),
    .Y(_05897_),
    .A2(_05896_),
    .A1(_05894_));
 sg13g2_nand2b_1 _15065_ (.Y(_05898_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][15] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _15066_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][15] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[15] ),
    .Y(_05899_));
 sg13g2_xnor2_1 _15067_ (.Y(_05900_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][15] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_xnor2_1 _15068_ (.Y(_00741_),
    .A(_05897_),
    .B(_05900_));
 sg13g2_nor2b_1 _15069_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[16] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][16] ),
    .Y(_05901_));
 sg13g2_nand2b_1 _15070_ (.Y(_05902_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[16] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][16] ));
 sg13g2_nand2b_1 _15071_ (.Y(_05903_),
    .B(_05902_),
    .A_N(_05901_));
 sg13g2_o21ai_1 _15072_ (.B1(_05898_),
    .Y(_05904_),
    .A1(_05897_),
    .A2(_05899_));
 sg13g2_xnor2_1 _15073_ (.Y(_00742_),
    .A(_05903_),
    .B(_05904_));
 sg13g2_a21oi_2 _15074_ (.B1(_05901_),
    .Y(_05905_),
    .A2(_05904_),
    .A1(_05902_));
 sg13g2_nand2b_1 _15075_ (.Y(_05906_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][17] ),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _15076_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][17] ),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[17] ),
    .Y(_05907_));
 sg13g2_xnor2_1 _15077_ (.Y(_05908_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][17] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _15078_ (.Y(_00743_),
    .A(_05905_),
    .B(_05908_));
 sg13g2_o21ai_1 _15079_ (.B1(_05906_),
    .Y(_05909_),
    .A1(_05905_),
    .A2(_05907_));
 sg13g2_xor2_1 _15080_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][18] ),
    .X(_05910_));
 sg13g2_xnor2_1 _15081_ (.Y(_00744_),
    .A(_05909_),
    .B(_05910_));
 sg13g2_nand2b_1 _15082_ (.Y(_05911_),
    .B(net4953),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_nor2b_1 _15083_ (.A(net4952),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[1] ),
    .Y(_05912_));
 sg13g2_xnor2_1 _15084_ (.Y(_05913_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[1] ),
    .B(net4952));
 sg13g2_xnor2_1 _15085_ (.Y(_00763_),
    .A(_01190_),
    .B(_05913_));
 sg13g2_xnor2_1 _15086_ (.Y(_05914_),
    .A(net4952),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_o21ai_1 _15087_ (.B1(_05911_),
    .Y(_05915_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[0] ),
    .A2(_05912_));
 sg13g2_nor2b_1 _15088_ (.A(_05915_),
    .B_N(_05914_),
    .Y(_05916_));
 sg13g2_xnor2_1 _15089_ (.Y(_00764_),
    .A(_05914_),
    .B(_05915_));
 sg13g2_a21oi_1 _15090_ (.A1(net4936),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[2] ),
    .Y(_05917_),
    .B1(_05916_));
 sg13g2_nor2_1 _15091_ (.A(net4936),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[3] ),
    .Y(_05918_));
 sg13g2_nand2_1 _15092_ (.Y(_05919_),
    .A(net4936),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_nor2b_1 _15093_ (.A(_05918_),
    .B_N(_05919_),
    .Y(_05920_));
 sg13g2_xnor2_1 _15094_ (.Y(_00765_),
    .A(_05917_),
    .B(_05920_));
 sg13g2_xor2_1 _15095_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[4] ),
    .A(net4952),
    .X(_05921_));
 sg13g2_a21oi_1 _15096_ (.A1(_05917_),
    .A2(_05919_),
    .Y(_05922_),
    .B1(_05918_));
 sg13g2_nor2b_1 _15097_ (.A(_05921_),
    .B_N(_05922_),
    .Y(_05923_));
 sg13g2_xnor2_1 _15098_ (.Y(_00766_),
    .A(_05921_),
    .B(_05922_));
 sg13g2_xnor2_1 _15099_ (.Y(_05924_),
    .A(net4952),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_a21oi_1 _15100_ (.A1(net4936),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[4] ),
    .Y(_05925_),
    .B1(_05923_));
 sg13g2_xnor2_1 _15101_ (.Y(_00767_),
    .A(_05924_),
    .B(_05925_));
 sg13g2_o21ai_1 _15102_ (.B1(net4936),
    .Y(_05926_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[4] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_and2_1 _15103_ (.A(_05923_),
    .B(_05924_),
    .X(_05927_));
 sg13g2_nor2b_1 _15104_ (.A(_05927_),
    .B_N(_05926_),
    .Y(_05928_));
 sg13g2_nand2_1 _15105_ (.Y(_05929_),
    .A(net4937),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_nor2_1 _15106_ (.A(net4936),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[6] ),
    .Y(_05930_));
 sg13g2_xnor2_1 _15107_ (.Y(_05931_),
    .A(net4952),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_xnor2_1 _15108_ (.Y(_00768_),
    .A(_05928_),
    .B(_05931_));
 sg13g2_nand2b_1 _15109_ (.Y(_05932_),
    .B(net4952),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_xor2_1 _15110_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[7] ),
    .A(net4952),
    .X(_05933_));
 sg13g2_o21ai_1 _15111_ (.B1(_05929_),
    .Y(_05934_),
    .A1(_05928_),
    .A2(_05930_));
 sg13g2_xnor2_1 _15112_ (.Y(_00769_),
    .A(_05933_),
    .B(_05934_));
 sg13g2_xnor2_1 _15113_ (.Y(_05935_),
    .A(net4953),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_o21ai_1 _15114_ (.B1(net4936),
    .Y(_05936_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_nand3_1 _15115_ (.B(_05931_),
    .C(_05932_),
    .A(_05927_),
    .Y(_05937_));
 sg13g2_and3_1 _15116_ (.X(_05938_),
    .A(_05926_),
    .B(_05936_),
    .C(_05937_));
 sg13g2_nand2b_1 _15117_ (.Y(_05939_),
    .B(_05935_),
    .A_N(_05938_));
 sg13g2_xnor2_1 _15118_ (.Y(_00770_),
    .A(_05935_),
    .B(_05938_));
 sg13g2_xor2_1 _15119_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[9] ),
    .A(net4953),
    .X(_05940_));
 sg13g2_o21ai_1 _15120_ (.B1(_05939_),
    .Y(_05941_),
    .A1(net4953),
    .A2(_02456_));
 sg13g2_xnor2_1 _15121_ (.Y(_00771_),
    .A(_05940_),
    .B(_05941_));
 sg13g2_o21ai_1 _15122_ (.B1(net4936),
    .Y(_05942_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[8] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_or2_1 _15123_ (.X(_05943_),
    .B(_05940_),
    .A(_05939_));
 sg13g2_nand2_1 _15124_ (.Y(_05944_),
    .A(_05942_),
    .B(_05943_));
 sg13g2_nor2b_1 _15125_ (.A(net4951),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[10] ),
    .Y(_05945_));
 sg13g2_xnor2_1 _15126_ (.Y(_05946_),
    .A(net4951),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_xor2_1 _15127_ (.B(_05946_),
    .A(_05944_),
    .X(_00754_));
 sg13g2_xnor2_1 _15128_ (.Y(_05947_),
    .A(net4951),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_a21oi_1 _15129_ (.A1(_05944_),
    .A2(_05946_),
    .Y(_05948_),
    .B1(_05945_));
 sg13g2_xnor2_1 _15130_ (.Y(_00755_),
    .A(_05947_),
    .B(_05948_));
 sg13g2_xnor2_1 _15131_ (.Y(_05949_),
    .A(net4951),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_nor2b_1 _15132_ (.A(_05943_),
    .B_N(_05946_),
    .Y(_05950_));
 sg13g2_o21ai_1 _15133_ (.B1(net4937),
    .Y(_05951_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[10] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_nand2_1 _15134_ (.Y(_05952_),
    .A(_05942_),
    .B(_05951_));
 sg13g2_a21oi_1 _15135_ (.A1(_05947_),
    .A2(_05950_),
    .Y(_05953_),
    .B1(_05952_));
 sg13g2_nand2b_1 _15136_ (.Y(_05954_),
    .B(_05949_),
    .A_N(_05953_));
 sg13g2_xnor2_1 _15137_ (.Y(_00756_),
    .A(_05949_),
    .B(_05953_));
 sg13g2_xor2_1 _15138_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[13] ),
    .A(net4951),
    .X(_05955_));
 sg13g2_o21ai_1 _15139_ (.B1(_05954_),
    .Y(_05956_),
    .A1(net4950),
    .A2(_02457_));
 sg13g2_xnor2_1 _15140_ (.Y(_00757_),
    .A(_05955_),
    .B(_05956_));
 sg13g2_o21ai_1 _15141_ (.B1(net4937),
    .Y(_05957_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[12] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_o21ai_1 _15142_ (.B1(_05957_),
    .Y(_05958_),
    .A1(_05954_),
    .A2(_05955_));
 sg13g2_nor2b_1 _15143_ (.A(net4950),
    .B_N(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[14] ),
    .Y(_05959_));
 sg13g2_nand2b_1 _15144_ (.Y(_05960_),
    .B(net4950),
    .A_N(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_nand2b_1 _15145_ (.Y(_05961_),
    .B(_05960_),
    .A_N(_05959_));
 sg13g2_xnor2_1 _15146_ (.Y(_00758_),
    .A(_05958_),
    .B(_05961_));
 sg13g2_xnor2_1 _15147_ (.Y(_05962_),
    .A(net4950),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_a21oi_1 _15148_ (.A1(_05958_),
    .A2(_05960_),
    .Y(_05963_),
    .B1(_05959_));
 sg13g2_xnor2_1 _15149_ (.Y(_00759_),
    .A(_05962_),
    .B(_05963_));
 sg13g2_xnor2_1 _15150_ (.Y(_05964_),
    .A(net4950),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_nand2b_1 _15151_ (.Y(_05965_),
    .B(_05962_),
    .A_N(_05961_));
 sg13g2_nor2_1 _15152_ (.A(_05955_),
    .B(_05965_),
    .Y(_05966_));
 sg13g2_and4_1 _15153_ (.A(_05947_),
    .B(_05949_),
    .C(_05950_),
    .D(_05966_),
    .X(_05967_));
 sg13g2_o21ai_1 _15154_ (.B1(net4937),
    .Y(_05968_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand2_1 _15155_ (.Y(_05969_),
    .A(_05957_),
    .B(_05968_));
 sg13g2_nor3_2 _15156_ (.A(_05952_),
    .B(_05967_),
    .C(_05969_),
    .Y(_05970_));
 sg13g2_nand2b_1 _15157_ (.Y(_05971_),
    .B(_05964_),
    .A_N(_05970_));
 sg13g2_xnor2_1 _15158_ (.Y(_00760_),
    .A(_05964_),
    .B(_05970_));
 sg13g2_xor2_1 _15159_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[17] ),
    .A(net4950),
    .X(_05972_));
 sg13g2_o21ai_1 _15160_ (.B1(_05971_),
    .Y(_05973_),
    .A1(net4950),
    .A2(_02458_));
 sg13g2_xnor2_1 _15161_ (.Y(_00761_),
    .A(_05972_),
    .B(_05973_));
 sg13g2_o21ai_1 _15162_ (.B1(net4937),
    .Y(_05974_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[16] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_o21ai_1 _15163_ (.B1(_05974_),
    .Y(_05975_),
    .A1(_05971_),
    .A2(_05972_));
 sg13g2_xor2_1 _15164_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[18] ),
    .A(net4950),
    .X(_05976_));
 sg13g2_xnor2_1 _15165_ (.Y(_00762_),
    .A(_05975_),
    .B(_05976_));
 sg13g2_nand2_1 _15166_ (.Y(_05977_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[0] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_xor2_1 _15167_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[0] ),
    .X(_00866_));
 sg13g2_nand2_1 _15168_ (.Y(_05978_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_nor2_1 _15169_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[1] ),
    .Y(_05979_));
 sg13g2_xor2_1 _15170_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[1] ),
    .X(_05980_));
 sg13g2_xnor2_1 _15171_ (.Y(_00876_),
    .A(_05977_),
    .B(_05980_));
 sg13g2_o21ai_1 _15172_ (.B1(_05978_),
    .Y(_05981_),
    .A1(_05977_),
    .A2(_05979_));
 sg13g2_xnor2_1 _15173_ (.Y(_05982_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[2] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_nor2b_1 _15174_ (.A(_05982_),
    .B_N(_05981_),
    .Y(_05983_));
 sg13g2_xnor2_1 _15175_ (.Y(_00877_),
    .A(_05981_),
    .B(_05982_));
 sg13g2_a21o_1 _15176_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[2] ),
    .B1(_05983_),
    .X(_05984_));
 sg13g2_xnor2_1 _15177_ (.Y(_05985_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[3] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_nor2b_1 _15178_ (.A(_05985_),
    .B_N(_05984_),
    .Y(_05986_));
 sg13g2_xnor2_1 _15179_ (.Y(_00878_),
    .A(_05984_),
    .B(_05985_));
 sg13g2_a21o_1 _15180_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[3] ),
    .B1(_05986_),
    .X(_05987_));
 sg13g2_xnor2_1 _15181_ (.Y(_05988_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[4] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_nor2b_1 _15182_ (.A(_05988_),
    .B_N(_05987_),
    .Y(_05989_));
 sg13g2_xnor2_1 _15183_ (.Y(_00879_),
    .A(_05987_),
    .B(_05988_));
 sg13g2_a21o_1 _15184_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[4] ),
    .B1(_05989_),
    .X(_05990_));
 sg13g2_nand2_1 _15185_ (.Y(_05991_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _15186_ (.Y(_05992_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _15187_ (.Y(_00880_),
    .A(_05990_),
    .B(_05992_));
 sg13g2_xnor2_1 _15188_ (.Y(_05993_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[6] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_o21ai_1 _15189_ (.B1(_05990_),
    .Y(_05994_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_a21oi_1 _15190_ (.A1(_05991_),
    .A2(_05994_),
    .Y(_05995_),
    .B1(_05993_));
 sg13g2_nand3_1 _15191_ (.B(_05993_),
    .C(_05994_),
    .A(_05991_),
    .Y(_05996_));
 sg13g2_nor2b_1 _15192_ (.A(_05995_),
    .B_N(_05996_),
    .Y(_00881_));
 sg13g2_a21oi_1 _15193_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[6] ),
    .Y(_05997_),
    .B1(_05995_));
 sg13g2_nand2_1 _15194_ (.Y(_05998_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_nor2_1 _15195_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[7] ),
    .Y(_05999_));
 sg13g2_xor2_1 _15196_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[7] ),
    .X(_06000_));
 sg13g2_xnor2_1 _15197_ (.Y(_00882_),
    .A(_05997_),
    .B(_06000_));
 sg13g2_o21ai_1 _15198_ (.B1(_05998_),
    .Y(_06001_),
    .A1(_05997_),
    .A2(_05999_));
 sg13g2_xnor2_1 _15199_ (.Y(_06002_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[8] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_nor2b_1 _15200_ (.A(_06002_),
    .B_N(_06001_),
    .Y(_06003_));
 sg13g2_xnor2_1 _15201_ (.Y(_00883_),
    .A(_06001_),
    .B(_06002_));
 sg13g2_a21o_1 _15202_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[8] ),
    .B1(_06003_),
    .X(_06004_));
 sg13g2_xnor2_1 _15203_ (.Y(_06005_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[9] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _15204_ (.Y(_00884_),
    .A(_06004_),
    .B(_06005_));
 sg13g2_nand2_1 _15205_ (.Y(_06006_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_nor2_1 _15206_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[10] ),
    .Y(_06007_));
 sg13g2_xor2_1 _15207_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[10] ),
    .X(_06008_));
 sg13g2_a21o_1 _15208_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[9] ),
    .B1(_06004_),
    .X(_06009_));
 sg13g2_o21ai_1 _15209_ (.B1(_06009_),
    .Y(_06010_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _15210_ (.Y(_00867_),
    .A(_06008_),
    .B(_06010_));
 sg13g2_o21ai_1 _15211_ (.B1(_06006_),
    .Y(_06011_),
    .A1(_06007_),
    .A2(_06010_));
 sg13g2_xnor2_1 _15212_ (.Y(_06012_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[11] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _15213_ (.Y(_00868_),
    .A(_06011_),
    .B(_06012_));
 sg13g2_xor2_1 _15214_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[12] ),
    .X(_06013_));
 sg13g2_a21o_1 _15215_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[11] ),
    .B1(_06011_),
    .X(_06014_));
 sg13g2_o21ai_1 _15216_ (.B1(_06014_),
    .Y(_06015_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_nand2b_1 _15217_ (.Y(_06016_),
    .B(_06013_),
    .A_N(_06015_));
 sg13g2_xnor2_1 _15218_ (.Y(_00869_),
    .A(_06013_),
    .B(_06015_));
 sg13g2_o21ai_1 _15219_ (.B1(_06016_),
    .Y(_06017_),
    .A1(_02448_),
    .A2(_02459_));
 sg13g2_xnor2_1 _15220_ (.Y(_06018_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[13] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_xnor2_1 _15221_ (.Y(_00870_),
    .A(_06017_),
    .B(_06018_));
 sg13g2_xnor2_1 _15222_ (.Y(_06019_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[14] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_a21o_1 _15223_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[13] ),
    .B1(_06017_),
    .X(_06020_));
 sg13g2_o21ai_1 _15224_ (.B1(_06020_),
    .Y(_06021_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_nor2_1 _15225_ (.A(_06019_),
    .B(_06021_),
    .Y(_06022_));
 sg13g2_xor2_1 _15226_ (.B(_06021_),
    .A(_06019_),
    .X(_00871_));
 sg13g2_a21oi_1 _15227_ (.A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[14] ),
    .Y(_06023_),
    .B1(_06022_));
 sg13g2_nand2_1 _15228_ (.Y(_06024_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_nor2_1 _15229_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[15] ),
    .Y(_06025_));
 sg13g2_xor2_1 _15230_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[15] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[15] ),
    .X(_06026_));
 sg13g2_xnor2_1 _15231_ (.Y(_00872_),
    .A(_06023_),
    .B(_06026_));
 sg13g2_and2_1 _15232_ (.A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[16] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[16] ),
    .X(_06027_));
 sg13g2_xor2_1 _15233_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[16] ),
    .X(_06028_));
 sg13g2_o21ai_1 _15234_ (.B1(_06024_),
    .Y(_06029_),
    .A1(_06023_),
    .A2(_06025_));
 sg13g2_xor2_1 _15235_ (.B(_06029_),
    .A(_06028_),
    .X(_00873_));
 sg13g2_a21o_1 _15236_ (.A2(_06029_),
    .A1(_06028_),
    .B1(_06027_),
    .X(_06030_));
 sg13g2_xnor2_1 _15237_ (.Y(_06031_),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[17] ),
    .B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xnor2_1 _15238_ (.Y(_00874_),
    .A(_06030_),
    .B(_06031_));
 sg13g2_a21o_1 _15239_ (.A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[17] ),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[17] ),
    .B1(_06030_),
    .X(_06032_));
 sg13g2_o21ai_1 _15240_ (.B1(_06032_),
    .Y(_06033_),
    .A1(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xor2_1 _15241_ (.B(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[18] ),
    .X(_06034_));
 sg13g2_xnor2_1 _15242_ (.Y(_00875_),
    .A(_06033_),
    .B(_06034_));
 sg13g2_and2_1 _15243_ (.A(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.u_mux_shift.sum_res ),
    .B(net4930),
    .X(_00223_));
 sg13g2_nor2b_1 _15244_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][1] ),
    .Y(_06035_));
 sg13g2_xnor2_1 _15245_ (.Y(_06036_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][1] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _15246_ (.B(_06036_),
    .A(_02515_),
    .X(_00933_));
 sg13g2_a21oi_1 _15247_ (.A1(_02515_),
    .A2(_06036_),
    .Y(_06037_),
    .B1(_06035_));
 sg13g2_xnor2_1 _15248_ (.Y(_06038_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][2] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _15249_ (.A(_06037_),
    .B_N(_06038_),
    .Y(_06039_));
 sg13g2_xnor2_1 _15250_ (.Y(_00934_),
    .A(_06037_),
    .B(_06038_));
 sg13g2_a21oi_1 _15251_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][2] ),
    .A2(_02460_),
    .Y(_06040_),
    .B1(_06039_));
 sg13g2_xnor2_1 _15252_ (.Y(_06041_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][3] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _15253_ (.A(_06040_),
    .B_N(_06041_),
    .Y(_06042_));
 sg13g2_xnor2_1 _15254_ (.Y(_00935_),
    .A(_06040_),
    .B(_06041_));
 sg13g2_a21oi_1 _15255_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][3] ),
    .A2(_02461_),
    .Y(_06043_),
    .B1(_06042_));
 sg13g2_xnor2_1 _15256_ (.Y(_06044_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][4] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _15257_ (.A(_06043_),
    .B_N(_06044_),
    .Y(_06045_));
 sg13g2_xnor2_1 _15258_ (.Y(_00936_),
    .A(_06043_),
    .B(_06044_));
 sg13g2_a21oi_1 _15259_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][4] ),
    .A2(_02462_),
    .Y(_06046_),
    .B1(_06045_));
 sg13g2_xnor2_1 _15260_ (.Y(_06047_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][5] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _15261_ (.A(_06046_),
    .B_N(_06047_),
    .Y(_06048_));
 sg13g2_xnor2_1 _15262_ (.Y(_00937_),
    .A(_06046_),
    .B(_06047_));
 sg13g2_a21oi_2 _15263_ (.B1(_06048_),
    .Y(_06049_),
    .A2(_02463_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][5] ));
 sg13g2_xnor2_1 _15264_ (.Y(_06050_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][6] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_nor2b_1 _15265_ (.A(_06049_),
    .B_N(_06050_),
    .Y(_06051_));
 sg13g2_xnor2_1 _15266_ (.Y(_00938_),
    .A(_06049_),
    .B(_06050_));
 sg13g2_a21oi_2 _15267_ (.B1(_06051_),
    .Y(_06052_),
    .A2(_02464_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][6] ));
 sg13g2_xnor2_1 _15268_ (.Y(_06053_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][7] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _15269_ (.A(_06052_),
    .B_N(_06053_),
    .Y(_06054_));
 sg13g2_xnor2_1 _15270_ (.Y(_00939_),
    .A(_06052_),
    .B(_06053_));
 sg13g2_a21oi_2 _15271_ (.B1(_06054_),
    .Y(_06055_),
    .A2(_02465_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][7] ));
 sg13g2_xnor2_1 _15272_ (.Y(_06056_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][8] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_nor2b_1 _15273_ (.A(_06055_),
    .B_N(_06056_),
    .Y(_06057_));
 sg13g2_xnor2_1 _15274_ (.Y(_00940_),
    .A(_06055_),
    .B(_06056_));
 sg13g2_a21oi_2 _15275_ (.B1(_06057_),
    .Y(_06058_),
    .A2(_02466_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][8] ));
 sg13g2_nor2b_1 _15276_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][9] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[9] ),
    .Y(_06059_));
 sg13g2_nand2b_1 _15277_ (.Y(_06060_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][9] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _15278_ (.A(_06059_),
    .B_N(_06060_),
    .Y(_06061_));
 sg13g2_xnor2_1 _15279_ (.Y(_00941_),
    .A(_06058_),
    .B(_06061_));
 sg13g2_nor2b_1 _15280_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][10] ),
    .Y(_06062_));
 sg13g2_nand2b_1 _15281_ (.Y(_06063_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][10] ));
 sg13g2_nand2b_1 _15282_ (.Y(_06064_),
    .B(_06063_),
    .A_N(_06062_));
 sg13g2_a21oi_1 _15283_ (.A1(_06058_),
    .A2(_06060_),
    .Y(_06065_),
    .B1(_06059_));
 sg13g2_xnor2_1 _15284_ (.Y(_00924_),
    .A(_06064_),
    .B(_06065_));
 sg13g2_a21oi_1 _15285_ (.A1(_06063_),
    .A2(_06065_),
    .Y(_06066_),
    .B1(_06062_));
 sg13g2_nor2b_1 _15286_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][11] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[11] ),
    .Y(_06067_));
 sg13g2_nand2b_1 _15287_ (.Y(_06068_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][11] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _15288_ (.A(_06067_),
    .B_N(_06068_),
    .Y(_06069_));
 sg13g2_xnor2_1 _15289_ (.Y(_00925_),
    .A(_06066_),
    .B(_06069_));
 sg13g2_nor2b_1 _15290_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][12] ),
    .Y(_06070_));
 sg13g2_nand2b_1 _15291_ (.Y(_06071_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][12] ));
 sg13g2_nand2b_1 _15292_ (.Y(_06072_),
    .B(_06071_),
    .A_N(_06070_));
 sg13g2_a21oi_1 _15293_ (.A1(_06066_),
    .A2(_06068_),
    .Y(_06073_),
    .B1(_06067_));
 sg13g2_xnor2_1 _15294_ (.Y(_00926_),
    .A(_06072_),
    .B(_06073_));
 sg13g2_a21oi_1 _15295_ (.A1(_06071_),
    .A2(_06073_),
    .Y(_06074_),
    .B1(_06070_));
 sg13g2_nor2b_1 _15296_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][13] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[13] ),
    .Y(_06075_));
 sg13g2_nand2b_1 _15297_ (.Y(_06076_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][13] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _15298_ (.A(_06075_),
    .B_N(_06076_),
    .Y(_06077_));
 sg13g2_xnor2_1 _15299_ (.Y(_00927_),
    .A(_06074_),
    .B(_06077_));
 sg13g2_nor2b_1 _15300_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][14] ),
    .Y(_06078_));
 sg13g2_nand2b_1 _15301_ (.Y(_06079_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][14] ));
 sg13g2_nand2b_1 _15302_ (.Y(_06080_),
    .B(_06079_),
    .A_N(_06078_));
 sg13g2_a21oi_1 _15303_ (.A1(_06074_),
    .A2(_06076_),
    .Y(_06081_),
    .B1(_06075_));
 sg13g2_xnor2_1 _15304_ (.Y(_00928_),
    .A(_06080_),
    .B(_06081_));
 sg13g2_a21oi_1 _15305_ (.A1(_06079_),
    .A2(_06081_),
    .Y(_06082_),
    .B1(_06078_));
 sg13g2_nor2b_1 _15306_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][15] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[15] ),
    .Y(_06083_));
 sg13g2_nand2b_1 _15307_ (.Y(_06084_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][15] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _15308_ (.A(_06083_),
    .B_N(_06084_),
    .Y(_06085_));
 sg13g2_xnor2_1 _15309_ (.Y(_00929_),
    .A(_06082_),
    .B(_06085_));
 sg13g2_xor2_1 _15310_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][16] ),
    .X(_06086_));
 sg13g2_a21oi_1 _15311_ (.A1(_06082_),
    .A2(_06084_),
    .Y(_06087_),
    .B1(_06083_));
 sg13g2_nor2b_1 _15312_ (.A(_06086_),
    .B_N(_06087_),
    .Y(_06088_));
 sg13g2_xnor2_1 _15313_ (.Y(_00930_),
    .A(_06086_),
    .B(_06087_));
 sg13g2_a21oi_2 _15314_ (.B1(_06088_),
    .Y(_06089_),
    .A2(_02467_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][16] ));
 sg13g2_nand2b_1 _15315_ (.Y(_06090_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][17] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _15316_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][17] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[17] ),
    .Y(_06091_));
 sg13g2_xnor2_1 _15317_ (.Y(_06092_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][17] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _15318_ (.Y(_00931_),
    .A(_06089_),
    .B(_06092_));
 sg13g2_o21ai_1 _15319_ (.B1(_06090_),
    .Y(_06093_),
    .A1(_06089_),
    .A2(_06091_));
 sg13g2_xor2_1 _15320_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][18] ),
    .X(_06094_));
 sg13g2_xnor2_1 _15321_ (.Y(_00932_),
    .A(_06093_),
    .B(_06094_));
 sg13g2_nand2_1 _15322_ (.Y(_06095_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[0] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_nand2_1 _15323_ (.Y(_06096_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_nor2_1 _15324_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[1] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[1] ),
    .Y(_06097_));
 sg13g2_xor2_1 _15325_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[1] ),
    .X(_06098_));
 sg13g2_xnor2_1 _15326_ (.Y(_00782_),
    .A(_06095_),
    .B(_06098_));
 sg13g2_o21ai_1 _15327_ (.B1(_06096_),
    .Y(_06099_),
    .A1(_06095_),
    .A2(_06097_));
 sg13g2_xnor2_1 _15328_ (.Y(_06100_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[2] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_nor2b_1 _15329_ (.A(_06100_),
    .B_N(_06099_),
    .Y(_06101_));
 sg13g2_xnor2_1 _15330_ (.Y(_00783_),
    .A(_06099_),
    .B(_06100_));
 sg13g2_a21o_1 _15331_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[2] ),
    .B1(_06101_),
    .X(_06102_));
 sg13g2_xnor2_1 _15332_ (.Y(_06103_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[3] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_nor2b_1 _15333_ (.A(_06103_),
    .B_N(_06102_),
    .Y(_06104_));
 sg13g2_xnor2_1 _15334_ (.Y(_00784_),
    .A(_06102_),
    .B(_06103_));
 sg13g2_a21o_1 _15335_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[3] ),
    .B1(_06104_),
    .X(_06105_));
 sg13g2_xnor2_1 _15336_ (.Y(_06106_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[4] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_nor2b_1 _15337_ (.A(_06106_),
    .B_N(_06105_),
    .Y(_06107_));
 sg13g2_xnor2_1 _15338_ (.Y(_00785_),
    .A(_06105_),
    .B(_06106_));
 sg13g2_a21o_1 _15339_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[4] ),
    .B1(_06107_),
    .X(_06108_));
 sg13g2_nand2_1 _15340_ (.Y(_06109_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _15341_ (.Y(_06110_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[5] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_xnor2_1 _15342_ (.Y(_00786_),
    .A(_06108_),
    .B(_06110_));
 sg13g2_xnor2_1 _15343_ (.Y(_06111_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[6] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_o21ai_1 _15344_ (.B1(_06108_),
    .Y(_06112_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_a21oi_1 _15345_ (.A1(_06109_),
    .A2(_06112_),
    .Y(_06113_),
    .B1(_06111_));
 sg13g2_nand3_1 _15346_ (.B(_06111_),
    .C(_06112_),
    .A(_06109_),
    .Y(_06114_));
 sg13g2_nor2b_1 _15347_ (.A(_06113_),
    .B_N(_06114_),
    .Y(_00787_));
 sg13g2_a21oi_1 _15348_ (.A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[6] ),
    .Y(_06115_),
    .B1(_06113_));
 sg13g2_nand2_1 _15349_ (.Y(_06116_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_nor2_1 _15350_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[7] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[7] ),
    .Y(_06117_));
 sg13g2_xor2_1 _15351_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[7] ),
    .X(_06118_));
 sg13g2_xnor2_1 _15352_ (.Y(_00788_),
    .A(_06115_),
    .B(_06118_));
 sg13g2_o21ai_1 _15353_ (.B1(_06116_),
    .Y(_06119_),
    .A1(_06115_),
    .A2(_06117_));
 sg13g2_xnor2_1 _15354_ (.Y(_06120_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[8] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_nor2b_1 _15355_ (.A(_06120_),
    .B_N(_06119_),
    .Y(_06121_));
 sg13g2_xnor2_1 _15356_ (.Y(_00789_),
    .A(_06119_),
    .B(_06120_));
 sg13g2_a21o_1 _15357_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[8] ),
    .B1(_06121_),
    .X(_06122_));
 sg13g2_xnor2_1 _15358_ (.Y(_06123_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[9] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _15359_ (.Y(_00790_),
    .A(_06122_),
    .B(_06123_));
 sg13g2_nand2_1 _15360_ (.Y(_06124_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_nor2_1 _15361_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[10] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[10] ),
    .Y(_06125_));
 sg13g2_xor2_1 _15362_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[10] ),
    .X(_06126_));
 sg13g2_a21o_1 _15363_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[9] ),
    .B1(_06122_),
    .X(_06127_));
 sg13g2_o21ai_1 _15364_ (.B1(_06127_),
    .Y(_06128_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_xnor2_1 _15365_ (.Y(_00773_),
    .A(_06126_),
    .B(_06128_));
 sg13g2_o21ai_1 _15366_ (.B1(_06124_),
    .Y(_06129_),
    .A1(_06125_),
    .A2(_06128_));
 sg13g2_xnor2_1 _15367_ (.Y(_06130_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[11] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _15368_ (.Y(_00774_),
    .A(_06129_),
    .B(_06130_));
 sg13g2_nand2_1 _15369_ (.Y(_06131_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[12] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_nor2_1 _15370_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[12] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[12] ),
    .Y(_06132_));
 sg13g2_xor2_1 _15371_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[12] ),
    .X(_06133_));
 sg13g2_a21o_1 _15372_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[11] ),
    .B1(_06129_),
    .X(_06134_));
 sg13g2_o21ai_1 _15373_ (.B1(_06134_),
    .Y(_06135_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_xnor2_1 _15374_ (.Y(_00775_),
    .A(_06133_),
    .B(_06135_));
 sg13g2_o21ai_1 _15375_ (.B1(_06131_),
    .Y(_06136_),
    .A1(_06132_),
    .A2(_06135_));
 sg13g2_xnor2_1 _15376_ (.Y(_06137_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[13] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_xnor2_1 _15377_ (.Y(_00776_),
    .A(_06136_),
    .B(_06137_));
 sg13g2_xor2_1 _15378_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[14] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[14] ),
    .X(_06138_));
 sg13g2_a21o_1 _15379_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[13] ),
    .B1(_06136_),
    .X(_06139_));
 sg13g2_o21ai_1 _15380_ (.B1(_06139_),
    .Y(_06140_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_nor2b_1 _15381_ (.A(_06140_),
    .B_N(_06138_),
    .Y(_06141_));
 sg13g2_xnor2_1 _15382_ (.Y(_00777_),
    .A(_06138_),
    .B(_06140_));
 sg13g2_a21o_1 _15383_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[14] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[14] ),
    .B1(_06141_),
    .X(_06142_));
 sg13g2_and2_1 _15384_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[15] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[15] ),
    .X(_06143_));
 sg13g2_or2_1 _15385_ (.X(_06144_),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[15] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand2b_1 _15386_ (.Y(_06145_),
    .B(_06144_),
    .A_N(_06143_));
 sg13g2_xnor2_1 _15387_ (.Y(_00778_),
    .A(_06142_),
    .B(_06145_));
 sg13g2_and2_1 _15388_ (.A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[16] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[16] ),
    .X(_06146_));
 sg13g2_xor2_1 _15389_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[16] ),
    .X(_06147_));
 sg13g2_a21o_1 _15390_ (.A2(_06144_),
    .A1(_06142_),
    .B1(_06143_),
    .X(_06148_));
 sg13g2_xor2_1 _15391_ (.B(_06148_),
    .A(_06147_),
    .X(_00779_));
 sg13g2_a21o_1 _15392_ (.A2(_06148_),
    .A1(_06147_),
    .B1(_06146_),
    .X(_06149_));
 sg13g2_xnor2_1 _15393_ (.Y(_06150_),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[17] ),
    .B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xnor2_1 _15394_ (.Y(_00780_),
    .A(_06149_),
    .B(_06150_));
 sg13g2_a21o_1 _15395_ (.A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[17] ),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[17] ),
    .B1(_06149_),
    .X(_06151_));
 sg13g2_o21ai_1 _15396_ (.B1(_06151_),
    .Y(_06152_),
    .A1(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_xor2_1 _15397_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[18] ),
    .X(_06153_));
 sg13g2_xnor2_1 _15398_ (.Y(_00781_),
    .A(_06152_),
    .B(_06153_));
 sg13g2_xor2_1 _15399_ (.B(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[0] ),
    .X(_00772_));
 sg13g2_nor2b_1 _15400_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][1] ),
    .Y(_06154_));
 sg13g2_xnor2_1 _15401_ (.Y(_06155_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][1] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _15402_ (.B(_06155_),
    .A(_02516_),
    .X(_01008_));
 sg13g2_a21oi_2 _15403_ (.B1(_06154_),
    .Y(_06156_),
    .A2(_06155_),
    .A1(_02516_));
 sg13g2_xnor2_1 _15404_ (.Y(_06157_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][2] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _15405_ (.A(_06156_),
    .B_N(_06157_),
    .Y(_06158_));
 sg13g2_xnor2_1 _15406_ (.Y(_01009_),
    .A(_06156_),
    .B(_06157_));
 sg13g2_a21oi_1 _15407_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][2] ),
    .A2(_02468_),
    .Y(_06159_),
    .B1(_06158_));
 sg13g2_xnor2_1 _15408_ (.Y(_06160_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][3] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _15409_ (.A(_06159_),
    .B_N(_06160_),
    .Y(_06161_));
 sg13g2_xnor2_1 _15410_ (.Y(_01010_),
    .A(_06159_),
    .B(_06160_));
 sg13g2_a21oi_1 _15411_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][3] ),
    .A2(_02469_),
    .Y(_06162_),
    .B1(_06161_));
 sg13g2_xnor2_1 _15412_ (.Y(_06163_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][4] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _15413_ (.A(_06162_),
    .B_N(_06163_),
    .Y(_06164_));
 sg13g2_xnor2_1 _15414_ (.Y(_01011_),
    .A(_06162_),
    .B(_06163_));
 sg13g2_a21oi_1 _15415_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][4] ),
    .A2(_02470_),
    .Y(_06165_),
    .B1(_06164_));
 sg13g2_nand2b_1 _15416_ (.Y(_06166_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][5] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _15417_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][5] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[5] ),
    .Y(_06167_));
 sg13g2_xnor2_1 _15418_ (.Y(_06168_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][5] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_xnor2_1 _15419_ (.Y(_01012_),
    .A(_06165_),
    .B(_06168_));
 sg13g2_nor2b_1 _15420_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[6] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][6] ),
    .Y(_06169_));
 sg13g2_nand2b_1 _15421_ (.Y(_06170_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[6] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][6] ));
 sg13g2_nand2b_1 _15422_ (.Y(_06171_),
    .B(_06170_),
    .A_N(_06169_));
 sg13g2_o21ai_1 _15423_ (.B1(_06166_),
    .Y(_06172_),
    .A1(_06165_),
    .A2(_06167_));
 sg13g2_xnor2_1 _15424_ (.Y(_01013_),
    .A(_06171_),
    .B(_06172_));
 sg13g2_a21oi_1 _15425_ (.A1(_06170_),
    .A2(_06172_),
    .Y(_06173_),
    .B1(_06169_));
 sg13g2_xnor2_1 _15426_ (.Y(_06174_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][7] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nand2b_1 _15427_ (.Y(_06175_),
    .B(_06174_),
    .A_N(_06173_));
 sg13g2_xnor2_1 _15428_ (.Y(_01014_),
    .A(_06173_),
    .B(_06174_));
 sg13g2_o21ai_1 _15429_ (.B1(_06175_),
    .Y(_06176_),
    .A1(_02471_),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _15430_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[8] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][8] ),
    .Y(_06177_));
 sg13g2_nand2b_1 _15431_ (.Y(_06178_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[8] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][8] ));
 sg13g2_nand2b_1 _15432_ (.Y(_06179_),
    .B(_06178_),
    .A_N(_06177_));
 sg13g2_xnor2_1 _15433_ (.Y(_01015_),
    .A(_06176_),
    .B(_06179_));
 sg13g2_a21oi_1 _15434_ (.A1(_06176_),
    .A2(_06178_),
    .Y(_06180_),
    .B1(_06177_));
 sg13g2_nand2b_1 _15435_ (.Y(_06181_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][9] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _15436_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][9] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[9] ),
    .Y(_06182_));
 sg13g2_xnor2_1 _15437_ (.Y(_06183_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][9] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_xnor2_1 _15438_ (.Y(_01016_),
    .A(_06180_),
    .B(_06183_));
 sg13g2_nor2b_1 _15439_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][10] ),
    .Y(_06184_));
 sg13g2_nand2b_1 _15440_ (.Y(_06185_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][10] ));
 sg13g2_nand2b_1 _15441_ (.Y(_06186_),
    .B(_06185_),
    .A_N(_06184_));
 sg13g2_a21oi_1 _15442_ (.A1(_06180_),
    .A2(_06181_),
    .Y(_06187_),
    .B1(_06182_));
 sg13g2_xnor2_1 _15443_ (.Y(_00999_),
    .A(_06186_),
    .B(_06187_));
 sg13g2_a21oi_1 _15444_ (.A1(_06185_),
    .A2(_06187_),
    .Y(_06188_),
    .B1(_06184_));
 sg13g2_nor2b_1 _15445_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][11] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[11] ),
    .Y(_06189_));
 sg13g2_nand2b_1 _15446_ (.Y(_06190_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][11] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _15447_ (.A(_06189_),
    .B_N(_06190_),
    .Y(_06191_));
 sg13g2_xnor2_1 _15448_ (.Y(_01000_),
    .A(_06188_),
    .B(_06191_));
 sg13g2_nor2b_1 _15449_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][12] ),
    .Y(_06192_));
 sg13g2_nand2b_1 _15450_ (.Y(_06193_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][12] ));
 sg13g2_nand2b_1 _15451_ (.Y(_06194_),
    .B(_06193_),
    .A_N(_06192_));
 sg13g2_a21oi_1 _15452_ (.A1(_06188_),
    .A2(_06190_),
    .Y(_06195_),
    .B1(_06189_));
 sg13g2_xnor2_1 _15453_ (.Y(_01001_),
    .A(_06194_),
    .B(_06195_));
 sg13g2_a21oi_1 _15454_ (.A1(_06193_),
    .A2(_06195_),
    .Y(_06196_),
    .B1(_06192_));
 sg13g2_nand2b_1 _15455_ (.Y(_06197_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][13] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _15456_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][13] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[13] ),
    .Y(_06198_));
 sg13g2_xnor2_1 _15457_ (.Y(_06199_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][13] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_xnor2_1 _15458_ (.Y(_01002_),
    .A(_06196_),
    .B(_06199_));
 sg13g2_nor2b_1 _15459_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][14] ),
    .Y(_06200_));
 sg13g2_nand2b_1 _15460_ (.Y(_06201_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][14] ));
 sg13g2_nand2b_1 _15461_ (.Y(_06202_),
    .B(_06201_),
    .A_N(_06200_));
 sg13g2_a21oi_1 _15462_ (.A1(_06196_),
    .A2(_06197_),
    .Y(_06203_),
    .B1(_06198_));
 sg13g2_xnor2_1 _15463_ (.Y(_01003_),
    .A(_06202_),
    .B(_06203_));
 sg13g2_a21oi_1 _15464_ (.A1(_06201_),
    .A2(_06203_),
    .Y(_06204_),
    .B1(_06200_));
 sg13g2_nand2b_1 _15465_ (.Y(_06205_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][15] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _15466_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][15] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[15] ),
    .Y(_06206_));
 sg13g2_xnor2_1 _15467_ (.Y(_06207_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][15] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_xnor2_1 _15468_ (.Y(_01004_),
    .A(_06204_),
    .B(_06207_));
 sg13g2_xor2_1 _15469_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][16] ),
    .X(_06208_));
 sg13g2_a21oi_1 _15470_ (.A1(_06204_),
    .A2(_06205_),
    .Y(_06209_),
    .B1(_06206_));
 sg13g2_nor2b_1 _15471_ (.A(_06208_),
    .B_N(_06209_),
    .Y(_06210_));
 sg13g2_xnor2_1 _15472_ (.Y(_01005_),
    .A(_06208_),
    .B(_06209_));
 sg13g2_a21oi_1 _15473_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][16] ),
    .A2(_02472_),
    .Y(_06211_),
    .B1(_06210_));
 sg13g2_nand2b_1 _15474_ (.Y(_06212_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][17] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _15475_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][17] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[17] ),
    .Y(_06213_));
 sg13g2_xnor2_1 _15476_ (.Y(_06214_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][17] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _15477_ (.Y(_01006_),
    .A(_06211_),
    .B(_06214_));
 sg13g2_o21ai_1 _15478_ (.B1(_06212_),
    .Y(_06215_),
    .A1(_06211_),
    .A2(_06213_));
 sg13g2_xor2_1 _15479_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][18] ),
    .X(_06216_));
 sg13g2_xnor2_1 _15480_ (.Y(_01007_),
    .A(_06215_),
    .B(_06216_));
 sg13g2_nand2_1 _15481_ (.Y(_06217_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[0] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_xor2_1 _15482_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[0] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[0] ),
    .X(_00979_));
 sg13g2_nand2_1 _15483_ (.Y(_06218_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[1] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_nor2_1 _15484_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[1] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[1] ),
    .Y(_06219_));
 sg13g2_xor2_1 _15485_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[1] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[1] ),
    .X(_06220_));
 sg13g2_xnor2_1 _15486_ (.Y(_00989_),
    .A(_06217_),
    .B(_06220_));
 sg13g2_o21ai_1 _15487_ (.B1(_06218_),
    .Y(_06221_),
    .A1(_06217_),
    .A2(_06219_));
 sg13g2_xnor2_1 _15488_ (.Y(_06222_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[2] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_nor2b_1 _15489_ (.A(_06222_),
    .B_N(_06221_),
    .Y(_06223_));
 sg13g2_xnor2_1 _15490_ (.Y(_00990_),
    .A(_06221_),
    .B(_06222_));
 sg13g2_a21o_1 _15491_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[2] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[2] ),
    .B1(_06223_),
    .X(_06224_));
 sg13g2_xnor2_1 _15492_ (.Y(_06225_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[3] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_nor2b_1 _15493_ (.A(_06225_),
    .B_N(_06224_),
    .Y(_06226_));
 sg13g2_xnor2_1 _15494_ (.Y(_00991_),
    .A(_06224_),
    .B(_06225_));
 sg13g2_a21o_1 _15495_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[3] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[3] ),
    .B1(_06226_),
    .X(_06227_));
 sg13g2_xnor2_1 _15496_ (.Y(_06228_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[4] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_nor2b_1 _15497_ (.A(_06228_),
    .B_N(_06227_),
    .Y(_06229_));
 sg13g2_xnor2_1 _15498_ (.Y(_00992_),
    .A(_06227_),
    .B(_06228_));
 sg13g2_a21o_1 _15499_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[4] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[4] ),
    .B1(_06229_),
    .X(_06230_));
 sg13g2_nand2_1 _15500_ (.Y(_06231_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[5] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_xnor2_1 _15501_ (.Y(_06232_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[5] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_xnor2_1 _15502_ (.Y(_00993_),
    .A(_06230_),
    .B(_06232_));
 sg13g2_xnor2_1 _15503_ (.Y(_06233_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[6] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_o21ai_1 _15504_ (.B1(_06230_),
    .Y(_06234_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[5] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_a21oi_1 _15505_ (.A1(_06231_),
    .A2(_06234_),
    .Y(_06235_),
    .B1(_06233_));
 sg13g2_nand3_1 _15506_ (.B(_06233_),
    .C(_06234_),
    .A(_06231_),
    .Y(_06236_));
 sg13g2_nor2b_1 _15507_ (.A(_06235_),
    .B_N(_06236_),
    .Y(_00994_));
 sg13g2_a21oi_2 _15508_ (.B1(_06235_),
    .Y(_06237_),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[6] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_nand2_1 _15509_ (.Y(_06238_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[7] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_nor2_1 _15510_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[7] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[7] ),
    .Y(_06239_));
 sg13g2_xor2_1 _15511_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[7] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[7] ),
    .X(_06240_));
 sg13g2_xnor2_1 _15512_ (.Y(_00995_),
    .A(_06237_),
    .B(_06240_));
 sg13g2_o21ai_1 _15513_ (.B1(_06238_),
    .Y(_06241_),
    .A1(_06237_),
    .A2(_06239_));
 sg13g2_xnor2_1 _15514_ (.Y(_06242_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[8] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_nor2b_1 _15515_ (.A(_06242_),
    .B_N(_06241_),
    .Y(_06243_));
 sg13g2_xnor2_1 _15516_ (.Y(_00996_),
    .A(_06241_),
    .B(_06242_));
 sg13g2_a21o_1 _15517_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[8] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[8] ),
    .B1(_06243_),
    .X(_06244_));
 sg13g2_xnor2_1 _15518_ (.Y(_06245_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[9] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_xnor2_1 _15519_ (.Y(_00997_),
    .A(_06244_),
    .B(_06245_));
 sg13g2_nand2_1 _15520_ (.Y(_06246_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[10] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_nor2_1 _15521_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[10] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[10] ),
    .Y(_06247_));
 sg13g2_xor2_1 _15522_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[10] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[10] ),
    .X(_06248_));
 sg13g2_a21o_1 _15523_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[9] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[9] ),
    .B1(_06244_),
    .X(_06249_));
 sg13g2_o21ai_1 _15524_ (.B1(_06249_),
    .Y(_06250_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[9] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_xnor2_1 _15525_ (.Y(_00980_),
    .A(_06248_),
    .B(_06250_));
 sg13g2_o21ai_1 _15526_ (.B1(_06246_),
    .Y(_01808_),
    .A1(_06247_),
    .A2(_06250_));
 sg13g2_xnor2_1 _15527_ (.Y(_01809_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[11] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_xnor2_1 _15528_ (.Y(_00981_),
    .A(_01808_),
    .B(_01809_));
 sg13g2_nand2_1 _15529_ (.Y(_01810_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[12] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_nor2_1 _15530_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[12] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[12] ),
    .Y(_01811_));
 sg13g2_xor2_1 _15531_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[12] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[12] ),
    .X(_01812_));
 sg13g2_a21o_1 _15532_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[11] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[11] ),
    .B1(_01808_),
    .X(_01813_));
 sg13g2_o21ai_1 _15533_ (.B1(_01813_),
    .Y(_01814_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[11] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_xnor2_1 _15534_ (.Y(_00982_),
    .A(_01812_),
    .B(_01814_));
 sg13g2_o21ai_1 _15535_ (.B1(_01810_),
    .Y(_01815_),
    .A1(_01811_),
    .A2(_01814_));
 sg13g2_xnor2_1 _15536_ (.Y(_01816_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[13] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_xnor2_1 _15537_ (.Y(_00983_),
    .A(_01815_),
    .B(_01816_));
 sg13g2_xnor2_1 _15538_ (.Y(_01817_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[14] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_a21o_1 _15539_ (.A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[13] ),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[13] ),
    .B1(_01815_),
    .X(_01818_));
 sg13g2_o21ai_1 _15540_ (.B1(_01818_),
    .Y(_01819_),
    .A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[13] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_nor2_1 _15541_ (.A(_01817_),
    .B(_01819_),
    .Y(_01820_));
 sg13g2_xor2_1 _15542_ (.B(_01819_),
    .A(_01817_),
    .X(_00984_));
 sg13g2_a21oi_1 _15543_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[14] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[14] ),
    .Y(_01821_),
    .B1(_01820_));
 sg13g2_nand2_1 _15544_ (.Y(_01822_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[15] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_nor2_1 _15545_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[15] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[15] ),
    .Y(_01823_));
 sg13g2_xor2_1 _15546_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[15] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[15] ),
    .X(_01824_));
 sg13g2_xnor2_1 _15547_ (.Y(_00985_),
    .A(_01821_),
    .B(_01824_));
 sg13g2_nand2_1 _15548_ (.Y(_01825_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[16] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_xor2_1 _15549_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[16] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[16] ),
    .X(_01826_));
 sg13g2_o21ai_1 _15550_ (.B1(_01822_),
    .Y(_01827_),
    .A1(_01821_),
    .A2(_01823_));
 sg13g2_nand2_1 _15551_ (.Y(_01828_),
    .A(_01826_),
    .B(_01827_));
 sg13g2_xor2_1 _15552_ (.B(_01827_),
    .A(_01826_),
    .X(_00986_));
 sg13g2_xnor2_1 _15553_ (.Y(_01829_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[17] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_a21oi_1 _15554_ (.A1(_01825_),
    .A2(_01828_),
    .Y(_01830_),
    .B1(_01829_));
 sg13g2_nand3_1 _15555_ (.B(_01828_),
    .C(_01829_),
    .A(_01825_),
    .Y(_01831_));
 sg13g2_nor2b_1 _15556_ (.A(_01830_),
    .B_N(_01831_),
    .Y(_00987_));
 sg13g2_a21oi_1 _15557_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[17] ),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[17] ),
    .Y(_01832_),
    .B1(_01830_));
 sg13g2_xor2_1 _15558_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[18] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[18] ),
    .X(_01833_));
 sg13g2_xnor2_1 _15559_ (.Y(_00988_),
    .A(_01832_),
    .B(_01833_));
 sg13g2_nand2_1 _15560_ (.Y(_01834_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[0] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_xor2_1 _15561_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[0] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[0] ),
    .X(_01073_));
 sg13g2_nand2_1 _15562_ (.Y(_01835_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[1] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_nor2_1 _15563_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[1] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[1] ),
    .Y(_01836_));
 sg13g2_xor2_1 _15564_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[1] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[1] ),
    .X(_01837_));
 sg13g2_xnor2_1 _15565_ (.Y(_01083_),
    .A(_01834_),
    .B(_01837_));
 sg13g2_o21ai_1 _15566_ (.B1(_01835_),
    .Y(_01838_),
    .A1(_01834_),
    .A2(_01836_));
 sg13g2_xnor2_1 _15567_ (.Y(_01839_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[2] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_nor2b_1 _15568_ (.A(_01839_),
    .B_N(_01838_),
    .Y(_01840_));
 sg13g2_xnor2_1 _15569_ (.Y(_01084_),
    .A(_01838_),
    .B(_01839_));
 sg13g2_a21o_1 _15570_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[2] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[2] ),
    .B1(_01840_),
    .X(_01841_));
 sg13g2_xnor2_1 _15571_ (.Y(_01842_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[3] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_nor2b_1 _15572_ (.A(_01842_),
    .B_N(_01841_),
    .Y(_01843_));
 sg13g2_xnor2_1 _15573_ (.Y(_01085_),
    .A(_01841_),
    .B(_01842_));
 sg13g2_a21o_1 _15574_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[3] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[3] ),
    .B1(_01843_),
    .X(_01844_));
 sg13g2_xnor2_1 _15575_ (.Y(_01845_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[4] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_nor2b_1 _15576_ (.A(_01845_),
    .B_N(_01844_),
    .Y(_01846_));
 sg13g2_xnor2_1 _15577_ (.Y(_01086_),
    .A(_01844_),
    .B(_01845_));
 sg13g2_a21o_1 _15578_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[4] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[4] ),
    .B1(_01846_),
    .X(_01847_));
 sg13g2_nand2_1 _15579_ (.Y(_01848_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[5] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_xnor2_1 _15580_ (.Y(_01849_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[5] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_xnor2_1 _15581_ (.Y(_01087_),
    .A(_01847_),
    .B(_01849_));
 sg13g2_xnor2_1 _15582_ (.Y(_01850_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[6] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_o21ai_1 _15583_ (.B1(_01847_),
    .Y(_01851_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[5] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_a21oi_1 _15584_ (.A1(_01848_),
    .A2(_01851_),
    .Y(_01852_),
    .B1(_01850_));
 sg13g2_nand3_1 _15585_ (.B(_01850_),
    .C(_01851_),
    .A(_01848_),
    .Y(_01853_));
 sg13g2_nor2b_1 _15586_ (.A(_01852_),
    .B_N(_01853_),
    .Y(_01088_));
 sg13g2_a21oi_2 _15587_ (.B1(_01852_),
    .Y(_01854_),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[6] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_nand2_1 _15588_ (.Y(_01855_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[7] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_nor2_1 _15589_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[7] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[7] ),
    .Y(_01856_));
 sg13g2_xor2_1 _15590_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[7] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[7] ),
    .X(_01857_));
 sg13g2_xnor2_1 _15591_ (.Y(_01089_),
    .A(_01854_),
    .B(_01857_));
 sg13g2_o21ai_1 _15592_ (.B1(_01855_),
    .Y(_01858_),
    .A1(_01854_),
    .A2(_01856_));
 sg13g2_xnor2_1 _15593_ (.Y(_01859_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[8] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_nor2b_1 _15594_ (.A(_01859_),
    .B_N(_01858_),
    .Y(_01860_));
 sg13g2_xnor2_1 _15595_ (.Y(_01090_),
    .A(_01858_),
    .B(_01859_));
 sg13g2_a21o_1 _15596_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[8] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[8] ),
    .B1(_01860_),
    .X(_01861_));
 sg13g2_xnor2_1 _15597_ (.Y(_01862_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[9] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_xnor2_1 _15598_ (.Y(_01091_),
    .A(_01861_),
    .B(_01862_));
 sg13g2_nand2_1 _15599_ (.Y(_01863_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[10] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_nor2_1 _15600_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[10] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[10] ),
    .Y(_01864_));
 sg13g2_xor2_1 _15601_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[10] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[10] ),
    .X(_01865_));
 sg13g2_a21o_1 _15602_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[9] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[9] ),
    .B1(_01861_),
    .X(_01866_));
 sg13g2_o21ai_1 _15603_ (.B1(_01866_),
    .Y(_01867_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[9] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_xnor2_1 _15604_ (.Y(_01074_),
    .A(_01865_),
    .B(_01867_));
 sg13g2_o21ai_1 _15605_ (.B1(_01863_),
    .Y(_01868_),
    .A1(_01864_),
    .A2(_01867_));
 sg13g2_xnor2_1 _15606_ (.Y(_01869_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[11] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_xnor2_1 _15607_ (.Y(_01075_),
    .A(_01868_),
    .B(_01869_));
 sg13g2_nand2_1 _15608_ (.Y(_01870_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[12] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_nor2_1 _15609_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[12] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[12] ),
    .Y(_01871_));
 sg13g2_xor2_1 _15610_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[12] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[12] ),
    .X(_01872_));
 sg13g2_a21o_1 _15611_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[11] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[11] ),
    .B1(_01868_),
    .X(_01873_));
 sg13g2_o21ai_1 _15612_ (.B1(_01873_),
    .Y(_01874_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[11] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_xnor2_1 _15613_ (.Y(_01076_),
    .A(_01872_),
    .B(_01874_));
 sg13g2_o21ai_1 _15614_ (.B1(_01870_),
    .Y(_01875_),
    .A1(_01871_),
    .A2(_01874_));
 sg13g2_xnor2_1 _15615_ (.Y(_01876_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[13] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_xnor2_1 _15616_ (.Y(_01077_),
    .A(_01875_),
    .B(_01876_));
 sg13g2_xor2_1 _15617_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[14] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[14] ),
    .X(_01877_));
 sg13g2_a21o_1 _15618_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[13] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[13] ),
    .B1(_01875_),
    .X(_01878_));
 sg13g2_o21ai_1 _15619_ (.B1(_01878_),
    .Y(_01879_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[13] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_nor2b_1 _15620_ (.A(_01879_),
    .B_N(_01877_),
    .Y(_01880_));
 sg13g2_xnor2_1 _15621_ (.Y(_01078_),
    .A(_01877_),
    .B(_01879_));
 sg13g2_a21o_1 _15622_ (.A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[14] ),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[14] ),
    .B1(_01880_),
    .X(_01881_));
 sg13g2_nand2_1 _15623_ (.Y(_01882_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[15] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_xnor2_1 _15624_ (.Y(_01883_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[15] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_xnor2_1 _15625_ (.Y(_01079_),
    .A(_01881_),
    .B(_01883_));
 sg13g2_nand2_1 _15626_ (.Y(_01884_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[16] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_xor2_1 _15627_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[16] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[16] ),
    .X(_01885_));
 sg13g2_o21ai_1 _15628_ (.B1(_01881_),
    .Y(_01886_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[15] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_nand2_1 _15629_ (.Y(_01887_),
    .A(_01882_),
    .B(_01886_));
 sg13g2_nand2_1 _15630_ (.Y(_01888_),
    .A(_01885_),
    .B(_01887_));
 sg13g2_xor2_1 _15631_ (.B(_01887_),
    .A(_01885_),
    .X(_01080_));
 sg13g2_xnor2_1 _15632_ (.Y(_01889_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[17] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_a21oi_1 _15633_ (.A1(_01884_),
    .A2(_01888_),
    .Y(_01890_),
    .B1(_01889_));
 sg13g2_nand3_1 _15634_ (.B(_01888_),
    .C(_01889_),
    .A(_01884_),
    .Y(_01891_));
 sg13g2_nor2b_1 _15635_ (.A(_01890_),
    .B_N(_01891_),
    .Y(_01081_));
 sg13g2_a21oi_1 _15636_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[17] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[17] ),
    .Y(_01892_),
    .B1(_01890_));
 sg13g2_xor2_1 _15637_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[18] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[18] ),
    .X(_01893_));
 sg13g2_xnor2_1 _15638_ (.Y(_01082_),
    .A(_01892_),
    .B(_01893_));
 sg13g2_nor2b_1 _15639_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][1] ),
    .Y(_01894_));
 sg13g2_xnor2_1 _15640_ (.Y(_01895_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][1] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _15641_ (.B(_01895_),
    .A(_02517_),
    .X(_00914_));
 sg13g2_a21oi_1 _15642_ (.A1(_02517_),
    .A2(_01895_),
    .Y(_01896_),
    .B1(_01894_));
 sg13g2_xnor2_1 _15643_ (.Y(_01897_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][2] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _15644_ (.A(_01896_),
    .B_N(_01897_),
    .Y(_01898_));
 sg13g2_xnor2_1 _15645_ (.Y(_00915_),
    .A(_01896_),
    .B(_01897_));
 sg13g2_a21oi_1 _15646_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][2] ),
    .A2(_02473_),
    .Y(_01899_),
    .B1(_01898_));
 sg13g2_xnor2_1 _15647_ (.Y(_01900_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][3] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _15648_ (.A(_01899_),
    .B_N(_01900_),
    .Y(_01901_));
 sg13g2_xnor2_1 _15649_ (.Y(_00916_),
    .A(_01899_),
    .B(_01900_));
 sg13g2_a21oi_1 _15650_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][3] ),
    .A2(_02474_),
    .Y(_01902_),
    .B1(_01901_));
 sg13g2_xnor2_1 _15651_ (.Y(_01903_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][4] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _15652_ (.A(_01902_),
    .B_N(_01903_),
    .Y(_01904_));
 sg13g2_xnor2_1 _15653_ (.Y(_00917_),
    .A(_01902_),
    .B(_01903_));
 sg13g2_a21oi_1 _15654_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][4] ),
    .A2(_02475_),
    .Y(_01905_),
    .B1(_01904_));
 sg13g2_nand2b_1 _15655_ (.Y(_01906_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][5] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _15656_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][5] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[5] ),
    .Y(_01907_));
 sg13g2_xnor2_1 _15657_ (.Y(_01908_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][5] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_xnor2_1 _15658_ (.Y(_00918_),
    .A(_01905_),
    .B(_01908_));
 sg13g2_nor2b_1 _15659_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[6] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][6] ),
    .Y(_01909_));
 sg13g2_nand2b_1 _15660_ (.Y(_01910_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[6] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][6] ));
 sg13g2_nand2b_1 _15661_ (.Y(_01911_),
    .B(_01910_),
    .A_N(_01909_));
 sg13g2_o21ai_1 _15662_ (.B1(_01906_),
    .Y(_01912_),
    .A1(_01905_),
    .A2(_01907_));
 sg13g2_xnor2_1 _15663_ (.Y(_00919_),
    .A(_01911_),
    .B(_01912_));
 sg13g2_a21oi_1 _15664_ (.A1(_01910_),
    .A2(_01912_),
    .Y(_01913_),
    .B1(_01909_));
 sg13g2_xnor2_1 _15665_ (.Y(_01914_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][7] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nand2b_1 _15666_ (.Y(_01915_),
    .B(_01914_),
    .A_N(_01913_));
 sg13g2_xnor2_1 _15667_ (.Y(_00920_),
    .A(_01913_),
    .B(_01914_));
 sg13g2_o21ai_1 _15668_ (.B1(_01915_),
    .Y(_01916_),
    .A1(_02476_),
    .A2(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _15669_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[8] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][8] ),
    .Y(_01917_));
 sg13g2_nand2b_1 _15670_ (.Y(_01918_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[8] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][8] ));
 sg13g2_nand2b_1 _15671_ (.Y(_01919_),
    .B(_01918_),
    .A_N(_01917_));
 sg13g2_xnor2_1 _15672_ (.Y(_00921_),
    .A(_01916_),
    .B(_01919_));
 sg13g2_a21oi_2 _15673_ (.B1(_01917_),
    .Y(_01920_),
    .A2(_01918_),
    .A1(_01916_));
 sg13g2_nor2b_1 _15674_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][9] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[9] ),
    .Y(_01921_));
 sg13g2_nand2b_1 _15675_ (.Y(_01922_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][9] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _15676_ (.A(_01921_),
    .B_N(_01922_),
    .Y(_01923_));
 sg13g2_xnor2_1 _15677_ (.Y(_00922_),
    .A(_01920_),
    .B(_01923_));
 sg13g2_nor2b_1 _15678_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][10] ),
    .Y(_01924_));
 sg13g2_nand2b_1 _15679_ (.Y(_01925_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][10] ));
 sg13g2_nand2b_1 _15680_ (.Y(_01926_),
    .B(_01925_),
    .A_N(_01924_));
 sg13g2_a21oi_2 _15681_ (.B1(_01921_),
    .Y(_01927_),
    .A2(_01922_),
    .A1(_01920_));
 sg13g2_xnor2_1 _15682_ (.Y(_00905_),
    .A(_01926_),
    .B(_01927_));
 sg13g2_a21oi_2 _15683_ (.B1(_01924_),
    .Y(_01928_),
    .A2(_01927_),
    .A1(_01925_));
 sg13g2_nor2b_1 _15684_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][11] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[11] ),
    .Y(_01929_));
 sg13g2_nand2b_1 _15685_ (.Y(_01930_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][11] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _15686_ (.A(_01929_),
    .B_N(_01930_),
    .Y(_01931_));
 sg13g2_xnor2_1 _15687_ (.Y(_00906_),
    .A(_01928_),
    .B(_01931_));
 sg13g2_nor2b_1 _15688_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][12] ),
    .Y(_01932_));
 sg13g2_nand2b_1 _15689_ (.Y(_01933_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][12] ));
 sg13g2_nand2b_1 _15690_ (.Y(_01934_),
    .B(_01933_),
    .A_N(_01932_));
 sg13g2_a21oi_2 _15691_ (.B1(_01929_),
    .Y(_01935_),
    .A2(_01930_),
    .A1(_01928_));
 sg13g2_xnor2_1 _15692_ (.Y(_00907_),
    .A(_01934_),
    .B(_01935_));
 sg13g2_a21oi_2 _15693_ (.B1(_01932_),
    .Y(_01936_),
    .A2(_01935_),
    .A1(_01933_));
 sg13g2_nor2b_1 _15694_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][13] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[13] ),
    .Y(_01937_));
 sg13g2_nand2b_1 _15695_ (.Y(_01938_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][13] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _15696_ (.A(_01937_),
    .B_N(_01938_),
    .Y(_01939_));
 sg13g2_xnor2_1 _15697_ (.Y(_00908_),
    .A(_01936_),
    .B(_01939_));
 sg13g2_nor2b_1 _15698_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][14] ),
    .Y(_01940_));
 sg13g2_nand2b_1 _15699_ (.Y(_01941_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][14] ));
 sg13g2_nand2b_1 _15700_ (.Y(_01942_),
    .B(_01941_),
    .A_N(_01940_));
 sg13g2_a21oi_2 _15701_ (.B1(_01937_),
    .Y(_01943_),
    .A2(_01938_),
    .A1(_01936_));
 sg13g2_xnor2_1 _15702_ (.Y(_00909_),
    .A(_01942_),
    .B(_01943_));
 sg13g2_a21oi_2 _15703_ (.B1(_01940_),
    .Y(_01944_),
    .A2(_01943_),
    .A1(_01941_));
 sg13g2_nor2b_1 _15704_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][15] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[15] ),
    .Y(_01945_));
 sg13g2_nand2b_1 _15705_ (.Y(_01946_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][15] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _15706_ (.A(_01945_),
    .B_N(_01946_),
    .Y(_01947_));
 sg13g2_xnor2_1 _15707_ (.Y(_00910_),
    .A(_01944_),
    .B(_01947_));
 sg13g2_xor2_1 _15708_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][16] ),
    .X(_01948_));
 sg13g2_a21oi_1 _15709_ (.A1(_01944_),
    .A2(_01946_),
    .Y(_01949_),
    .B1(_01945_));
 sg13g2_nor2b_1 _15710_ (.A(_01948_),
    .B_N(_01949_),
    .Y(_01950_));
 sg13g2_xnor2_1 _15711_ (.Y(_00911_),
    .A(_01948_),
    .B(_01949_));
 sg13g2_a21oi_1 _15712_ (.A1(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][16] ),
    .A2(_02477_),
    .Y(_01951_),
    .B1(_01950_));
 sg13g2_nand2b_1 _15713_ (.Y(_01952_),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][17] ),
    .A_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _15714_ (.A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][17] ),
    .B_N(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[17] ),
    .Y(_01953_));
 sg13g2_xnor2_1 _15715_ (.Y(_01954_),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][17] ),
    .B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _15716_ (.Y(_00912_),
    .A(_01951_),
    .B(_01954_));
 sg13g2_o21ai_1 _15717_ (.B1(_01952_),
    .Y(_01955_),
    .A1(_01951_),
    .A2(_01953_));
 sg13g2_xor2_1 _15718_ (.B(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][18] ),
    .X(_01956_));
 sg13g2_xnor2_1 _15719_ (.Y(_00913_),
    .A(_01955_),
    .B(_01956_));
 sg13g2_nor2b_1 _15720_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][1] ),
    .Y(_01957_));
 sg13g2_xnor2_1 _15721_ (.Y(_01958_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][1] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _15722_ (.B(_01958_),
    .A(_02518_),
    .X(_01121_));
 sg13g2_a21oi_2 _15723_ (.B1(_01957_),
    .Y(_01959_),
    .A2(_01958_),
    .A1(_02518_));
 sg13g2_xnor2_1 _15724_ (.Y(_01960_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][2] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _15725_ (.A(_01959_),
    .B_N(_01960_),
    .Y(_01961_));
 sg13g2_xnor2_1 _15726_ (.Y(_01122_),
    .A(_01959_),
    .B(_01960_));
 sg13g2_a21oi_1 _15727_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][2] ),
    .A2(_02478_),
    .Y(_01962_),
    .B1(_01961_));
 sg13g2_xnor2_1 _15728_ (.Y(_01963_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][3] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _15729_ (.A(_01962_),
    .B_N(_01963_),
    .Y(_01964_));
 sg13g2_xnor2_1 _15730_ (.Y(_01123_),
    .A(_01962_),
    .B(_01963_));
 sg13g2_a21oi_2 _15731_ (.B1(_01964_),
    .Y(_01965_),
    .A2(_02479_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][3] ));
 sg13g2_xnor2_1 _15732_ (.Y(_01966_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][4] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _15733_ (.A(_01965_),
    .B_N(_01966_),
    .Y(_01967_));
 sg13g2_xnor2_1 _15734_ (.Y(_01124_),
    .A(_01965_),
    .B(_01966_));
 sg13g2_a21oi_2 _15735_ (.B1(_01967_),
    .Y(_01968_),
    .A2(_02480_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][4] ));
 sg13g2_nand2b_1 _15736_ (.Y(_01969_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][5] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _15737_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][5] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[5] ),
    .Y(_01970_));
 sg13g2_xnor2_1 _15738_ (.Y(_01971_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][5] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_xnor2_1 _15739_ (.Y(_01125_),
    .A(_01968_),
    .B(_01971_));
 sg13g2_nor2b_1 _15740_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][6] ),
    .Y(_01972_));
 sg13g2_nand2b_1 _15741_ (.Y(_01973_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][6] ));
 sg13g2_nand2b_1 _15742_ (.Y(_01974_),
    .B(_01973_),
    .A_N(_01972_));
 sg13g2_o21ai_1 _15743_ (.B1(_01969_),
    .Y(_01975_),
    .A1(_01968_),
    .A2(_01970_));
 sg13g2_xnor2_1 _15744_ (.Y(_01126_),
    .A(_01974_),
    .B(_01975_));
 sg13g2_a21oi_1 _15745_ (.A1(_01973_),
    .A2(_01975_),
    .Y(_01976_),
    .B1(_01972_));
 sg13g2_xnor2_1 _15746_ (.Y(_01977_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][7] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nand2b_1 _15747_ (.Y(_01978_),
    .B(_01977_),
    .A_N(_01976_));
 sg13g2_xnor2_1 _15748_ (.Y(_01127_),
    .A(_01976_),
    .B(_01977_));
 sg13g2_o21ai_1 _15749_ (.B1(_01978_),
    .Y(_01979_),
    .A1(_02481_),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _15750_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][8] ),
    .Y(_01980_));
 sg13g2_nand2b_1 _15751_ (.Y(_01981_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][8] ));
 sg13g2_nand2b_1 _15752_ (.Y(_01982_),
    .B(_01981_),
    .A_N(_01980_));
 sg13g2_xnor2_1 _15753_ (.Y(_01128_),
    .A(_01979_),
    .B(_01982_));
 sg13g2_nand2b_1 _15754_ (.Y(_01983_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][9] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _15755_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][9] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[9] ),
    .Y(_01984_));
 sg13g2_xnor2_1 _15756_ (.Y(_01985_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][9] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_a21oi_1 _15757_ (.A1(_01979_),
    .A2(_01981_),
    .Y(_01986_),
    .B1(_01980_));
 sg13g2_xnor2_1 _15758_ (.Y(_01129_),
    .A(_01985_),
    .B(_01986_));
 sg13g2_nor2b_1 _15759_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][10] ),
    .Y(_01987_));
 sg13g2_nand2b_1 _15760_ (.Y(_01988_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][10] ));
 sg13g2_nand2b_1 _15761_ (.Y(_01989_),
    .B(_01988_),
    .A_N(_01987_));
 sg13g2_o21ai_1 _15762_ (.B1(_01983_),
    .Y(_01990_),
    .A1(_01984_),
    .A2(_01986_));
 sg13g2_xnor2_1 _15763_ (.Y(_01112_),
    .A(_01989_),
    .B(_01990_));
 sg13g2_nand2b_1 _15764_ (.Y(_01991_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][11] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _15765_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][11] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[11] ),
    .Y(_01992_));
 sg13g2_xnor2_1 _15766_ (.Y(_01993_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][11] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_a21oi_2 _15767_ (.B1(_01987_),
    .Y(_01994_),
    .A2(_01990_),
    .A1(_01988_));
 sg13g2_xnor2_1 _15768_ (.Y(_01113_),
    .A(_01993_),
    .B(_01994_));
 sg13g2_nor2b_1 _15769_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][12] ),
    .Y(_01995_));
 sg13g2_nand2b_1 _15770_ (.Y(_01996_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][12] ));
 sg13g2_nand2b_1 _15771_ (.Y(_01997_),
    .B(_01996_),
    .A_N(_01995_));
 sg13g2_o21ai_1 _15772_ (.B1(_01991_),
    .Y(_01998_),
    .A1(_01992_),
    .A2(_01994_));
 sg13g2_xnor2_1 _15773_ (.Y(_01114_),
    .A(_01997_),
    .B(_01998_));
 sg13g2_nand2b_1 _15774_ (.Y(_01999_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][13] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _15775_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][13] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[13] ),
    .Y(_02000_));
 sg13g2_xnor2_1 _15776_ (.Y(_02001_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][13] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_a21oi_2 _15777_ (.B1(_01995_),
    .Y(_02002_),
    .A2(_01998_),
    .A1(_01996_));
 sg13g2_xnor2_1 _15778_ (.Y(_01115_),
    .A(_02001_),
    .B(_02002_));
 sg13g2_nor2b_1 _15779_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][14] ),
    .Y(_02003_));
 sg13g2_nand2b_1 _15780_ (.Y(_02004_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][14] ));
 sg13g2_nand2b_1 _15781_ (.Y(_02005_),
    .B(_02004_),
    .A_N(_02003_));
 sg13g2_o21ai_1 _15782_ (.B1(_01999_),
    .Y(_02006_),
    .A1(_02000_),
    .A2(_02002_));
 sg13g2_xnor2_1 _15783_ (.Y(_01116_),
    .A(_02005_),
    .B(_02006_));
 sg13g2_nand2b_1 _15784_ (.Y(_02007_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][15] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _15785_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][15] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[15] ),
    .Y(_02008_));
 sg13g2_xnor2_1 _15786_ (.Y(_02009_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][15] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_a21oi_2 _15787_ (.B1(_02003_),
    .Y(_02010_),
    .A2(_02006_),
    .A1(_02004_));
 sg13g2_xnor2_1 _15788_ (.Y(_01117_),
    .A(_02009_),
    .B(_02010_));
 sg13g2_xor2_1 _15789_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][16] ),
    .X(_02011_));
 sg13g2_o21ai_1 _15790_ (.B1(_02007_),
    .Y(_02012_),
    .A1(_02008_),
    .A2(_02010_));
 sg13g2_nor2b_1 _15791_ (.A(_02011_),
    .B_N(_02012_),
    .Y(_02013_));
 sg13g2_xnor2_1 _15792_ (.Y(_01118_),
    .A(_02011_),
    .B(_02012_));
 sg13g2_a21oi_2 _15793_ (.B1(_02013_),
    .Y(_02014_),
    .A2(_02482_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][16] ));
 sg13g2_nand2b_1 _15794_ (.Y(_02015_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][17] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _15795_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][17] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[17] ),
    .Y(_02016_));
 sg13g2_xnor2_1 _15796_ (.Y(_02017_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][17] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _15797_ (.Y(_01119_),
    .A(_02014_),
    .B(_02017_));
 sg13g2_o21ai_1 _15798_ (.B1(_02015_),
    .Y(_02018_),
    .A1(_02014_),
    .A2(_02016_));
 sg13g2_xor2_1 _15799_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][18] ),
    .X(_02019_));
 sg13g2_xnor2_1 _15800_ (.Y(_01120_),
    .A(_02018_),
    .B(_02019_));
 sg13g2_nor2b_1 _15801_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][1] ),
    .Y(_02020_));
 sg13g2_xnor2_1 _15802_ (.Y(_02021_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][1] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _15803_ (.B(_02021_),
    .A(_02519_),
    .X(_01102_));
 sg13g2_a21oi_2 _15804_ (.B1(_02020_),
    .Y(_02022_),
    .A2(_02021_),
    .A1(_02519_));
 sg13g2_xnor2_1 _15805_ (.Y(_02023_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][2] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _15806_ (.A(_02022_),
    .B_N(_02023_),
    .Y(_02024_));
 sg13g2_xnor2_1 _15807_ (.Y(_01103_),
    .A(_02022_),
    .B(_02023_));
 sg13g2_a21oi_2 _15808_ (.B1(_02024_),
    .Y(_02025_),
    .A2(_02483_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][2] ));
 sg13g2_xnor2_1 _15809_ (.Y(_02026_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][3] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _15810_ (.A(_02025_),
    .B_N(_02026_),
    .Y(_02027_));
 sg13g2_xnor2_1 _15811_ (.Y(_01104_),
    .A(_02025_),
    .B(_02026_));
 sg13g2_a21oi_2 _15812_ (.B1(_02027_),
    .Y(_02028_),
    .A2(_02484_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][3] ));
 sg13g2_xnor2_1 _15813_ (.Y(_02029_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][4] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _15814_ (.A(_02028_),
    .B_N(_02029_),
    .Y(_02030_));
 sg13g2_xnor2_1 _15815_ (.Y(_01105_),
    .A(_02028_),
    .B(_02029_));
 sg13g2_a21oi_2 _15816_ (.B1(_02030_),
    .Y(_02031_),
    .A2(_02485_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][4] ));
 sg13g2_xnor2_1 _15817_ (.Y(_02032_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][5] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _15818_ (.A(_02031_),
    .B_N(_02032_),
    .Y(_02033_));
 sg13g2_xnor2_1 _15819_ (.Y(_01106_),
    .A(_02031_),
    .B(_02032_));
 sg13g2_a21oi_1 _15820_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][5] ),
    .A2(_02486_),
    .Y(_02034_),
    .B1(_02033_));
 sg13g2_xnor2_1 _15821_ (.Y(_02035_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][6] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_nor2b_1 _15822_ (.A(_02034_),
    .B_N(_02035_),
    .Y(_02036_));
 sg13g2_xnor2_1 _15823_ (.Y(_01107_),
    .A(_02034_),
    .B(_02035_));
 sg13g2_a21oi_1 _15824_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][6] ),
    .A2(_02487_),
    .Y(_02037_),
    .B1(_02036_));
 sg13g2_xnor2_1 _15825_ (.Y(_02038_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][7] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _15826_ (.A(_02037_),
    .B_N(_02038_),
    .Y(_02039_));
 sg13g2_xnor2_1 _15827_ (.Y(_01108_),
    .A(_02037_),
    .B(_02038_));
 sg13g2_a21oi_1 _15828_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][7] ),
    .A2(_02488_),
    .Y(_02040_),
    .B1(_02039_));
 sg13g2_xnor2_1 _15829_ (.Y(_02041_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][8] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_nor2b_1 _15830_ (.A(_02040_),
    .B_N(_02041_),
    .Y(_02042_));
 sg13g2_xnor2_1 _15831_ (.Y(_01109_),
    .A(_02040_),
    .B(_02041_));
 sg13g2_a21oi_2 _15832_ (.B1(_02042_),
    .Y(_02043_),
    .A2(_02489_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][8] ));
 sg13g2_nor2b_1 _15833_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][9] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[9] ),
    .Y(_02044_));
 sg13g2_nand2b_1 _15834_ (.Y(_02045_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][9] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _15835_ (.A(_02044_),
    .B_N(_02045_),
    .Y(_02046_));
 sg13g2_xnor2_1 _15836_ (.Y(_01110_),
    .A(_02043_),
    .B(_02046_));
 sg13g2_nor2b_1 _15837_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][10] ),
    .Y(_02047_));
 sg13g2_nand2b_1 _15838_ (.Y(_02048_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][10] ));
 sg13g2_nand2b_1 _15839_ (.Y(_02049_),
    .B(_02048_),
    .A_N(_02047_));
 sg13g2_a21oi_2 _15840_ (.B1(_02044_),
    .Y(_02050_),
    .A2(_02045_),
    .A1(_02043_));
 sg13g2_xnor2_1 _15841_ (.Y(_01093_),
    .A(_02049_),
    .B(_02050_));
 sg13g2_a21oi_2 _15842_ (.B1(_02047_),
    .Y(_02051_),
    .A2(_02050_),
    .A1(_02048_));
 sg13g2_nand2b_1 _15843_ (.Y(_02052_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][11] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _15844_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][11] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[11] ),
    .Y(_02053_));
 sg13g2_xnor2_1 _15845_ (.Y(_02054_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][11] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_xnor2_1 _15846_ (.Y(_01094_),
    .A(_02051_),
    .B(_02054_));
 sg13g2_nor2b_1 _15847_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][12] ),
    .Y(_02055_));
 sg13g2_nand2b_1 _15848_ (.Y(_02056_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][12] ));
 sg13g2_nand2b_1 _15849_ (.Y(_02057_),
    .B(_02056_),
    .A_N(_02055_));
 sg13g2_a21oi_2 _15850_ (.B1(_02053_),
    .Y(_02058_),
    .A2(_02052_),
    .A1(_02051_));
 sg13g2_xnor2_1 _15851_ (.Y(_01095_),
    .A(_02057_),
    .B(_02058_));
 sg13g2_a21oi_2 _15852_ (.B1(_02055_),
    .Y(_02059_),
    .A2(_02058_),
    .A1(_02056_));
 sg13g2_nor2b_1 _15853_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][13] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[13] ),
    .Y(_02060_));
 sg13g2_nand2b_1 _15854_ (.Y(_02061_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][13] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _15855_ (.A(_02060_),
    .B_N(_02061_),
    .Y(_02062_));
 sg13g2_xnor2_1 _15856_ (.Y(_01096_),
    .A(_02059_),
    .B(_02062_));
 sg13g2_nor2b_1 _15857_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][14] ),
    .Y(_02063_));
 sg13g2_nand2b_1 _15858_ (.Y(_02064_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][14] ));
 sg13g2_nand2b_1 _15859_ (.Y(_02065_),
    .B(_02064_),
    .A_N(_02063_));
 sg13g2_a21oi_1 _15860_ (.A1(_02059_),
    .A2(_02061_),
    .Y(_02066_),
    .B1(_02060_));
 sg13g2_xnor2_1 _15861_ (.Y(_01097_),
    .A(_02065_),
    .B(_02066_));
 sg13g2_a21oi_1 _15862_ (.A1(_02064_),
    .A2(_02066_),
    .Y(_02067_),
    .B1(_02063_));
 sg13g2_nor2b_1 _15863_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][15] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[15] ),
    .Y(_02068_));
 sg13g2_nand2b_1 _15864_ (.Y(_02069_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][15] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _15865_ (.A(_02068_),
    .B_N(_02069_),
    .Y(_02070_));
 sg13g2_xnor2_1 _15866_ (.Y(_01098_),
    .A(_02067_),
    .B(_02070_));
 sg13g2_xor2_1 _15867_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][16] ),
    .X(_02071_));
 sg13g2_a21oi_1 _15868_ (.A1(_02067_),
    .A2(_02069_),
    .Y(_02072_),
    .B1(_02068_));
 sg13g2_nor2b_1 _15869_ (.A(_02071_),
    .B_N(_02072_),
    .Y(_02073_));
 sg13g2_xnor2_1 _15870_ (.Y(_01099_),
    .A(_02071_),
    .B(_02072_));
 sg13g2_a21oi_1 _15871_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][16] ),
    .A2(_02490_),
    .Y(_02074_),
    .B1(_02073_));
 sg13g2_nand2b_1 _15872_ (.Y(_02075_),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][17] ),
    .A_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _15873_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][17] ),
    .B_N(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[17] ),
    .Y(_02076_));
 sg13g2_xnor2_1 _15874_ (.Y(_02077_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][17] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _15875_ (.Y(_01100_),
    .A(_02074_),
    .B(_02077_));
 sg13g2_o21ai_1 _15876_ (.B1(_02075_),
    .Y(_02078_),
    .A1(_02074_),
    .A2(_02076_));
 sg13g2_xor2_1 _15877_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][18] ),
    .X(_02079_));
 sg13g2_xnor2_1 _15878_ (.Y(_01101_),
    .A(_02078_),
    .B(_02079_));
 sg13g2_and2_1 _15879_ (.A(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.u_mux_shift.sum_res ),
    .B(net4927),
    .X(_00191_));
 sg13g2_and2_1 _15880_ (.A(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ),
    .B(net4928),
    .X(_00159_));
 sg13g2_and2_1 _15881_ (.A(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.u_mux_shift.sum_res ),
    .B(net4932),
    .X(_00127_));
 sg13g2_and2_1 _15882_ (.A(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.u_mux_shift.sum_res ),
    .B(net4929),
    .X(_00095_));
 sg13g2_and2_1 _15883_ (.A(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.u_mux_shift.sum_res ),
    .B(net4927),
    .X(_00063_));
 sg13g2_and2_1 _15884_ (.A(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.u_mux_shift.sum_res ),
    .B(net4928),
    .X(_00031_));
 sg13g2_nand2_1 _15885_ (.Y(_02080_),
    .A(net4929),
    .B(_02846_));
 sg13g2_a21oi_1 _15886_ (.A1(_02755_),
    .A2(_02844_),
    .Y(_00287_),
    .B1(_02080_));
 sg13g2_nor2b_1 _15887_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][1] ),
    .Y(_02081_));
 sg13g2_xnor2_1 _15888_ (.Y(_02082_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][1] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _15889_ (.B(_02082_),
    .A(_02505_),
    .X(_00444_));
 sg13g2_a21oi_1 _15890_ (.A1(_02505_),
    .A2(_02082_),
    .Y(_02083_),
    .B1(_02081_));
 sg13g2_xnor2_1 _15891_ (.Y(_02084_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][2] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _15892_ (.A(_02083_),
    .B_N(_02084_),
    .Y(_02085_));
 sg13g2_xnor2_1 _15893_ (.Y(_00445_),
    .A(_02083_),
    .B(_02084_));
 sg13g2_a21oi_1 _15894_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][2] ),
    .A2(_02491_),
    .Y(_02086_),
    .B1(_02085_));
 sg13g2_xnor2_1 _15895_ (.Y(_02087_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][3] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _15896_ (.A(_02086_),
    .B_N(_02087_),
    .Y(_02088_));
 sg13g2_xnor2_1 _15897_ (.Y(_00446_),
    .A(_02086_),
    .B(_02087_));
 sg13g2_a21oi_1 _15898_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][3] ),
    .A2(_02492_),
    .Y(_02089_),
    .B1(_02088_));
 sg13g2_xnor2_1 _15899_ (.Y(_02090_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][4] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _15900_ (.A(_02089_),
    .B_N(_02090_),
    .Y(_02091_));
 sg13g2_xnor2_1 _15901_ (.Y(_00447_),
    .A(_02089_),
    .B(_02090_));
 sg13g2_a21oi_1 _15902_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][4] ),
    .A2(_02493_),
    .Y(_02092_),
    .B1(_02091_));
 sg13g2_xnor2_1 _15903_ (.Y(_02093_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][5] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _15904_ (.A(_02092_),
    .B_N(_02093_),
    .Y(_02094_));
 sg13g2_xnor2_1 _15905_ (.Y(_00448_),
    .A(_02092_),
    .B(_02093_));
 sg13g2_a21oi_1 _15906_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][5] ),
    .A2(_02494_),
    .Y(_02095_),
    .B1(_02094_));
 sg13g2_xnor2_1 _15907_ (.Y(_02096_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][6] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_nor2b_1 _15908_ (.A(_02095_),
    .B_N(_02096_),
    .Y(_02097_));
 sg13g2_xnor2_1 _15909_ (.Y(_00449_),
    .A(_02095_),
    .B(_02096_));
 sg13g2_a21oi_1 _15910_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][6] ),
    .A2(_02495_),
    .Y(_02098_),
    .B1(_02097_));
 sg13g2_xnor2_1 _15911_ (.Y(_02099_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][7] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _15912_ (.A(_02098_),
    .B_N(_02099_),
    .Y(_02100_));
 sg13g2_xnor2_1 _15913_ (.Y(_00450_),
    .A(_02098_),
    .B(_02099_));
 sg13g2_a21oi_1 _15914_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][7] ),
    .A2(_02496_),
    .Y(_02101_),
    .B1(_02100_));
 sg13g2_xnor2_1 _15915_ (.Y(_02102_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][8] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_nor2b_1 _15916_ (.A(_02101_),
    .B_N(_02102_),
    .Y(_02103_));
 sg13g2_xnor2_1 _15917_ (.Y(_00451_),
    .A(_02101_),
    .B(_02102_));
 sg13g2_nand2b_1 _15918_ (.Y(_02104_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][9] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _15919_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][9] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[9] ),
    .Y(_02105_));
 sg13g2_xnor2_1 _15920_ (.Y(_02106_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][9] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_a21oi_2 _15921_ (.B1(_02103_),
    .Y(_02107_),
    .A2(_02497_),
    .A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][8] ));
 sg13g2_xnor2_1 _15922_ (.Y(_00452_),
    .A(_02106_),
    .B(_02107_));
 sg13g2_nor2b_1 _15923_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][10] ),
    .Y(_02108_));
 sg13g2_nand2b_1 _15924_ (.Y(_02109_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][10] ));
 sg13g2_nand2b_1 _15925_ (.Y(_02110_),
    .B(_02109_),
    .A_N(_02108_));
 sg13g2_o21ai_1 _15926_ (.B1(_02104_),
    .Y(_02111_),
    .A1(_02105_),
    .A2(_02107_));
 sg13g2_xnor2_1 _15927_ (.Y(_00435_),
    .A(_02110_),
    .B(_02111_));
 sg13g2_nand2b_1 _15928_ (.Y(_02112_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][11] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _15929_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][11] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[11] ),
    .Y(_02113_));
 sg13g2_xnor2_1 _15930_ (.Y(_02114_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][11] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_a21oi_1 _15931_ (.A1(_02109_),
    .A2(_02111_),
    .Y(_02115_),
    .B1(_02108_));
 sg13g2_xnor2_1 _15932_ (.Y(_00436_),
    .A(_02114_),
    .B(_02115_));
 sg13g2_nor2b_1 _15933_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][12] ),
    .Y(_02116_));
 sg13g2_nand2b_1 _15934_ (.Y(_02117_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][12] ));
 sg13g2_nand2b_1 _15935_ (.Y(_02118_),
    .B(_02117_),
    .A_N(_02116_));
 sg13g2_o21ai_1 _15936_ (.B1(_02112_),
    .Y(_02119_),
    .A1(_02113_),
    .A2(_02115_));
 sg13g2_xnor2_1 _15937_ (.Y(_00437_),
    .A(_02118_),
    .B(_02119_));
 sg13g2_a21oi_1 _15938_ (.A1(_02117_),
    .A2(_02119_),
    .Y(_02120_),
    .B1(_02116_));
 sg13g2_nor2b_1 _15939_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][13] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[13] ),
    .Y(_02121_));
 sg13g2_nand2b_1 _15940_ (.Y(_02122_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][13] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _15941_ (.A(_02121_),
    .B_N(_02122_),
    .Y(_02123_));
 sg13g2_xnor2_1 _15942_ (.Y(_00438_),
    .A(_02120_),
    .B(_02123_));
 sg13g2_nor2b_1 _15943_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][14] ),
    .Y(_02124_));
 sg13g2_nand2b_1 _15944_ (.Y(_02125_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][14] ));
 sg13g2_nand2b_1 _15945_ (.Y(_02126_),
    .B(_02125_),
    .A_N(_02124_));
 sg13g2_a21oi_1 _15946_ (.A1(_02120_),
    .A2(_02122_),
    .Y(_02127_),
    .B1(_02121_));
 sg13g2_xnor2_1 _15947_ (.Y(_00439_),
    .A(_02126_),
    .B(_02127_));
 sg13g2_a21oi_1 _15948_ (.A1(_02125_),
    .A2(_02127_),
    .Y(_02128_),
    .B1(_02124_));
 sg13g2_nor2b_1 _15949_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][15] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[15] ),
    .Y(_02129_));
 sg13g2_nand2b_1 _15950_ (.Y(_02130_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][15] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _15951_ (.A(_02129_),
    .B_N(_02130_),
    .Y(_02131_));
 sg13g2_xnor2_1 _15952_ (.Y(_00440_),
    .A(_02128_),
    .B(_02131_));
 sg13g2_xor2_1 _15953_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][16] ),
    .X(_02132_));
 sg13g2_a21oi_1 _15954_ (.A1(_02128_),
    .A2(_02130_),
    .Y(_02133_),
    .B1(_02129_));
 sg13g2_nor2b_1 _15955_ (.A(_02132_),
    .B_N(_02133_),
    .Y(_02134_));
 sg13g2_xnor2_1 _15956_ (.Y(_00441_),
    .A(_02132_),
    .B(_02133_));
 sg13g2_a21oi_1 _15957_ (.A1(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][16] ),
    .A2(_02498_),
    .Y(_02135_),
    .B1(_02134_));
 sg13g2_nand2b_1 _15958_ (.Y(_02136_),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][17] ),
    .A_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _15959_ (.A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][17] ),
    .B_N(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[17] ),
    .Y(_02137_));
 sg13g2_xnor2_1 _15960_ (.Y(_02138_),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][17] ),
    .B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _15961_ (.Y(_00442_),
    .A(_02135_),
    .B(_02138_));
 sg13g2_o21ai_1 _15962_ (.B1(_02136_),
    .Y(_02139_),
    .A1(_02135_),
    .A2(_02137_));
 sg13g2_xor2_1 _15963_ (.B(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][18] ),
    .X(_02140_));
 sg13g2_xnor2_1 _15964_ (.Y(_00443_),
    .A(_02139_),
    .B(_02140_));
 sg13g2_nand2b_1 _15965_ (.Y(_02141_),
    .B(net4965),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_nor2b_1 _15966_ (.A(net4965),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[1] ),
    .Y(_02142_));
 sg13g2_xnor2_1 _15967_ (.Y(_02143_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[1] ),
    .B(net4965));
 sg13g2_xnor2_1 _15968_ (.Y(_01045_),
    .A(_01187_),
    .B(_02143_));
 sg13g2_xnor2_1 _15969_ (.Y(_02144_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[2] ),
    .B(net4965));
 sg13g2_o21ai_1 _15970_ (.B1(_02141_),
    .Y(_02145_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[0] ),
    .A2(_02142_));
 sg13g2_nor2b_1 _15971_ (.A(_02145_),
    .B_N(_02144_),
    .Y(_02146_));
 sg13g2_xnor2_1 _15972_ (.Y(_01046_),
    .A(_02144_),
    .B(_02145_));
 sg13g2_a21oi_1 _15973_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[2] ),
    .A2(net4935),
    .Y(_02147_),
    .B1(_02146_));
 sg13g2_nor2_1 _15974_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4935),
    .Y(_02148_));
 sg13g2_nand2_1 _15975_ (.Y(_02149_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[3] ),
    .B(net4935));
 sg13g2_nor2b_1 _15976_ (.A(_02148_),
    .B_N(_02149_),
    .Y(_02150_));
 sg13g2_xnor2_1 _15977_ (.Y(_01047_),
    .A(_02147_),
    .B(_02150_));
 sg13g2_xnor2_1 _15978_ (.Y(_02151_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[4] ),
    .B(net4966));
 sg13g2_o21ai_1 _15979_ (.B1(_02149_),
    .Y(_02152_),
    .A1(_02147_),
    .A2(_02148_));
 sg13g2_and2_1 _15980_ (.A(_02151_),
    .B(_02152_),
    .X(_02153_));
 sg13g2_xor2_1 _15981_ (.B(_02152_),
    .A(_02151_),
    .X(_01048_));
 sg13g2_xnor2_1 _15982_ (.Y(_02154_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[5] ),
    .B(net4965));
 sg13g2_a21oi_1 _15983_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[4] ),
    .A2(net4935),
    .Y(_02155_),
    .B1(_02153_));
 sg13g2_xnor2_1 _15984_ (.Y(_01049_),
    .A(_02154_),
    .B(_02155_));
 sg13g2_o21ai_1 _15985_ (.B1(net4935),
    .Y(_02156_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[4] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_and2_1 _15986_ (.A(_02153_),
    .B(_02154_),
    .X(_02157_));
 sg13g2_nor2b_1 _15987_ (.A(_02157_),
    .B_N(_02156_),
    .Y(_02158_));
 sg13g2_nand2_1 _15988_ (.Y(_02159_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4935));
 sg13g2_nor2_1 _15989_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4935),
    .Y(_02160_));
 sg13g2_xnor2_1 _15990_ (.Y(_02161_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[6] ),
    .B(net4965));
 sg13g2_xnor2_1 _15991_ (.Y(_01050_),
    .A(_02158_),
    .B(_02161_));
 sg13g2_nand2b_1 _15992_ (.Y(_02162_),
    .B(net4965),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_xor2_1 _15993_ (.B(net4965),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[7] ),
    .X(_02163_));
 sg13g2_o21ai_1 _15994_ (.B1(_02159_),
    .Y(_02164_),
    .A1(_02158_),
    .A2(_02160_));
 sg13g2_xnor2_1 _15995_ (.Y(_01051_),
    .A(_02163_),
    .B(_02164_));
 sg13g2_xnor2_1 _15996_ (.Y(_02165_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[8] ),
    .B(net4966));
 sg13g2_o21ai_1 _15997_ (.B1(net4934),
    .Y(_02166_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_nand3_1 _15998_ (.B(_02161_),
    .C(_02162_),
    .A(_02157_),
    .Y(_02167_));
 sg13g2_and3_1 _15999_ (.X(_02168_),
    .A(_02156_),
    .B(_02166_),
    .C(_02167_));
 sg13g2_nand2b_1 _16000_ (.Y(_02169_),
    .B(_02165_),
    .A_N(_02168_));
 sg13g2_xnor2_1 _16001_ (.Y(_01052_),
    .A(_02165_),
    .B(_02168_));
 sg13g2_xor2_1 _16002_ (.B(net4966),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[9] ),
    .X(_02170_));
 sg13g2_o21ai_1 _16003_ (.B1(_02169_),
    .Y(_02171_),
    .A1(_02389_),
    .A2(net4966));
 sg13g2_xnor2_1 _16004_ (.Y(_01053_),
    .A(_02170_),
    .B(_02171_));
 sg13g2_o21ai_1 _16005_ (.B1(net4934),
    .Y(_02172_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[8] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_nor2_1 _16006_ (.A(_02169_),
    .B(_02170_),
    .Y(_02173_));
 sg13g2_nor2b_1 _16007_ (.A(_02173_),
    .B_N(_02172_),
    .Y(_02174_));
 sg13g2_nand2_1 _16008_ (.Y(_02175_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4934));
 sg13g2_nor2_1 _16009_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4934),
    .Y(_02176_));
 sg13g2_xnor2_1 _16010_ (.Y(_02177_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[10] ),
    .B(net4964));
 sg13g2_xnor2_1 _16011_ (.Y(_01036_),
    .A(_02174_),
    .B(_02177_));
 sg13g2_xor2_1 _16012_ (.B(net4963),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[11] ),
    .X(_02178_));
 sg13g2_o21ai_1 _16013_ (.B1(_02175_),
    .Y(_02179_),
    .A1(_02174_),
    .A2(_02176_));
 sg13g2_xnor2_1 _16014_ (.Y(_01037_),
    .A(_02178_),
    .B(_02179_));
 sg13g2_xnor2_1 _16015_ (.Y(_02180_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[12] ),
    .B(net4963));
 sg13g2_nand2_1 _16016_ (.Y(_02181_),
    .A(_02173_),
    .B(_02177_));
 sg13g2_nor2_1 _16017_ (.A(_02178_),
    .B(_02181_),
    .Y(_02182_));
 sg13g2_o21ai_1 _16018_ (.B1(net4934),
    .Y(_02183_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[10] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_nand2_1 _16019_ (.Y(_02184_),
    .A(_02172_),
    .B(_02183_));
 sg13g2_inv_1 _16020_ (.Y(_02185_),
    .A(_02184_));
 sg13g2_o21ai_1 _16021_ (.B1(_02180_),
    .Y(_02186_),
    .A1(_02182_),
    .A2(_02184_));
 sg13g2_or3_1 _16022_ (.A(_02180_),
    .B(_02182_),
    .C(_02184_),
    .X(_02187_));
 sg13g2_and2_1 _16023_ (.A(_02186_),
    .B(_02187_),
    .X(_01038_));
 sg13g2_nand2_1 _16024_ (.Y(_02188_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[13] ),
    .B(net4934));
 sg13g2_nand2_1 _16025_ (.Y(_02189_),
    .A(_02391_),
    .B(net4963));
 sg13g2_nand2_1 _16026_ (.Y(_02190_),
    .A(_02188_),
    .B(_02189_));
 sg13g2_o21ai_1 _16027_ (.B1(_02186_),
    .Y(_02191_),
    .A1(_02390_),
    .A2(net4963));
 sg13g2_xnor2_1 _16028_ (.Y(_01039_),
    .A(_02190_),
    .B(_02191_));
 sg13g2_nor2b_1 _16029_ (.A(net4963),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[14] ),
    .Y(_02192_));
 sg13g2_xnor2_1 _16030_ (.Y(_02193_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[14] ),
    .B(net4963));
 sg13g2_o21ai_1 _16031_ (.B1(net4934),
    .Y(_02194_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[12] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_a22oi_1 _16032_ (.Y(_02195_),
    .B1(_02186_),
    .B2(_02194_),
    .A2(net4963),
    .A1(_02391_));
 sg13g2_xor2_1 _16033_ (.B(_02195_),
    .A(_02193_),
    .X(_01040_));
 sg13g2_xnor2_1 _16034_ (.Y(_02196_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[15] ),
    .B(net4964));
 sg13g2_a21oi_1 _16035_ (.A1(_02193_),
    .A2(_02195_),
    .Y(_02197_),
    .B1(_02192_));
 sg13g2_xnor2_1 _16036_ (.Y(_01041_),
    .A(_02196_),
    .B(_02197_));
 sg13g2_and4_1 _16037_ (.A(_02180_),
    .B(_02188_),
    .C(_02189_),
    .D(_02193_),
    .X(_02198_));
 sg13g2_nand3_1 _16038_ (.B(_02196_),
    .C(_02198_),
    .A(_02182_),
    .Y(_02199_));
 sg13g2_o21ai_1 _16039_ (.B1(net4934),
    .Y(_02200_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[14] ),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_nand4_1 _16040_ (.B(_02194_),
    .C(_02199_),
    .A(_02185_),
    .Y(_02201_),
    .D(_02200_));
 sg13g2_nor2b_1 _16041_ (.A(net4964),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[16] ),
    .Y(_02202_));
 sg13g2_xnor2_1 _16042_ (.Y(_02203_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[16] ),
    .B(net4964));
 sg13g2_xor2_1 _16043_ (.B(_02203_),
    .A(_02201_),
    .X(_01042_));
 sg13g2_a21o_1 _16044_ (.A2(_02203_),
    .A1(_02201_),
    .B1(_02202_),
    .X(_02204_));
 sg13g2_xor2_1 _16045_ (.B(net4964),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[17] ),
    .X(_02205_));
 sg13g2_xnor2_1 _16046_ (.Y(_01043_),
    .A(_02204_),
    .B(_02205_));
 sg13g2_nor3_1 _16047_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[17] ),
    .B(net4964),
    .C(_02204_),
    .Y(_02206_));
 sg13g2_nand3_1 _16048_ (.B(net4964),
    .C(_02204_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[17] ),
    .Y(_02207_));
 sg13g2_nor2b_1 _16049_ (.A(_02206_),
    .B_N(_02207_),
    .Y(_02208_));
 sg13g2_xnor2_1 _16050_ (.Y(_01044_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[18] ),
    .B(_02208_));
 sg13g2_nor2b_1 _16051_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[1] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][1] ),
    .Y(_02209_));
 sg13g2_xnor2_1 _16052_ (.Y(_02210_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][1] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_xor2_1 _16053_ (.B(_02210_),
    .A(_02506_),
    .X(_01027_));
 sg13g2_a21oi_2 _16054_ (.B1(_02209_),
    .Y(_02211_),
    .A2(_02210_),
    .A1(_02506_));
 sg13g2_xnor2_1 _16055_ (.Y(_02212_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][2] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_nor2b_1 _16056_ (.A(_02211_),
    .B_N(_02212_),
    .Y(_02213_));
 sg13g2_xnor2_1 _16057_ (.Y(_01028_),
    .A(_02211_),
    .B(_02212_));
 sg13g2_a21oi_2 _16058_ (.B1(_02213_),
    .Y(_02214_),
    .A2(_02500_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][2] ));
 sg13g2_xnor2_1 _16059_ (.Y(_02215_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][3] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_nor2b_1 _16060_ (.A(_02214_),
    .B_N(_02215_),
    .Y(_02216_));
 sg13g2_xnor2_1 _16061_ (.Y(_01029_),
    .A(_02214_),
    .B(_02215_));
 sg13g2_a21oi_2 _16062_ (.B1(_02216_),
    .Y(_02217_),
    .A2(_02501_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][3] ));
 sg13g2_xnor2_1 _16063_ (.Y(_02218_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][4] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_nor2b_1 _16064_ (.A(_02217_),
    .B_N(_02218_),
    .Y(_02219_));
 sg13g2_xnor2_1 _16065_ (.Y(_01030_),
    .A(_02217_),
    .B(_02218_));
 sg13g2_a21oi_1 _16066_ (.A1(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][4] ),
    .A2(_02502_),
    .Y(_02220_),
    .B1(_02219_));
 sg13g2_nand2b_1 _16067_ (.Y(_02221_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][5] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_nor2b_1 _16068_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][5] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[5] ),
    .Y(_02222_));
 sg13g2_xnor2_1 _16069_ (.Y(_02223_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][5] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_xnor2_1 _16070_ (.Y(_01031_),
    .A(_02220_),
    .B(_02223_));
 sg13g2_nor2b_1 _16071_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][6] ),
    .Y(_02224_));
 sg13g2_nand2b_1 _16072_ (.Y(_02225_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[6] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][6] ));
 sg13g2_nand2b_1 _16073_ (.Y(_02226_),
    .B(_02225_),
    .A_N(_02224_));
 sg13g2_o21ai_1 _16074_ (.B1(_02221_),
    .Y(_02227_),
    .A1(_02220_),
    .A2(_02222_));
 sg13g2_xnor2_1 _16075_ (.Y(_01032_),
    .A(_02226_),
    .B(_02227_));
 sg13g2_a21oi_2 _16076_ (.B1(_02224_),
    .Y(_02228_),
    .A2(_02227_),
    .A1(_02225_));
 sg13g2_xnor2_1 _16077_ (.Y(_02229_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][7] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nand2b_1 _16078_ (.Y(_02230_),
    .B(_02229_),
    .A_N(_02228_));
 sg13g2_xnor2_1 _16079_ (.Y(_01033_),
    .A(_02228_),
    .B(_02229_));
 sg13g2_o21ai_1 _16080_ (.B1(_02230_),
    .Y(_02231_),
    .A1(_02503_),
    .A2(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_nor2b_1 _16081_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][8] ),
    .Y(_02232_));
 sg13g2_nand2b_1 _16082_ (.Y(_02233_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[8] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][8] ));
 sg13g2_nand2b_1 _16083_ (.Y(_02234_),
    .B(_02233_),
    .A_N(_02232_));
 sg13g2_xnor2_1 _16084_ (.Y(_01034_),
    .A(_02231_),
    .B(_02234_));
 sg13g2_a21oi_2 _16085_ (.B1(_02232_),
    .Y(_02235_),
    .A2(_02233_),
    .A1(_02231_));
 sg13g2_nor2b_1 _16086_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][9] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[9] ),
    .Y(_02236_));
 sg13g2_nand2b_1 _16087_ (.Y(_02237_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][9] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_nor2b_1 _16088_ (.A(_02236_),
    .B_N(_02237_),
    .Y(_02238_));
 sg13g2_xnor2_1 _16089_ (.Y(_01035_),
    .A(_02235_),
    .B(_02238_));
 sg13g2_nor2b_1 _16090_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][10] ),
    .Y(_02239_));
 sg13g2_nand2b_1 _16091_ (.Y(_02240_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[10] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][10] ));
 sg13g2_nand2b_1 _16092_ (.Y(_02241_),
    .B(_02240_),
    .A_N(_02239_));
 sg13g2_a21oi_1 _16093_ (.A1(_02235_),
    .A2(_02237_),
    .Y(_02242_),
    .B1(_02236_));
 sg13g2_xnor2_1 _16094_ (.Y(_01018_),
    .A(_02241_),
    .B(_02242_));
 sg13g2_a21oi_1 _16095_ (.A1(_02240_),
    .A2(_02242_),
    .Y(_02243_),
    .B1(_02239_));
 sg13g2_nor2b_1 _16096_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][11] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[11] ),
    .Y(_02244_));
 sg13g2_nand2b_1 _16097_ (.Y(_02245_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][11] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_nor2b_1 _16098_ (.A(_02244_),
    .B_N(_02245_),
    .Y(_02246_));
 sg13g2_xnor2_1 _16099_ (.Y(_01019_),
    .A(_02243_),
    .B(_02246_));
 sg13g2_nor2b_1 _16100_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][12] ),
    .Y(_02247_));
 sg13g2_nand2b_1 _16101_ (.Y(_02248_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[12] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][12] ));
 sg13g2_nand2b_1 _16102_ (.Y(_02249_),
    .B(_02248_),
    .A_N(_02247_));
 sg13g2_a21oi_1 _16103_ (.A1(_02243_),
    .A2(_02245_),
    .Y(_02250_),
    .B1(_02244_));
 sg13g2_xnor2_1 _16104_ (.Y(_01020_),
    .A(_02249_),
    .B(_02250_));
 sg13g2_a21oi_1 _16105_ (.A1(_02248_),
    .A2(_02250_),
    .Y(_02251_),
    .B1(_02247_));
 sg13g2_nand2b_1 _16106_ (.Y(_02252_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][13] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_nor2b_1 _16107_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][13] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[13] ),
    .Y(_02253_));
 sg13g2_xnor2_1 _16108_ (.Y(_02254_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][13] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_xnor2_1 _16109_ (.Y(_01021_),
    .A(_02251_),
    .B(_02254_));
 sg13g2_nor2b_1 _16110_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][14] ),
    .Y(_02255_));
 sg13g2_nand2b_1 _16111_ (.Y(_02256_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[14] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][14] ));
 sg13g2_nand2b_1 _16112_ (.Y(_02257_),
    .B(_02256_),
    .A_N(_02255_));
 sg13g2_a21oi_1 _16113_ (.A1(_02251_),
    .A2(_02252_),
    .Y(_02258_),
    .B1(_02253_));
 sg13g2_xnor2_1 _16114_ (.Y(_01022_),
    .A(_02257_),
    .B(_02258_));
 sg13g2_a21oi_1 _16115_ (.A1(_02256_),
    .A2(_02258_),
    .Y(_02259_),
    .B1(_02255_));
 sg13g2_nor2b_1 _16116_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][15] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[15] ),
    .Y(_02260_));
 sg13g2_nand2b_1 _16117_ (.Y(_02261_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][15] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_nor2b_1 _16118_ (.A(_02260_),
    .B_N(_02261_),
    .Y(_02262_));
 sg13g2_xnor2_1 _16119_ (.Y(_01023_),
    .A(_02259_),
    .B(_02262_));
 sg13g2_xor2_1 _16120_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[16] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][16] ),
    .X(_02263_));
 sg13g2_a21oi_1 _16121_ (.A1(_02259_),
    .A2(_02261_),
    .Y(_02264_),
    .B1(_02260_));
 sg13g2_nor2b_1 _16122_ (.A(_02263_),
    .B_N(_02264_),
    .Y(_02265_));
 sg13g2_xnor2_1 _16123_ (.Y(_01024_),
    .A(_02263_),
    .B(_02264_));
 sg13g2_a21oi_2 _16124_ (.B1(_02265_),
    .Y(_02266_),
    .A2(_02504_),
    .A1(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][16] ));
 sg13g2_nand2b_1 _16125_ (.Y(_02267_),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][17] ),
    .A_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_nor2b_1 _16126_ (.A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][17] ),
    .B_N(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[17] ),
    .Y(_02268_));
 sg13g2_xnor2_1 _16127_ (.Y(_02269_),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][17] ),
    .B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_xnor2_1 _16128_ (.Y(_01025_),
    .A(_02266_),
    .B(_02269_));
 sg13g2_o21ai_1 _16129_ (.B1(_02267_),
    .Y(_02270_),
    .A1(_02266_),
    .A2(_02268_));
 sg13g2_xor2_1 _16130_ (.B(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[18] ),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][18] ),
    .X(_02271_));
 sg13g2_xnor2_1 _16131_ (.Y(_01026_),
    .A(_02270_),
    .B(_02271_));
 sg13g2_nand2_1 _16132_ (.Y(_02272_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[0] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_nand2_1 _16133_ (.Y(_02273_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_nor2_1 _16134_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[1] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[1] ),
    .Y(_02274_));
 sg13g2_xor2_1 _16135_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[1] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[1] ),
    .X(_02275_));
 sg13g2_xnor2_1 _16136_ (.Y(_01177_),
    .A(_02272_),
    .B(_02275_));
 sg13g2_o21ai_1 _16137_ (.B1(_02273_),
    .Y(_02276_),
    .A1(_02272_),
    .A2(_02274_));
 sg13g2_xnor2_1 _16138_ (.Y(_02277_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[2] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_nor2b_1 _16139_ (.A(_02277_),
    .B_N(_02276_),
    .Y(_02278_));
 sg13g2_xnor2_1 _16140_ (.Y(_01178_),
    .A(_02276_),
    .B(_02277_));
 sg13g2_a21o_1 _16141_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[2] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[2] ),
    .B1(_02278_),
    .X(_02279_));
 sg13g2_xnor2_1 _16142_ (.Y(_02280_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[3] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_nor2b_1 _16143_ (.A(_02280_),
    .B_N(_02279_),
    .Y(_02281_));
 sg13g2_xnor2_1 _16144_ (.Y(_01179_),
    .A(_02279_),
    .B(_02280_));
 sg13g2_a21o_1 _16145_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[3] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[3] ),
    .B1(_02281_),
    .X(_02282_));
 sg13g2_xnor2_1 _16146_ (.Y(_02283_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[4] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_nor2b_1 _16147_ (.A(_02283_),
    .B_N(_02282_),
    .Y(_02284_));
 sg13g2_xnor2_1 _16148_ (.Y(_01180_),
    .A(_02282_),
    .B(_02283_));
 sg13g2_a21o_1 _16149_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[4] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[4] ),
    .B1(_02284_),
    .X(_02285_));
 sg13g2_nand2_1 _16150_ (.Y(_02286_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[5] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_xnor2_1 _16151_ (.Y(_02287_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[5] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_xnor2_1 _16152_ (.Y(_01181_),
    .A(_02285_),
    .B(_02287_));
 sg13g2_xnor2_1 _16153_ (.Y(_02288_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[6] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_o21ai_1 _16154_ (.B1(_02285_),
    .Y(_02289_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[5] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_a21oi_1 _16155_ (.A1(_02286_),
    .A2(_02289_),
    .Y(_02290_),
    .B1(_02288_));
 sg13g2_nand3_1 _16156_ (.B(_02288_),
    .C(_02289_),
    .A(_02286_),
    .Y(_02291_));
 sg13g2_nor2b_1 _16157_ (.A(_02290_),
    .B_N(_02291_),
    .Y(_01182_));
 sg13g2_a21oi_1 _16158_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[6] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[6] ),
    .Y(_02292_),
    .B1(_02290_));
 sg13g2_nand2_1 _16159_ (.Y(_02293_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[7] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_nor2_1 _16160_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[7] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[7] ),
    .Y(_02294_));
 sg13g2_xor2_1 _16161_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[7] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[7] ),
    .X(_02295_));
 sg13g2_xnor2_1 _16162_ (.Y(_01183_),
    .A(_02292_),
    .B(_02295_));
 sg13g2_o21ai_1 _16163_ (.B1(_02293_),
    .Y(_02296_),
    .A1(_02292_),
    .A2(_02294_));
 sg13g2_xnor2_1 _16164_ (.Y(_02297_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[8] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_nor2b_1 _16165_ (.A(_02297_),
    .B_N(_02296_),
    .Y(_02298_));
 sg13g2_xnor2_1 _16166_ (.Y(_01184_),
    .A(_02296_),
    .B(_02297_));
 sg13g2_xnor2_1 _16167_ (.Y(_02299_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[9] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_a21o_1 _16168_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[8] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[8] ),
    .B1(_02298_),
    .X(_02300_));
 sg13g2_xnor2_1 _16169_ (.Y(_01185_),
    .A(_02299_),
    .B(_02300_));
 sg13g2_nand2_1 _16170_ (.Y(_02301_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[10] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_nor2_1 _16171_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[10] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[10] ),
    .Y(_02302_));
 sg13g2_xor2_1 _16172_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[10] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[10] ),
    .X(_02303_));
 sg13g2_a21o_1 _16173_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[9] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[9] ),
    .B1(_02300_),
    .X(_02304_));
 sg13g2_o21ai_1 _16174_ (.B1(_02304_),
    .Y(_02305_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[9] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_xnor2_1 _16175_ (.Y(_01168_),
    .A(_02303_),
    .B(_02305_));
 sg13g2_xnor2_1 _16176_ (.Y(_02306_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[11] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_o21ai_1 _16177_ (.B1(_02301_),
    .Y(_02307_),
    .A1(_02302_),
    .A2(_02305_));
 sg13g2_xnor2_1 _16178_ (.Y(_01169_),
    .A(_02306_),
    .B(_02307_));
 sg13g2_nand2_1 _16179_ (.Y(_02308_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[12] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_nor2_1 _16180_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[12] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[12] ),
    .Y(_02309_));
 sg13g2_xor2_1 _16181_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[12] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[12] ),
    .X(_02310_));
 sg13g2_a21o_1 _16182_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[11] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[11] ),
    .B1(_02307_),
    .X(_02311_));
 sg13g2_o21ai_1 _16183_ (.B1(_02311_),
    .Y(_02312_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[11] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_xnor2_1 _16184_ (.Y(_01170_),
    .A(_02310_),
    .B(_02312_));
 sg13g2_o21ai_1 _16185_ (.B1(_02308_),
    .Y(_02313_),
    .A1(_02309_),
    .A2(_02312_));
 sg13g2_xnor2_1 _16186_ (.Y(_02314_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[13] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_xnor2_1 _16187_ (.Y(_01171_),
    .A(_02313_),
    .B(_02314_));
 sg13g2_xnor2_1 _16188_ (.Y(_02315_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[14] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_a21o_1 _16189_ (.A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[13] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[13] ),
    .B1(_02313_),
    .X(_02316_));
 sg13g2_o21ai_1 _16190_ (.B1(_02316_),
    .Y(_02317_),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[13] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_nor2_1 _16191_ (.A(_02315_),
    .B(_02317_),
    .Y(_02318_));
 sg13g2_xor2_1 _16192_ (.B(_02317_),
    .A(_02315_),
    .X(_01172_));
 sg13g2_a21oi_2 _16193_ (.B1(_02318_),
    .Y(_02319_),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[14] ),
    .A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_nand2_1 _16194_ (.Y(_02320_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_nor2_1 _16195_ (.A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[15] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[15] ),
    .Y(_02321_));
 sg13g2_xor2_1 _16196_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[15] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[15] ),
    .X(_02322_));
 sg13g2_xnor2_1 _16197_ (.Y(_01173_),
    .A(_02319_),
    .B(_02322_));
 sg13g2_nand2_1 _16198_ (.Y(_02323_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[16] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_xor2_1 _16199_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[16] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[16] ),
    .X(_02324_));
 sg13g2_o21ai_1 _16200_ (.B1(_02320_),
    .Y(_02325_),
    .A1(_02319_),
    .A2(_02321_));
 sg13g2_nand2_1 _16201_ (.Y(_02326_),
    .A(_02324_),
    .B(_02325_));
 sg13g2_xor2_1 _16202_ (.B(_02325_),
    .A(_02324_),
    .X(_01174_));
 sg13g2_xnor2_1 _16203_ (.Y(_02327_),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[17] ),
    .B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_a21oi_1 _16204_ (.A1(_02323_),
    .A2(_02326_),
    .Y(_02328_),
    .B1(_02327_));
 sg13g2_nand3_1 _16205_ (.B(_02326_),
    .C(_02327_),
    .A(_02323_),
    .Y(_02329_));
 sg13g2_nor2b_1 _16206_ (.A(_02328_),
    .B_N(_02329_),
    .Y(_01175_));
 sg13g2_a21oi_1 _16207_ (.A1(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[17] ),
    .A2(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[17] ),
    .Y(_02330_),
    .B1(_02328_));
 sg13g2_xor2_1 _16208_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[18] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[18] ),
    .X(_02331_));
 sg13g2_xnor2_1 _16209_ (.Y(_01176_),
    .A(_02330_),
    .B(_02331_));
 sg13g2_xor2_1 _16210_ (.B(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[0] ),
    .A(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[0] ),
    .X(_01167_));
 sg13g2_inv_1 _16211_ (.Y(_01195_),
    .A(net5214));
 sg13g2_inv_1 _16212_ (.Y(_01196_),
    .A(net5593));
 sg13g2_inv_1 _16213_ (.Y(_01197_),
    .A(net5593));
 sg13g2_inv_1 _16214_ (.Y(_01198_),
    .A(net5631));
 sg13g2_inv_1 _16215_ (.Y(_01199_),
    .A(net5633));
 sg13g2_inv_1 _16216_ (.Y(_01200_),
    .A(net5643));
 sg13g2_inv_1 _16217_ (.Y(_01201_),
    .A(net5648));
 sg13g2_inv_1 _16218_ (.Y(_01202_),
    .A(net5644));
 sg13g2_inv_1 _16219_ (.Y(_01203_),
    .A(net5644));
 sg13g2_inv_1 _16220_ (.Y(_01204_),
    .A(net5663));
 sg13g2_inv_1 _16221_ (.Y(_01205_),
    .A(net5663));
 sg13g2_inv_1 _16222_ (.Y(_01206_),
    .A(net5663));
 sg13g2_inv_1 _16223_ (.Y(_01207_),
    .A(net5666));
 sg13g2_inv_1 _16224_ (.Y(_01208_),
    .A(net5661));
 sg13g2_inv_1 _16225_ (.Y(_01209_),
    .A(net5661));
 sg13g2_inv_1 _16226_ (.Y(_01210_),
    .A(net5651));
 sg13g2_inv_1 _16227_ (.Y(_01211_),
    .A(net5651));
 sg13g2_inv_1 _16228_ (.Y(_01212_),
    .A(net5618));
 sg13g2_inv_1 _16229_ (.Y(_01213_),
    .A(net5589));
 sg13g2_inv_1 _16230_ (.Y(_01214_),
    .A(net5592));
 sg13g2_inv_1 _16231_ (.Y(_01215_),
    .A(net5491));
 sg13g2_inv_1 _16232_ (.Y(_01216_),
    .A(net5488));
 sg13g2_inv_1 _16233_ (.Y(_01217_),
    .A(net5428));
 sg13g2_inv_1 _16234_ (.Y(_01218_),
    .A(net5351));
 sg13g2_inv_1 _16235_ (.Y(_01219_),
    .A(net5351));
 sg13g2_inv_1 _16236_ (.Y(_01220_),
    .A(net5369));
 sg13g2_inv_1 _16237_ (.Y(_01221_),
    .A(net5369));
 sg13g2_inv_1 _16238_ (.Y(_01222_),
    .A(net5352));
 sg13g2_inv_1 _16239_ (.Y(_01223_),
    .A(net5351));
 sg13g2_inv_1 _16240_ (.Y(_01224_),
    .A(net5351));
 sg13g2_inv_1 _16241_ (.Y(_01225_),
    .A(net5356));
 sg13g2_inv_1 _16242_ (.Y(_01226_),
    .A(net5365));
 sg13g2_inv_1 _16243_ (.Y(_01227_),
    .A(net5205));
 sg13g2_inv_1 _16244_ (.Y(_01228_),
    .A(net5209));
 sg13g2_inv_1 _16245_ (.Y(_01229_),
    .A(net5440));
 sg13g2_inv_1 _16246_ (.Y(_01230_),
    .A(net5456));
 sg13g2_inv_1 _16247_ (.Y(_01231_),
    .A(net5461));
 sg13g2_inv_1 _16248_ (.Y(_01232_),
    .A(net5502));
 sg13g2_inv_1 _16249_ (.Y(_01233_),
    .A(net5502));
 sg13g2_inv_1 _16250_ (.Y(_01234_),
    .A(net5480));
 sg13g2_inv_1 _16251_ (.Y(_01235_),
    .A(net5479));
 sg13g2_inv_1 _16252_ (.Y(_01236_),
    .A(net5456));
 sg13g2_inv_1 _16253_ (.Y(_01237_),
    .A(net5439));
 sg13g2_inv_1 _16254_ (.Y(_01238_),
    .A(net5440));
 sg13g2_inv_1 _16255_ (.Y(_01239_),
    .A(net5443));
 sg13g2_inv_1 _16256_ (.Y(_01240_),
    .A(net5443));
 sg13g2_inv_1 _16257_ (.Y(_01241_),
    .A(net5406));
 sg13g2_inv_1 _16258_ (.Y(_01242_),
    .A(net5406));
 sg13g2_inv_1 _16259_ (.Y(_01243_),
    .A(net5407));
 sg13g2_inv_1 _16260_ (.Y(_01244_),
    .A(net5379));
 sg13g2_inv_1 _16261_ (.Y(_01245_),
    .A(net5379));
 sg13g2_inv_1 _16262_ (.Y(_01246_),
    .A(net5379));
 sg13g2_inv_1 _16263_ (.Y(_01247_),
    .A(net5355));
 sg13g2_inv_1 _16264_ (.Y(_01248_),
    .A(net5350));
 sg13g2_inv_1 _16265_ (.Y(_01249_),
    .A(net5345));
 sg13g2_inv_1 _16266_ (.Y(_01250_),
    .A(net5343));
 sg13g2_inv_1 _16267_ (.Y(_01251_),
    .A(net5342));
 sg13g2_inv_1 _16268_ (.Y(_01252_),
    .A(net5300));
 sg13g2_inv_1 _16269_ (.Y(_01253_),
    .A(net5342));
 sg13g2_inv_1 _16270_ (.Y(_01254_),
    .A(net5343));
 sg13g2_inv_1 _16271_ (.Y(_01255_),
    .A(net5349));
 sg13g2_inv_1 _16272_ (.Y(_01256_),
    .A(net5354));
 sg13g2_inv_1 _16273_ (.Y(_01257_),
    .A(net5354));
 sg13g2_inv_1 _16274_ (.Y(_01258_),
    .A(net5355));
 sg13g2_inv_1 _16275_ (.Y(_01259_),
    .A(net5348));
 sg13g2_inv_1 _16276_ (.Y(_01260_),
    .A(net5218));
 sg13g2_inv_1 _16277_ (.Y(_01261_),
    .A(net5210));
 sg13g2_inv_1 _16278_ (.Y(_01262_),
    .A(net5408));
 sg13g2_inv_1 _16279_ (.Y(_01263_),
    .A(net5411));
 sg13g2_inv_1 _16280_ (.Y(_01264_),
    .A(net5411));
 sg13g2_inv_1 _16281_ (.Y(_01265_),
    .A(net5412));
 sg13g2_inv_1 _16282_ (.Y(_01266_),
    .A(net5412));
 sg13g2_inv_1 _16283_ (.Y(_01267_),
    .A(net5409));
 sg13g2_inv_1 _16284_ (.Y(_01268_),
    .A(net5398));
 sg13g2_inv_1 _16285_ (.Y(_01269_),
    .A(net5398));
 sg13g2_inv_1 _16286_ (.Y(_01270_),
    .A(net5397));
 sg13g2_inv_1 _16287_ (.Y(_01271_),
    .A(net5337));
 sg13g2_inv_1 _16288_ (.Y(_01272_),
    .A(net5332));
 sg13g2_inv_1 _16289_ (.Y(_01273_),
    .A(net5332));
 sg13g2_inv_1 _16290_ (.Y(_01274_),
    .A(net5326));
 sg13g2_inv_1 _16291_ (.Y(_01275_),
    .A(net5326));
 sg13g2_inv_1 _16292_ (.Y(_01276_),
    .A(net5326));
 sg13g2_inv_1 _16293_ (.Y(_01277_),
    .A(net5326));
 sg13g2_inv_1 _16294_ (.Y(_01278_),
    .A(net5327));
 sg13g2_inv_1 _16295_ (.Y(_01279_),
    .A(net5322));
 sg13g2_inv_1 _16296_ (.Y(_01280_),
    .A(net5275));
 sg13g2_inv_1 _16297_ (.Y(_01281_),
    .A(net5273));
 sg13g2_inv_1 _16298_ (.Y(_01282_),
    .A(net5262));
 sg13g2_inv_1 _16299_ (.Y(_01283_),
    .A(net5219));
 sg13g2_inv_1 _16300_ (.Y(_01284_),
    .A(net5213));
 sg13g2_inv_1 _16301_ (.Y(_01285_),
    .A(net5213));
 sg13g2_inv_1 _16302_ (.Y(_01286_),
    .A(net5209));
 sg13g2_inv_1 _16303_ (.Y(_01287_),
    .A(net5211));
 sg13g2_inv_1 _16304_ (.Y(_01288_),
    .A(net5211));
 sg13g2_inv_1 _16305_ (.Y(_01289_),
    .A(net5212));
 sg13g2_inv_1 _16306_ (.Y(_01290_),
    .A(net5212));
 sg13g2_inv_1 _16307_ (.Y(_01291_),
    .A(net5210));
 sg13g2_inv_1 _16308_ (.Y(_01292_),
    .A(net5210));
 sg13g2_inv_1 _16309_ (.Y(_01293_),
    .A(net5209));
 sg13g2_inv_1 _16310_ (.Y(_01294_),
    .A(net5218));
 sg13g2_inv_1 _16311_ (.Y(_01295_),
    .A(net5258));
 sg13g2_inv_1 _16312_ (.Y(_01296_),
    .A(net5260));
 sg13g2_inv_1 _16313_ (.Y(_01297_),
    .A(net5260));
 sg13g2_inv_1 _16314_ (.Y(_01298_),
    .A(net5233));
 sg13g2_inv_1 _16315_ (.Y(_01299_),
    .A(net5233));
 sg13g2_inv_1 _16316_ (.Y(_01300_),
    .A(net5232));
 sg13g2_inv_1 _16317_ (.Y(_01301_),
    .A(net5232));
 sg13g2_inv_1 _16318_ (.Y(_01302_),
    .A(net5232));
 sg13g2_inv_1 _16319_ (.Y(_01303_),
    .A(net5230));
 sg13g2_inv_1 _16320_ (.Y(_01304_),
    .A(net5230));
 sg13g2_inv_1 _16321_ (.Y(_01305_),
    .A(net5230));
 sg13g2_inv_1 _16322_ (.Y(_01306_),
    .A(net5234));
 sg13g2_inv_1 _16323_ (.Y(_01307_),
    .A(net5234));
 sg13g2_inv_1 _16324_ (.Y(_01308_),
    .A(net5234));
 sg13g2_inv_1 _16325_ (.Y(_01309_),
    .A(net5234));
 sg13g2_inv_1 _16326_ (.Y(_01310_),
    .A(net5231));
 sg13g2_inv_1 _16327_ (.Y(_01311_),
    .A(net5236));
 sg13g2_inv_1 _16328_ (.Y(_01312_),
    .A(net5233));
 sg13g2_inv_1 _16329_ (.Y(_01313_),
    .A(net5198));
 sg13g2_inv_1 _16330_ (.Y(_01314_),
    .A(net5198));
 sg13g2_inv_1 _16331_ (.Y(_01315_),
    .A(net5215));
 sg13g2_inv_1 _16332_ (.Y(_01316_),
    .A(net5215));
 sg13g2_inv_1 _16333_ (.Y(_01317_),
    .A(net5204));
 sg13g2_inv_1 _16334_ (.Y(_01318_),
    .A(net5205));
 sg13g2_inv_1 _16335_ (.Y(_01319_),
    .A(net5205));
 sg13g2_inv_1 _16336_ (.Y(_01320_),
    .A(net5206));
 sg13g2_inv_1 _16337_ (.Y(_01321_),
    .A(net5206));
 sg13g2_inv_1 _16338_ (.Y(_01322_),
    .A(net5213));
 sg13g2_inv_1 _16339_ (.Y(_01323_),
    .A(net5212));
 sg13g2_inv_1 _16340_ (.Y(_01324_),
    .A(net5213));
 sg13g2_inv_1 _16341_ (.Y(_01325_),
    .A(net5212));
 sg13g2_inv_1 _16342_ (.Y(_01326_),
    .A(net5214));
 sg13g2_inv_1 _16343_ (.Y(_01327_),
    .A(net5219));
 sg13g2_inv_1 _16344_ (.Y(_01328_),
    .A(net5566));
 sg13g2_inv_1 _16345_ (.Y(_01329_),
    .A(net5566));
 sg13g2_inv_1 _16346_ (.Y(_01330_),
    .A(net5571));
 sg13g2_inv_1 _16347_ (.Y(_01331_),
    .A(net5580));
 sg13g2_inv_1 _16348_ (.Y(_01332_),
    .A(net5580));
 sg13g2_inv_1 _16349_ (.Y(_01333_),
    .A(net5581));
 sg13g2_inv_1 _16350_ (.Y(_01334_),
    .A(net5581));
 sg13g2_inv_1 _16351_ (.Y(_01335_),
    .A(net5624));
 sg13g2_inv_1 _16352_ (.Y(_01336_),
    .A(net5624));
 sg13g2_inv_1 _16353_ (.Y(_01337_),
    .A(net5592));
 sg13g2_inv_1 _16354_ (.Y(_01338_),
    .A(net5592));
 sg13g2_inv_1 _16355_ (.Y(_01339_),
    .A(net5593));
 sg13g2_inv_1 _16356_ (.Y(_01340_),
    .A(net5591));
 sg13g2_inv_1 _16357_ (.Y(_01341_),
    .A(net5603));
 sg13g2_inv_1 _16358_ (.Y(_01342_),
    .A(net5569));
 sg13g2_inv_1 _16359_ (.Y(_01343_),
    .A(net5495));
 sg13g2_inv_1 _16360_ (.Y(_01344_),
    .A(net5483));
 sg13g2_inv_1 _16361_ (.Y(_01345_),
    .A(net5476));
 sg13g2_inv_1 _16362_ (.Y(_01346_),
    .A(net5429));
 sg13g2_inv_1 _16363_ (.Y(_01347_),
    .A(net5431));
 sg13g2_inv_1 _16364_ (.Y(_01348_),
    .A(net5417));
 sg13g2_inv_1 _16365_ (.Y(_01349_),
    .A(net5353));
 sg13g2_inv_1 _16366_ (.Y(_01350_),
    .A(net5350));
 sg13g2_inv_1 _16367_ (.Y(_01351_),
    .A(net5350));
 sg13g2_inv_1 _16368_ (.Y(_01352_),
    .A(net5345));
 sg13g2_inv_1 _16369_ (.Y(_01353_),
    .A(net5344));
 sg13g2_inv_1 _16370_ (.Y(_01354_),
    .A(net5344));
 sg13g2_inv_1 _16371_ (.Y(_01355_),
    .A(net5344));
 sg13g2_inv_1 _16372_ (.Y(_01356_),
    .A(net5300));
 sg13g2_inv_1 _16373_ (.Y(_01357_),
    .A(net5300));
 sg13g2_inv_1 _16374_ (.Y(_01358_),
    .A(net5303));
 sg13g2_inv_1 _16375_ (.Y(_01359_),
    .A(net5215));
 sg13g2_inv_1 _16376_ (.Y(_01360_),
    .A(net5214));
 sg13g2_inv_1 _16377_ (.Y(_01361_),
    .A(net5471));
 sg13g2_inv_1 _16378_ (.Y(_01362_),
    .A(net5466));
 sg13g2_inv_1 _16379_ (.Y(_01363_),
    .A(net5515));
 sg13g2_inv_1 _16380_ (.Y(_01364_),
    .A(net5515));
 sg13g2_inv_1 _16381_ (.Y(_01365_),
    .A(net5517));
 sg13g2_inv_1 _16382_ (.Y(_01366_),
    .A(net5519));
 sg13g2_inv_1 _16383_ (.Y(_01367_),
    .A(net5511));
 sg13g2_inv_1 _16384_ (.Y(_01368_),
    .A(net5505));
 sg13g2_inv_1 _16385_ (.Y(_01369_),
    .A(net5471));
 sg13g2_inv_1 _16386_ (.Y(_01370_),
    .A(net5471));
 sg13g2_inv_1 _16387_ (.Y(_01371_),
    .A(net5471));
 sg13g2_inv_1 _16388_ (.Y(_01372_),
    .A(net5451));
 sg13g2_inv_1 _16389_ (.Y(_01373_),
    .A(net5450));
 sg13g2_inv_1 _16390_ (.Y(_01374_),
    .A(net5452));
 sg13g2_inv_1 _16391_ (.Y(_01375_),
    .A(net5452));
 sg13g2_inv_1 _16392_ (.Y(_01376_),
    .A(net5452));
 sg13g2_inv_1 _16393_ (.Y(_01377_),
    .A(net5453));
 sg13g2_inv_1 _16394_ (.Y(_01378_),
    .A(net5443));
 sg13g2_inv_1 _16395_ (.Y(_01379_),
    .A(net5407));
 sg13g2_inv_1 _16396_ (.Y(_01380_),
    .A(net5379));
 sg13g2_inv_1 _16397_ (.Y(_01381_),
    .A(net5373));
 sg13g2_inv_1 _16398_ (.Y(_01382_),
    .A(net5356));
 sg13g2_inv_1 _16399_ (.Y(_01383_),
    .A(net5350));
 sg13g2_inv_1 _16400_ (.Y(_01384_),
    .A(net5345));
 sg13g2_inv_1 _16401_ (.Y(_01385_),
    .A(net5300));
 sg13g2_inv_1 _16402_ (.Y(_01386_),
    .A(net5299));
 sg13g2_inv_1 _16403_ (.Y(_01387_),
    .A(net5299));
 sg13g2_inv_1 _16404_ (.Y(_01388_),
    .A(net5284));
 sg13g2_inv_1 _16405_ (.Y(_01389_),
    .A(net5284));
 sg13g2_inv_1 _16406_ (.Y(_01390_),
    .A(net5283));
 sg13g2_inv_1 _16407_ (.Y(_01391_),
    .A(net5340));
 sg13g2_inv_1 _16408_ (.Y(_01392_),
    .A(net5220));
 sg13g2_inv_1 _16409_ (.Y(_01393_),
    .A(net5209));
 sg13g2_inv_1 _16410_ (.Y(_01394_),
    .A(net5325));
 sg13g2_inv_1 _16411_ (.Y(_01395_),
    .A(net5325));
 sg13g2_inv_1 _16412_ (.Y(_01396_),
    .A(net5325));
 sg13g2_inv_1 _16413_ (.Y(_01397_),
    .A(net5324));
 sg13g2_inv_1 _16414_ (.Y(_01398_),
    .A(net5324));
 sg13g2_inv_1 _16415_ (.Y(_01399_),
    .A(net5324));
 sg13g2_inv_1 _16416_ (.Y(_01400_),
    .A(net5293));
 sg13g2_inv_1 _16417_ (.Y(_01401_),
    .A(net5293));
 sg13g2_inv_1 _16418_ (.Y(_01402_),
    .A(net5293));
 sg13g2_inv_1 _16419_ (.Y(_01403_),
    .A(net5292));
 sg13g2_inv_1 _16420_ (.Y(_01404_),
    .A(net5292));
 sg13g2_inv_1 _16421_ (.Y(_01405_),
    .A(net5289));
 sg13g2_inv_1 _16422_ (.Y(_01406_),
    .A(net5289));
 sg13g2_inv_1 _16423_ (.Y(_01407_),
    .A(net5289));
 sg13g2_inv_1 _16424_ (.Y(_01408_),
    .A(net5289));
 sg13g2_inv_1 _16425_ (.Y(_01409_),
    .A(net5294));
 sg13g2_inv_1 _16426_ (.Y(_01410_),
    .A(net5295));
 sg13g2_inv_1 _16427_ (.Y(_01411_),
    .A(net5269));
 sg13g2_inv_1 _16428_ (.Y(_01412_),
    .A(net5260));
 sg13g2_inv_1 _16429_ (.Y(_01413_),
    .A(net5258));
 sg13g2_inv_1 _16430_ (.Y(_01414_),
    .A(net5255));
 sg13g2_inv_1 _16431_ (.Y(_01415_),
    .A(net5255));
 sg13g2_inv_1 _16432_ (.Y(_01416_),
    .A(net5216));
 sg13g2_inv_1 _16433_ (.Y(_01417_),
    .A(net5216));
 sg13g2_inv_1 _16434_ (.Y(_01418_),
    .A(net5216));
 sg13g2_inv_1 _16435_ (.Y(_01419_),
    .A(net5216));
 sg13g2_inv_1 _16436_ (.Y(_01420_),
    .A(net5215));
 sg13g2_inv_1 _16437_ (.Y(_01421_),
    .A(net5218));
 sg13g2_inv_1 _16438_ (.Y(_01422_),
    .A(net5218));
 sg13g2_inv_1 _16439_ (.Y(_01423_),
    .A(net5218));
 sg13g2_inv_1 _16440_ (.Y(_01424_),
    .A(net5219));
 sg13g2_inv_1 _16441_ (.Y(_01425_),
    .A(net5219));
 sg13g2_inv_1 _16442_ (.Y(_01426_),
    .A(net5283));
 sg13g2_inv_1 _16443_ (.Y(_01427_),
    .A(net5282));
 sg13g2_inv_1 _16444_ (.Y(_01428_),
    .A(net5281));
 sg13g2_inv_1 _16445_ (.Y(_01429_),
    .A(net5281));
 sg13g2_inv_1 _16446_ (.Y(_01430_),
    .A(net5281));
 sg13g2_inv_1 _16447_ (.Y(_01431_),
    .A(net5282));
 sg13g2_inv_1 _16448_ (.Y(_01432_),
    .A(net5282));
 sg13g2_inv_1 _16449_ (.Y(_01433_),
    .A(net5283));
 sg13g2_inv_1 _16450_ (.Y(_01434_),
    .A(net5284));
 sg13g2_inv_1 _16451_ (.Y(_01435_),
    .A(net5298));
 sg13g2_inv_1 _16452_ (.Y(_01436_),
    .A(net5297));
 sg13g2_inv_1 _16453_ (.Y(_01437_),
    .A(net5301));
 sg13g2_inv_1 _16454_ (.Y(_01438_),
    .A(net5342));
 sg13g2_inv_1 _16455_ (.Y(_01439_),
    .A(net5343));
 sg13g2_inv_1 _16456_ (.Y(_01440_),
    .A(net5343));
 sg13g2_inv_1 _16457_ (.Y(_01441_),
    .A(net5303));
 sg13g2_inv_1 _16458_ (.Y(_01442_),
    .A(net5297));
 sg13g2_inv_1 _16459_ (.Y(_01443_),
    .A(net5297));
 sg13g2_inv_1 _16460_ (.Y(_01444_),
    .A(net5238));
 sg13g2_inv_1 _16461_ (.Y(_01445_),
    .A(net5237));
 sg13g2_inv_1 _16462_ (.Y(_01446_),
    .A(net5229));
 sg13g2_inv_1 _16463_ (.Y(_01447_),
    .A(net5225));
 sg13g2_inv_1 _16464_ (.Y(_01448_),
    .A(net5196));
 sg13g2_inv_1 _16465_ (.Y(_01449_),
    .A(net5191));
 sg13g2_inv_1 _16466_ (.Y(_01450_),
    .A(net5177));
 sg13g2_inv_1 _16467_ (.Y(_01451_),
    .A(net5188));
 sg13g2_inv_1 _16468_ (.Y(_01452_),
    .A(net5177));
 sg13g2_inv_1 _16469_ (.Y(_01453_),
    .A(net5177));
 sg13g2_inv_1 _16470_ (.Y(_01454_),
    .A(net5177));
 sg13g2_inv_1 _16471_ (.Y(_01455_),
    .A(net5180));
 sg13g2_inv_1 _16472_ (.Y(_01456_),
    .A(net5180));
 sg13g2_inv_1 _16473_ (.Y(_01457_),
    .A(net5201));
 sg13g2_inv_1 _16474_ (.Y(_01459_),
    .A(net5161));
 sg13g2_inv_1 _16475_ (.Y(_01460_),
    .A(net5165));
 sg13g2_inv_1 _16476_ (.Y(_01461_),
    .A(net5166));
 sg13g2_inv_1 _16477_ (.Y(_01462_),
    .A(net5171));
 sg13g2_inv_1 _16478_ (.Y(_01463_),
    .A(net5168));
 sg13g2_inv_1 _16479_ (.Y(_01464_),
    .A(net5168));
 sg13g2_inv_1 _16480_ (.Y(_01465_),
    .A(net5168));
 sg13g2_inv_1 _16481_ (.Y(_01466_),
    .A(net5168));
 sg13g2_inv_1 _16482_ (.Y(_01467_),
    .A(net5168));
 sg13g2_inv_1 _16483_ (.Y(_01468_),
    .A(net5171));
 sg13g2_inv_1 _16484_ (.Y(_01469_),
    .A(net5166));
 sg13g2_inv_1 _16485_ (.Y(_01470_),
    .A(net5165));
 sg13g2_inv_1 _16486_ (.Y(_01471_),
    .A(net5161));
 sg13g2_inv_1 _16487_ (.Y(_01472_),
    .A(net5160));
 sg13g2_inv_1 _16488_ (.Y(_01473_),
    .A(net5157));
 sg13g2_inv_1 _16489_ (.Y(_01474_),
    .A(net5157));
 sg13g2_inv_1 _16490_ (.Y(_01475_),
    .A(net5157));
 sg13g2_inv_1 _16491_ (.Y(_01476_),
    .A(net5164));
 sg13g2_inv_1 _16492_ (.Y(_01477_),
    .A(net5151));
 sg13g2_inv_1 _16493_ (.Y(_01478_),
    .A(net5157));
 sg13g2_inv_1 _16494_ (.Y(_01479_),
    .A(net5160));
 sg13g2_inv_1 _16495_ (.Y(_01480_),
    .A(net5160));
 sg13g2_inv_1 _16496_ (.Y(_01481_),
    .A(net5165));
 sg13g2_inv_1 _16497_ (.Y(_01482_),
    .A(net5171));
 sg13g2_inv_1 _16498_ (.Y(_01483_),
    .A(net5169));
 sg13g2_inv_1 _16499_ (.Y(_01484_),
    .A(net5169));
 sg13g2_inv_1 _16500_ (.Y(_01485_),
    .A(net5169));
 sg13g2_inv_1 _16501_ (.Y(_01486_),
    .A(net5172));
 sg13g2_inv_1 _16502_ (.Y(_01487_),
    .A(net5173));
 sg13g2_inv_1 _16503_ (.Y(_01488_),
    .A(net5166));
 sg13g2_inv_1 _16504_ (.Y(_01489_),
    .A(net5167));
 sg13g2_inv_1 _16505_ (.Y(_01490_),
    .A(net5162));
 sg13g2_inv_1 _16506_ (.Y(_01491_),
    .A(net5162));
 sg13g2_inv_1 _16507_ (.Y(_01492_),
    .A(net5159));
 sg13g2_inv_1 _16508_ (.Y(_01493_),
    .A(net5159));
 sg13g2_inv_1 _16509_ (.Y(_01494_),
    .A(net5151));
 sg13g2_inv_1 _16510_ (.Y(_01495_),
    .A(net5152));
 sg13g2_inv_1 _16511_ (.Y(_01496_),
    .A(net5106));
 sg13g2_inv_1 _16512_ (.Y(_01497_),
    .A(net5106));
 sg13g2_inv_1 _16513_ (.Y(_01498_),
    .A(net5105));
 sg13g2_inv_1 _16514_ (.Y(_01499_),
    .A(net5117));
 sg13g2_inv_1 _16515_ (.Y(_01500_),
    .A(net5117));
 sg13g2_inv_1 _16516_ (.Y(_01501_),
    .A(net5117));
 sg13g2_inv_1 _16517_ (.Y(_01502_),
    .A(net5111));
 sg13g2_inv_1 _16518_ (.Y(_01503_),
    .A(net5105));
 sg13g2_inv_1 _16519_ (.Y(_01504_),
    .A(net5105));
 sg13g2_inv_1 _16520_ (.Y(_01505_),
    .A(net5086));
 sg13g2_inv_1 _16521_ (.Y(_01506_),
    .A(net5091));
 sg13g2_inv_1 _16522_ (.Y(_01507_),
    .A(net5089));
 sg13g2_inv_1 _16523_ (.Y(_01508_),
    .A(net5086));
 sg13g2_inv_1 _16524_ (.Y(_01509_),
    .A(net5086));
 sg13g2_inv_1 _16525_ (.Y(_01510_),
    .A(net5086));
 sg13g2_inv_1 _16526_ (.Y(_01511_),
    .A(net5085));
 sg13g2_inv_1 _16527_ (.Y(_01512_),
    .A(net5085));
 sg13g2_inv_1 _16528_ (.Y(_01513_),
    .A(net5084));
 sg13g2_inv_1 _16529_ (.Y(_01514_),
    .A(net5084));
 sg13g2_inv_1 _16530_ (.Y(_01515_),
    .A(net5109));
 sg13g2_inv_1 _16531_ (.Y(_01516_),
    .A(net5109));
 sg13g2_inv_1 _16532_ (.Y(_01517_),
    .A(net5114));
 sg13g2_inv_1 _16533_ (.Y(_01518_),
    .A(net5113));
 sg13g2_inv_1 _16534_ (.Y(_01519_),
    .A(net5115));
 sg13g2_inv_1 _16535_ (.Y(_01520_),
    .A(net5115));
 sg13g2_inv_1 _16536_ (.Y(_01521_),
    .A(net5115));
 sg13g2_inv_1 _16537_ (.Y(_01522_),
    .A(net5112));
 sg13g2_inv_1 _16538_ (.Y(_01523_),
    .A(net5107));
 sg13g2_inv_1 _16539_ (.Y(_01524_),
    .A(net5106));
 sg13g2_inv_1 _16540_ (.Y(_01525_),
    .A(net5090));
 sg13g2_inv_1 _16541_ (.Y(_01526_),
    .A(net5090));
 sg13g2_inv_1 _16542_ (.Y(_01527_),
    .A(net5091));
 sg13g2_inv_1 _16543_ (.Y(_01528_),
    .A(net5090));
 sg13g2_inv_1 _16544_ (.Y(_01529_),
    .A(net5088));
 sg13g2_inv_1 _16545_ (.Y(_01530_),
    .A(net5088));
 sg13g2_inv_1 _16546_ (.Y(_01531_),
    .A(net5088));
 sg13g2_inv_1 _16547_ (.Y(_01532_),
    .A(net5092));
 sg13g2_inv_1 _16548_ (.Y(_01533_),
    .A(net5085));
 sg13g2_inv_1 _16549_ (.Y(_01534_),
    .A(net5096));
 sg13g2_inv_1 _16550_ (.Y(_01535_),
    .A(net5094));
 sg13g2_inv_1 _16551_ (.Y(_01536_),
    .A(net5094));
 sg13g2_inv_1 _16552_ (.Y(_01537_),
    .A(net5095));
 sg13g2_inv_1 _16553_ (.Y(_01538_),
    .A(net5095));
 sg13g2_inv_1 _16554_ (.Y(_01539_),
    .A(net5094));
 sg13g2_inv_1 _16555_ (.Y(_01540_),
    .A(net5093));
 sg13g2_inv_1 _16556_ (.Y(_01541_),
    .A(net5103));
 sg13g2_inv_1 _16557_ (.Y(_01542_),
    .A(net5082));
 sg13g2_inv_1 _16558_ (.Y(_01543_),
    .A(net5081));
 sg13g2_inv_1 _16559_ (.Y(_01544_),
    .A(net5082));
 sg13g2_inv_1 _16560_ (.Y(_01545_),
    .A(net5080));
 sg13g2_inv_1 _16561_ (.Y(_01546_),
    .A(net5077));
 sg13g2_inv_1 _16562_ (.Y(_01547_),
    .A(net5077));
 sg13g2_inv_1 _16563_ (.Y(_01548_),
    .A(net5077));
 sg13g2_inv_1 _16564_ (.Y(_01549_),
    .A(net5076));
 sg13g2_inv_1 _16565_ (.Y(_01550_),
    .A(net5070));
 sg13g2_inv_1 _16566_ (.Y(_01551_),
    .A(net5076));
 sg13g2_inv_1 _16567_ (.Y(_01552_),
    .A(net5054));
 sg13g2_inv_1 _16568_ (.Y(_01553_),
    .A(net5097));
 sg13g2_inv_1 _16569_ (.Y(_01554_),
    .A(net5100));
 sg13g2_inv_1 _16570_ (.Y(_01555_),
    .A(net5101));
 sg13g2_inv_1 _16571_ (.Y(_01556_),
    .A(net5101));
 sg13g2_inv_1 _16572_ (.Y(_01557_),
    .A(net5101));
 sg13g2_inv_1 _16573_ (.Y(_01558_),
    .A(net5099));
 sg13g2_inv_1 _16574_ (.Y(_01559_),
    .A(net5098));
 sg13g2_inv_1 _16575_ (.Y(_01560_),
    .A(net5094));
 sg13g2_inv_1 _16576_ (.Y(_01561_),
    .A(net5093));
 sg13g2_inv_1 _16577_ (.Y(_01562_),
    .A(net5081));
 sg13g2_inv_1 _16578_ (.Y(_01563_),
    .A(net5081));
 sg13g2_inv_1 _16579_ (.Y(_01564_),
    .A(net5080));
 sg13g2_inv_1 _16580_ (.Y(_01565_),
    .A(net5079));
 sg13g2_inv_1 _16581_ (.Y(_01566_),
    .A(net5078));
 sg13g2_inv_1 _16582_ (.Y(_01567_),
    .A(net5078));
 sg13g2_inv_1 _16583_ (.Y(_01568_),
    .A(net5073));
 sg13g2_inv_1 _16584_ (.Y(_01569_),
    .A(net5073));
 sg13g2_inv_1 _16585_ (.Y(_01570_),
    .A(net5072));
 sg13g2_inv_1 _16586_ (.Y(_01571_),
    .A(net5076));
 sg13g2_inv_1 _16587_ (.Y(_01572_),
    .A(net5027));
 sg13g2_inv_1 _16588_ (.Y(_01573_),
    .A(net5027));
 sg13g2_inv_1 _16589_ (.Y(_01574_),
    .A(net5029));
 sg13g2_inv_1 _16590_ (.Y(_01575_),
    .A(net5025));
 sg13g2_inv_1 _16591_ (.Y(_01576_),
    .A(net5025));
 sg13g2_inv_1 _16592_ (.Y(_01577_),
    .A(net5025));
 sg13g2_inv_1 _16593_ (.Y(_01578_),
    .A(net5013));
 sg13g2_inv_1 _16594_ (.Y(_01579_),
    .A(net5012));
 sg13g2_inv_1 _16595_ (.Y(_01580_),
    .A(net5012));
 sg13g2_inv_1 _16596_ (.Y(_01581_),
    .A(net5012));
 sg13g2_inv_1 _16597_ (.Y(_01582_),
    .A(net5012));
 sg13g2_inv_1 _16598_ (.Y(_01583_),
    .A(net5011));
 sg13g2_inv_1 _16599_ (.Y(_01584_),
    .A(net5011));
 sg13g2_inv_1 _16600_ (.Y(_01585_),
    .A(net5011));
 sg13g2_inv_1 _16601_ (.Y(_01586_),
    .A(net5014));
 sg13g2_inv_1 _16602_ (.Y(_01587_),
    .A(net5014));
 sg13g2_inv_1 _16603_ (.Y(_01588_),
    .A(net5014));
 sg13g2_inv_1 _16604_ (.Y(_01589_),
    .A(net5015));
 sg13g2_inv_1 _16605_ (.Y(_01590_),
    .A(net5014));
 sg13g2_inv_1 _16606_ (.Y(_01591_),
    .A(net5028));
 sg13g2_inv_1 _16607_ (.Y(_01592_),
    .A(net5028));
 sg13g2_inv_1 _16608_ (.Y(_01593_),
    .A(net5026));
 sg13g2_inv_1 _16609_ (.Y(_01594_),
    .A(net5026));
 sg13g2_inv_1 _16610_ (.Y(_01595_),
    .A(net5026));
 sg13g2_inv_1 _16611_ (.Y(_01596_),
    .A(net5023));
 sg13g2_inv_1 _16612_ (.Y(_01597_),
    .A(net5023));
 sg13g2_inv_1 _16613_ (.Y(_01598_),
    .A(net5023));
 sg13g2_inv_1 _16614_ (.Y(_01599_),
    .A(net5023));
 sg13g2_inv_1 _16615_ (.Y(_01600_),
    .A(net5020));
 sg13g2_inv_1 _16616_ (.Y(_01601_),
    .A(net5017));
 sg13g2_inv_1 _16617_ (.Y(_01602_),
    .A(net5017));
 sg13g2_inv_1 _16618_ (.Y(_01603_),
    .A(net5016));
 sg13g2_inv_1 _16619_ (.Y(_01604_),
    .A(net5022));
 sg13g2_inv_1 _16620_ (.Y(_01605_),
    .A(net5016));
 sg13g2_inv_1 _16621_ (.Y(_01606_),
    .A(net5024));
 sg13g2_inv_1 _16622_ (.Y(_01607_),
    .A(net5016));
 sg13g2_inv_1 _16623_ (.Y(_01608_),
    .A(net5016));
 sg13g2_inv_1 _16624_ (.Y(_01609_),
    .A(net5018));
 sg13g2_inv_1 _16625_ (.Y(_01610_),
    .A(net5143));
 sg13g2_inv_1 _16626_ (.Y(_01611_),
    .A(net5143));
 sg13g2_inv_1 _16627_ (.Y(_01612_),
    .A(net5146));
 sg13g2_inv_1 _16628_ (.Y(_01613_),
    .A(net5146));
 sg13g2_inv_1 _16629_ (.Y(_01614_),
    .A(net5149));
 sg13g2_inv_1 _16630_ (.Y(_01615_),
    .A(net5149));
 sg13g2_inv_1 _16631_ (.Y(_01616_),
    .A(net5154));
 sg13g2_inv_1 _16632_ (.Y(_01617_),
    .A(net5154));
 sg13g2_inv_1 _16633_ (.Y(_01618_),
    .A(net5148));
 sg13g2_inv_1 _16634_ (.Y(_01619_),
    .A(net5148));
 sg13g2_inv_1 _16635_ (.Y(_01620_),
    .A(net5146));
 sg13g2_inv_1 _16636_ (.Y(_01621_),
    .A(net5141));
 sg13g2_inv_1 _16637_ (.Y(_01622_),
    .A(net5135));
 sg13g2_inv_1 _16638_ (.Y(_01623_),
    .A(net5135));
 sg13g2_inv_1 _16639_ (.Y(_01624_),
    .A(net5134));
 sg13g2_inv_1 _16640_ (.Y(_01625_),
    .A(net5134));
 sg13g2_inv_1 _16641_ (.Y(_01626_),
    .A(net5134));
 sg13g2_inv_1 _16642_ (.Y(_01627_),
    .A(net5134));
 sg13g2_inv_1 _16643_ (.Y(_01628_),
    .A(net5134));
 sg13g2_inv_1 _16644_ (.Y(_01629_),
    .A(net5142));
 sg13g2_inv_1 _16645_ (.Y(_01630_),
    .A(net5142));
 sg13g2_inv_1 _16646_ (.Y(_01631_),
    .A(net5144));
 sg13g2_inv_1 _16647_ (.Y(_01632_),
    .A(net5146));
 sg13g2_inv_1 _16648_ (.Y(_01633_),
    .A(net5148));
 sg13g2_inv_1 _16649_ (.Y(_01634_),
    .A(net5154));
 sg13g2_inv_1 _16650_ (.Y(_01635_),
    .A(net5155));
 sg13g2_inv_1 _16651_ (.Y(_01636_),
    .A(net5155));
 sg13g2_inv_1 _16652_ (.Y(_01637_),
    .A(net5155));
 sg13g2_inv_1 _16653_ (.Y(_01638_),
    .A(net5150));
 sg13g2_inv_1 _16654_ (.Y(_01639_),
    .A(net5150));
 sg13g2_inv_1 _16655_ (.Y(_01640_),
    .A(net5147));
 sg13g2_inv_1 _16656_ (.Y(_01641_),
    .A(net5142));
 sg13g2_inv_1 _16657_ (.Y(_01642_),
    .A(net5145));
 sg13g2_inv_1 _16658_ (.Y(_01643_),
    .A(net5136));
 sg13g2_inv_1 _16659_ (.Y(_01644_),
    .A(net5136));
 sg13g2_inv_1 _16660_ (.Y(_01645_),
    .A(net5136));
 sg13g2_inv_1 _16661_ (.Y(_01646_),
    .A(net5133));
 sg13g2_inv_1 _16662_ (.Y(_01647_),
    .A(net5130));
 sg13g2_inv_1 _16663_ (.Y(_01648_),
    .A(net5113));
 sg13g2_inv_1 _16664_ (.Y(_01649_),
    .A(net5115));
 sg13g2_inv_1 _16665_ (.Y(_01650_),
    .A(net5115));
 sg13g2_inv_1 _16666_ (.Y(_01651_),
    .A(net5131));
 sg13g2_inv_1 _16667_ (.Y(_01652_),
    .A(net5130));
 sg13g2_inv_1 _16668_ (.Y(_01653_),
    .A(net5130));
 sg13g2_inv_1 _16669_ (.Y(_01654_),
    .A(net5131));
 sg13g2_inv_1 _16670_ (.Y(_01655_),
    .A(net5116));
 sg13g2_inv_1 _16671_ (.Y(_01656_),
    .A(net5113));
 sg13g2_inv_1 _16672_ (.Y(_01657_),
    .A(net5112));
 sg13g2_inv_1 _16673_ (.Y(_01658_),
    .A(net5112));
 sg13g2_inv_1 _16674_ (.Y(_01659_),
    .A(net5108));
 sg13g2_inv_1 _16675_ (.Y(_01660_),
    .A(net5108));
 sg13g2_inv_1 _16676_ (.Y(_01661_),
    .A(net5109));
 sg13g2_inv_1 _16677_ (.Y(_01662_),
    .A(net5107));
 sg13g2_inv_1 _16678_ (.Y(_01663_),
    .A(net5106));
 sg13g2_inv_1 _16679_ (.Y(_01664_),
    .A(net5107));
 sg13g2_inv_1 _16680_ (.Y(_01665_),
    .A(net5107));
 sg13g2_inv_1 _16681_ (.Y(_01666_),
    .A(net5112));
 sg13g2_inv_1 _16682_ (.Y(_01667_),
    .A(net5125));
 sg13g2_inv_1 _16683_ (.Y(_01668_),
    .A(net5125));
 sg13g2_inv_1 _16684_ (.Y(_01669_),
    .A(net5125));
 sg13g2_inv_1 _16685_ (.Y(_01670_),
    .A(net5127));
 sg13g2_inv_1 _16686_ (.Y(_01671_),
    .A(net5139));
 sg13g2_inv_1 _16687_ (.Y(_01672_),
    .A(net5139));
 sg13g2_inv_1 _16688_ (.Y(_01673_),
    .A(net5139));
 sg13g2_inv_1 _16689_ (.Y(_01674_),
    .A(net5127));
 sg13g2_inv_1 _16690_ (.Y(_01675_),
    .A(net5126));
 sg13g2_inv_1 _16691_ (.Y(_01676_),
    .A(net5120));
 sg13g2_inv_1 _16692_ (.Y(_01677_),
    .A(net5124));
 sg13g2_inv_1 _16693_ (.Y(_01678_),
    .A(net5122));
 sg13g2_inv_1 _16694_ (.Y(_01679_),
    .A(net5122));
 sg13g2_inv_1 _16695_ (.Y(_01680_),
    .A(net5123));
 sg13g2_inv_1 _16696_ (.Y(_01681_),
    .A(net5122));
 sg13g2_inv_1 _16697_ (.Y(_01682_),
    .A(net5122));
 sg13g2_inv_1 _16698_ (.Y(_01683_),
    .A(net5121));
 sg13g2_inv_1 _16699_ (.Y(_01684_),
    .A(net5120));
 sg13g2_inv_1 _16700_ (.Y(_01685_),
    .A(net5120));
 sg13g2_inv_1 _16701_ (.Y(_01686_),
    .A(net5075));
 sg13g2_inv_1 _16702_ (.Y(_01687_),
    .A(net5052));
 sg13g2_inv_1 _16703_ (.Y(_01688_),
    .A(net5075));
 sg13g2_inv_1 _16704_ (.Y(_01689_),
    .A(net5052));
 sg13g2_inv_1 _16705_ (.Y(_01690_),
    .A(net5052));
 sg13g2_inv_1 _16706_ (.Y(_01691_),
    .A(net5051));
 sg13g2_inv_1 _16707_ (.Y(_01692_),
    .A(net5050));
 sg13g2_inv_1 _16708_ (.Y(_01693_),
    .A(net5050));
 sg13g2_inv_1 _16709_ (.Y(_01694_),
    .A(net5053));
 sg13g2_inv_1 _16710_ (.Y(_01695_),
    .A(net5049));
 sg13g2_inv_1 _16711_ (.Y(_01696_),
    .A(net5048));
 sg13g2_inv_1 _16712_ (.Y(_01697_),
    .A(net5049));
 sg13g2_inv_1 _16713_ (.Y(_01698_),
    .A(net5049));
 sg13g2_inv_1 _16714_ (.Y(_01699_),
    .A(net5046));
 sg13g2_inv_1 _16715_ (.Y(_01700_),
    .A(net5045));
 sg13g2_inv_1 _16716_ (.Y(_01701_),
    .A(net5045));
 sg13g2_inv_1 _16717_ (.Y(_01702_),
    .A(net5045));
 sg13g2_inv_1 _16718_ (.Y(_01703_),
    .A(net5047));
 sg13g2_inv_1 _16719_ (.Y(_01704_),
    .A(net5047));
 sg13g2_inv_1 _16720_ (.Y(_01705_),
    .A(net5074));
 sg13g2_inv_1 _16721_ (.Y(_01706_),
    .A(net5074));
 sg13g2_inv_1 _16722_ (.Y(_01707_),
    .A(net5071));
 sg13g2_inv_1 _16723_ (.Y(_01708_),
    .A(net5071));
 sg13g2_inv_1 _16724_ (.Y(_01709_),
    .A(net5071));
 sg13g2_inv_1 _16725_ (.Y(_01710_),
    .A(net5069));
 sg13g2_inv_1 _16726_ (.Y(_01711_),
    .A(net5069));
 sg13g2_inv_1 _16727_ (.Y(_01712_),
    .A(net5069));
 sg13g2_inv_1 _16728_ (.Y(_01713_),
    .A(net5068));
 sg13g2_inv_1 _16729_ (.Y(_01714_),
    .A(net5068));
 sg13g2_inv_1 _16730_ (.Y(_01715_),
    .A(net5068));
 sg13g2_inv_1 _16731_ (.Y(_01716_),
    .A(net5061));
 sg13g2_inv_1 _16732_ (.Y(_01717_),
    .A(net5061));
 sg13g2_inv_1 _16733_ (.Y(_01718_),
    .A(net5042));
 sg13g2_inv_1 _16734_ (.Y(_01719_),
    .A(net5042));
 sg13g2_inv_1 _16735_ (.Y(_01720_),
    .A(net5042));
 sg13g2_inv_1 _16736_ (.Y(_01721_),
    .A(net5050));
 sg13g2_inv_1 _16737_ (.Y(_01722_),
    .A(net5049));
 sg13g2_inv_1 _16738_ (.Y(_01723_),
    .A(net5046));
 sg13g2_inv_1 _16739_ (.Y(_01724_),
    .A(net5033));
 sg13g2_inv_1 _16740_ (.Y(_01725_),
    .A(net5031));
 sg13g2_inv_1 _16741_ (.Y(_01726_),
    .A(net5031));
 sg13g2_inv_1 _16742_ (.Y(_01727_),
    .A(net5030));
 sg13g2_inv_1 _16743_ (.Y(_01728_),
    .A(net5030));
 sg13g2_inv_1 _16744_ (.Y(_01729_),
    .A(net5030));
 sg13g2_inv_1 _16745_ (.Y(_01730_),
    .A(net5032));
 sg13g2_inv_1 _16746_ (.Y(_01731_),
    .A(net5032));
 sg13g2_inv_1 _16747_ (.Y(_01732_),
    .A(net5035));
 sg13g2_inv_1 _16748_ (.Y(_01733_),
    .A(net5035));
 sg13g2_inv_1 _16749_ (.Y(_01734_),
    .A(net5035));
 sg13g2_inv_1 _16750_ (.Y(_01735_),
    .A(net5039));
 sg13g2_inv_1 _16751_ (.Y(_01736_),
    .A(net5038));
 sg13g2_inv_1 _16752_ (.Y(_01737_),
    .A(net5057));
 sg13g2_inv_1 _16753_ (.Y(_01738_),
    .A(net5057));
 sg13g2_inv_1 _16754_ (.Y(_01739_),
    .A(net5057));
 sg13g2_inv_1 _16755_ (.Y(_01740_),
    .A(net5038));
 sg13g2_inv_1 _16756_ (.Y(_01741_),
    .A(net5039));
 sg13g2_inv_1 _16757_ (.Y(_01742_),
    .A(net5037));
 sg13g2_inv_1 _16758_ (.Y(_01743_),
    .A(net5040));
 sg13g2_inv_1 _16759_ (.Y(_01744_),
    .A(net5040));
 sg13g2_inv_1 _16760_ (.Y(_01745_),
    .A(net5037));
 sg13g2_inv_1 _16761_ (.Y(_01746_),
    .A(net5036));
 sg13g2_inv_1 _16762_ (.Y(_01747_),
    .A(net5036));
 sg13g2_inv_1 _16763_ (.Y(_01748_),
    .A(net5040));
 sg13g2_inv_1 _16764_ (.Y(_01749_),
    .A(net5040));
 sg13g2_inv_1 _16765_ (.Y(_01750_),
    .A(net5038));
 sg13g2_inv_1 _16766_ (.Y(_01751_),
    .A(net5057));
 sg13g2_inv_1 _16767_ (.Y(_01752_),
    .A(net5058));
 sg13g2_inv_1 _16768_ (.Y(_01753_),
    .A(net5059));
 sg13g2_inv_1 _16769_ (.Y(_01754_),
    .A(net5064));
 sg13g2_inv_1 _16770_ (.Y(_01755_),
    .A(net5065));
 sg13g2_inv_1 _16771_ (.Y(_01756_),
    .A(net5065));
 sg13g2_inv_1 _16772_ (.Y(_01757_),
    .A(net5067));
 sg13g2_inv_1 _16773_ (.Y(_01758_),
    .A(net5064));
 sg13g2_inv_1 _16774_ (.Y(_01759_),
    .A(net5059));
 sg13g2_inv_1 _16775_ (.Y(_01760_),
    .A(net5059));
 sg13g2_inv_1 _16776_ (.Y(_01761_),
    .A(net5058));
 sg13g2_inv_1 _16777_ (.Y(_01762_),
    .A(net5211));
 sg13g2_inv_1 _16778_ (.Y(_01763_),
    .A(net5461));
 sg13g2_inv_1 _16779_ (.Y(_01764_),
    .A(net5502));
 sg13g2_inv_1 _16780_ (.Y(_01765_),
    .A(net5506));
 sg13g2_inv_1 _16781_ (.Y(_01766_),
    .A(net5506));
 sg13g2_inv_1 _16782_ (.Y(_01767_),
    .A(net5508));
 sg13g2_inv_1 _16783_ (.Y(_01768_),
    .A(net5508));
 sg13g2_inv_1 _16784_ (.Y(_01769_),
    .A(net5528));
 sg13g2_inv_1 _16785_ (.Y(_01770_),
    .A(net5507));
 sg13g2_inv_1 _16786_ (.Y(_01771_),
    .A(net5479));
 sg13g2_inv_1 _16787_ (.Y(_01772_),
    .A(net5435));
 sg13g2_inv_1 _16788_ (.Y(_01773_),
    .A(net5439));
 sg13g2_inv_1 _16789_ (.Y(_01774_),
    .A(net5443));
 sg13g2_inv_1 _16790_ (.Y(_01775_),
    .A(net5443));
 sg13g2_inv_1 _16791_ (.Y(_01776_),
    .A(net5407));
 sg13g2_inv_1 _16792_ (.Y(_01777_),
    .A(net5401));
 sg13g2_inv_1 _16793_ (.Y(_01778_),
    .A(net5401));
 sg13g2_inv_1 _16794_ (.Y(_01779_),
    .A(net5400));
 sg13g2_inv_1 _16795_ (.Y(_01780_),
    .A(net5400));
 sg13g2_inv_1 _16796_ (.Y(_01781_),
    .A(net5366));
 sg13g2_inv_1 _16797_ (.Y(_01782_),
    .A(net5366));
 sg13g2_inv_1 _16798_ (.Y(_01783_),
    .A(net5364));
 sg13g2_inv_1 _16799_ (.Y(_01784_),
    .A(net5346));
 sg13g2_inv_1 _16800_ (.Y(_01785_),
    .A(net5346));
 sg13g2_inv_1 _16801_ (.Y(_01786_),
    .A(net5355));
 sg13g2_inv_1 _16802_ (.Y(_01787_),
    .A(net5355));
 sg13g2_inv_1 _16803_ (.Y(_01788_),
    .A(net5346));
 sg13g2_inv_1 _16804_ (.Y(_01789_),
    .A(net5302));
 sg13g2_inv_1 _16805_ (.Y(_01790_),
    .A(net5302));
 sg13g2_inv_1 _16806_ (.Y(_01791_),
    .A(net5297));
 sg13g2_inv_1 _16807_ (.Y(_01792_),
    .A(net5298));
 sg13g2_inv_1 _16808_ (.Y(_01793_),
    .A(net5307));
 sg13g2_inv_1 _16809_ (.Y(_01794_),
    .A(net5220));
 sg13g2_inv_1 _16810_ (.Y(_01795_),
    .A(net5267));
 sg13g2_inv_1 _16811_ (.Y(_01796_),
    .A(net5376));
 sg13g2_inv_1 _16812_ (.Y(_01797_),
    .A(net5624));
 sg13g2_inv_1 _16813_ (.Y(_01798_),
    .A(net5185));
 sg13g2_dfrbp_1 _16814_ (.CLK(_01194_),
    .RESET_B(net19),
    .D(_01799_),
    .Q_N(_06855_),
    .Q(\u_supermic_top_module.i2s_out ));
 sg13g2_dfrbp_1 _16815_ (.CLK(_01195_),
    .RESET_B(net20),
    .D(_01800_),
    .Q_N(_06856_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.out ));
 sg13g2_dfrbp_1 _16816_ (.CLK(net5591),
    .RESET_B(net6100),
    .D(_00255_),
    .Q_N(_06854_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _16817_ (.CLK(_01196_),
    .RESET_B(net6102),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.u_mux_shift.data ),
    .Q_N(_06857_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _16818_ (.CLK(net5593),
    .RESET_B(net6102),
    .D(_00234_),
    .Q_N(_06853_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16819_ (.CLK(_01197_),
    .RESET_B(net6102),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_06858_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16820_ (.CLK(net5630),
    .RESET_B(net6139),
    .D(_00245_),
    .Q_N(_06852_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16821_ (.CLK(_01198_),
    .RESET_B(net6139),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_06859_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16822_ (.CLK(net5630),
    .RESET_B(net6140),
    .D(_00248_),
    .Q_N(_06851_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16823_ (.CLK(_01199_),
    .RESET_B(net6142),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_06860_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16824_ (.CLK(net5632),
    .RESET_B(net6141),
    .D(_00249_),
    .Q_N(_06850_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16825_ (.CLK(_01200_),
    .RESET_B(net6152),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_06861_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16826_ (.CLK(net5643),
    .RESET_B(net6152),
    .D(_00250_),
    .Q_N(_06849_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16827_ (.CLK(_01201_),
    .RESET_B(net6157),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_06862_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16828_ (.CLK(net5644),
    .RESET_B(net6153),
    .D(_00251_),
    .Q_N(_06848_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16829_ (.CLK(_01202_),
    .RESET_B(net6153),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_06863_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16830_ (.CLK(net5645),
    .RESET_B(net6154),
    .D(_00252_),
    .Q_N(_06847_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16831_ (.CLK(_01203_),
    .RESET_B(net6153),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_06864_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16832_ (.CLK(net5663),
    .RESET_B(net6173),
    .D(_00253_),
    .Q_N(_06846_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16833_ (.CLK(_01204_),
    .RESET_B(net6173),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_06865_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16834_ (.CLK(net5683),
    .RESET_B(net6193),
    .D(_00254_),
    .Q_N(_06845_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16835_ (.CLK(_01205_),
    .RESET_B(net6173),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_06866_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _16836_ (.CLK(net5663),
    .RESET_B(net6173),
    .D(_00224_),
    .Q_N(_06844_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16837_ (.CLK(_01206_),
    .RESET_B(net6173),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_06867_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16838_ (.CLK(net5666),
    .RESET_B(net6176),
    .D(_00225_),
    .Q_N(_06843_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16839_ (.CLK(_01207_),
    .RESET_B(net6176),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_06868_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16840_ (.CLK(net5662),
    .RESET_B(net6172),
    .D(_00226_),
    .Q_N(_06842_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16841_ (.CLK(_01208_),
    .RESET_B(net6171),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_06869_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16842_ (.CLK(net5661),
    .RESET_B(net6171),
    .D(_00227_),
    .Q_N(_06841_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16843_ (.CLK(_01209_),
    .RESET_B(net6171),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_06870_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16844_ (.CLK(net5657),
    .RESET_B(net6161),
    .D(_00228_),
    .Q_N(_06840_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16845_ (.CLK(_01210_),
    .RESET_B(net6161),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_06871_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16846_ (.CLK(net5651),
    .RESET_B(net6160),
    .D(_00229_),
    .Q_N(_06839_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16847_ (.CLK(_01211_),
    .RESET_B(net6160),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_06872_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16848_ (.CLK(net5618),
    .RESET_B(net6127),
    .D(_00230_),
    .Q_N(_06838_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16849_ (.CLK(_01212_),
    .RESET_B(net6127),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_06873_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16850_ (.CLK(net5591),
    .RESET_B(net6100),
    .D(_00231_),
    .Q_N(_06837_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16851_ (.CLK(_01213_),
    .RESET_B(net6100),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_06874_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16852_ (.CLK(net5592),
    .RESET_B(net6101),
    .D(_00232_),
    .Q_N(_06836_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16853_ (.CLK(_01214_),
    .RESET_B(net6101),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_06875_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16854_ (.CLK(net5500),
    .RESET_B(net6009),
    .D(_00233_),
    .Q_N(_06835_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16855_ (.CLK(_01215_),
    .RESET_B(net6000),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_06876_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16856_ (.CLK(net5488),
    .RESET_B(net5997),
    .D(_00235_),
    .Q_N(_06834_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16857_ (.CLK(_01216_),
    .RESET_B(net5997),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_06877_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16858_ (.CLK(net5431),
    .RESET_B(net5940),
    .D(_00236_),
    .Q_N(_06833_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16859_ (.CLK(_01217_),
    .RESET_B(net5937),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_06878_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16860_ (.CLK(net5353),
    .RESET_B(net5861),
    .D(_00237_),
    .Q_N(_06832_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16861_ (.CLK(_01218_),
    .RESET_B(net5861),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_06879_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16862_ (.CLK(net5351),
    .RESET_B(net5859),
    .D(_00238_),
    .Q_N(_06831_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16863_ (.CLK(_01219_),
    .RESET_B(net5859),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_06880_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16864_ (.CLK(net5351),
    .RESET_B(net5859),
    .D(_00239_),
    .Q_N(_06830_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16865_ (.CLK(_01220_),
    .RESET_B(net5878),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_06881_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16866_ (.CLK(net5352),
    .RESET_B(net5859),
    .D(_00240_),
    .Q_N(_06829_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16867_ (.CLK(_01221_),
    .RESET_B(net5878),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_06882_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16868_ (.CLK(net5352),
    .RESET_B(net5860),
    .D(_00241_),
    .Q_N(_06828_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16869_ (.CLK(_01222_),
    .RESET_B(net5860),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_06883_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16870_ (.CLK(net5351),
    .RESET_B(net5859),
    .D(_00242_),
    .Q_N(_06827_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16871_ (.CLK(_01223_),
    .RESET_B(net5859),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_06884_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16872_ (.CLK(net5351),
    .RESET_B(net5859),
    .D(_00243_),
    .Q_N(_06826_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16873_ (.CLK(_01224_),
    .RESET_B(net5859),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_06885_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16874_ (.CLK(net5353),
    .RESET_B(net5861),
    .D(_00244_),
    .Q_N(_06825_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16875_ (.CLK(_01225_),
    .RESET_B(net5864),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_06886_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16876_ (.CLK(net5356),
    .RESET_B(net5864),
    .D(_00246_),
    .Q_N(_06824_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16877_ (.CLK(_01226_),
    .RESET_B(net5874),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_06887_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16878_ (.CLK(net5186),
    .RESET_B(net5696),
    .D(_00247_),
    .Q_N(_06823_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16879_ (.CLK(_01227_),
    .RESET_B(net5715),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_06822_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16880_ (.CLK(_01228_),
    .RESET_B(net21),
    .D(_01801_),
    .Q_N(_06888_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.out ));
 sg13g2_dfrbp_1 _16881_ (.CLK(net5440),
    .RESET_B(net5949),
    .D(_00223_),
    .Q_N(_06821_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _16882_ (.CLK(_01229_),
    .RESET_B(net5965),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.u_mux_shift.data ),
    .Q_N(_06889_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _16883_ (.CLK(net5456),
    .RESET_B(net5965),
    .D(_00202_),
    .Q_N(_06820_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16884_ (.CLK(_01230_),
    .RESET_B(net5965),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_06890_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16885_ (.CLK(net5461),
    .RESET_B(net5969),
    .D(_00213_),
    .Q_N(_06819_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16886_ (.CLK(_01231_),
    .RESET_B(net5969),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_06891_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16887_ (.CLK(net5502),
    .RESET_B(net6011),
    .D(_00216_),
    .Q_N(_06818_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16888_ (.CLK(_01232_),
    .RESET_B(net6011),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_06892_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16889_ (.CLK(net5502),
    .RESET_B(net6011),
    .D(_00217_),
    .Q_N(_06817_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16890_ (.CLK(_01233_),
    .RESET_B(net6011),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_06893_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16891_ (.CLK(net5480),
    .RESET_B(net5989),
    .D(_00218_),
    .Q_N(_06816_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16892_ (.CLK(_01234_),
    .RESET_B(net5989),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_06894_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16893_ (.CLK(net5479),
    .RESET_B(net5988),
    .D(_00219_),
    .Q_N(_06815_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16894_ (.CLK(_01235_),
    .RESET_B(net5988),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_06895_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16895_ (.CLK(net5437),
    .RESET_B(net5946),
    .D(_00220_),
    .Q_N(_06814_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16896_ (.CLK(_01236_),
    .RESET_B(net5965),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_06896_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16897_ (.CLK(net5439),
    .RESET_B(net5948),
    .D(_00221_),
    .Q_N(_06813_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16898_ (.CLK(_01237_),
    .RESET_B(net5948),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_06897_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16899_ (.CLK(net5440),
    .RESET_B(net5949),
    .D(_00222_),
    .Q_N(_06812_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16900_ (.CLK(_01238_),
    .RESET_B(net5949),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_06898_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _16901_ (.CLK(net5443),
    .RESET_B(net5952),
    .D(_00192_),
    .Q_N(_06811_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16902_ (.CLK(_01239_),
    .RESET_B(net5952),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_06899_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16903_ (.CLK(net5443),
    .RESET_B(net5952),
    .D(_00193_),
    .Q_N(_06810_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16904_ (.CLK(_01240_),
    .RESET_B(net5952),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_06900_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16905_ (.CLK(net5406),
    .RESET_B(net5915),
    .D(_00194_),
    .Q_N(_06809_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16906_ (.CLK(_01241_),
    .RESET_B(net5915),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_06901_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16907_ (.CLK(net5406),
    .RESET_B(net5915),
    .D(_00195_),
    .Q_N(_06808_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16908_ (.CLK(_01242_),
    .RESET_B(net5915),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_06902_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16909_ (.CLK(net5406),
    .RESET_B(net5915),
    .D(_00196_),
    .Q_N(_06807_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16910_ (.CLK(_01243_),
    .RESET_B(net5916),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_06903_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16911_ (.CLK(net5407),
    .RESET_B(net5916),
    .D(_00197_),
    .Q_N(_06806_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16912_ (.CLK(_01244_),
    .RESET_B(net5888),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_06904_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16913_ (.CLK(net5379),
    .RESET_B(net5888),
    .D(_00198_),
    .Q_N(_06805_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16914_ (.CLK(_01245_),
    .RESET_B(net5888),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_06905_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16915_ (.CLK(net5379),
    .RESET_B(net5888),
    .D(_00199_),
    .Q_N(_06804_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16916_ (.CLK(_01246_),
    .RESET_B(net5888),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_06906_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16917_ (.CLK(net5355),
    .RESET_B(net5863),
    .D(_00200_),
    .Q_N(_06803_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16918_ (.CLK(_01247_),
    .RESET_B(net5863),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_06907_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16919_ (.CLK(net5347),
    .RESET_B(net5855),
    .D(_00201_),
    .Q_N(_06802_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16920_ (.CLK(_01248_),
    .RESET_B(net5858),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_06908_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16921_ (.CLK(net5345),
    .RESET_B(net5854),
    .D(_00203_),
    .Q_N(_06801_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16922_ (.CLK(_01249_),
    .RESET_B(net5854),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_06909_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16923_ (.CLK(net5342),
    .RESET_B(net5852),
    .D(_00204_),
    .Q_N(_06800_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16924_ (.CLK(_01250_),
    .RESET_B(net5852),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_06910_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16925_ (.CLK(net5342),
    .RESET_B(net5851),
    .D(_00205_),
    .Q_N(_06799_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16926_ (.CLK(_01251_),
    .RESET_B(net5851),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_06911_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16927_ (.CLK(net5300),
    .RESET_B(net5810),
    .D(_00206_),
    .Q_N(_06798_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16928_ (.CLK(_01252_),
    .RESET_B(net5851),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_06912_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16929_ (.CLK(net5301),
    .RESET_B(net5810),
    .D(_00207_),
    .Q_N(_06797_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16930_ (.CLK(_01253_),
    .RESET_B(net5851),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_06913_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16931_ (.CLK(net5342),
    .RESET_B(net5851),
    .D(_00208_),
    .Q_N(_06796_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16932_ (.CLK(_01254_),
    .RESET_B(net5852),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_06914_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16933_ (.CLK(net5345),
    .RESET_B(net5854),
    .D(_00209_),
    .Q_N(_06795_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16934_ (.CLK(_01255_),
    .RESET_B(net5857),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_06915_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16935_ (.CLK(net5345),
    .RESET_B(net5854),
    .D(_00210_),
    .Q_N(_06794_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16936_ (.CLK(_01256_),
    .RESET_B(net5862),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_06916_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16937_ (.CLK(net5350),
    .RESET_B(net5862),
    .D(_00211_),
    .Q_N(_06793_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16938_ (.CLK(_01257_),
    .RESET_B(net5858),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_06917_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16939_ (.CLK(net5354),
    .RESET_B(net5862),
    .D(_00212_),
    .Q_N(_06792_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16940_ (.CLK(_01258_),
    .RESET_B(net5863),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_06918_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16941_ (.CLK(net5347),
    .RESET_B(net5855),
    .D(_00214_),
    .Q_N(_06791_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16942_ (.CLK(_01259_),
    .RESET_B(net5856),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_06919_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16943_ (.CLK(net5221),
    .RESET_B(net5727),
    .D(_00215_),
    .Q_N(_06790_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16944_ (.CLK(_01260_),
    .RESET_B(net5729),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_06789_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16945_ (.CLK(_01261_),
    .RESET_B(net22),
    .D(_01802_),
    .Q_N(_06920_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.out ));
 sg13g2_dfrbp_1 _16946_ (.CLK(net5403),
    .RESET_B(net5912),
    .D(_00191_),
    .Q_N(_06788_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _16947_ (.CLK(_01262_),
    .RESET_B(net5917),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.u_mux_shift.data ),
    .Q_N(_06921_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _16948_ (.CLK(net5408),
    .RESET_B(net5917),
    .D(_00170_),
    .Q_N(_06787_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16949_ (.CLK(_01263_),
    .RESET_B(net5920),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_06922_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16950_ (.CLK(net5411),
    .RESET_B(net5920),
    .D(_00181_),
    .Q_N(_06786_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16951_ (.CLK(_01264_),
    .RESET_B(net5920),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_06923_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16952_ (.CLK(net5412),
    .RESET_B(net5921),
    .D(_00184_),
    .Q_N(_06785_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16953_ (.CLK(_01265_),
    .RESET_B(net5921),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_06924_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16954_ (.CLK(net5412),
    .RESET_B(net5921),
    .D(_00185_),
    .Q_N(_06784_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16955_ (.CLK(_01266_),
    .RESET_B(net5921),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_06925_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16956_ (.CLK(net5413),
    .RESET_B(net5922),
    .D(_00186_),
    .Q_N(_06783_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16957_ (.CLK(_01267_),
    .RESET_B(net5918),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_06926_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16958_ (.CLK(net5409),
    .RESET_B(net5918),
    .D(_00187_),
    .Q_N(_06782_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16959_ (.CLK(_01268_),
    .RESET_B(net5907),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_06927_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16960_ (.CLK(net5398),
    .RESET_B(net5907),
    .D(_00188_),
    .Q_N(_06781_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16961_ (.CLK(_01269_),
    .RESET_B(net5907),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_06928_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16962_ (.CLK(net5397),
    .RESET_B(net5906),
    .D(_00189_),
    .Q_N(_06780_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16963_ (.CLK(_01270_),
    .RESET_B(net5906),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_06929_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16964_ (.CLK(net5337),
    .RESET_B(net5847),
    .D(_00190_),
    .Q_N(_06779_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16965_ (.CLK(_01271_),
    .RESET_B(net5847),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_06930_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _16966_ (.CLK(net5332),
    .RESET_B(net5842),
    .D(_00160_),
    .Q_N(_06778_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16967_ (.CLK(_01272_),
    .RESET_B(net5842),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_06931_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16968_ (.CLK(net5332),
    .RESET_B(net5842),
    .D(_00161_),
    .Q_N(_06777_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16969_ (.CLK(_01273_),
    .RESET_B(net5842),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_06932_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16970_ (.CLK(net5326),
    .RESET_B(net5836),
    .D(_00162_),
    .Q_N(_06776_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16971_ (.CLK(_01274_),
    .RESET_B(net5836),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_06933_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16972_ (.CLK(net5326),
    .RESET_B(net5836),
    .D(_00163_),
    .Q_N(_06775_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16973_ (.CLK(_01275_),
    .RESET_B(net5836),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_06934_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16974_ (.CLK(net5326),
    .RESET_B(net5836),
    .D(_00164_),
    .Q_N(_06774_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16975_ (.CLK(_01276_),
    .RESET_B(net5836),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_06935_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16976_ (.CLK(net5326),
    .RESET_B(net5836),
    .D(_00165_),
    .Q_N(_06773_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16977_ (.CLK(_01277_),
    .RESET_B(net5836),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_06936_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16978_ (.CLK(net5327),
    .RESET_B(net5837),
    .D(_00166_),
    .Q_N(_06772_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16979_ (.CLK(_01278_),
    .RESET_B(net5837),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_06937_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16980_ (.CLK(net5322),
    .RESET_B(net5832),
    .D(_00167_),
    .Q_N(_06771_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16981_ (.CLK(_01279_),
    .RESET_B(net5832),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_06938_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16982_ (.CLK(net5319),
    .RESET_B(net5829),
    .D(_00168_),
    .Q_N(_06770_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16983_ (.CLK(_01280_),
    .RESET_B(net5785),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_06939_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16984_ (.CLK(net5274),
    .RESET_B(net5784),
    .D(_00169_),
    .Q_N(_06769_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16985_ (.CLK(_01281_),
    .RESET_B(net5783),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_06940_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16986_ (.CLK(net5262),
    .RESET_B(net5772),
    .D(_00171_),
    .Q_N(_06768_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16987_ (.CLK(_01282_),
    .RESET_B(net5772),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_06941_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16988_ (.CLK(net5219),
    .RESET_B(net5729),
    .D(_00172_),
    .Q_N(_06767_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16989_ (.CLK(_01283_),
    .RESET_B(net5729),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_06942_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16990_ (.CLK(net5213),
    .RESET_B(net5723),
    .D(_00173_),
    .Q_N(_06766_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16991_ (.CLK(_01284_),
    .RESET_B(net5723),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_06943_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16992_ (.CLK(net5213),
    .RESET_B(net5723),
    .D(_00174_),
    .Q_N(_06765_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16993_ (.CLK(_01285_),
    .RESET_B(net5723),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_06944_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16994_ (.CLK(net5209),
    .RESET_B(net5719),
    .D(_00175_),
    .Q_N(_06764_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16995_ (.CLK(_01286_),
    .RESET_B(net5723),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_06945_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16996_ (.CLK(net5209),
    .RESET_B(net5719),
    .D(_00176_),
    .Q_N(_06763_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16997_ (.CLK(_01287_),
    .RESET_B(net5720),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_06946_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _16998_ (.CLK(net5211),
    .RESET_B(net5720),
    .D(_00177_),
    .Q_N(_06762_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _16999_ (.CLK(_01288_),
    .RESET_B(net5720),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_06947_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17000_ (.CLK(net5211),
    .RESET_B(net5720),
    .D(_00178_),
    .Q_N(_06761_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17001_ (.CLK(_01289_),
    .RESET_B(net5721),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_06948_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17002_ (.CLK(net5211),
    .RESET_B(net5720),
    .D(_00179_),
    .Q_N(_06760_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17003_ (.CLK(_01290_),
    .RESET_B(net5721),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_06949_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17004_ (.CLK(net5209),
    .RESET_B(net5719),
    .D(_00180_),
    .Q_N(_06759_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17005_ (.CLK(_01291_),
    .RESET_B(net5719),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_06950_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17006_ (.CLK(net5210),
    .RESET_B(net5719),
    .D(_00182_),
    .Q_N(_06758_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17007_ (.CLK(_01292_),
    .RESET_B(net5724),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_06951_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17008_ (.CLK(net5209),
    .RESET_B(net5719),
    .D(_00183_),
    .Q_N(_06757_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17009_ (.CLK(_01293_),
    .RESET_B(net5719),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_06756_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17010_ (.CLK(_01294_),
    .RESET_B(net23),
    .D(_01803_),
    .Q_N(_06952_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.out ));
 sg13g2_dfrbp_1 _17011_ (.CLK(net5258),
    .RESET_B(net5768),
    .D(_00159_),
    .Q_N(_06755_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _17012_ (.CLK(_01295_),
    .RESET_B(net5768),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.data ),
    .Q_N(_06953_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17013_ (.CLK(net5258),
    .RESET_B(net5768),
    .D(_00138_),
    .Q_N(_06754_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17014_ (.CLK(_01296_),
    .RESET_B(net5770),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_06954_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17015_ (.CLK(net5258),
    .RESET_B(net5768),
    .D(_00149_),
    .Q_N(_06753_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17016_ (.CLK(_01297_),
    .RESET_B(net5770),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_06955_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17017_ (.CLK(net5232),
    .RESET_B(net5743),
    .D(_00152_),
    .Q_N(_06752_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17018_ (.CLK(_01298_),
    .RESET_B(net5742),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_06956_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17019_ (.CLK(net5232),
    .RESET_B(net5743),
    .D(_00153_),
    .Q_N(_06751_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17020_ (.CLK(_01299_),
    .RESET_B(net5742),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_06957_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17021_ (.CLK(net5232),
    .RESET_B(net5742),
    .D(_00154_),
    .Q_N(_06750_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17022_ (.CLK(_01300_),
    .RESET_B(net5742),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_06958_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17023_ (.CLK(net5232),
    .RESET_B(net5742),
    .D(_00155_),
    .Q_N(_06749_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17024_ (.CLK(_01301_),
    .RESET_B(net5742),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_06959_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17025_ (.CLK(net5232),
    .RESET_B(net5742),
    .D(_00156_),
    .Q_N(_06748_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17026_ (.CLK(_01302_),
    .RESET_B(net5742),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_06960_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17027_ (.CLK(net5230),
    .RESET_B(net5740),
    .D(_00157_),
    .Q_N(_06747_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17028_ (.CLK(_01303_),
    .RESET_B(net5740),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_06961_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17029_ (.CLK(net5231),
    .RESET_B(net5740),
    .D(_00158_),
    .Q_N(_06746_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17030_ (.CLK(_01304_),
    .RESET_B(net5740),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_06962_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17031_ (.CLK(net5230),
    .RESET_B(net5740),
    .D(_00128_),
    .Q_N(_06745_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17032_ (.CLK(_01305_),
    .RESET_B(net5740),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_06963_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17033_ (.CLK(net5230),
    .RESET_B(net5740),
    .D(_00129_),
    .Q_N(_06744_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17034_ (.CLK(_01306_),
    .RESET_B(net5744),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_06964_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17035_ (.CLK(net5230),
    .RESET_B(net5741),
    .D(_00130_),
    .Q_N(_06743_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17036_ (.CLK(_01307_),
    .RESET_B(net5744),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_06965_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17037_ (.CLK(net5234),
    .RESET_B(net5744),
    .D(_00131_),
    .Q_N(_06742_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17038_ (.CLK(_01308_),
    .RESET_B(net5744),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_06966_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17039_ (.CLK(net5234),
    .RESET_B(net5744),
    .D(_00132_),
    .Q_N(_06741_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17040_ (.CLK(_01309_),
    .RESET_B(net5744),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_06967_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17041_ (.CLK(net5231),
    .RESET_B(net5741),
    .D(_00133_),
    .Q_N(_06740_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17042_ (.CLK(_01310_),
    .RESET_B(net5741),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_06968_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17043_ (.CLK(net5230),
    .RESET_B(net5740),
    .D(_00134_),
    .Q_N(_06739_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17044_ (.CLK(_01311_),
    .RESET_B(net5746),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_06969_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17045_ (.CLK(net5233),
    .RESET_B(net5743),
    .D(_00135_),
    .Q_N(_06738_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17046_ (.CLK(_01312_),
    .RESET_B(net5743),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_06970_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17047_ (.CLK(net5198),
    .RESET_B(net5708),
    .D(_00136_),
    .Q_N(_06737_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17048_ (.CLK(_01313_),
    .RESET_B(net5708),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_06971_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17049_ (.CLK(net5198),
    .RESET_B(net5708),
    .D(_00137_),
    .Q_N(_06736_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17050_ (.CLK(_01314_),
    .RESET_B(net5708),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_06972_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17051_ (.CLK(net5215),
    .RESET_B(net5727),
    .D(_00139_),
    .Q_N(_06735_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17052_ (.CLK(_01315_),
    .RESET_B(net5727),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_06973_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17053_ (.CLK(net5215),
    .RESET_B(net5727),
    .D(_00140_),
    .Q_N(_06734_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17054_ (.CLK(_01316_),
    .RESET_B(net5727),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_06974_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17055_ (.CLK(net5208),
    .RESET_B(net5718),
    .D(_00141_),
    .Q_N(_06733_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17056_ (.CLK(_01317_),
    .RESET_B(net5714),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_06975_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17057_ (.CLK(net5208),
    .RESET_B(net5718),
    .D(_00142_),
    .Q_N(_06732_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17058_ (.CLK(_01318_),
    .RESET_B(net5715),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_06976_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17059_ (.CLK(net5205),
    .RESET_B(net5715),
    .D(_00143_),
    .Q_N(_06731_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17060_ (.CLK(_01319_),
    .RESET_B(net5715),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_06977_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17061_ (.CLK(net5205),
    .RESET_B(net5715),
    .D(_00144_),
    .Q_N(_06730_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17062_ (.CLK(_01320_),
    .RESET_B(net5716),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_06978_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17063_ (.CLK(net5206),
    .RESET_B(net5716),
    .D(_00145_),
    .Q_N(_06729_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17064_ (.CLK(_01321_),
    .RESET_B(net5716),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_06979_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17065_ (.CLK(net5213),
    .RESET_B(net5722),
    .D(_00146_),
    .Q_N(_06728_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17066_ (.CLK(_01322_),
    .RESET_B(net5722),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_06980_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17067_ (.CLK(net5212),
    .RESET_B(net5722),
    .D(_00147_),
    .Q_N(_06727_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17068_ (.CLK(_01323_),
    .RESET_B(net5721),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_06981_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17069_ (.CLK(net5212),
    .RESET_B(net5721),
    .D(_00148_),
    .Q_N(_06726_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17070_ (.CLK(_01324_),
    .RESET_B(net5721),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_06982_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17071_ (.CLK(net5212),
    .RESET_B(net5721),
    .D(_00150_),
    .Q_N(_06725_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17072_ (.CLK(_01325_),
    .RESET_B(net5722),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_06983_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17073_ (.CLK(net5212),
    .RESET_B(net5721),
    .D(_00151_),
    .Q_N(_06724_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17074_ (.CLK(_01326_),
    .RESET_B(net5724),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_06723_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17075_ (.CLK(_01327_),
    .RESET_B(net53),
    .D(_01804_),
    .Q_N(_06984_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.out ));
 sg13g2_dfrbp_1 _17076_ (.CLK(net5566),
    .RESET_B(net6075),
    .D(_00127_),
    .Q_N(_06722_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _17077_ (.CLK(_01328_),
    .RESET_B(net6075),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.u_mux_shift.data ),
    .Q_N(_06985_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17078_ (.CLK(net5566),
    .RESET_B(net6075),
    .D(_00106_),
    .Q_N(_06721_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17079_ (.CLK(_01329_),
    .RESET_B(net6075),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_06986_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17080_ (.CLK(net5565),
    .RESET_B(net6074),
    .D(_00117_),
    .Q_N(_06720_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17081_ (.CLK(_01330_),
    .RESET_B(net6080),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_06987_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17082_ (.CLK(net5562),
    .RESET_B(net6071),
    .D(_00120_),
    .Q_N(_06719_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17083_ (.CLK(_01331_),
    .RESET_B(net6089),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_06988_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17084_ (.CLK(net5580),
    .RESET_B(net6089),
    .D(_00121_),
    .Q_N(_06718_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17085_ (.CLK(_01332_),
    .RESET_B(net6089),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_06989_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17086_ (.CLK(net5581),
    .RESET_B(net6090),
    .D(_00122_),
    .Q_N(_06717_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17087_ (.CLK(_01333_),
    .RESET_B(net6090),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_06990_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17088_ (.CLK(net5581),
    .RESET_B(net6090),
    .D(_00123_),
    .Q_N(_06716_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17089_ (.CLK(_01334_),
    .RESET_B(net6090),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_06991_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17090_ (.CLK(net5581),
    .RESET_B(net6090),
    .D(_00124_),
    .Q_N(_06715_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17091_ (.CLK(_01335_),
    .RESET_B(net6133),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_06992_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17092_ (.CLK(net5624),
    .RESET_B(net6133),
    .D(_00125_),
    .Q_N(_06714_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17093_ (.CLK(_01336_),
    .RESET_B(net6133),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_06993_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17094_ (.CLK(net5581),
    .RESET_B(net6090),
    .D(_00126_),
    .Q_N(_06713_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17095_ (.CLK(_01337_),
    .RESET_B(net6101),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_06994_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17096_ (.CLK(net5592),
    .RESET_B(net6101),
    .D(_00096_),
    .Q_N(_06712_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17097_ (.CLK(_01338_),
    .RESET_B(net6101),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_06995_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17098_ (.CLK(net5593),
    .RESET_B(net6102),
    .D(_00097_),
    .Q_N(_06711_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17099_ (.CLK(_01339_),
    .RESET_B(net6102),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_06996_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17100_ (.CLK(net5591),
    .RESET_B(net6099),
    .D(_00098_),
    .Q_N(_06710_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17101_ (.CLK(_01340_),
    .RESET_B(net6099),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_06997_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17102_ (.CLK(net5602),
    .RESET_B(net6111),
    .D(_00099_),
    .Q_N(_06709_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17103_ (.CLK(_01341_),
    .RESET_B(net6112),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_06998_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17104_ (.CLK(net5598),
    .RESET_B(net6107),
    .D(_00100_),
    .Q_N(_06708_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17105_ (.CLK(_01342_),
    .RESET_B(net6078),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_06999_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17106_ (.CLK(net5494),
    .RESET_B(net6003),
    .D(_00101_),
    .Q_N(_06707_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17107_ (.CLK(_01343_),
    .RESET_B(net6004),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_07000_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17108_ (.CLK(net5483),
    .RESET_B(net5992),
    .D(_00102_),
    .Q_N(_06706_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17109_ (.CLK(_01344_),
    .RESET_B(net5992),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_07001_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17110_ (.CLK(net5480),
    .RESET_B(net5989),
    .D(_00103_),
    .Q_N(_06705_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17111_ (.CLK(_01345_),
    .RESET_B(net5985),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_07002_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17112_ (.CLK(net5429),
    .RESET_B(net5938),
    .D(_00104_),
    .Q_N(_06704_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17113_ (.CLK(_01346_),
    .RESET_B(net5938),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_07003_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17114_ (.CLK(net5429),
    .RESET_B(net5938),
    .D(_00105_),
    .Q_N(_06703_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17115_ (.CLK(_01347_),
    .RESET_B(net5940),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_07004_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17116_ (.CLK(net5419),
    .RESET_B(net5928),
    .D(_00107_),
    .Q_N(_06702_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17117_ (.CLK(_01348_),
    .RESET_B(net5926),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_07005_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17118_ (.CLK(net5353),
    .RESET_B(net5861),
    .D(_00108_),
    .Q_N(_06701_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17119_ (.CLK(_01349_),
    .RESET_B(net5861),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_07006_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17120_ (.CLK(net5350),
    .RESET_B(net5858),
    .D(_00109_),
    .Q_N(_06700_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17121_ (.CLK(_01350_),
    .RESET_B(net5858),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_07007_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17122_ (.CLK(net5350),
    .RESET_B(net5858),
    .D(_00110_),
    .Q_N(_06699_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17123_ (.CLK(_01351_),
    .RESET_B(net5858),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_07008_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17124_ (.CLK(net5345),
    .RESET_B(net5854),
    .D(_00111_),
    .Q_N(_06698_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17125_ (.CLK(_01352_),
    .RESET_B(net5854),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_07009_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17126_ (.CLK(net5344),
    .RESET_B(net5853),
    .D(_00112_),
    .Q_N(_06697_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17127_ (.CLK(_01353_),
    .RESET_B(net5853),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_07010_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17128_ (.CLK(net5344),
    .RESET_B(net5853),
    .D(_00113_),
    .Q_N(_06696_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17129_ (.CLK(_01354_),
    .RESET_B(net5853),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_07011_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17130_ (.CLK(net5344),
    .RESET_B(net5853),
    .D(_00114_),
    .Q_N(_06695_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17131_ (.CLK(_01355_),
    .RESET_B(net5853),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_07012_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17132_ (.CLK(net5300),
    .RESET_B(net5810),
    .D(_00115_),
    .Q_N(_06694_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17133_ (.CLK(_01356_),
    .RESET_B(net5810),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_07013_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17134_ (.CLK(net5300),
    .RESET_B(net5810),
    .D(_00116_),
    .Q_N(_06693_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17135_ (.CLK(_01357_),
    .RESET_B(net5810),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_07014_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17136_ (.CLK(net5303),
    .RESET_B(net5812),
    .D(_00118_),
    .Q_N(_06692_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17137_ (.CLK(_01358_),
    .RESET_B(net5812),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_07015_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17138_ (.CLK(net5198),
    .RESET_B(net5708),
    .D(_00119_),
    .Q_N(_06691_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17139_ (.CLK(_01359_),
    .RESET_B(net5727),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_06690_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17140_ (.CLK(_01360_),
    .RESET_B(net87),
    .D(_01805_),
    .Q_N(_07016_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.out ));
 sg13g2_dfrbp_1 _17141_ (.CLK(net5471),
    .RESET_B(net5980),
    .D(_00095_),
    .Q_N(_06689_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _17142_ (.CLK(_01361_),
    .RESET_B(net5980),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.u_mux_shift.data ),
    .Q_N(_07017_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17143_ (.CLK(net5466),
    .RESET_B(net5975),
    .D(_00074_),
    .Q_N(_06688_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17144_ (.CLK(_01362_),
    .RESET_B(net5975),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_07018_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17145_ (.CLK(net5466),
    .RESET_B(net5975),
    .D(_00085_),
    .Q_N(_06687_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17146_ (.CLK(_01363_),
    .RESET_B(net6024),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_07019_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17147_ (.CLK(net5515),
    .RESET_B(net6024),
    .D(_00088_),
    .Q_N(_06686_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17148_ (.CLK(_01364_),
    .RESET_B(net6024),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_07020_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17149_ (.CLK(net5517),
    .RESET_B(net6026),
    .D(_00089_),
    .Q_N(_06685_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17150_ (.CLK(_01365_),
    .RESET_B(net6026),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_07021_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17151_ (.CLK(net5519),
    .RESET_B(net6028),
    .D(_00090_),
    .Q_N(_06684_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17152_ (.CLK(_01366_),
    .RESET_B(net6028),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_07022_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17153_ (.CLK(net5511),
    .RESET_B(net6020),
    .D(_00091_),
    .Q_N(_06683_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17154_ (.CLK(_01367_),
    .RESET_B(net6020),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_07023_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17155_ (.CLK(net5505),
    .RESET_B(net6014),
    .D(_00092_),
    .Q_N(_06682_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17156_ (.CLK(_01368_),
    .RESET_B(net6024),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_07024_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17157_ (.CLK(net5466),
    .RESET_B(net5975),
    .D(_00093_),
    .Q_N(_06681_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17158_ (.CLK(_01369_),
    .RESET_B(net5980),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_07025_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17159_ (.CLK(net5471),
    .RESET_B(net5980),
    .D(_00094_),
    .Q_N(_06680_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17160_ (.CLK(_01370_),
    .RESET_B(net5980),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_07026_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17161_ (.CLK(net5471),
    .RESET_B(net5980),
    .D(_00064_),
    .Q_N(_06679_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17162_ (.CLK(_01371_),
    .RESET_B(net5980),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_07027_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17163_ (.CLK(net5449),
    .RESET_B(net5958),
    .D(_00065_),
    .Q_N(_06678_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17164_ (.CLK(_01372_),
    .RESET_B(net5960),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_07028_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17165_ (.CLK(net5450),
    .RESET_B(net5959),
    .D(_00066_),
    .Q_N(_06677_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17166_ (.CLK(_01373_),
    .RESET_B(net5959),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_07029_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17167_ (.CLK(net5452),
    .RESET_B(net5961),
    .D(_00067_),
    .Q_N(_06676_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17168_ (.CLK(_01374_),
    .RESET_B(net5961),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_07030_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17169_ (.CLK(net5452),
    .RESET_B(net5961),
    .D(_00068_),
    .Q_N(_06675_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17170_ (.CLK(_01375_),
    .RESET_B(net5961),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_07031_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17171_ (.CLK(net5453),
    .RESET_B(net5962),
    .D(_00069_),
    .Q_N(_06674_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17172_ (.CLK(_01376_),
    .RESET_B(net5961),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_07032_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17173_ (.CLK(net5453),
    .RESET_B(net5962),
    .D(_00070_),
    .Q_N(_06673_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17174_ (.CLK(_01377_),
    .RESET_B(net5962),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_07033_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17175_ (.CLK(net5453),
    .RESET_B(net5962),
    .D(_00071_),
    .Q_N(_06672_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17176_ (.CLK(_01378_),
    .RESET_B(net5952),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_07034_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17177_ (.CLK(net5407),
    .RESET_B(net5916),
    .D(_00072_),
    .Q_N(_06671_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17178_ (.CLK(_01379_),
    .RESET_B(net5916),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_07035_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17179_ (.CLK(net5379),
    .RESET_B(net5888),
    .D(_00073_),
    .Q_N(_06670_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17180_ (.CLK(_01380_),
    .RESET_B(net5889),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_07036_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17181_ (.CLK(net5380),
    .RESET_B(net5888),
    .D(_00075_),
    .Q_N(_06669_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17182_ (.CLK(_01381_),
    .RESET_B(net5882),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_07037_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17183_ (.CLK(net5355),
    .RESET_B(net5864),
    .D(_00076_),
    .Q_N(_06668_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17184_ (.CLK(_01382_),
    .RESET_B(net5864),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_07038_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17185_ (.CLK(net5350),
    .RESET_B(net5858),
    .D(_00077_),
    .Q_N(_06667_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17186_ (.CLK(_01383_),
    .RESET_B(net5858),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_07039_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17187_ (.CLK(net5345),
    .RESET_B(net5854),
    .D(_00078_),
    .Q_N(_06666_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17188_ (.CLK(_01384_),
    .RESET_B(net5854),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_07040_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17189_ (.CLK(net5300),
    .RESET_B(net5810),
    .D(_00079_),
    .Q_N(_06665_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17190_ (.CLK(_01385_),
    .RESET_B(net5810),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_07041_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17191_ (.CLK(net5299),
    .RESET_B(net5809),
    .D(_00080_),
    .Q_N(_06664_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17192_ (.CLK(_01386_),
    .RESET_B(net5809),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_07042_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17193_ (.CLK(net5299),
    .RESET_B(net5809),
    .D(_00081_),
    .Q_N(_06663_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17194_ (.CLK(_01387_),
    .RESET_B(net5809),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_07043_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17195_ (.CLK(net5284),
    .RESET_B(net5794),
    .D(_00082_),
    .Q_N(_06662_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17196_ (.CLK(_01388_),
    .RESET_B(net5794),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_07044_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17197_ (.CLK(net5284),
    .RESET_B(net5794),
    .D(_00083_),
    .Q_N(_06661_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17198_ (.CLK(_01389_),
    .RESET_B(net5794),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_07045_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17199_ (.CLK(net5283),
    .RESET_B(net5793),
    .D(_00084_),
    .Q_N(_06660_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17200_ (.CLK(_01390_),
    .RESET_B(net5793),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_07046_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17201_ (.CLK(net5294),
    .RESET_B(net5804),
    .D(_00086_),
    .Q_N(_06659_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17202_ (.CLK(_01391_),
    .RESET_B(net5850),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_07047_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17203_ (.CLK(net5220),
    .RESET_B(net5730),
    .D(_00087_),
    .Q_N(_06658_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17204_ (.CLK(_01392_),
    .RESET_B(net5730),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_06657_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17205_ (.CLK(_01393_),
    .RESET_B(net121),
    .D(_01806_),
    .Q_N(_07048_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.out ));
 sg13g2_dfrbp_1 _17206_ (.CLK(net5324),
    .RESET_B(net5834),
    .D(_00063_),
    .Q_N(_06656_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _17207_ (.CLK(_01394_),
    .RESET_B(net5834),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.u_mux_shift.data ),
    .Q_N(_07049_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17208_ (.CLK(net5324),
    .RESET_B(net5835),
    .D(_00042_),
    .Q_N(_06655_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17209_ (.CLK(_01395_),
    .RESET_B(net5835),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_07050_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17210_ (.CLK(net5325),
    .RESET_B(net5835),
    .D(_00053_),
    .Q_N(_06654_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17211_ (.CLK(_01396_),
    .RESET_B(net5835),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_07051_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17212_ (.CLK(net5324),
    .RESET_B(net5834),
    .D(_00056_),
    .Q_N(_06653_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17213_ (.CLK(_01397_),
    .RESET_B(net5834),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_07052_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17214_ (.CLK(net5324),
    .RESET_B(net5834),
    .D(_00057_),
    .Q_N(_06652_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17215_ (.CLK(_01398_),
    .RESET_B(net5834),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_07053_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17216_ (.CLK(net5324),
    .RESET_B(net5834),
    .D(_00058_),
    .Q_N(_06651_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17217_ (.CLK(_01399_),
    .RESET_B(net5834),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_07054_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17218_ (.CLK(net5340),
    .RESET_B(net5850),
    .D(_00059_),
    .Q_N(_06650_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17219_ (.CLK(_01400_),
    .RESET_B(net5803),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_07055_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17220_ (.CLK(net5292),
    .RESET_B(net5802),
    .D(_00060_),
    .Q_N(_06649_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17221_ (.CLK(_01401_),
    .RESET_B(net5803),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_07056_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17222_ (.CLK(net5293),
    .RESET_B(net5803),
    .D(_00061_),
    .Q_N(_06648_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17223_ (.CLK(_01402_),
    .RESET_B(net5803),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_07057_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17224_ (.CLK(net5292),
    .RESET_B(net5802),
    .D(_00062_),
    .Q_N(_06647_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17225_ (.CLK(_01403_),
    .RESET_B(net5802),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_07058_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17226_ (.CLK(net5292),
    .RESET_B(net5802),
    .D(_00032_),
    .Q_N(_06646_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17227_ (.CLK(_01404_),
    .RESET_B(net5802),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_07059_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17228_ (.CLK(net5289),
    .RESET_B(net5799),
    .D(_00033_),
    .Q_N(_06645_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17229_ (.CLK(_01405_),
    .RESET_B(net5799),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_07060_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17230_ (.CLK(net5289),
    .RESET_B(net5799),
    .D(_00034_),
    .Q_N(_06644_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17231_ (.CLK(_01406_),
    .RESET_B(net5799),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_07061_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17232_ (.CLK(net5289),
    .RESET_B(net5799),
    .D(_00035_),
    .Q_N(_06643_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17233_ (.CLK(_01407_),
    .RESET_B(net5799),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_07062_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17234_ (.CLK(net5289),
    .RESET_B(net5799),
    .D(_00036_),
    .Q_N(_06642_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17235_ (.CLK(_01408_),
    .RESET_B(net5799),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_07063_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17236_ (.CLK(net5294),
    .RESET_B(net5804),
    .D(_00037_),
    .Q_N(_06641_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17237_ (.CLK(_01409_),
    .RESET_B(net5804),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_07064_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17238_ (.CLK(net5295),
    .RESET_B(net5805),
    .D(_00038_),
    .Q_N(_06640_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17239_ (.CLK(_01410_),
    .RESET_B(net5805),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_07065_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17240_ (.CLK(net5269),
    .RESET_B(net5779),
    .D(_00039_),
    .Q_N(_06639_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17241_ (.CLK(_01411_),
    .RESET_B(net5779),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_07066_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17242_ (.CLK(net5260),
    .RESET_B(net5770),
    .D(_00040_),
    .Q_N(_06638_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17243_ (.CLK(_01412_),
    .RESET_B(net5770),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_07067_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17244_ (.CLK(net5258),
    .RESET_B(net5768),
    .D(_00041_),
    .Q_N(_06637_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17245_ (.CLK(_01413_),
    .RESET_B(net5768),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_07068_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17246_ (.CLK(net5258),
    .RESET_B(net5768),
    .D(_00043_),
    .Q_N(_06636_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17247_ (.CLK(_01414_),
    .RESET_B(net5765),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_07069_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17248_ (.CLK(net5216),
    .RESET_B(net5725),
    .D(_00044_),
    .Q_N(_06635_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17249_ (.CLK(_01415_),
    .RESET_B(net5765),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_07070_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17250_ (.CLK(net5217),
    .RESET_B(net5726),
    .D(_00045_),
    .Q_N(_06634_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17251_ (.CLK(_01416_),
    .RESET_B(net5725),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_07071_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17252_ (.CLK(net5216),
    .RESET_B(net5726),
    .D(_00046_),
    .Q_N(_06633_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17253_ (.CLK(_01417_),
    .RESET_B(net5725),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_07072_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17254_ (.CLK(net5216),
    .RESET_B(net5725),
    .D(_00047_),
    .Q_N(_06632_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17255_ (.CLK(_01418_),
    .RESET_B(net5725),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_07073_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17256_ (.CLK(net5216),
    .RESET_B(net5725),
    .D(_00048_),
    .Q_N(_06631_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17257_ (.CLK(_01419_),
    .RESET_B(net5725),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_07074_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17258_ (.CLK(net5215),
    .RESET_B(net5727),
    .D(_00049_),
    .Q_N(_06630_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17259_ (.CLK(_01420_),
    .RESET_B(net5725),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_07075_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17260_ (.CLK(net5215),
    .RESET_B(net5727),
    .D(_00050_),
    .Q_N(_06629_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17261_ (.CLK(_01421_),
    .RESET_B(net5728),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_07076_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17262_ (.CLK(net5218),
    .RESET_B(net5728),
    .D(_00051_),
    .Q_N(_06628_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17263_ (.CLK(_01422_),
    .RESET_B(net5728),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_07077_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17264_ (.CLK(net5218),
    .RESET_B(net5728),
    .D(_00052_),
    .Q_N(_06627_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17265_ (.CLK(_01423_),
    .RESET_B(net5728),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_07078_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17266_ (.CLK(net5218),
    .RESET_B(net5728),
    .D(_00054_),
    .Q_N(_06626_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17267_ (.CLK(_01424_),
    .RESET_B(net5728),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_07079_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17268_ (.CLK(net5219),
    .RESET_B(net5729),
    .D(_00055_),
    .Q_N(_06625_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17269_ (.CLK(_01425_),
    .RESET_B(net5729),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_07080_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17270_ (.CLK(net5283),
    .RESET_B(net5793),
    .D(_00031_),
    .Q_N(_06624_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _17271_ (.CLK(_01426_),
    .RESET_B(net5793),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.u_mux_shift.data ),
    .Q_N(_07081_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17272_ (.CLK(net5281),
    .RESET_B(net5792),
    .D(_00010_),
    .Q_N(_06623_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17273_ (.CLK(_01427_),
    .RESET_B(net5791),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_07082_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17274_ (.CLK(net5286),
    .RESET_B(net5796),
    .D(_00021_),
    .Q_N(_06622_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17275_ (.CLK(_01428_),
    .RESET_B(net5791),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_07083_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17276_ (.CLK(net5281),
    .RESET_B(net5791),
    .D(_00024_),
    .Q_N(_06621_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17277_ (.CLK(_01429_),
    .RESET_B(net5791),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_07084_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17278_ (.CLK(net5281),
    .RESET_B(net5791),
    .D(_00025_),
    .Q_N(_06620_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17279_ (.CLK(_01430_),
    .RESET_B(net5791),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_07085_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17280_ (.CLK(net5281),
    .RESET_B(net5791),
    .D(_00026_),
    .Q_N(_06619_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17281_ (.CLK(_01431_),
    .RESET_B(net5792),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_07086_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17282_ (.CLK(net5282),
    .RESET_B(net5792),
    .D(_00027_),
    .Q_N(_06618_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17283_ (.CLK(_01432_),
    .RESET_B(net5792),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_07087_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17284_ (.CLK(net5283),
    .RESET_B(net5793),
    .D(_00028_),
    .Q_N(_06617_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17285_ (.CLK(_01433_),
    .RESET_B(net5793),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_07088_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17286_ (.CLK(net5283),
    .RESET_B(net5794),
    .D(_00029_),
    .Q_N(_06616_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17287_ (.CLK(_01434_),
    .RESET_B(net5793),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_07089_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17288_ (.CLK(net5298),
    .RESET_B(net5808),
    .D(_00030_),
    .Q_N(_06615_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17289_ (.CLK(_01435_),
    .RESET_B(net5808),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_07090_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _17290_ (.CLK(net5297),
    .RESET_B(net5807),
    .D(_00000_),
    .Q_N(_06614_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17291_ (.CLK(_01436_),
    .RESET_B(net5807),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_07091_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17292_ (.CLK(net5592),
    .RESET_B(net6101),
    .D(net5151),
    .Q_N(_07092_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ));
 sg13g2_dfrbp_1 _17293_ (.CLK(net5302),
    .RESET_B(net5811),
    .D(_00001_),
    .Q_N(_06613_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17294_ (.CLK(_01437_),
    .RESET_B(net5813),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_07093_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17295_ (.CLK(net5301),
    .RESET_B(net5813),
    .D(_00002_),
    .Q_N(_06612_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17296_ (.CLK(_01438_),
    .RESET_B(net5851),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_07094_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17297_ (.CLK(net5342),
    .RESET_B(net5851),
    .D(_00003_),
    .Q_N(_06611_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17298_ (.CLK(_01439_),
    .RESET_B(net5852),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_07095_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17299_ (.CLK(net5342),
    .RESET_B(net5851),
    .D(_00004_),
    .Q_N(_06610_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17300_ (.CLK(_01440_),
    .RESET_B(net5852),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_07096_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17301_ (.CLK(net5303),
    .RESET_B(net5812),
    .D(_00005_),
    .Q_N(_06609_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17302_ (.CLK(_01441_),
    .RESET_B(net5812),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_07097_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17303_ (.CLK(net5302),
    .RESET_B(net5811),
    .D(_00006_),
    .Q_N(_06608_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17304_ (.CLK(_01442_),
    .RESET_B(net5807),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_07098_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17305_ (.CLK(net5299),
    .RESET_B(net5809),
    .D(_00007_),
    .Q_N(_06607_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17306_ (.CLK(_01443_),
    .RESET_B(net5807),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_07099_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17307_ (.CLK(net5238),
    .RESET_B(net5748),
    .D(_00008_),
    .Q_N(_06606_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17308_ (.CLK(_01444_),
    .RESET_B(net5748),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_07100_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17309_ (.CLK(net5237),
    .RESET_B(net5747),
    .D(_00009_),
    .Q_N(_06605_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17310_ (.CLK(_01445_),
    .RESET_B(net5747),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_07101_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17311_ (.CLK(net5229),
    .RESET_B(net5739),
    .D(_00011_),
    .Q_N(_06604_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17312_ (.CLK(_01446_),
    .RESET_B(net5739),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_07102_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17313_ (.CLK(net5225),
    .RESET_B(net5735),
    .D(_00012_),
    .Q_N(_06603_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17314_ (.CLK(_01447_),
    .RESET_B(net5735),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_07103_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17315_ (.CLK(net5196),
    .RESET_B(net5706),
    .D(_00013_),
    .Q_N(_06602_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17316_ (.CLK(_01448_),
    .RESET_B(net5706),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_07104_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17317_ (.CLK(net5191),
    .RESET_B(net5701),
    .D(_00014_),
    .Q_N(_06601_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17318_ (.CLK(_01449_),
    .RESET_B(net5701),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_07105_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17319_ (.CLK(net5177),
    .RESET_B(net5687),
    .D(_00015_),
    .Q_N(_06600_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17320_ (.CLK(_01450_),
    .RESET_B(net5698),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_07106_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17321_ (.CLK(net5188),
    .RESET_B(net5687),
    .D(_00016_),
    .Q_N(_06599_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17322_ (.CLK(_01451_),
    .RESET_B(net5698),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_07107_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17323_ (.CLK(net5177),
    .RESET_B(net5687),
    .D(_00017_),
    .Q_N(_06598_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17324_ (.CLK(_01452_),
    .RESET_B(net5687),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_07108_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17325_ (.CLK(net5177),
    .RESET_B(net5687),
    .D(_00018_),
    .Q_N(_06597_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17326_ (.CLK(_01453_),
    .RESET_B(net5687),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_07109_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17327_ (.CLK(net5177),
    .RESET_B(net5687),
    .D(_00019_),
    .Q_N(_06596_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17328_ (.CLK(_01454_),
    .RESET_B(net5687),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_07110_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17329_ (.CLK(net5180),
    .RESET_B(net5690),
    .D(_00020_),
    .Q_N(_06595_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17330_ (.CLK(_01455_),
    .RESET_B(net5690),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_07111_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17331_ (.CLK(net5180),
    .RESET_B(net5690),
    .D(_00022_),
    .Q_N(_06594_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17332_ (.CLK(_01456_),
    .RESET_B(net5690),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_07112_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17333_ (.CLK(net5199),
    .RESET_B(net5709),
    .D(_00023_),
    .Q_N(_06593_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _17334_ (.CLK(_01457_),
    .RESET_B(net5711),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_07113_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _17335_ (.CLK(net5632),
    .RESET_B(net6141),
    .D(_01167_),
    .Q_N(_07114_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_dfrbp_1 _17336_ (.CLK(net5632),
    .RESET_B(net6141),
    .D(_01177_),
    .Q_N(_07115_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_dfrbp_1 _17337_ (.CLK(net5635),
    .RESET_B(net6144),
    .D(_01178_),
    .Q_N(_07116_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_dfrbp_1 _17338_ (.CLK(net5636),
    .RESET_B(net6145),
    .D(_01179_),
    .Q_N(_07117_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_dfrbp_1 _17339_ (.CLK(net5640),
    .RESET_B(net6149),
    .D(_01180_),
    .Q_N(_07118_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_dfrbp_1 _17340_ (.CLK(net5640),
    .RESET_B(net6149),
    .D(_01181_),
    .Q_N(_07119_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_dfrbp_1 _17341_ (.CLK(net5640),
    .RESET_B(net6149),
    .D(_01182_),
    .Q_N(_07120_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_dfrbp_1 _17342_ (.CLK(net5641),
    .RESET_B(net6150),
    .D(_01183_),
    .Q_N(_07121_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_dfrbp_1 _17343_ (.CLK(net5640),
    .RESET_B(net6149),
    .D(_01184_),
    .Q_N(_07122_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_dfrbp_1 _17344_ (.CLK(net5636),
    .RESET_B(net6145),
    .D(_01185_),
    .Q_N(_07123_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_dfrbp_1 _17345_ (.CLK(net5635),
    .RESET_B(net6144),
    .D(_01168_),
    .Q_N(_07124_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_dfrbp_1 _17346_ (.CLK(net5635),
    .RESET_B(net6144),
    .D(_01169_),
    .Q_N(_07125_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_dfrbp_1 _17347_ (.CLK(net5628),
    .RESET_B(net6137),
    .D(_01170_),
    .Q_N(_07126_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_dfrbp_1 _17348_ (.CLK(net5627),
    .RESET_B(net6136),
    .D(_01171_),
    .Q_N(_07127_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_dfrbp_1 _17349_ (.CLK(net5627),
    .RESET_B(net6136),
    .D(_01172_),
    .Q_N(_07128_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_dfrbp_1 _17350_ (.CLK(net5624),
    .RESET_B(net6133),
    .D(_01173_),
    .Q_N(_07129_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_dfrbp_1 _17351_ (.CLK(net5629),
    .RESET_B(net6138),
    .D(_01174_),
    .Q_N(_07130_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_dfrbp_1 _17352_ (.CLK(net5624),
    .RESET_B(net6133),
    .D(_01175_),
    .Q_N(_07131_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_dfrbp_1 _17353_ (.CLK(net5627),
    .RESET_B(net6136),
    .D(_01176_),
    .Q_N(_07132_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u3.reg_value[18] ));
 sg13g2_dfrbp_1 _17354_ (.CLK(net5631),
    .RESET_B(net6140),
    .D(_01167_),
    .Q_N(_07133_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][0] ));
 sg13g2_dfrbp_1 _17355_ (.CLK(net5632),
    .RESET_B(net6141),
    .D(_01177_),
    .Q_N(_07134_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][1] ));
 sg13g2_dfrbp_1 _17356_ (.CLK(net5632),
    .RESET_B(net6141),
    .D(_01178_),
    .Q_N(_07135_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][2] ));
 sg13g2_dfrbp_1 _17357_ (.CLK(net5643),
    .RESET_B(net6152),
    .D(_01179_),
    .Q_N(_07136_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][3] ));
 sg13g2_dfrbp_1 _17358_ (.CLK(net5636),
    .RESET_B(net6145),
    .D(_01180_),
    .Q_N(_07137_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][4] ));
 sg13g2_dfrbp_1 _17359_ (.CLK(net5640),
    .RESET_B(net6149),
    .D(_01181_),
    .Q_N(_07138_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][5] ));
 sg13g2_dfrbp_1 _17360_ (.CLK(net5641),
    .RESET_B(net6150),
    .D(_01182_),
    .Q_N(_07139_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][6] ));
 sg13g2_dfrbp_1 _17361_ (.CLK(net5641),
    .RESET_B(net6150),
    .D(_01183_),
    .Q_N(_07140_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][7] ));
 sg13g2_dfrbp_1 _17362_ (.CLK(net5639),
    .RESET_B(net6148),
    .D(_01184_),
    .Q_N(_07141_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][8] ));
 sg13g2_dfrbp_1 _17363_ (.CLK(net5639),
    .RESET_B(net6148),
    .D(_01185_),
    .Q_N(_07142_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][9] ));
 sg13g2_dfrbp_1 _17364_ (.CLK(net5643),
    .RESET_B(net6152),
    .D(_01168_),
    .Q_N(_07143_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][10] ));
 sg13g2_dfrbp_1 _17365_ (.CLK(net5643),
    .RESET_B(net6152),
    .D(_01169_),
    .Q_N(_07144_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][11] ));
 sg13g2_dfrbp_1 _17366_ (.CLK(net5632),
    .RESET_B(net6141),
    .D(_01170_),
    .Q_N(_07145_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][12] ));
 sg13g2_dfrbp_1 _17367_ (.CLK(net5632),
    .RESET_B(net6141),
    .D(_01171_),
    .Q_N(_07146_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][13] ));
 sg13g2_dfrbp_1 _17368_ (.CLK(net5632),
    .RESET_B(net6141),
    .D(_01172_),
    .Q_N(_07147_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][14] ));
 sg13g2_dfrbp_1 _17369_ (.CLK(net5631),
    .RESET_B(net6140),
    .D(_01173_),
    .Q_N(_07148_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][15] ));
 sg13g2_dfrbp_1 _17370_ (.CLK(net5631),
    .RESET_B(net6140),
    .D(_01174_),
    .Q_N(_07149_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][16] ));
 sg13g2_dfrbp_1 _17371_ (.CLK(net5629),
    .RESET_B(net6138),
    .D(_01175_),
    .Q_N(_07150_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][17] ));
 sg13g2_dfrbp_1 _17372_ (.CLK(net5624),
    .RESET_B(net6133),
    .D(_01176_),
    .Q_N(_07151_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][18] ));
 sg13g2_dfrbp_1 _17373_ (.CLK(net5637),
    .RESET_B(net6146),
    .D(_01148_),
    .Q_N(_07152_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_dfrbp_1 _17374_ (.CLK(net5635),
    .RESET_B(net6144),
    .D(_01158_),
    .Q_N(_07153_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_dfrbp_1 _17375_ (.CLK(net5636),
    .RESET_B(net6145),
    .D(_01159_),
    .Q_N(_07154_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_dfrbp_1 _17376_ (.CLK(net5636),
    .RESET_B(net6145),
    .D(_01160_),
    .Q_N(_07155_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_dfrbp_1 _17377_ (.CLK(net5639),
    .RESET_B(net6148),
    .D(_01161_),
    .Q_N(_07156_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_dfrbp_1 _17378_ (.CLK(net5642),
    .RESET_B(net6151),
    .D(_01162_),
    .Q_N(_07157_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_dfrbp_1 _17379_ (.CLK(net5642),
    .RESET_B(net6151),
    .D(_01163_),
    .Q_N(_07158_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_dfrbp_1 _17380_ (.CLK(net5642),
    .RESET_B(net6151),
    .D(_01164_),
    .Q_N(_07159_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_dfrbp_1 _17381_ (.CLK(net5634),
    .RESET_B(net6143),
    .D(_01165_),
    .Q_N(_07160_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_dfrbp_1 _17382_ (.CLK(net5634),
    .RESET_B(net6143),
    .D(_01166_),
    .Q_N(_07161_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_dfrbp_1 _17383_ (.CLK(net5634),
    .RESET_B(net6143),
    .D(_01149_),
    .Q_N(_07162_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_dfrbp_1 _17384_ (.CLK(net5628),
    .RESET_B(net6137),
    .D(_01150_),
    .Q_N(_07163_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_dfrbp_1 _17385_ (.CLK(net5628),
    .RESET_B(net6137),
    .D(_01151_),
    .Q_N(_07164_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_dfrbp_1 _17386_ (.CLK(net5628),
    .RESET_B(net6137),
    .D(_01152_),
    .Q_N(_07165_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_dfrbp_1 _17387_ (.CLK(net5626),
    .RESET_B(net6136),
    .D(_01153_),
    .Q_N(_07166_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_dfrbp_1 _17388_ (.CLK(net5626),
    .RESET_B(net6135),
    .D(_01154_),
    .Q_N(_07167_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_dfrbp_1 _17389_ (.CLK(net5627),
    .RESET_B(net6136),
    .D(_01155_),
    .Q_N(_07168_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[16] ));
 sg13g2_dfrbp_1 _17390_ (.CLK(net5627),
    .RESET_B(net6135),
    .D(_01156_),
    .Q_N(_07169_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_dfrbp_1 _17391_ (.CLK(net5625),
    .RESET_B(net6134),
    .D(_01157_),
    .Q_N(_07170_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.u2.reg_value[18] ));
 sg13g2_dfrbp_1 _17392_ (.CLK(net5628),
    .RESET_B(net6137),
    .D(_01148_),
    .Q_N(_07171_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_dfrbp_1 _17393_ (.CLK(net5635),
    .RESET_B(net6144),
    .D(_01158_),
    .Q_N(_07172_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_dfrbp_1 _17394_ (.CLK(net5637),
    .RESET_B(net6146),
    .D(_01159_),
    .Q_N(_07173_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_dfrbp_1 _17395_ (.CLK(net5637),
    .RESET_B(net6146),
    .D(_01160_),
    .Q_N(_07174_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_dfrbp_1 _17396_ (.CLK(net5639),
    .RESET_B(net6148),
    .D(_01161_),
    .Q_N(_07175_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_dfrbp_1 _17397_ (.CLK(net5639),
    .RESET_B(net6148),
    .D(_01162_),
    .Q_N(_07176_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_dfrbp_1 _17398_ (.CLK(net5639),
    .RESET_B(net6148),
    .D(_01163_),
    .Q_N(_07177_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_dfrbp_1 _17399_ (.CLK(net5639),
    .RESET_B(net6148),
    .D(_01164_),
    .Q_N(_07178_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_dfrbp_1 _17400_ (.CLK(net5639),
    .RESET_B(net6148),
    .D(_01165_),
    .Q_N(_07179_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_dfrbp_1 _17401_ (.CLK(net5636),
    .RESET_B(net6145),
    .D(_01166_),
    .Q_N(_07180_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_dfrbp_1 _17402_ (.CLK(net5635),
    .RESET_B(net6144),
    .D(_01149_),
    .Q_N(_07181_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_dfrbp_1 _17403_ (.CLK(net5628),
    .RESET_B(net6137),
    .D(_01150_),
    .Q_N(_07182_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_dfrbp_1 _17404_ (.CLK(net5628),
    .RESET_B(net6137),
    .D(_01151_),
    .Q_N(_07183_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_dfrbp_1 _17405_ (.CLK(net5626),
    .RESET_B(net6135),
    .D(_01152_),
    .Q_N(_07184_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_dfrbp_1 _17406_ (.CLK(net5626),
    .RESET_B(net6135),
    .D(_01153_),
    .Q_N(_07185_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_dfrbp_1 _17407_ (.CLK(net5626),
    .RESET_B(net6135),
    .D(_01154_),
    .Q_N(_07186_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_dfrbp_1 _17408_ (.CLK(net5626),
    .RESET_B(net6135),
    .D(_01155_),
    .Q_N(_07187_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_dfrbp_1 _17409_ (.CLK(net5626),
    .RESET_B(net6135),
    .D(_01156_),
    .Q_N(_07188_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_dfrbp_1 _17410_ (.CLK(net5626),
    .RESET_B(net6135),
    .D(_01157_),
    .Q_N(_07189_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator2_out[18] ));
 sg13g2_dfrbp_1 _17411_ (.CLK(net5635),
    .RESET_B(net6144),
    .D(_01186_),
    .Q_N(_01186_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[0] ));
 sg13g2_dfrbp_1 _17412_ (.CLK(net5635),
    .RESET_B(net6144),
    .D(_01139_),
    .Q_N(_07190_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_dfrbp_1 _17413_ (.CLK(net5636),
    .RESET_B(net6145),
    .D(_01140_),
    .Q_N(_07191_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_dfrbp_1 _17414_ (.CLK(net5636),
    .RESET_B(net6145),
    .D(_01141_),
    .Q_N(_07192_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_dfrbp_1 _17415_ (.CLK(net5634),
    .RESET_B(net6143),
    .D(_01142_),
    .Q_N(_07193_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[4] ));
 sg13g2_dfrbp_1 _17416_ (.CLK(net5638),
    .RESET_B(net6143),
    .D(_01143_),
    .Q_N(_07194_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_dfrbp_1 _17417_ (.CLK(net5634),
    .RESET_B(net6147),
    .D(_01144_),
    .Q_N(_07195_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_dfrbp_1 _17418_ (.CLK(net5634),
    .RESET_B(net6147),
    .D(_01145_),
    .Q_N(_07196_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_dfrbp_1 _17419_ (.CLK(net5638),
    .RESET_B(net6143),
    .D(_01146_),
    .Q_N(_07197_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_dfrbp_1 _17420_ (.CLK(net5634),
    .RESET_B(net6143),
    .D(_01147_),
    .Q_N(_07198_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_dfrbp_1 _17421_ (.CLK(net5634),
    .RESET_B(net6143),
    .D(_01130_),
    .Q_N(_07199_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_dfrbp_1 _17422_ (.CLK(net5625),
    .RESET_B(net6134),
    .D(_01131_),
    .Q_N(_07200_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_dfrbp_1 _17423_ (.CLK(net5625),
    .RESET_B(net6134),
    .D(_01132_),
    .Q_N(_07201_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_dfrbp_1 _17424_ (.CLK(net5625),
    .RESET_B(net6134),
    .D(_01133_),
    .Q_N(_07202_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_dfrbp_1 _17425_ (.CLK(net5625),
    .RESET_B(net6134),
    .D(_01134_),
    .Q_N(_07203_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_dfrbp_1 _17426_ (.CLK(net5625),
    .RESET_B(net6134),
    .D(_01135_),
    .Q_N(_07204_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_dfrbp_1 _17427_ (.CLK(net5625),
    .RESET_B(net6138),
    .D(_01136_),
    .Q_N(_07205_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_dfrbp_1 _17428_ (.CLK(net5629),
    .RESET_B(net6134),
    .D(_01137_),
    .Q_N(_07206_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_dfrbp_1 _17429_ (.CLK(net5625),
    .RESET_B(net6134),
    .D(_01138_),
    .Q_N(_07207_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.u_top_module.integrator1_out[18] ));
 sg13g2_dfrbp_1 _17430_ (.CLK(net5158),
    .RESET_B(net185),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][0] ),
    .Q_N(_07208_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _17431_ (.CLK(net5160),
    .RESET_B(net186),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][1] ),
    .Q_N(_07209_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _17432_ (.CLK(net5161),
    .RESET_B(net187),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][2] ),
    .Q_N(_07210_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _17433_ (.CLK(net5166),
    .RESET_B(net188),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][3] ),
    .Q_N(_07211_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _17434_ (.CLK(net5171),
    .RESET_B(net189),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][4] ),
    .Q_N(_07212_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _17435_ (.CLK(net5170),
    .RESET_B(net190),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][5] ),
    .Q_N(_07213_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _17436_ (.CLK(net5168),
    .RESET_B(net191),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][6] ),
    .Q_N(_07214_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _17437_ (.CLK(net5168),
    .RESET_B(net192),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][7] ),
    .Q_N(_07215_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _17438_ (.CLK(net5168),
    .RESET_B(net193),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][8] ),
    .Q_N(_07216_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _17439_ (.CLK(net5171),
    .RESET_B(net194),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][9] ),
    .Q_N(_07217_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _17440_ (.CLK(net5171),
    .RESET_B(net195),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][10] ),
    .Q_N(_07218_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _17441_ (.CLK(net5165),
    .RESET_B(net196),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][11] ),
    .Q_N(_07219_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _17442_ (.CLK(net5165),
    .RESET_B(net197),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][12] ),
    .Q_N(_07220_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _17443_ (.CLK(net5161),
    .RESET_B(net198),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][13] ),
    .Q_N(_07221_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _17444_ (.CLK(net5160),
    .RESET_B(net199),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][14] ),
    .Q_N(_07222_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _17445_ (.CLK(net5157),
    .RESET_B(net200),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][15] ),
    .Q_N(_07223_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _17446_ (.CLK(net5157),
    .RESET_B(net201),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][16] ),
    .Q_N(_07224_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _17447_ (.CLK(net5157),
    .RESET_B(net202),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][17] ),
    .Q_N(_07225_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _17448_ (.CLK(net5164),
    .RESET_B(net203),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[0][18] ),
    .Q_N(_07226_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _17449_ (.CLK(net5158),
    .RESET_B(net204),
    .D(_01092_),
    .Q_N(_07227_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][0] ));
 sg13g2_dfrbp_1 _17450_ (.CLK(net5158),
    .RESET_B(net205),
    .D(_01102_),
    .Q_N(_07228_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][1] ));
 sg13g2_dfrbp_1 _17451_ (.CLK(net5160),
    .RESET_B(net206),
    .D(_01103_),
    .Q_N(_07229_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][2] ));
 sg13g2_dfrbp_1 _17452_ (.CLK(net5161),
    .RESET_B(net207),
    .D(_01104_),
    .Q_N(_07230_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][3] ));
 sg13g2_dfrbp_1 _17453_ (.CLK(net5165),
    .RESET_B(net208),
    .D(_01105_),
    .Q_N(_07231_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][4] ));
 sg13g2_dfrbp_1 _17454_ (.CLK(net5171),
    .RESET_B(net209),
    .D(_01106_),
    .Q_N(_07232_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][5] ));
 sg13g2_dfrbp_1 _17455_ (.CLK(net5169),
    .RESET_B(net210),
    .D(_01107_),
    .Q_N(_07233_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][6] ));
 sg13g2_dfrbp_1 _17456_ (.CLK(net5170),
    .RESET_B(net211),
    .D(_01108_),
    .Q_N(_07234_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][7] ));
 sg13g2_dfrbp_1 _17457_ (.CLK(net5170),
    .RESET_B(net212),
    .D(_01109_),
    .Q_N(_07235_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][8] ));
 sg13g2_dfrbp_1 _17458_ (.CLK(net5169),
    .RESET_B(net213),
    .D(_01110_),
    .Q_N(_07236_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][9] ));
 sg13g2_dfrbp_1 _17459_ (.CLK(net5165),
    .RESET_B(net214),
    .D(_01093_),
    .Q_N(_07237_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][10] ));
 sg13g2_dfrbp_1 _17460_ (.CLK(net5167),
    .RESET_B(net215),
    .D(_01094_),
    .Q_N(_07238_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][11] ));
 sg13g2_dfrbp_1 _17461_ (.CLK(net5167),
    .RESET_B(net216),
    .D(_01095_),
    .Q_N(_07239_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][12] ));
 sg13g2_dfrbp_1 _17462_ (.CLK(net5163),
    .RESET_B(net217),
    .D(_01096_),
    .Q_N(_07240_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][13] ));
 sg13g2_dfrbp_1 _17463_ (.CLK(net5163),
    .RESET_B(net218),
    .D(_01097_),
    .Q_N(_07241_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][14] ));
 sg13g2_dfrbp_1 _17464_ (.CLK(net5159),
    .RESET_B(net219),
    .D(_01098_),
    .Q_N(_07242_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][15] ));
 sg13g2_dfrbp_1 _17465_ (.CLK(net5158),
    .RESET_B(net220),
    .D(_01099_),
    .Q_N(_07243_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][16] ));
 sg13g2_dfrbp_1 _17466_ (.CLK(net5158),
    .RESET_B(net240),
    .D(_01100_),
    .Q_N(_07244_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][17] ));
 sg13g2_dfrbp_1 _17467_ (.CLK(net5158),
    .RESET_B(net633),
    .D(_01101_),
    .Q_N(_06592_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][18] ));
 sg13g2_dfrbp_1 _17468_ (.CLK(_01458_),
    .RESET_B(net632),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[0] ),
    .Q_N(_06591_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _17469_ (.CLK(_01459_),
    .RESET_B(net631),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[1] ),
    .Q_N(_06590_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _17470_ (.CLK(_01460_),
    .RESET_B(net630),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[2] ),
    .Q_N(_06589_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _17471_ (.CLK(_01461_),
    .RESET_B(net629),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[3] ),
    .Q_N(_06588_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _17472_ (.CLK(_01462_),
    .RESET_B(net628),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[4] ),
    .Q_N(_06587_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _17473_ (.CLK(_01463_),
    .RESET_B(net627),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[5] ),
    .Q_N(_06586_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _17474_ (.CLK(_01464_),
    .RESET_B(net626),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[6] ),
    .Q_N(_06585_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _17475_ (.CLK(_01465_),
    .RESET_B(net625),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[7] ),
    .Q_N(_06584_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _17476_ (.CLK(_01466_),
    .RESET_B(net624),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[8] ),
    .Q_N(_06583_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _17477_ (.CLK(_01467_),
    .RESET_B(net623),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[9] ),
    .Q_N(_06582_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _17478_ (.CLK(_01468_),
    .RESET_B(net622),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[10] ),
    .Q_N(_06581_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _17479_ (.CLK(_01469_),
    .RESET_B(net621),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[11] ),
    .Q_N(_06580_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _17480_ (.CLK(_01470_),
    .RESET_B(net620),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[12] ),
    .Q_N(_06579_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _17481_ (.CLK(_01471_),
    .RESET_B(net581),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[13] ),
    .Q_N(_06578_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _17482_ (.CLK(_01472_),
    .RESET_B(net580),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[14] ),
    .Q_N(_06577_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _17483_ (.CLK(_01473_),
    .RESET_B(net579),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[15] ),
    .Q_N(_06576_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _17484_ (.CLK(_01474_),
    .RESET_B(net578),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[16] ),
    .Q_N(_06575_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _17485_ (.CLK(_01475_),
    .RESET_B(net577),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[17] ),
    .Q_N(_06574_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _17486_ (.CLK(_01476_),
    .RESET_B(net241),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.temp_delay[18] ),
    .Q_N(_07245_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[1].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _17487_ (.CLK(net5151),
    .RESET_B(net242),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][0] ),
    .Q_N(_07246_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _17488_ (.CLK(net5157),
    .RESET_B(net243),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][1] ),
    .Q_N(_07247_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _17489_ (.CLK(net5160),
    .RESET_B(net244),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][2] ),
    .Q_N(_07248_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _17490_ (.CLK(net5160),
    .RESET_B(net245),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][3] ),
    .Q_N(_07249_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _17491_ (.CLK(net5165),
    .RESET_B(net246),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][4] ),
    .Q_N(_07250_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _17492_ (.CLK(net5171),
    .RESET_B(net247),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][5] ),
    .Q_N(_07251_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _17493_ (.CLK(net5169),
    .RESET_B(net248),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][6] ),
    .Q_N(_07252_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _17494_ (.CLK(net5169),
    .RESET_B(net249),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][7] ),
    .Q_N(_07253_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _17495_ (.CLK(net5169),
    .RESET_B(net250),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][8] ),
    .Q_N(_07254_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _17496_ (.CLK(net5172),
    .RESET_B(net251),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][9] ),
    .Q_N(_07255_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _17497_ (.CLK(net5167),
    .RESET_B(net252),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][10] ),
    .Q_N(_07256_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _17498_ (.CLK(net5166),
    .RESET_B(net253),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][11] ),
    .Q_N(_07257_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _17499_ (.CLK(net5166),
    .RESET_B(net254),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][12] ),
    .Q_N(_07258_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _17500_ (.CLK(net5162),
    .RESET_B(net255),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][13] ),
    .Q_N(_07259_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _17501_ (.CLK(net5162),
    .RESET_B(net256),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][14] ),
    .Q_N(_07260_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _17502_ (.CLK(net5159),
    .RESET_B(net257),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][15] ),
    .Q_N(_07261_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _17503_ (.CLK(net5152),
    .RESET_B(net258),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][16] ),
    .Q_N(_07262_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _17504_ (.CLK(net5152),
    .RESET_B(net259),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][17] ),
    .Q_N(_07263_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _17505_ (.CLK(net5151),
    .RESET_B(net260),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.comb_data[1][18] ),
    .Q_N(_07264_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _17506_ (.CLK(net5152),
    .RESET_B(net261),
    .D(_01111_),
    .Q_N(_07265_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17507_ (.CLK(net5152),
    .RESET_B(net262),
    .D(_01121_),
    .Q_N(_07266_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17508_ (.CLK(net5159),
    .RESET_B(net263),
    .D(_01122_),
    .Q_N(_07267_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17509_ (.CLK(net5162),
    .RESET_B(net264),
    .D(_01123_),
    .Q_N(_07268_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17510_ (.CLK(net5162),
    .RESET_B(net265),
    .D(_01124_),
    .Q_N(_07269_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17511_ (.CLK(net5166),
    .RESET_B(net266),
    .D(_01125_),
    .Q_N(_07270_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17512_ (.CLK(net5172),
    .RESET_B(net267),
    .D(_01126_),
    .Q_N(_07271_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17513_ (.CLK(net5172),
    .RESET_B(net268),
    .D(_01127_),
    .Q_N(_07272_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17514_ (.CLK(net5172),
    .RESET_B(net269),
    .D(_01128_),
    .Q_N(_07273_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17515_ (.CLK(net5172),
    .RESET_B(net270),
    .D(_01129_),
    .Q_N(_07274_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17516_ (.CLK(net5174),
    .RESET_B(net271),
    .D(_01112_),
    .Q_N(_07275_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17517_ (.CLK(net5174),
    .RESET_B(net272),
    .D(_01113_),
    .Q_N(_07276_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17518_ (.CLK(net5174),
    .RESET_B(net273),
    .D(_01114_),
    .Q_N(_07277_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17519_ (.CLK(net5174),
    .RESET_B(net274),
    .D(_01115_),
    .Q_N(_07278_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17520_ (.CLK(net5174),
    .RESET_B(net275),
    .D(_01116_),
    .Q_N(_07279_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17521_ (.CLK(net5174),
    .RESET_B(net276),
    .D(_01117_),
    .Q_N(_07280_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17522_ (.CLK(net5175),
    .RESET_B(net277),
    .D(_01118_),
    .Q_N(_07281_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17523_ (.CLK(net5152),
    .RESET_B(net297),
    .D(_01119_),
    .Q_N(_07282_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17524_ (.CLK(net5151),
    .RESET_B(net576),
    .D(_01120_),
    .Q_N(_06573_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17525_ (.CLK(_01477_),
    .RESET_B(net575),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[0] ),
    .Q_N(_06572_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _17526_ (.CLK(_01478_),
    .RESET_B(net574),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[1] ),
    .Q_N(_06571_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _17527_ (.CLK(_01479_),
    .RESET_B(net573),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[2] ),
    .Q_N(_06570_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _17528_ (.CLK(_01480_),
    .RESET_B(net572),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[3] ),
    .Q_N(_06569_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _17529_ (.CLK(_01481_),
    .RESET_B(net571),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[4] ),
    .Q_N(_06568_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _17530_ (.CLK(_01482_),
    .RESET_B(net570),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[5] ),
    .Q_N(_06567_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _17531_ (.CLK(_01483_),
    .RESET_B(net569),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[6] ),
    .Q_N(_06566_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _17532_ (.CLK(_01484_),
    .RESET_B(net568),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[7] ),
    .Q_N(_06565_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _17533_ (.CLK(_01485_),
    .RESET_B(net567),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[8] ),
    .Q_N(_06564_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _17534_ (.CLK(_01486_),
    .RESET_B(net566),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[9] ),
    .Q_N(_06563_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _17535_ (.CLK(_01487_),
    .RESET_B(net565),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[10] ),
    .Q_N(_06562_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _17536_ (.CLK(_01488_),
    .RESET_B(net564),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[11] ),
    .Q_N(_06561_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _17537_ (.CLK(_01489_),
    .RESET_B(net563),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[12] ),
    .Q_N(_06560_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _17538_ (.CLK(_01490_),
    .RESET_B(net524),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[13] ),
    .Q_N(_06559_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _17539_ (.CLK(_01491_),
    .RESET_B(net523),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[14] ),
    .Q_N(_06558_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _17540_ (.CLK(_01492_),
    .RESET_B(net522),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[15] ),
    .Q_N(_06557_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _17541_ (.CLK(_01493_),
    .RESET_B(net521),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[16] ),
    .Q_N(_06556_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _17542_ (.CLK(_01494_),
    .RESET_B(net520),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[17] ),
    .Q_N(_06555_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _17543_ (.CLK(_01495_),
    .RESET_B(net298),
    .D(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.temp_delay[18] ),
    .Q_N(_07283_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.genblk1[2].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _17544_ (.CLK(net5418),
    .RESET_B(net5927),
    .D(_01073_),
    .Q_N(_07284_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_dfrbp_1 _17545_ (.CLK(net5418),
    .RESET_B(net5927),
    .D(_01083_),
    .Q_N(_07285_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_dfrbp_1 _17546_ (.CLK(net5421),
    .RESET_B(net5930),
    .D(_01084_),
    .Q_N(_07286_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_dfrbp_1 _17547_ (.CLK(net5419),
    .RESET_B(net5928),
    .D(_01085_),
    .Q_N(_07287_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_dfrbp_1 _17548_ (.CLK(net5420),
    .RESET_B(net5929),
    .D(_01086_),
    .Q_N(_07288_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_dfrbp_1 _17549_ (.CLK(net5420),
    .RESET_B(net5929),
    .D(_01087_),
    .Q_N(_07289_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_dfrbp_1 _17550_ (.CLK(net5419),
    .RESET_B(net5928),
    .D(_01088_),
    .Q_N(_07290_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_dfrbp_1 _17551_ (.CLK(net5416),
    .RESET_B(net5925),
    .D(_01089_),
    .Q_N(_07291_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_dfrbp_1 _17552_ (.CLK(net5422),
    .RESET_B(net5927),
    .D(_01090_),
    .Q_N(_07292_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_dfrbp_1 _17553_ (.CLK(net5377),
    .RESET_B(net5886),
    .D(_01091_),
    .Q_N(_07293_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_dfrbp_1 _17554_ (.CLK(net5377),
    .RESET_B(net5886),
    .D(_01074_),
    .Q_N(_07294_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_dfrbp_1 _17555_ (.CLK(net5376),
    .RESET_B(net5885),
    .D(_01075_),
    .Q_N(_07295_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_dfrbp_1 _17556_ (.CLK(net5376),
    .RESET_B(net5885),
    .D(_01076_),
    .Q_N(_07296_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_dfrbp_1 _17557_ (.CLK(net5376),
    .RESET_B(net5885),
    .D(_01077_),
    .Q_N(_07297_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_dfrbp_1 _17558_ (.CLK(net5373),
    .RESET_B(net5882),
    .D(_01078_),
    .Q_N(_07298_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_dfrbp_1 _17559_ (.CLK(net5371),
    .RESET_B(net5880),
    .D(_01079_),
    .Q_N(_07299_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_dfrbp_1 _17560_ (.CLK(net5369),
    .RESET_B(net5878),
    .D(_01080_),
    .Q_N(_07300_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_dfrbp_1 _17561_ (.CLK(net5370),
    .RESET_B(net5879),
    .D(_01081_),
    .Q_N(_07301_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_dfrbp_1 _17562_ (.CLK(net5369),
    .RESET_B(net5878),
    .D(_01082_),
    .Q_N(_07302_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u3.reg_value[18] ));
 sg13g2_dfrbp_1 _17563_ (.CLK(net5425),
    .RESET_B(net5934),
    .D(_01073_),
    .Q_N(_07303_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][0] ));
 sg13g2_dfrbp_1 _17564_ (.CLK(net5418),
    .RESET_B(net5927),
    .D(_01083_),
    .Q_N(_07304_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][1] ));
 sg13g2_dfrbp_1 _17565_ (.CLK(net5421),
    .RESET_B(net5930),
    .D(_01084_),
    .Q_N(_07305_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][2] ));
 sg13g2_dfrbp_1 _17566_ (.CLK(net5421),
    .RESET_B(net5930),
    .D(_01085_),
    .Q_N(_07306_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][3] ));
 sg13g2_dfrbp_1 _17567_ (.CLK(net5420),
    .RESET_B(net5928),
    .D(_01086_),
    .Q_N(_07307_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][4] ));
 sg13g2_dfrbp_1 _17568_ (.CLK(net5419),
    .RESET_B(net5929),
    .D(_01087_),
    .Q_N(_07308_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][5] ));
 sg13g2_dfrbp_1 _17569_ (.CLK(net5420),
    .RESET_B(net5929),
    .D(_01088_),
    .Q_N(_07309_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][6] ));
 sg13g2_dfrbp_1 _17570_ (.CLK(net5421),
    .RESET_B(net5930),
    .D(_01089_),
    .Q_N(_07310_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][7] ));
 sg13g2_dfrbp_1 _17571_ (.CLK(net5418),
    .RESET_B(net5927),
    .D(_01090_),
    .Q_N(_07311_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][8] ));
 sg13g2_dfrbp_1 _17572_ (.CLK(net5376),
    .RESET_B(net5885),
    .D(_01091_),
    .Q_N(_07312_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][9] ));
 sg13g2_dfrbp_1 _17573_ (.CLK(net5377),
    .RESET_B(net5886),
    .D(_01074_),
    .Q_N(_07313_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][10] ));
 sg13g2_dfrbp_1 _17574_ (.CLK(net5377),
    .RESET_B(net5886),
    .D(_01075_),
    .Q_N(_07314_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][11] ));
 sg13g2_dfrbp_1 _17575_ (.CLK(net5376),
    .RESET_B(net5885),
    .D(_01076_),
    .Q_N(_07315_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][12] ));
 sg13g2_dfrbp_1 _17576_ (.CLK(net5376),
    .RESET_B(net5885),
    .D(_01077_),
    .Q_N(_07316_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][13] ));
 sg13g2_dfrbp_1 _17577_ (.CLK(net5373),
    .RESET_B(net5882),
    .D(_01078_),
    .Q_N(_07317_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][14] ));
 sg13g2_dfrbp_1 _17578_ (.CLK(net5373),
    .RESET_B(net5882),
    .D(_01079_),
    .Q_N(_07318_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][15] ));
 sg13g2_dfrbp_1 _17579_ (.CLK(net5373),
    .RESET_B(net5882),
    .D(_01080_),
    .Q_N(_07319_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][16] ));
 sg13g2_dfrbp_1 _17580_ (.CLK(net5373),
    .RESET_B(net5882),
    .D(_01081_),
    .Q_N(_07320_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][17] ));
 sg13g2_dfrbp_1 _17581_ (.CLK(net5370),
    .RESET_B(net5879),
    .D(_01082_),
    .Q_N(_07321_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][18] ));
 sg13g2_dfrbp_1 _17582_ (.CLK(net5417),
    .RESET_B(net5926),
    .D(_01054_),
    .Q_N(_07322_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_dfrbp_1 _17583_ (.CLK(net5416),
    .RESET_B(net5925),
    .D(_01064_),
    .Q_N(_07323_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_dfrbp_1 _17584_ (.CLK(net5416),
    .RESET_B(net5925),
    .D(_01065_),
    .Q_N(_07324_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_dfrbp_1 _17585_ (.CLK(net5416),
    .RESET_B(net5925),
    .D(_01066_),
    .Q_N(_07325_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_dfrbp_1 _17586_ (.CLK(net5419),
    .RESET_B(net5928),
    .D(_01067_),
    .Q_N(_07326_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_dfrbp_1 _17587_ (.CLK(net5415),
    .RESET_B(net5924),
    .D(_01068_),
    .Q_N(_07327_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_dfrbp_1 _17588_ (.CLK(net5415),
    .RESET_B(net5924),
    .D(_01069_),
    .Q_N(_07328_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_dfrbp_1 _17589_ (.CLK(net5417),
    .RESET_B(net5926),
    .D(_01070_),
    .Q_N(_07329_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_dfrbp_1 _17590_ (.CLK(net5375),
    .RESET_B(net5884),
    .D(_01071_),
    .Q_N(_07330_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_dfrbp_1 _17591_ (.CLK(net5375),
    .RESET_B(net5884),
    .D(_01072_),
    .Q_N(_07331_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_dfrbp_1 _17592_ (.CLK(net5374),
    .RESET_B(net5883),
    .D(_01055_),
    .Q_N(_07332_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_dfrbp_1 _17593_ (.CLK(net5374),
    .RESET_B(net5883),
    .D(_01056_),
    .Q_N(_07333_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_dfrbp_1 _17594_ (.CLK(net5375),
    .RESET_B(net5884),
    .D(_01057_),
    .Q_N(_07334_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_dfrbp_1 _17595_ (.CLK(net5371),
    .RESET_B(net5880),
    .D(_01058_),
    .Q_N(_07335_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_dfrbp_1 _17596_ (.CLK(net5371),
    .RESET_B(net5880),
    .D(_01059_),
    .Q_N(_07336_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_dfrbp_1 _17597_ (.CLK(net5371),
    .RESET_B(net5880),
    .D(_01060_),
    .Q_N(_07337_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_dfrbp_1 _17598_ (.CLK(net5369),
    .RESET_B(net5878),
    .D(_01061_),
    .Q_N(_07338_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[16] ));
 sg13g2_dfrbp_1 _17599_ (.CLK(net5369),
    .RESET_B(net5878),
    .D(_01062_),
    .Q_N(_07339_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_dfrbp_1 _17600_ (.CLK(net5352),
    .RESET_B(net5860),
    .D(_01063_),
    .Q_N(_07340_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.u2.reg_value[18] ));
 sg13g2_dfrbp_1 _17601_ (.CLK(net5418),
    .RESET_B(net5927),
    .D(_01054_),
    .Q_N(_07341_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_dfrbp_1 _17602_ (.CLK(net5418),
    .RESET_B(net5931),
    .D(_01064_),
    .Q_N(_07342_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_dfrbp_1 _17603_ (.CLK(net5416),
    .RESET_B(net5925),
    .D(_01065_),
    .Q_N(_07343_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_dfrbp_1 _17604_ (.CLK(net5419),
    .RESET_B(net5928),
    .D(_01066_),
    .Q_N(_07344_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_dfrbp_1 _17605_ (.CLK(net5419),
    .RESET_B(net5928),
    .D(_01067_),
    .Q_N(_07345_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_dfrbp_1 _17606_ (.CLK(net5419),
    .RESET_B(net5928),
    .D(_01068_),
    .Q_N(_07346_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_dfrbp_1 _17607_ (.CLK(net5415),
    .RESET_B(net5924),
    .D(_01069_),
    .Q_N(_07347_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_dfrbp_1 _17608_ (.CLK(net5415),
    .RESET_B(net5924),
    .D(_01070_),
    .Q_N(_07348_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_dfrbp_1 _17609_ (.CLK(net5417),
    .RESET_B(net5926),
    .D(_01071_),
    .Q_N(_07349_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_dfrbp_1 _17610_ (.CLK(net5375),
    .RESET_B(net5884),
    .D(_01072_),
    .Q_N(_07350_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_dfrbp_1 _17611_ (.CLK(net5375),
    .RESET_B(net5884),
    .D(_01055_),
    .Q_N(_07351_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_dfrbp_1 _17612_ (.CLK(net5374),
    .RESET_B(net5883),
    .D(_01056_),
    .Q_N(_07352_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_dfrbp_1 _17613_ (.CLK(net5374),
    .RESET_B(net5883),
    .D(_01057_),
    .Q_N(_07353_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_dfrbp_1 _17614_ (.CLK(net5374),
    .RESET_B(net5883),
    .D(_01058_),
    .Q_N(_07354_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_dfrbp_1 _17615_ (.CLK(net5371),
    .RESET_B(net5880),
    .D(_01059_),
    .Q_N(_07355_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_dfrbp_1 _17616_ (.CLK(net5372),
    .RESET_B(net5881),
    .D(_01060_),
    .Q_N(_07356_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_dfrbp_1 _17617_ (.CLK(net5370),
    .RESET_B(net5879),
    .D(_01061_),
    .Q_N(_07357_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_dfrbp_1 _17618_ (.CLK(net5370),
    .RESET_B(net5879),
    .D(_01062_),
    .Q_N(_07358_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_dfrbp_1 _17619_ (.CLK(net5353),
    .RESET_B(net5861),
    .D(_01063_),
    .Q_N(_07359_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator2_out[18] ));
 sg13g2_dfrbp_1 _17620_ (.CLK(net5417),
    .RESET_B(net5926),
    .D(_01187_),
    .Q_N(_01187_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[0] ));
 sg13g2_dfrbp_1 _17621_ (.CLK(net5417),
    .RESET_B(net5926),
    .D(_01045_),
    .Q_N(_07360_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_dfrbp_1 _17622_ (.CLK(net5415),
    .RESET_B(net5924),
    .D(_01046_),
    .Q_N(_07361_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_dfrbp_1 _17623_ (.CLK(net5415),
    .RESET_B(net5924),
    .D(_01047_),
    .Q_N(_07362_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_dfrbp_1 _17624_ (.CLK(net5415),
    .RESET_B(net5924),
    .D(_01048_),
    .Q_N(_07363_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[4] ));
 sg13g2_dfrbp_1 _17625_ (.CLK(net5415),
    .RESET_B(net5924),
    .D(_01049_),
    .Q_N(_07364_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_dfrbp_1 _17626_ (.CLK(net5417),
    .RESET_B(net5926),
    .D(_01050_),
    .Q_N(_07365_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_dfrbp_1 _17627_ (.CLK(net5417),
    .RESET_B(net5926),
    .D(_01051_),
    .Q_N(_07366_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_dfrbp_1 _17628_ (.CLK(net5375),
    .RESET_B(net5884),
    .D(_01052_),
    .Q_N(_07367_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_dfrbp_1 _17629_ (.CLK(net5375),
    .RESET_B(net5884),
    .D(_01053_),
    .Q_N(_07368_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_dfrbp_1 _17630_ (.CLK(net5374),
    .RESET_B(net5883),
    .D(_01036_),
    .Q_N(_07369_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_dfrbp_1 _17631_ (.CLK(net5374),
    .RESET_B(net5883),
    .D(_01037_),
    .Q_N(_07370_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_dfrbp_1 _17632_ (.CLK(net5374),
    .RESET_B(net5883),
    .D(_01038_),
    .Q_N(_07371_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_dfrbp_1 _17633_ (.CLK(net5371),
    .RESET_B(net5880),
    .D(_01039_),
    .Q_N(_07372_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_dfrbp_1 _17634_ (.CLK(net5371),
    .RESET_B(net5880),
    .D(_01040_),
    .Q_N(_07373_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_dfrbp_1 _17635_ (.CLK(net5371),
    .RESET_B(net5880),
    .D(_01041_),
    .Q_N(_07374_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_dfrbp_1 _17636_ (.CLK(net5369),
    .RESET_B(net5878),
    .D(_01042_),
    .Q_N(_07375_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_dfrbp_1 _17637_ (.CLK(net5369),
    .RESET_B(net5878),
    .D(_01043_),
    .Q_N(_07376_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_dfrbp_1 _17638_ (.CLK(net5352),
    .RESET_B(net5860),
    .D(_01044_),
    .Q_N(_07377_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.u_top_module.integrator1_out[18] ));
 sg13g2_dfrbp_1 _17639_ (.CLK(net5106),
    .RESET_B(net299),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][0] ),
    .Q_N(_07378_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _17640_ (.CLK(net5106),
    .RESET_B(net300),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][1] ),
    .Q_N(_07379_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _17641_ (.CLK(net5105),
    .RESET_B(net301),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][2] ),
    .Q_N(_07380_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _17642_ (.CLK(net5105),
    .RESET_B(net302),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][3] ),
    .Q_N(_07381_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _17643_ (.CLK(net5117),
    .RESET_B(net303),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][4] ),
    .Q_N(_07382_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _17644_ (.CLK(net5117),
    .RESET_B(net304),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][5] ),
    .Q_N(_07383_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _17645_ (.CLK(net5105),
    .RESET_B(net305),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][6] ),
    .Q_N(_07384_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _17646_ (.CLK(net5105),
    .RESET_B(net306),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][7] ),
    .Q_N(_07385_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _17647_ (.CLK(net5105),
    .RESET_B(net307),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][8] ),
    .Q_N(_07386_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _17648_ (.CLK(net5086),
    .RESET_B(net308),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][9] ),
    .Q_N(_07387_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _17649_ (.CLK(net5089),
    .RESET_B(net309),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][10] ),
    .Q_N(_07388_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _17650_ (.CLK(net5087),
    .RESET_B(net310),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][11] ),
    .Q_N(_07389_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _17651_ (.CLK(net5086),
    .RESET_B(net311),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][12] ),
    .Q_N(_07390_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _17652_ (.CLK(net5086),
    .RESET_B(net312),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][13] ),
    .Q_N(_07391_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _17653_ (.CLK(net5086),
    .RESET_B(net313),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][14] ),
    .Q_N(_07392_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _17654_ (.CLK(net5085),
    .RESET_B(net314),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][15] ),
    .Q_N(_07393_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _17655_ (.CLK(net5084),
    .RESET_B(net315),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][16] ),
    .Q_N(_07394_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _17656_ (.CLK(net5084),
    .RESET_B(net316),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][17] ),
    .Q_N(_07395_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _17657_ (.CLK(net5084),
    .RESET_B(net317),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[0][18] ),
    .Q_N(_07396_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _17658_ (.CLK(net5109),
    .RESET_B(net318),
    .D(_00998_),
    .Q_N(_07397_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][0] ));
 sg13g2_dfrbp_1 _17659_ (.CLK(net5109),
    .RESET_B(net319),
    .D(_01008_),
    .Q_N(_07398_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][1] ));
 sg13g2_dfrbp_1 _17660_ (.CLK(net5108),
    .RESET_B(net320),
    .D(_01009_),
    .Q_N(_07399_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][2] ));
 sg13g2_dfrbp_1 _17661_ (.CLK(net5112),
    .RESET_B(net321),
    .D(_01010_),
    .Q_N(_07400_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][3] ));
 sg13g2_dfrbp_1 _17662_ (.CLK(net5117),
    .RESET_B(net322),
    .D(_01011_),
    .Q_N(_07401_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][4] ));
 sg13g2_dfrbp_1 _17663_ (.CLK(net5117),
    .RESET_B(net323),
    .D(_01012_),
    .Q_N(_07402_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][5] ));
 sg13g2_dfrbp_1 _17664_ (.CLK(net5117),
    .RESET_B(net324),
    .D(_01013_),
    .Q_N(_07403_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][6] ));
 sg13g2_dfrbp_1 _17665_ (.CLK(net5108),
    .RESET_B(net325),
    .D(_01014_),
    .Q_N(_07404_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][7] ));
 sg13g2_dfrbp_1 _17666_ (.CLK(net5107),
    .RESET_B(net326),
    .D(_01015_),
    .Q_N(_07405_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][8] ));
 sg13g2_dfrbp_1 _17667_ (.CLK(net5106),
    .RESET_B(net327),
    .D(_01016_),
    .Q_N(_07406_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][9] ));
 sg13g2_dfrbp_1 _17668_ (.CLK(net5089),
    .RESET_B(net328),
    .D(_00999_),
    .Q_N(_07407_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][10] ));
 sg13g2_dfrbp_1 _17669_ (.CLK(net5089),
    .RESET_B(net329),
    .D(_01000_),
    .Q_N(_07408_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][11] ));
 sg13g2_dfrbp_1 _17670_ (.CLK(net5089),
    .RESET_B(net330),
    .D(_01001_),
    .Q_N(_07409_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][12] ));
 sg13g2_dfrbp_1 _17671_ (.CLK(net5089),
    .RESET_B(net331),
    .D(_01002_),
    .Q_N(_07410_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][13] ));
 sg13g2_dfrbp_1 _17672_ (.CLK(net5088),
    .RESET_B(net332),
    .D(_01003_),
    .Q_N(_07411_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][14] ));
 sg13g2_dfrbp_1 _17673_ (.CLK(net5088),
    .RESET_B(net333),
    .D(_01004_),
    .Q_N(_07412_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][15] ));
 sg13g2_dfrbp_1 _17674_ (.CLK(net5085),
    .RESET_B(net334),
    .D(_01005_),
    .Q_N(_07413_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][16] ));
 sg13g2_dfrbp_1 _17675_ (.CLK(net5085),
    .RESET_B(net354),
    .D(_01006_),
    .Q_N(_07414_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][17] ));
 sg13g2_dfrbp_1 _17676_ (.CLK(net5084),
    .RESET_B(net519),
    .D(_01007_),
    .Q_N(_06554_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][18] ));
 sg13g2_dfrbp_1 _17677_ (.CLK(_01496_),
    .RESET_B(net518),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[0] ),
    .Q_N(_06553_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _17678_ (.CLK(_01497_),
    .RESET_B(net517),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[1] ),
    .Q_N(_06552_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _17679_ (.CLK(_01498_),
    .RESET_B(net516),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[2] ),
    .Q_N(_06551_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _17680_ (.CLK(_01499_),
    .RESET_B(net515),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[3] ),
    .Q_N(_06550_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _17681_ (.CLK(_01500_),
    .RESET_B(net514),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[4] ),
    .Q_N(_06549_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _17682_ (.CLK(_01501_),
    .RESET_B(net513),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[5] ),
    .Q_N(_06548_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _17683_ (.CLK(_01502_),
    .RESET_B(net512),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[6] ),
    .Q_N(_06547_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _17684_ (.CLK(_01503_),
    .RESET_B(net511),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[7] ),
    .Q_N(_06546_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _17685_ (.CLK(_01504_),
    .RESET_B(net510),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[8] ),
    .Q_N(_06545_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _17686_ (.CLK(_01505_),
    .RESET_B(net509),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[9] ),
    .Q_N(_06544_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _17687_ (.CLK(_01506_),
    .RESET_B(net508),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[10] ),
    .Q_N(_06543_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _17688_ (.CLK(_01507_),
    .RESET_B(net507),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[11] ),
    .Q_N(_06542_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _17689_ (.CLK(_01508_),
    .RESET_B(net506),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[12] ),
    .Q_N(_06541_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _17690_ (.CLK(_01509_),
    .RESET_B(net467),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[13] ),
    .Q_N(_06540_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _17691_ (.CLK(_01510_),
    .RESET_B(net466),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[14] ),
    .Q_N(_06539_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _17692_ (.CLK(_01511_),
    .RESET_B(net465),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[15] ),
    .Q_N(_06538_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _17693_ (.CLK(_01512_),
    .RESET_B(net464),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[16] ),
    .Q_N(_06537_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _17694_ (.CLK(_01513_),
    .RESET_B(net463),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[17] ),
    .Q_N(_06536_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _17695_ (.CLK(_01514_),
    .RESET_B(net355),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.temp_delay[18] ),
    .Q_N(_07415_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[1].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _17696_ (.CLK(net5109),
    .RESET_B(net356),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][0] ),
    .Q_N(_07416_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _17697_ (.CLK(net5110),
    .RESET_B(net357),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][1] ),
    .Q_N(_07417_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _17698_ (.CLK(net5114),
    .RESET_B(net358),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][2] ),
    .Q_N(_07418_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _17699_ (.CLK(net5113),
    .RESET_B(net359),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][3] ),
    .Q_N(_07419_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _17700_ (.CLK(net5115),
    .RESET_B(net360),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][4] ),
    .Q_N(_07420_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _17701_ (.CLK(net5115),
    .RESET_B(net361),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][5] ),
    .Q_N(_07421_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _17702_ (.CLK(net5113),
    .RESET_B(net362),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][6] ),
    .Q_N(_07422_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _17703_ (.CLK(net5112),
    .RESET_B(net363),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][7] ),
    .Q_N(_07423_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _17704_ (.CLK(net5107),
    .RESET_B(net364),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][8] ),
    .Q_N(_07424_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _17705_ (.CLK(net5106),
    .RESET_B(net365),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][9] ),
    .Q_N(_07425_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _17706_ (.CLK(net5090),
    .RESET_B(net366),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][10] ),
    .Q_N(_07426_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _17707_ (.CLK(net5091),
    .RESET_B(net367),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][11] ),
    .Q_N(_07427_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _17708_ (.CLK(net5090),
    .RESET_B(net368),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][12] ),
    .Q_N(_07428_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _17709_ (.CLK(net5090),
    .RESET_B(net369),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][13] ),
    .Q_N(_07429_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _17710_ (.CLK(net5089),
    .RESET_B(net370),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][14] ),
    .Q_N(_07430_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _17711_ (.CLK(net5088),
    .RESET_B(net371),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][15] ),
    .Q_N(_07431_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _17712_ (.CLK(net5088),
    .RESET_B(net372),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][16] ),
    .Q_N(_07432_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _17713_ (.CLK(net5092),
    .RESET_B(net373),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][17] ),
    .Q_N(_07433_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _17714_ (.CLK(net5084),
    .RESET_B(net374),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.comb_data[1][18] ),
    .Q_N(_07434_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _17715_ (.CLK(net5119),
    .RESET_B(net375),
    .D(_01017_),
    .Q_N(_07435_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17716_ (.CLK(net5126),
    .RESET_B(net376),
    .D(_01027_),
    .Q_N(_07436_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17717_ (.CLK(net5126),
    .RESET_B(net377),
    .D(_01028_),
    .Q_N(_07437_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17718_ (.CLK(net5116),
    .RESET_B(net378),
    .D(_01029_),
    .Q_N(_07438_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17719_ (.CLK(net5131),
    .RESET_B(net379),
    .D(_01030_),
    .Q_N(_07439_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17720_ (.CLK(net5131),
    .RESET_B(net380),
    .D(_01031_),
    .Q_N(_07440_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17721_ (.CLK(net5131),
    .RESET_B(net381),
    .D(_01032_),
    .Q_N(_07441_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17722_ (.CLK(net5116),
    .RESET_B(net382),
    .D(_01033_),
    .Q_N(_07442_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17723_ (.CLK(net5114),
    .RESET_B(net383),
    .D(_01034_),
    .Q_N(_07443_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17724_ (.CLK(net5109),
    .RESET_B(net384),
    .D(_01035_),
    .Q_N(_07444_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17725_ (.CLK(net5119),
    .RESET_B(net385),
    .D(_01018_),
    .Q_N(_07445_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17726_ (.CLK(net5119),
    .RESET_B(net386),
    .D(_01019_),
    .Q_N(_07446_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17727_ (.CLK(net5102),
    .RESET_B(net387),
    .D(_01020_),
    .Q_N(_07447_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17728_ (.CLK(net5102),
    .RESET_B(net388),
    .D(_01021_),
    .Q_N(_07448_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17729_ (.CLK(net5102),
    .RESET_B(net389),
    .D(_01022_),
    .Q_N(_07449_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17730_ (.CLK(net5090),
    .RESET_B(net390),
    .D(_01023_),
    .Q_N(_07450_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17731_ (.CLK(net5090),
    .RESET_B(net391),
    .D(_01024_),
    .Q_N(_07451_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17732_ (.CLK(net5088),
    .RESET_B(net411),
    .D(_01025_),
    .Q_N(_07452_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17733_ (.CLK(net5084),
    .RESET_B(net462),
    .D(_01026_),
    .Q_N(_06535_),
    .Q(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17734_ (.CLK(_01515_),
    .RESET_B(net461),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[0] ),
    .Q_N(_06534_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _17735_ (.CLK(_01516_),
    .RESET_B(net460),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[1] ),
    .Q_N(_06533_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _17736_ (.CLK(_01517_),
    .RESET_B(net459),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[2] ),
    .Q_N(_06532_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _17737_ (.CLK(_01518_),
    .RESET_B(net458),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[3] ),
    .Q_N(_06531_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _17738_ (.CLK(_01519_),
    .RESET_B(net457),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[4] ),
    .Q_N(_06530_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _17739_ (.CLK(_01520_),
    .RESET_B(net456),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[5] ),
    .Q_N(_06529_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _17740_ (.CLK(_01521_),
    .RESET_B(net455),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[6] ),
    .Q_N(_06528_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _17741_ (.CLK(_01522_),
    .RESET_B(net454),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[7] ),
    .Q_N(_06527_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _17742_ (.CLK(_01523_),
    .RESET_B(net453),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[8] ),
    .Q_N(_06526_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _17743_ (.CLK(_01524_),
    .RESET_B(net452),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[9] ),
    .Q_N(_06525_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _17744_ (.CLK(_01525_),
    .RESET_B(net451),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[10] ),
    .Q_N(_06524_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _17745_ (.CLK(_01526_),
    .RESET_B(net450),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[11] ),
    .Q_N(_06523_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _17746_ (.CLK(_01527_),
    .RESET_B(net449),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[12] ),
    .Q_N(_06522_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _17747_ (.CLK(_01528_),
    .RESET_B(net410),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[13] ),
    .Q_N(_06521_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _17748_ (.CLK(_01529_),
    .RESET_B(net409),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[14] ),
    .Q_N(_06520_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _17749_ (.CLK(_01530_),
    .RESET_B(net408),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[15] ),
    .Q_N(_06519_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _17750_ (.CLK(_01531_),
    .RESET_B(net407),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[16] ),
    .Q_N(_06518_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _17751_ (.CLK(_01532_),
    .RESET_B(net406),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[17] ),
    .Q_N(_06517_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _17752_ (.CLK(_01533_),
    .RESET_B(net412),
    .D(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.temp_delay[18] ),
    .Q_N(_07453_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.genblk1[2].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _17753_ (.CLK(net5395),
    .RESET_B(net5904),
    .D(_00979_),
    .Q_N(_07454_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_dfrbp_1 _17754_ (.CLK(net5395),
    .RESET_B(net5904),
    .D(_00989_),
    .Q_N(_07455_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_dfrbp_1 _17755_ (.CLK(net5395),
    .RESET_B(net5904),
    .D(_00990_),
    .Q_N(_07456_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_dfrbp_1 _17756_ (.CLK(net5395),
    .RESET_B(net5904),
    .D(_00991_),
    .Q_N(_07457_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_dfrbp_1 _17757_ (.CLK(net5395),
    .RESET_B(net5904),
    .D(_00992_),
    .Q_N(_07458_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_dfrbp_1 _17758_ (.CLK(net5395),
    .RESET_B(net5904),
    .D(_00993_),
    .Q_N(_07459_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_dfrbp_1 _17759_ (.CLK(net5336),
    .RESET_B(net5846),
    .D(_00994_),
    .Q_N(_07460_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_dfrbp_1 _17760_ (.CLK(net5335),
    .RESET_B(net5845),
    .D(_00995_),
    .Q_N(_07461_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_dfrbp_1 _17761_ (.CLK(net5333),
    .RESET_B(net5843),
    .D(_00996_),
    .Q_N(_07462_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_dfrbp_1 _17762_ (.CLK(net5334),
    .RESET_B(net5844),
    .D(_00997_),
    .Q_N(_07463_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_dfrbp_1 _17763_ (.CLK(net5321),
    .RESET_B(net5831),
    .D(_00980_),
    .Q_N(_07464_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_dfrbp_1 _17764_ (.CLK(net5322),
    .RESET_B(net5832),
    .D(_00981_),
    .Q_N(_07465_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_dfrbp_1 _17765_ (.CLK(net5322),
    .RESET_B(net5832),
    .D(_00982_),
    .Q_N(_07466_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_dfrbp_1 _17766_ (.CLK(net5322),
    .RESET_B(net5832),
    .D(_00983_),
    .Q_N(_07467_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_dfrbp_1 _17767_ (.CLK(net5319),
    .RESET_B(net5829),
    .D(_00984_),
    .Q_N(_07468_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_dfrbp_1 _17768_ (.CLK(net5319),
    .RESET_B(net5829),
    .D(_00985_),
    .Q_N(_07469_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_dfrbp_1 _17769_ (.CLK(net5275),
    .RESET_B(net5785),
    .D(_00986_),
    .Q_N(_07470_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_dfrbp_1 _17770_ (.CLK(net5275),
    .RESET_B(net5785),
    .D(_00987_),
    .Q_N(_07471_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_dfrbp_1 _17771_ (.CLK(net5275),
    .RESET_B(net5785),
    .D(_00988_),
    .Q_N(_07472_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u3.reg_value[18] ));
 sg13g2_dfrbp_1 _17772_ (.CLK(net5396),
    .RESET_B(net5905),
    .D(_00979_),
    .Q_N(_07473_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][0] ));
 sg13g2_dfrbp_1 _17773_ (.CLK(net5395),
    .RESET_B(net5904),
    .D(_00989_),
    .Q_N(_07474_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][1] ));
 sg13g2_dfrbp_1 _17774_ (.CLK(net5396),
    .RESET_B(net5905),
    .D(_00990_),
    .Q_N(_07475_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][2] ));
 sg13g2_dfrbp_1 _17775_ (.CLK(net5396),
    .RESET_B(net5905),
    .D(_00991_),
    .Q_N(_07476_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][3] ));
 sg13g2_dfrbp_1 _17776_ (.CLK(net5396),
    .RESET_B(net5905),
    .D(_00992_),
    .Q_N(_07477_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][4] ));
 sg13g2_dfrbp_1 _17777_ (.CLK(net5396),
    .RESET_B(net5905),
    .D(_00993_),
    .Q_N(_07478_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][5] ));
 sg13g2_dfrbp_1 _17778_ (.CLK(net5395),
    .RESET_B(net5904),
    .D(_00994_),
    .Q_N(_07479_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][6] ));
 sg13g2_dfrbp_1 _17779_ (.CLK(net5336),
    .RESET_B(net5846),
    .D(_00995_),
    .Q_N(_07480_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][7] ));
 sg13g2_dfrbp_1 _17780_ (.CLK(net5335),
    .RESET_B(net5845),
    .D(_00996_),
    .Q_N(_07481_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][8] ));
 sg13g2_dfrbp_1 _17781_ (.CLK(net5333),
    .RESET_B(net5843),
    .D(_00997_),
    .Q_N(_07482_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][9] ));
 sg13g2_dfrbp_1 _17782_ (.CLK(net5338),
    .RESET_B(net5848),
    .D(_00980_),
    .Q_N(_07483_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][10] ));
 sg13g2_dfrbp_1 _17783_ (.CLK(net5322),
    .RESET_B(net5832),
    .D(_00981_),
    .Q_N(_07484_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][11] ));
 sg13g2_dfrbp_1 _17784_ (.CLK(net5322),
    .RESET_B(net5832),
    .D(_00982_),
    .Q_N(_07485_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][12] ));
 sg13g2_dfrbp_1 _17785_ (.CLK(net5322),
    .RESET_B(net5832),
    .D(_00983_),
    .Q_N(_07486_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][13] ));
 sg13g2_dfrbp_1 _17786_ (.CLK(net5319),
    .RESET_B(net5829),
    .D(_00984_),
    .Q_N(_07487_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][14] ));
 sg13g2_dfrbp_1 _17787_ (.CLK(net5319),
    .RESET_B(net5829),
    .D(_00985_),
    .Q_N(_07488_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][15] ));
 sg13g2_dfrbp_1 _17788_ (.CLK(net5319),
    .RESET_B(net5829),
    .D(_00986_),
    .Q_N(_07489_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][16] ));
 sg13g2_dfrbp_1 _17789_ (.CLK(net5275),
    .RESET_B(net5785),
    .D(_00987_),
    .Q_N(_07490_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][17] ));
 sg13g2_dfrbp_1 _17790_ (.CLK(net5275),
    .RESET_B(net5786),
    .D(_00988_),
    .Q_N(_07491_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][18] ));
 sg13g2_dfrbp_1 _17791_ (.CLK(net5335),
    .RESET_B(net5845),
    .D(_00960_),
    .Q_N(_07492_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_dfrbp_1 _17792_ (.CLK(net5335),
    .RESET_B(net5845),
    .D(_00970_),
    .Q_N(_07493_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_dfrbp_1 _17793_ (.CLK(net5335),
    .RESET_B(net5845),
    .D(_00971_),
    .Q_N(_07494_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_dfrbp_1 _17794_ (.CLK(net5335),
    .RESET_B(net5845),
    .D(_00972_),
    .Q_N(_07495_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_dfrbp_1 _17795_ (.CLK(net5336),
    .RESET_B(net5846),
    .D(_00973_),
    .Q_N(_07496_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_dfrbp_1 _17796_ (.CLK(net5338),
    .RESET_B(net5848),
    .D(_00974_),
    .Q_N(_07497_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_dfrbp_1 _17797_ (.CLK(net5333),
    .RESET_B(net5843),
    .D(_00975_),
    .Q_N(_07498_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_dfrbp_1 _17798_ (.CLK(net5334),
    .RESET_B(net5844),
    .D(_00976_),
    .Q_N(_07499_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_dfrbp_1 _17799_ (.CLK(net5321),
    .RESET_B(net5833),
    .D(_00977_),
    .Q_N(_07500_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_dfrbp_1 _17800_ (.CLK(net5323),
    .RESET_B(net5831),
    .D(_00978_),
    .Q_N(_07501_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_dfrbp_1 _17801_ (.CLK(net5321),
    .RESET_B(net5831),
    .D(_00961_),
    .Q_N(_07502_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_dfrbp_1 _17802_ (.CLK(net5320),
    .RESET_B(net5828),
    .D(_00962_),
    .Q_N(_07503_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_dfrbp_1 _17803_ (.CLK(net5318),
    .RESET_B(net5828),
    .D(_00963_),
    .Q_N(_07504_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_dfrbp_1 _17804_ (.CLK(net5318),
    .RESET_B(net5828),
    .D(_00964_),
    .Q_N(_07505_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_dfrbp_1 _17805_ (.CLK(net5318),
    .RESET_B(net5828),
    .D(_00965_),
    .Q_N(_07506_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_dfrbp_1 _17806_ (.CLK(net5276),
    .RESET_B(net5787),
    .D(_00966_),
    .Q_N(_07507_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_dfrbp_1 _17807_ (.CLK(net5276),
    .RESET_B(net5786),
    .D(_00967_),
    .Q_N(_07508_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[16] ));
 sg13g2_dfrbp_1 _17808_ (.CLK(net5275),
    .RESET_B(net5785),
    .D(_00968_),
    .Q_N(_07509_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_dfrbp_1 _17809_ (.CLK(net5277),
    .RESET_B(net5787),
    .D(_00969_),
    .Q_N(_07510_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.u2.reg_value[18] ));
 sg13g2_dfrbp_1 _17810_ (.CLK(net5336),
    .RESET_B(net5846),
    .D(_00960_),
    .Q_N(_07511_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_dfrbp_1 _17811_ (.CLK(net5337),
    .RESET_B(net5846),
    .D(_00970_),
    .Q_N(_07512_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_dfrbp_1 _17812_ (.CLK(net5336),
    .RESET_B(net5847),
    .D(_00971_),
    .Q_N(_07513_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_dfrbp_1 _17813_ (.CLK(net5336),
    .RESET_B(net5846),
    .D(_00972_),
    .Q_N(_07514_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_dfrbp_1 _17814_ (.CLK(net5336),
    .RESET_B(net5846),
    .D(_00973_),
    .Q_N(_07515_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_dfrbp_1 _17815_ (.CLK(net5335),
    .RESET_B(net5845),
    .D(_00974_),
    .Q_N(_07516_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_dfrbp_1 _17816_ (.CLK(net5335),
    .RESET_B(net5845),
    .D(_00975_),
    .Q_N(_07517_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_dfrbp_1 _17817_ (.CLK(net5333),
    .RESET_B(net5843),
    .D(_00976_),
    .Q_N(_07518_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_dfrbp_1 _17818_ (.CLK(net5334),
    .RESET_B(net5844),
    .D(_00977_),
    .Q_N(_07519_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_dfrbp_1 _17819_ (.CLK(net5321),
    .RESET_B(net5831),
    .D(_00978_),
    .Q_N(_07520_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_dfrbp_1 _17820_ (.CLK(net5321),
    .RESET_B(net5831),
    .D(_00961_),
    .Q_N(_07521_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_dfrbp_1 _17821_ (.CLK(net5321),
    .RESET_B(net5831),
    .D(_00962_),
    .Q_N(_07522_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_dfrbp_1 _17822_ (.CLK(net5320),
    .RESET_B(net5828),
    .D(_00963_),
    .Q_N(_07523_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_dfrbp_1 _17823_ (.CLK(net5320),
    .RESET_B(net5830),
    .D(_00964_),
    .Q_N(_07524_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_dfrbp_1 _17824_ (.CLK(net5319),
    .RESET_B(net5829),
    .D(_00965_),
    .Q_N(_07525_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_dfrbp_1 _17825_ (.CLK(net5319),
    .RESET_B(net5829),
    .D(_00966_),
    .Q_N(_07526_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_dfrbp_1 _17826_ (.CLK(net5276),
    .RESET_B(net5786),
    .D(_00967_),
    .Q_N(_07527_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_dfrbp_1 _17827_ (.CLK(net5276),
    .RESET_B(net5785),
    .D(_00968_),
    .Q_N(_07528_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_dfrbp_1 _17828_ (.CLK(net5275),
    .RESET_B(net5785),
    .D(_00969_),
    .Q_N(_07529_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator2_out[18] ));
 sg13g2_dfrbp_1 _17829_ (.CLK(net5333),
    .RESET_B(net5843),
    .D(_01188_),
    .Q_N(_01188_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[0] ));
 sg13g2_dfrbp_1 _17830_ (.CLK(net5333),
    .RESET_B(net5843),
    .D(_00951_),
    .Q_N(_07530_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_dfrbp_1 _17831_ (.CLK(net5333),
    .RESET_B(net5843),
    .D(_00952_),
    .Q_N(_07531_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_dfrbp_1 _17832_ (.CLK(net5333),
    .RESET_B(net5843),
    .D(_00953_),
    .Q_N(_07532_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_dfrbp_1 _17833_ (.CLK(net5334),
    .RESET_B(net5844),
    .D(_00954_),
    .Q_N(_07533_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[4] ));
 sg13g2_dfrbp_1 _17834_ (.CLK(net5334),
    .RESET_B(net5844),
    .D(_00955_),
    .Q_N(_07534_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_dfrbp_1 _17835_ (.CLK(net5334),
    .RESET_B(net5844),
    .D(_00956_),
    .Q_N(_07535_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_dfrbp_1 _17836_ (.CLK(net5334),
    .RESET_B(net5844),
    .D(_00957_),
    .Q_N(_07536_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_dfrbp_1 _17837_ (.CLK(net5321),
    .RESET_B(net5831),
    .D(_00958_),
    .Q_N(_07537_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_dfrbp_1 _17838_ (.CLK(net5321),
    .RESET_B(net5831),
    .D(_00959_),
    .Q_N(_07538_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_dfrbp_1 _17839_ (.CLK(net5318),
    .RESET_B(net5830),
    .D(_00942_),
    .Q_N(_07539_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_dfrbp_1 _17840_ (.CLK(net5318),
    .RESET_B(net5830),
    .D(_00943_),
    .Q_N(_07540_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_dfrbp_1 _17841_ (.CLK(net5318),
    .RESET_B(net5828),
    .D(_00944_),
    .Q_N(_07541_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_dfrbp_1 _17842_ (.CLK(net5318),
    .RESET_B(net5828),
    .D(_00945_),
    .Q_N(_07542_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_dfrbp_1 _17843_ (.CLK(net5318),
    .RESET_B(net5828),
    .D(_00946_),
    .Q_N(_07543_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_dfrbp_1 _17844_ (.CLK(net5276),
    .RESET_B(net5786),
    .D(_00947_),
    .Q_N(_07544_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_dfrbp_1 _17845_ (.CLK(net5276),
    .RESET_B(net5786),
    .D(_00948_),
    .Q_N(_07545_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_dfrbp_1 _17846_ (.CLK(net5277),
    .RESET_B(net5786),
    .D(_00949_),
    .Q_N(_07546_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_dfrbp_1 _17847_ (.CLK(net5276),
    .RESET_B(net5786),
    .D(_00950_),
    .Q_N(_07547_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.u_top_module.integrator1_out[18] ));
 sg13g2_dfrbp_1 _17848_ (.CLK(net5096),
    .RESET_B(net413),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][0] ),
    .Q_N(_07548_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _17849_ (.CLK(net5093),
    .RESET_B(net414),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][1] ),
    .Q_N(_07549_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _17850_ (.CLK(net5094),
    .RESET_B(net415),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][2] ),
    .Q_N(_07550_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _17851_ (.CLK(net5094),
    .RESET_B(net416),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][3] ),
    .Q_N(_07551_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _17852_ (.CLK(net5095),
    .RESET_B(net417),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][4] ),
    .Q_N(_07552_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _17853_ (.CLK(net5095),
    .RESET_B(net418),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][5] ),
    .Q_N(_07553_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _17854_ (.CLK(net5093),
    .RESET_B(net419),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][6] ),
    .Q_N(_07554_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _17855_ (.CLK(net5093),
    .RESET_B(net420),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][7] ),
    .Q_N(_07555_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _17856_ (.CLK(net5081),
    .RESET_B(net421),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][8] ),
    .Q_N(_07556_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _17857_ (.CLK(net5082),
    .RESET_B(net422),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][9] ),
    .Q_N(_07557_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _17858_ (.CLK(net5080),
    .RESET_B(net423),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][10] ),
    .Q_N(_07558_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _17859_ (.CLK(net5080),
    .RESET_B(net424),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][11] ),
    .Q_N(_07559_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _17860_ (.CLK(net5077),
    .RESET_B(net425),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][12] ),
    .Q_N(_07560_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _17861_ (.CLK(net5077),
    .RESET_B(net426),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][13] ),
    .Q_N(_07561_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _17862_ (.CLK(net5076),
    .RESET_B(net427),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][14] ),
    .Q_N(_07562_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _17863_ (.CLK(net5076),
    .RESET_B(net428),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][15] ),
    .Q_N(_07563_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _17864_ (.CLK(net5076),
    .RESET_B(net429),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][16] ),
    .Q_N(_07564_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _17865_ (.CLK(net5054),
    .RESET_B(net430),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][17] ),
    .Q_N(_07565_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _17866_ (.CLK(net5054),
    .RESET_B(net431),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[0][18] ),
    .Q_N(_07566_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _17867_ (.CLK(net5096),
    .RESET_B(net432),
    .D(_00904_),
    .Q_N(_07567_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][0] ));
 sg13g2_dfrbp_1 _17868_ (.CLK(net5097),
    .RESET_B(net433),
    .D(_00914_),
    .Q_N(_07568_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][1] ));
 sg13g2_dfrbp_1 _17869_ (.CLK(net5098),
    .RESET_B(net434),
    .D(_00915_),
    .Q_N(_07569_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][2] ));
 sg13g2_dfrbp_1 _17870_ (.CLK(net5098),
    .RESET_B(net435),
    .D(_00916_),
    .Q_N(_07570_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][3] ));
 sg13g2_dfrbp_1 _17871_ (.CLK(net5098),
    .RESET_B(net436),
    .D(_00917_),
    .Q_N(_07571_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][4] ));
 sg13g2_dfrbp_1 _17872_ (.CLK(net5098),
    .RESET_B(net437),
    .D(_00918_),
    .Q_N(_07572_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][5] ));
 sg13g2_dfrbp_1 _17873_ (.CLK(net5095),
    .RESET_B(net438),
    .D(_00919_),
    .Q_N(_07573_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][6] ));
 sg13g2_dfrbp_1 _17874_ (.CLK(net5094),
    .RESET_B(net439),
    .D(_00920_),
    .Q_N(_07574_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][7] ));
 sg13g2_dfrbp_1 _17875_ (.CLK(net5093),
    .RESET_B(net440),
    .D(_00921_),
    .Q_N(_07575_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][8] ));
 sg13g2_dfrbp_1 _17876_ (.CLK(net5081),
    .RESET_B(net441),
    .D(_00922_),
    .Q_N(_07576_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][9] ));
 sg13g2_dfrbp_1 _17877_ (.CLK(net5080),
    .RESET_B(net442),
    .D(_00905_),
    .Q_N(_07577_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][10] ));
 sg13g2_dfrbp_1 _17878_ (.CLK(net5080),
    .RESET_B(net443),
    .D(_00906_),
    .Q_N(_07578_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][11] ));
 sg13g2_dfrbp_1 _17879_ (.CLK(net5080),
    .RESET_B(net444),
    .D(_00907_),
    .Q_N(_07579_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][12] ));
 sg13g2_dfrbp_1 _17880_ (.CLK(net5073),
    .RESET_B(net445),
    .D(_00908_),
    .Q_N(_07580_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][13] ));
 sg13g2_dfrbp_1 _17881_ (.CLK(net5073),
    .RESET_B(net446),
    .D(_00909_),
    .Q_N(_07581_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][14] ));
 sg13g2_dfrbp_1 _17882_ (.CLK(net5072),
    .RESET_B(net447),
    .D(_00910_),
    .Q_N(_07582_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][15] ));
 sg13g2_dfrbp_1 _17883_ (.CLK(net5072),
    .RESET_B(net448),
    .D(_00911_),
    .Q_N(_07583_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][16] ));
 sg13g2_dfrbp_1 _17884_ (.CLK(net5070),
    .RESET_B(net468),
    .D(_00912_),
    .Q_N(_07584_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][17] ));
 sg13g2_dfrbp_1 _17885_ (.CLK(net5076),
    .RESET_B(net405),
    .D(_00913_),
    .Q_N(_06516_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][18] ));
 sg13g2_dfrbp_1 _17886_ (.CLK(_01534_),
    .RESET_B(net404),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[0] ),
    .Q_N(_06515_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _17887_ (.CLK(_01535_),
    .RESET_B(net403),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[1] ),
    .Q_N(_06514_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _17888_ (.CLK(_01536_),
    .RESET_B(net402),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[2] ),
    .Q_N(_06513_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _17889_ (.CLK(_01537_),
    .RESET_B(net401),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[3] ),
    .Q_N(_06512_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _17890_ (.CLK(_01538_),
    .RESET_B(net400),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[4] ),
    .Q_N(_06511_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _17891_ (.CLK(_01539_),
    .RESET_B(net399),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[5] ),
    .Q_N(_06510_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _17892_ (.CLK(_01540_),
    .RESET_B(net398),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[6] ),
    .Q_N(_06509_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _17893_ (.CLK(_01541_),
    .RESET_B(net397),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[7] ),
    .Q_N(_06508_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _17894_ (.CLK(_01542_),
    .RESET_B(net396),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[8] ),
    .Q_N(_06507_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _17895_ (.CLK(_01543_),
    .RESET_B(net395),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[9] ),
    .Q_N(_06506_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _17896_ (.CLK(_01544_),
    .RESET_B(net394),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[10] ),
    .Q_N(_06505_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _17897_ (.CLK(_01545_),
    .RESET_B(net393),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[11] ),
    .Q_N(_06504_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _17898_ (.CLK(_01546_),
    .RESET_B(net392),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[12] ),
    .Q_N(_06503_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _17899_ (.CLK(_01547_),
    .RESET_B(net353),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[13] ),
    .Q_N(_06502_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _17900_ (.CLK(_01548_),
    .RESET_B(net352),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[14] ),
    .Q_N(_06501_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _17901_ (.CLK(_01549_),
    .RESET_B(net351),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[15] ),
    .Q_N(_06500_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _17902_ (.CLK(_01550_),
    .RESET_B(net350),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[16] ),
    .Q_N(_06499_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _17903_ (.CLK(_01551_),
    .RESET_B(net349),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[17] ),
    .Q_N(_06498_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _17904_ (.CLK(_01552_),
    .RESET_B(net469),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.temp_delay[18] ),
    .Q_N(_07585_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[1].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _17905_ (.CLK(net5097),
    .RESET_B(net470),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][0] ),
    .Q_N(_07586_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _17906_ (.CLK(net5097),
    .RESET_B(net471),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][1] ),
    .Q_N(_07587_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _17907_ (.CLK(net5099),
    .RESET_B(net472),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][2] ),
    .Q_N(_07588_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _17908_ (.CLK(net5099),
    .RESET_B(net473),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][3] ),
    .Q_N(_07589_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _17909_ (.CLK(net5098),
    .RESET_B(net474),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][4] ),
    .Q_N(_07590_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _17910_ (.CLK(net5098),
    .RESET_B(net475),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][5] ),
    .Q_N(_07591_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _17911_ (.CLK(net5098),
    .RESET_B(net476),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][6] ),
    .Q_N(_07592_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _17912_ (.CLK(net5094),
    .RESET_B(net477),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][7] ),
    .Q_N(_07593_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _17913_ (.CLK(net5093),
    .RESET_B(net478),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][8] ),
    .Q_N(_07594_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _17914_ (.CLK(net5081),
    .RESET_B(net479),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][9] ),
    .Q_N(_07595_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _17915_ (.CLK(net5081),
    .RESET_B(net480),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][10] ),
    .Q_N(_07596_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _17916_ (.CLK(net5080),
    .RESET_B(net481),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][11] ),
    .Q_N(_07597_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _17917_ (.CLK(net5078),
    .RESET_B(net482),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][12] ),
    .Q_N(_07598_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _17918_ (.CLK(net5078),
    .RESET_B(net483),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][13] ),
    .Q_N(_07599_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _17919_ (.CLK(net5073),
    .RESET_B(net484),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][14] ),
    .Q_N(_07600_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _17920_ (.CLK(net5073),
    .RESET_B(net485),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][15] ),
    .Q_N(_07601_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _17921_ (.CLK(net5072),
    .RESET_B(net486),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][16] ),
    .Q_N(_07602_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _17922_ (.CLK(net5072),
    .RESET_B(net487),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][17] ),
    .Q_N(_07603_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _17923_ (.CLK(net5076),
    .RESET_B(net488),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.comb_data[1][18] ),
    .Q_N(_07604_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _17924_ (.CLK(net5102),
    .RESET_B(net489),
    .D(_00923_),
    .Q_N(_07605_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17925_ (.CLK(net5097),
    .RESET_B(net490),
    .D(_00933_),
    .Q_N(_07606_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17926_ (.CLK(net5097),
    .RESET_B(net491),
    .D(_00934_),
    .Q_N(_07607_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17927_ (.CLK(net5097),
    .RESET_B(net492),
    .D(_00935_),
    .Q_N(_07608_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17928_ (.CLK(net5099),
    .RESET_B(net493),
    .D(_00936_),
    .Q_N(_07609_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17929_ (.CLK(net5099),
    .RESET_B(net494),
    .D(_00937_),
    .Q_N(_07610_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17930_ (.CLK(net5097),
    .RESET_B(net495),
    .D(_00938_),
    .Q_N(_07611_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17931_ (.CLK(net5096),
    .RESET_B(net496),
    .D(_00939_),
    .Q_N(_07612_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17932_ (.CLK(net5093),
    .RESET_B(net497),
    .D(_00940_),
    .Q_N(_07613_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17933_ (.CLK(net5081),
    .RESET_B(net498),
    .D(_00941_),
    .Q_N(_07614_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17934_ (.CLK(net5083),
    .RESET_B(net499),
    .D(_00924_),
    .Q_N(_07615_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17935_ (.CLK(net5078),
    .RESET_B(net500),
    .D(_00925_),
    .Q_N(_07616_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17936_ (.CLK(net5079),
    .RESET_B(net501),
    .D(_00926_),
    .Q_N(_07617_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17937_ (.CLK(net5079),
    .RESET_B(net502),
    .D(_00927_),
    .Q_N(_07618_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17938_ (.CLK(net5078),
    .RESET_B(net503),
    .D(_00928_),
    .Q_N(_07619_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17939_ (.CLK(net5078),
    .RESET_B(net504),
    .D(_00929_),
    .Q_N(_07620_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17940_ (.CLK(net5078),
    .RESET_B(net505),
    .D(_00930_),
    .Q_N(_07621_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17941_ (.CLK(net5073),
    .RESET_B(net525),
    .D(_00931_),
    .Q_N(_07622_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17942_ (.CLK(net5072),
    .RESET_B(net348),
    .D(_00932_),
    .Q_N(_06497_),
    .Q(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _17943_ (.CLK(_01553_),
    .RESET_B(net347),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[0] ),
    .Q_N(_06496_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _17944_ (.CLK(_01554_),
    .RESET_B(net346),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[1] ),
    .Q_N(_06495_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _17945_ (.CLK(_01555_),
    .RESET_B(net345),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[2] ),
    .Q_N(_06494_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _17946_ (.CLK(_01556_),
    .RESET_B(net344),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[3] ),
    .Q_N(_06493_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _17947_ (.CLK(_01557_),
    .RESET_B(net343),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[4] ),
    .Q_N(_06492_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _17948_ (.CLK(_01558_),
    .RESET_B(net342),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[5] ),
    .Q_N(_06491_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _17949_ (.CLK(_01559_),
    .RESET_B(net341),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[6] ),
    .Q_N(_06490_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _17950_ (.CLK(_01560_),
    .RESET_B(net340),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[7] ),
    .Q_N(_06489_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _17951_ (.CLK(_01561_),
    .RESET_B(net339),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[8] ),
    .Q_N(_06488_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _17952_ (.CLK(_01562_),
    .RESET_B(net338),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[9] ),
    .Q_N(_06487_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _17953_ (.CLK(_01563_),
    .RESET_B(net337),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[10] ),
    .Q_N(_06486_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _17954_ (.CLK(_01564_),
    .RESET_B(net336),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[11] ),
    .Q_N(_06485_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _17955_ (.CLK(_01565_),
    .RESET_B(net335),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[12] ),
    .Q_N(_06484_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _17956_ (.CLK(_01566_),
    .RESET_B(net296),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[13] ),
    .Q_N(_06483_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _17957_ (.CLK(_01567_),
    .RESET_B(net295),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[14] ),
    .Q_N(_06482_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _17958_ (.CLK(_01568_),
    .RESET_B(net294),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[15] ),
    .Q_N(_06481_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _17959_ (.CLK(_01569_),
    .RESET_B(net293),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[16] ),
    .Q_N(_06480_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _17960_ (.CLK(_01570_),
    .RESET_B(net292),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[17] ),
    .Q_N(_06479_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _17961_ (.CLK(_01571_),
    .RESET_B(net526),
    .D(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.temp_delay[18] ),
    .Q_N(_07623_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.genblk1[2].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _17962_ (.CLK(net5207),
    .RESET_B(net5717),
    .D(_00885_),
    .Q_N(_07624_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_dfrbp_1 _17963_ (.CLK(net5207),
    .RESET_B(net5717),
    .D(_00895_),
    .Q_N(_07625_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_dfrbp_1 _17964_ (.CLK(net5207),
    .RESET_B(net5717),
    .D(_00896_),
    .Q_N(_07626_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_dfrbp_1 _17965_ (.CLK(net5207),
    .RESET_B(net5717),
    .D(_00897_),
    .Q_N(_07627_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_dfrbp_1 _17966_ (.CLK(net5204),
    .RESET_B(net5714),
    .D(_00898_),
    .Q_N(_07628_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_dfrbp_1 _17967_ (.CLK(net5204),
    .RESET_B(net5714),
    .D(_00899_),
    .Q_N(_07629_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_dfrbp_1 _17968_ (.CLK(net5204),
    .RESET_B(net5714),
    .D(_00900_),
    .Q_N(_07630_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_dfrbp_1 _17969_ (.CLK(net5204),
    .RESET_B(net5714),
    .D(_00901_),
    .Q_N(_07631_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_dfrbp_1 _17970_ (.CLK(net5186),
    .RESET_B(net5696),
    .D(_00902_),
    .Q_N(_07632_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_dfrbp_1 _17971_ (.CLK(net5185),
    .RESET_B(net5695),
    .D(_00903_),
    .Q_N(_07633_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_dfrbp_1 _17972_ (.CLK(net5184),
    .RESET_B(net5694),
    .D(_00886_),
    .Q_N(_07634_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_dfrbp_1 _17973_ (.CLK(net5187),
    .RESET_B(net5697),
    .D(_00887_),
    .Q_N(_07635_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_dfrbp_1 _17974_ (.CLK(net5184),
    .RESET_B(net5694),
    .D(_00888_),
    .Q_N(_07636_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_dfrbp_1 _17975_ (.CLK(net5181),
    .RESET_B(net5691),
    .D(_00889_),
    .Q_N(_07637_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_dfrbp_1 _17976_ (.CLK(net5181),
    .RESET_B(net5691),
    .D(_00890_),
    .Q_N(_07638_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_dfrbp_1 _17977_ (.CLK(net5178),
    .RESET_B(net5688),
    .D(_00891_),
    .Q_N(_07639_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_dfrbp_1 _17978_ (.CLK(net5179),
    .RESET_B(net5689),
    .D(_00892_),
    .Q_N(_07640_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_dfrbp_1 _17979_ (.CLK(net5179),
    .RESET_B(net5689),
    .D(_00893_),
    .Q_N(_07641_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_dfrbp_1 _17980_ (.CLK(net5179),
    .RESET_B(net5689),
    .D(_00894_),
    .Q_N(_07642_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u3.reg_value[18] ));
 sg13g2_dfrbp_1 _17981_ (.CLK(net5205),
    .RESET_B(net5715),
    .D(_00885_),
    .Q_N(_07643_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][0] ));
 sg13g2_dfrbp_1 _17982_ (.CLK(net5206),
    .RESET_B(net5716),
    .D(_00895_),
    .Q_N(_07644_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][1] ));
 sg13g2_dfrbp_1 _17983_ (.CLK(net5205),
    .RESET_B(net5715),
    .D(_00896_),
    .Q_N(_07645_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][2] ));
 sg13g2_dfrbp_1 _17984_ (.CLK(net5205),
    .RESET_B(net5715),
    .D(_00897_),
    .Q_N(_07646_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][3] ));
 sg13g2_dfrbp_1 _17985_ (.CLK(net5204),
    .RESET_B(net5714),
    .D(_00898_),
    .Q_N(_07647_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][4] ));
 sg13g2_dfrbp_1 _17986_ (.CLK(net5204),
    .RESET_B(net5714),
    .D(_00899_),
    .Q_N(_07648_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][5] ));
 sg13g2_dfrbp_1 _17987_ (.CLK(net5204),
    .RESET_B(net5714),
    .D(_00900_),
    .Q_N(_07649_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][6] ));
 sg13g2_dfrbp_1 _17988_ (.CLK(net5185),
    .RESET_B(net5695),
    .D(_00901_),
    .Q_N(_07650_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][7] ));
 sg13g2_dfrbp_1 _17989_ (.CLK(net5185),
    .RESET_B(net5695),
    .D(_00902_),
    .Q_N(_07651_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][8] ));
 sg13g2_dfrbp_1 _17990_ (.CLK(net5185),
    .RESET_B(net5695),
    .D(_00903_),
    .Q_N(_07652_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][9] ));
 sg13g2_dfrbp_1 _17991_ (.CLK(net5185),
    .RESET_B(net5695),
    .D(_00886_),
    .Q_N(_07653_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][10] ));
 sg13g2_dfrbp_1 _17992_ (.CLK(net5185),
    .RESET_B(net5695),
    .D(_00887_),
    .Q_N(_07654_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][11] ));
 sg13g2_dfrbp_1 _17993_ (.CLK(net5186),
    .RESET_B(net5696),
    .D(_00888_),
    .Q_N(_07655_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][12] ));
 sg13g2_dfrbp_1 _17994_ (.CLK(net5186),
    .RESET_B(net5696),
    .D(_00889_),
    .Q_N(_07656_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][13] ));
 sg13g2_dfrbp_1 _17995_ (.CLK(net5181),
    .RESET_B(net5691),
    .D(_00890_),
    .Q_N(_07657_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][14] ));
 sg13g2_dfrbp_1 _17996_ (.CLK(net5180),
    .RESET_B(net5690),
    .D(_00891_),
    .Q_N(_07658_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][15] ));
 sg13g2_dfrbp_1 _17997_ (.CLK(net5180),
    .RESET_B(net5690),
    .D(_00892_),
    .Q_N(_07659_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][16] ));
 sg13g2_dfrbp_1 _17998_ (.CLK(net5180),
    .RESET_B(net5690),
    .D(_00893_),
    .Q_N(_07660_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][17] ));
 sg13g2_dfrbp_1 _17999_ (.CLK(net5180),
    .RESET_B(net5690),
    .D(_00894_),
    .Q_N(_07661_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][18] ));
 sg13g2_dfrbp_1 _18000_ (.CLK(net5202),
    .RESET_B(net5711),
    .D(_00866_),
    .Q_N(_07662_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_dfrbp_1 _18001_ (.CLK(net5202),
    .RESET_B(net5712),
    .D(_00876_),
    .Q_N(_07663_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_dfrbp_1 _18002_ (.CLK(net5202),
    .RESET_B(net5712),
    .D(_00877_),
    .Q_N(_07664_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_dfrbp_1 _18003_ (.CLK(net5202),
    .RESET_B(net5712),
    .D(_00878_),
    .Q_N(_07665_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_dfrbp_1 _18004_ (.CLK(net5203),
    .RESET_B(net5713),
    .D(_00879_),
    .Q_N(_07666_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_dfrbp_1 _18005_ (.CLK(net5203),
    .RESET_B(net5710),
    .D(_00880_),
    .Q_N(_07667_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_dfrbp_1 _18006_ (.CLK(net5200),
    .RESET_B(net5713),
    .D(_00881_),
    .Q_N(_07668_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_dfrbp_1 _18007_ (.CLK(net5199),
    .RESET_B(net5709),
    .D(_00882_),
    .Q_N(_07669_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_dfrbp_1 _18008_ (.CLK(net5199),
    .RESET_B(net5709),
    .D(_00883_),
    .Q_N(_07670_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_dfrbp_1 _18009_ (.CLK(net5199),
    .RESET_B(net5709),
    .D(_00884_),
    .Q_N(_07671_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_dfrbp_1 _18010_ (.CLK(net5183),
    .RESET_B(net5693),
    .D(_00867_),
    .Q_N(_07672_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_dfrbp_1 _18011_ (.CLK(net5183),
    .RESET_B(net5693),
    .D(_00868_),
    .Q_N(_07673_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_dfrbp_1 _18012_ (.CLK(net5183),
    .RESET_B(net5693),
    .D(_00869_),
    .Q_N(_07674_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_dfrbp_1 _18013_ (.CLK(net5183),
    .RESET_B(net5693),
    .D(_00870_),
    .Q_N(_07675_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_dfrbp_1 _18014_ (.CLK(net5182),
    .RESET_B(net5692),
    .D(_00871_),
    .Q_N(_07676_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_dfrbp_1 _18015_ (.CLK(net5182),
    .RESET_B(net5692),
    .D(_00872_),
    .Q_N(_07677_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_dfrbp_1 _18016_ (.CLK(net5178),
    .RESET_B(net5688),
    .D(_00873_),
    .Q_N(_07678_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[16] ));
 sg13g2_dfrbp_1 _18017_ (.CLK(net5178),
    .RESET_B(net5688),
    .D(_00874_),
    .Q_N(_07679_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_dfrbp_1 _18018_ (.CLK(net5178),
    .RESET_B(net5688),
    .D(_00875_),
    .Q_N(_07680_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.u2.reg_value[18] ));
 sg13g2_dfrbp_1 _18019_ (.CLK(net5201),
    .RESET_B(net5712),
    .D(_00866_),
    .Q_N(_07681_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_dfrbp_1 _18020_ (.CLK(net5202),
    .RESET_B(net5712),
    .D(_00876_),
    .Q_N(_07682_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_dfrbp_1 _18021_ (.CLK(net5201),
    .RESET_B(net5711),
    .D(_00877_),
    .Q_N(_07683_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_dfrbp_1 _18022_ (.CLK(net5201),
    .RESET_B(net5711),
    .D(_00878_),
    .Q_N(_07684_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_dfrbp_1 _18023_ (.CLK(net5200),
    .RESET_B(net5710),
    .D(_00879_),
    .Q_N(_07685_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_dfrbp_1 _18024_ (.CLK(net5200),
    .RESET_B(net5710),
    .D(_00880_),
    .Q_N(_07686_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_dfrbp_1 _18025_ (.CLK(net5200),
    .RESET_B(net5710),
    .D(_00881_),
    .Q_N(_07687_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_dfrbp_1 _18026_ (.CLK(net5200),
    .RESET_B(net5710),
    .D(_00882_),
    .Q_N(_07688_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_dfrbp_1 _18027_ (.CLK(net5203),
    .RESET_B(net5713),
    .D(_00883_),
    .Q_N(_07689_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_dfrbp_1 _18028_ (.CLK(net5184),
    .RESET_B(net5694),
    .D(_00884_),
    .Q_N(_07690_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_dfrbp_1 _18029_ (.CLK(net5184),
    .RESET_B(net5694),
    .D(_00867_),
    .Q_N(_07691_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_dfrbp_1 _18030_ (.CLK(net5184),
    .RESET_B(net5694),
    .D(_00868_),
    .Q_N(_07692_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_dfrbp_1 _18031_ (.CLK(net5184),
    .RESET_B(net5694),
    .D(_00869_),
    .Q_N(_07693_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_dfrbp_1 _18032_ (.CLK(net5183),
    .RESET_B(net5692),
    .D(_00870_),
    .Q_N(_07694_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_dfrbp_1 _18033_ (.CLK(net5182),
    .RESET_B(net5693),
    .D(_00871_),
    .Q_N(_07695_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_dfrbp_1 _18034_ (.CLK(net5179),
    .RESET_B(net5689),
    .D(_00872_),
    .Q_N(_07696_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_dfrbp_1 _18035_ (.CLK(net5178),
    .RESET_B(net5688),
    .D(_00873_),
    .Q_N(_07697_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_dfrbp_1 _18036_ (.CLK(net5178),
    .RESET_B(net5688),
    .D(_00874_),
    .Q_N(_07698_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_dfrbp_1 _18037_ (.CLK(net5178),
    .RESET_B(net5688),
    .D(_00875_),
    .Q_N(_07699_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator2_out[18] ));
 sg13g2_dfrbp_1 _18038_ (.CLK(net5201),
    .RESET_B(net5711),
    .D(_01189_),
    .Q_N(_01189_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[0] ));
 sg13g2_dfrbp_1 _18039_ (.CLK(net5201),
    .RESET_B(net5711),
    .D(_00857_),
    .Q_N(_07700_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_dfrbp_1 _18040_ (.CLK(net5201),
    .RESET_B(net5711),
    .D(_00858_),
    .Q_N(_07701_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_dfrbp_1 _18041_ (.CLK(net5201),
    .RESET_B(net5711),
    .D(_00859_),
    .Q_N(_07702_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_dfrbp_1 _18042_ (.CLK(net5200),
    .RESET_B(net5710),
    .D(_00860_),
    .Q_N(_07703_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[4] ));
 sg13g2_dfrbp_1 _18043_ (.CLK(net5200),
    .RESET_B(net5710),
    .D(_00861_),
    .Q_N(_07704_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_dfrbp_1 _18044_ (.CLK(net5199),
    .RESET_B(net5709),
    .D(_00862_),
    .Q_N(_07705_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_dfrbp_1 _18045_ (.CLK(net5199),
    .RESET_B(net5709),
    .D(_00863_),
    .Q_N(_07706_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_dfrbp_1 _18046_ (.CLK(net5199),
    .RESET_B(net5709),
    .D(_00864_),
    .Q_N(_07707_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_dfrbp_1 _18047_ (.CLK(net5199),
    .RESET_B(net5709),
    .D(_00865_),
    .Q_N(_07708_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_dfrbp_1 _18048_ (.CLK(net5184),
    .RESET_B(net5694),
    .D(_00848_),
    .Q_N(_07709_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_dfrbp_1 _18049_ (.CLK(net5183),
    .RESET_B(net5693),
    .D(_00849_),
    .Q_N(_07710_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_dfrbp_1 _18050_ (.CLK(net5183),
    .RESET_B(net5693),
    .D(_00850_),
    .Q_N(_07711_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_dfrbp_1 _18051_ (.CLK(net5182),
    .RESET_B(net5692),
    .D(_00851_),
    .Q_N(_07712_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_dfrbp_1 _18052_ (.CLK(net5182),
    .RESET_B(net5692),
    .D(_00852_),
    .Q_N(_07713_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_dfrbp_1 _18053_ (.CLK(net5182),
    .RESET_B(net5692),
    .D(_00853_),
    .Q_N(_07714_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_dfrbp_1 _18054_ (.CLK(net5182),
    .RESET_B(net5692),
    .D(_00854_),
    .Q_N(_07715_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_dfrbp_1 _18055_ (.CLK(net5182),
    .RESET_B(net5692),
    .D(_00855_),
    .Q_N(_07716_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_dfrbp_1 _18056_ (.CLK(net5178),
    .RESET_B(net5688),
    .D(_00856_),
    .Q_N(_07717_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.u_top_module.integrator1_out[18] ));
 sg13g2_dfrbp_1 _18057_ (.CLK(net5027),
    .RESET_B(net527),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][0] ),
    .Q_N(_07718_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18058_ (.CLK(net5025),
    .RESET_B(net528),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][1] ),
    .Q_N(_07719_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18059_ (.CLK(net5025),
    .RESET_B(net529),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][2] ),
    .Q_N(_07720_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18060_ (.CLK(net5025),
    .RESET_B(net530),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][3] ),
    .Q_N(_07721_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18061_ (.CLK(net5025),
    .RESET_B(net531),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][4] ),
    .Q_N(_07722_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18062_ (.CLK(net5025),
    .RESET_B(net532),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][5] ),
    .Q_N(_07723_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18063_ (.CLK(net5012),
    .RESET_B(net533),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][6] ),
    .Q_N(_07724_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18064_ (.CLK(net5013),
    .RESET_B(net534),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][7] ),
    .Q_N(_07725_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18065_ (.CLK(net5012),
    .RESET_B(net535),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][8] ),
    .Q_N(_07726_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18066_ (.CLK(net5012),
    .RESET_B(net536),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][9] ),
    .Q_N(_07727_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18067_ (.CLK(net5012),
    .RESET_B(net537),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][10] ),
    .Q_N(_07728_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18068_ (.CLK(net5011),
    .RESET_B(net538),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][11] ),
    .Q_N(_07729_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18069_ (.CLK(net5011),
    .RESET_B(net539),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][12] ),
    .Q_N(_07730_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18070_ (.CLK(net5011),
    .RESET_B(net540),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][13] ),
    .Q_N(_07731_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18071_ (.CLK(net5014),
    .RESET_B(net541),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][14] ),
    .Q_N(_07732_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18072_ (.CLK(net5014),
    .RESET_B(net542),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][15] ),
    .Q_N(_07733_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18073_ (.CLK(net5014),
    .RESET_B(net543),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][16] ),
    .Q_N(_07734_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18074_ (.CLK(net5015),
    .RESET_B(net544),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][17] ),
    .Q_N(_07735_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18075_ (.CLK(net5015),
    .RESET_B(net545),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[0][18] ),
    .Q_N(_07736_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18076_ (.CLK(net5027),
    .RESET_B(net546),
    .D(_00810_),
    .Q_N(_07737_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][0] ));
 sg13g2_dfrbp_1 _18077_ (.CLK(net5027),
    .RESET_B(net547),
    .D(_00820_),
    .Q_N(_07738_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][1] ));
 sg13g2_dfrbp_1 _18078_ (.CLK(net5027),
    .RESET_B(net548),
    .D(_00821_),
    .Q_N(_07739_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][2] ));
 sg13g2_dfrbp_1 _18079_ (.CLK(net5027),
    .RESET_B(net549),
    .D(_00822_),
    .Q_N(_07740_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][3] ));
 sg13g2_dfrbp_1 _18080_ (.CLK(net5027),
    .RESET_B(net550),
    .D(_00823_),
    .Q_N(_07741_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][4] ));
 sg13g2_dfrbp_1 _18081_ (.CLK(net5019),
    .RESET_B(net551),
    .D(_00824_),
    .Q_N(_07742_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][5] ));
 sg13g2_dfrbp_1 _18082_ (.CLK(net5019),
    .RESET_B(net552),
    .D(_00825_),
    .Q_N(_07743_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][6] ));
 sg13g2_dfrbp_1 _18083_ (.CLK(net5019),
    .RESET_B(net553),
    .D(_00826_),
    .Q_N(_07744_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][7] ));
 sg13g2_dfrbp_1 _18084_ (.CLK(net5019),
    .RESET_B(net554),
    .D(_00827_),
    .Q_N(_07745_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][8] ));
 sg13g2_dfrbp_1 _18085_ (.CLK(net5019),
    .RESET_B(net555),
    .D(_00828_),
    .Q_N(_07746_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][9] ));
 sg13g2_dfrbp_1 _18086_ (.CLK(net5018),
    .RESET_B(net556),
    .D(_00811_),
    .Q_N(_07747_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][10] ));
 sg13g2_dfrbp_1 _18087_ (.CLK(net5018),
    .RESET_B(net557),
    .D(_00812_),
    .Q_N(_07748_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][11] ));
 sg13g2_dfrbp_1 _18088_ (.CLK(net5018),
    .RESET_B(net558),
    .D(_00813_),
    .Q_N(_07749_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][12] ));
 sg13g2_dfrbp_1 _18089_ (.CLK(net5018),
    .RESET_B(net559),
    .D(_00814_),
    .Q_N(_07750_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][13] ));
 sg13g2_dfrbp_1 _18090_ (.CLK(net5018),
    .RESET_B(net560),
    .D(_00815_),
    .Q_N(_07751_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][14] ));
 sg13g2_dfrbp_1 _18091_ (.CLK(net5013),
    .RESET_B(net561),
    .D(_00816_),
    .Q_N(_07752_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][15] ));
 sg13g2_dfrbp_1 _18092_ (.CLK(net5011),
    .RESET_B(net562),
    .D(_00817_),
    .Q_N(_07753_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][16] ));
 sg13g2_dfrbp_1 _18093_ (.CLK(net5011),
    .RESET_B(net582),
    .D(_00818_),
    .Q_N(_07754_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][17] ));
 sg13g2_dfrbp_1 _18094_ (.CLK(net5013),
    .RESET_B(net291),
    .D(_00819_),
    .Q_N(_06478_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][18] ));
 sg13g2_dfrbp_1 _18095_ (.CLK(_01572_),
    .RESET_B(net290),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[0] ),
    .Q_N(_06477_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18096_ (.CLK(_01573_),
    .RESET_B(net289),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[1] ),
    .Q_N(_06476_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18097_ (.CLK(_01574_),
    .RESET_B(net288),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[2] ),
    .Q_N(_06475_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18098_ (.CLK(_01575_),
    .RESET_B(net287),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[3] ),
    .Q_N(_06474_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18099_ (.CLK(_01576_),
    .RESET_B(net286),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[4] ),
    .Q_N(_06473_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18100_ (.CLK(_01577_),
    .RESET_B(net285),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[5] ),
    .Q_N(_06472_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18101_ (.CLK(_01578_),
    .RESET_B(net284),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[6] ),
    .Q_N(_06471_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18102_ (.CLK(_01579_),
    .RESET_B(net283),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[7] ),
    .Q_N(_06470_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18103_ (.CLK(_01580_),
    .RESET_B(net282),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[8] ),
    .Q_N(_06469_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18104_ (.CLK(_01581_),
    .RESET_B(net281),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[9] ),
    .Q_N(_06468_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18105_ (.CLK(_01582_),
    .RESET_B(net280),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[10] ),
    .Q_N(_06467_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18106_ (.CLK(_01583_),
    .RESET_B(net279),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[11] ),
    .Q_N(_06466_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _18107_ (.CLK(_01584_),
    .RESET_B(net278),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[12] ),
    .Q_N(_06465_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _18108_ (.CLK(_01585_),
    .RESET_B(net239),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[13] ),
    .Q_N(_06464_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _18109_ (.CLK(_01586_),
    .RESET_B(net238),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[14] ),
    .Q_N(_06463_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _18110_ (.CLK(_01587_),
    .RESET_B(net237),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[15] ),
    .Q_N(_06462_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _18111_ (.CLK(_01588_),
    .RESET_B(net236),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[16] ),
    .Q_N(_06461_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _18112_ (.CLK(_01589_),
    .RESET_B(net235),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[17] ),
    .Q_N(_06460_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _18113_ (.CLK(_01590_),
    .RESET_B(net583),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.temp_delay[18] ),
    .Q_N(_07755_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[1].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _18114_ (.CLK(net5026),
    .RESET_B(net584),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][0] ),
    .Q_N(_07756_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18115_ (.CLK(net5026),
    .RESET_B(net585),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][1] ),
    .Q_N(_07757_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18116_ (.CLK(net5026),
    .RESET_B(net586),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][2] ),
    .Q_N(_07758_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18117_ (.CLK(net5026),
    .RESET_B(net587),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][3] ),
    .Q_N(_07759_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18118_ (.CLK(net5026),
    .RESET_B(net588),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][4] ),
    .Q_N(_07760_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18119_ (.CLK(net5023),
    .RESET_B(net589),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][5] ),
    .Q_N(_07761_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18120_ (.CLK(net5023),
    .RESET_B(net590),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][6] ),
    .Q_N(_07762_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18121_ (.CLK(net5019),
    .RESET_B(net591),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][7] ),
    .Q_N(_07763_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18122_ (.CLK(net5019),
    .RESET_B(net592),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][8] ),
    .Q_N(_07764_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18123_ (.CLK(net5019),
    .RESET_B(net593),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][9] ),
    .Q_N(_07765_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18124_ (.CLK(net5017),
    .RESET_B(net594),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][10] ),
    .Q_N(_07766_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18125_ (.CLK(net5016),
    .RESET_B(net595),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][11] ),
    .Q_N(_07767_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18126_ (.CLK(net5017),
    .RESET_B(net596),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][12] ),
    .Q_N(_07768_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18127_ (.CLK(net5016),
    .RESET_B(net597),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][13] ),
    .Q_N(_07769_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18128_ (.CLK(net5016),
    .RESET_B(net598),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][14] ),
    .Q_N(_07770_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18129_ (.CLK(net5024),
    .RESET_B(net599),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][15] ),
    .Q_N(_07771_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18130_ (.CLK(net5016),
    .RESET_B(net600),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][16] ),
    .Q_N(_07772_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18131_ (.CLK(net5018),
    .RESET_B(net601),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][17] ),
    .Q_N(_07773_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18132_ (.CLK(net5018),
    .RESET_B(net602),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.comb_data[1][18] ),
    .Q_N(_07774_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18133_ (.CLK(net5047),
    .RESET_B(net603),
    .D(_00829_),
    .Q_N(_07775_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18134_ (.CLK(net5047),
    .RESET_B(net604),
    .D(_00839_),
    .Q_N(_07776_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18135_ (.CLK(net5047),
    .RESET_B(net605),
    .D(_00840_),
    .Q_N(_07777_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18136_ (.CLK(net5034),
    .RESET_B(net606),
    .D(_00841_),
    .Q_N(_07778_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18137_ (.CLK(net5034),
    .RESET_B(net607),
    .D(_00842_),
    .Q_N(_07779_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18138_ (.CLK(net5023),
    .RESET_B(net608),
    .D(_00843_),
    .Q_N(_07780_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18139_ (.CLK(net5034),
    .RESET_B(net609),
    .D(_00844_),
    .Q_N(_07781_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18140_ (.CLK(net5034),
    .RESET_B(net610),
    .D(_00845_),
    .Q_N(_07782_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18141_ (.CLK(net5022),
    .RESET_B(net611),
    .D(_00846_),
    .Q_N(_07783_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18142_ (.CLK(net5021),
    .RESET_B(net612),
    .D(_00847_),
    .Q_N(_07784_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18143_ (.CLK(net5021),
    .RESET_B(net613),
    .D(_00830_),
    .Q_N(_07785_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18144_ (.CLK(net5021),
    .RESET_B(net614),
    .D(_00831_),
    .Q_N(_07786_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18145_ (.CLK(net5021),
    .RESET_B(net615),
    .D(_00832_),
    .Q_N(_07787_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18146_ (.CLK(net5022),
    .RESET_B(net616),
    .D(_00833_),
    .Q_N(_07788_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18147_ (.CLK(net5021),
    .RESET_B(net617),
    .D(_00834_),
    .Q_N(_07789_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18148_ (.CLK(net5021),
    .RESET_B(net618),
    .D(_00835_),
    .Q_N(_07790_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18149_ (.CLK(net5021),
    .RESET_B(net619),
    .D(_00836_),
    .Q_N(_07791_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18150_ (.CLK(net5021),
    .RESET_B(net634),
    .D(_00837_),
    .Q_N(_07792_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18151_ (.CLK(net5022),
    .RESET_B(net234),
    .D(_00838_),
    .Q_N(_06459_),
    .Q(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18152_ (.CLK(_01591_),
    .RESET_B(net233),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[0] ),
    .Q_N(_06458_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18153_ (.CLK(_01592_),
    .RESET_B(net232),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[1] ),
    .Q_N(_06457_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18154_ (.CLK(_01593_),
    .RESET_B(net231),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[2] ),
    .Q_N(_06456_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18155_ (.CLK(_01594_),
    .RESET_B(net230),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[3] ),
    .Q_N(_06455_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18156_ (.CLK(_01595_),
    .RESET_B(net229),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[4] ),
    .Q_N(_06454_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18157_ (.CLK(_01596_),
    .RESET_B(net228),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[5] ),
    .Q_N(_06453_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18158_ (.CLK(_01597_),
    .RESET_B(net227),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[6] ),
    .Q_N(_06452_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18159_ (.CLK(_01598_),
    .RESET_B(net226),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[7] ),
    .Q_N(_06451_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18160_ (.CLK(_01599_),
    .RESET_B(net225),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[8] ),
    .Q_N(_06450_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18161_ (.CLK(_01600_),
    .RESET_B(net224),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[9] ),
    .Q_N(_06449_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18162_ (.CLK(_01601_),
    .RESET_B(net223),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[10] ),
    .Q_N(_06448_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18163_ (.CLK(_01602_),
    .RESET_B(net222),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[11] ),
    .Q_N(_06447_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _18164_ (.CLK(_01603_),
    .RESET_B(net221),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[12] ),
    .Q_N(_06446_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _18165_ (.CLK(_01604_),
    .RESET_B(net184),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[13] ),
    .Q_N(_06445_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _18166_ (.CLK(_01605_),
    .RESET_B(net183),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[14] ),
    .Q_N(_06444_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _18167_ (.CLK(_01606_),
    .RESET_B(net182),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[15] ),
    .Q_N(_06443_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _18168_ (.CLK(_01607_),
    .RESET_B(net181),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[16] ),
    .Q_N(_06442_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _18169_ (.CLK(_01608_),
    .RESET_B(net180),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[17] ),
    .Q_N(_06441_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _18170_ (.CLK(_01609_),
    .RESET_B(net635),
    .D(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.temp_delay[18] ),
    .Q_N(_07793_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.genblk1[2].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _18171_ (.CLK(net5558),
    .RESET_B(net6067),
    .D(_00791_),
    .Q_N(_07794_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_dfrbp_1 _18172_ (.CLK(net5561),
    .RESET_B(net6070),
    .D(_00801_),
    .Q_N(_07795_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_dfrbp_1 _18173_ (.CLK(net5561),
    .RESET_B(net6070),
    .D(_00802_),
    .Q_N(_07796_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_dfrbp_1 _18174_ (.CLK(net5561),
    .RESET_B(net6070),
    .D(_00803_),
    .Q_N(_07797_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_dfrbp_1 _18175_ (.CLK(net5579),
    .RESET_B(net6088),
    .D(_00804_),
    .Q_N(_07798_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_dfrbp_1 _18176_ (.CLK(net5579),
    .RESET_B(net6088),
    .D(_00805_),
    .Q_N(_07799_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_dfrbp_1 _18177_ (.CLK(net5579),
    .RESET_B(net6088),
    .D(_00806_),
    .Q_N(_07800_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_dfrbp_1 _18178_ (.CLK(net5579),
    .RESET_B(net6088),
    .D(_00807_),
    .Q_N(_07801_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_dfrbp_1 _18179_ (.CLK(net5561),
    .RESET_B(net6071),
    .D(_00808_),
    .Q_N(_07802_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_dfrbp_1 _18180_ (.CLK(net5561),
    .RESET_B(net6070),
    .D(_00809_),
    .Q_N(_07803_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_dfrbp_1 _18181_ (.CLK(net5558),
    .RESET_B(net6067),
    .D(_00792_),
    .Q_N(_07804_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_dfrbp_1 _18182_ (.CLK(net5489),
    .RESET_B(net5998),
    .D(_00793_),
    .Q_N(_07805_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_dfrbp_1 _18183_ (.CLK(net5491),
    .RESET_B(net6000),
    .D(_00794_),
    .Q_N(_07806_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_dfrbp_1 _18184_ (.CLK(net5491),
    .RESET_B(net6000),
    .D(_00795_),
    .Q_N(_07807_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_dfrbp_1 _18185_ (.CLK(net5488),
    .RESET_B(net5997),
    .D(_00796_),
    .Q_N(_07808_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_dfrbp_1 _18186_ (.CLK(net5487),
    .RESET_B(net5996),
    .D(_00797_),
    .Q_N(_07809_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_dfrbp_1 _18187_ (.CLK(net5487),
    .RESET_B(net5996),
    .D(_00798_),
    .Q_N(_07810_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_dfrbp_1 _18188_ (.CLK(net5487),
    .RESET_B(net5996),
    .D(_00799_),
    .Q_N(_07811_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_dfrbp_1 _18189_ (.CLK(net5487),
    .RESET_B(net5996),
    .D(_00800_),
    .Q_N(_07812_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u3.reg_value[18] ));
 sg13g2_dfrbp_1 _18190_ (.CLK(net5560),
    .RESET_B(net6069),
    .D(_00791_),
    .Q_N(_07813_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][0] ));
 sg13g2_dfrbp_1 _18191_ (.CLK(net5560),
    .RESET_B(net6069),
    .D(_00801_),
    .Q_N(_07814_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][1] ));
 sg13g2_dfrbp_1 _18192_ (.CLK(net5561),
    .RESET_B(net6070),
    .D(_00802_),
    .Q_N(_07815_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][2] ));
 sg13g2_dfrbp_1 _18193_ (.CLK(net5579),
    .RESET_B(net6088),
    .D(_00803_),
    .Q_N(_07816_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][3] ));
 sg13g2_dfrbp_1 _18194_ (.CLK(net5579),
    .RESET_B(net6088),
    .D(_00804_),
    .Q_N(_07817_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][4] ));
 sg13g2_dfrbp_1 _18195_ (.CLK(net5580),
    .RESET_B(net6088),
    .D(_00805_),
    .Q_N(_07818_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][5] ));
 sg13g2_dfrbp_1 _18196_ (.CLK(net5581),
    .RESET_B(net6090),
    .D(_00806_),
    .Q_N(_07819_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][6] ));
 sg13g2_dfrbp_1 _18197_ (.CLK(net5579),
    .RESET_B(net6089),
    .D(_00807_),
    .Q_N(_07820_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][7] ));
 sg13g2_dfrbp_1 _18198_ (.CLK(net5580),
    .RESET_B(net6089),
    .D(_00808_),
    .Q_N(_07821_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][8] ));
 sg13g2_dfrbp_1 _18199_ (.CLK(net5579),
    .RESET_B(net6088),
    .D(_00809_),
    .Q_N(_07822_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][9] ));
 sg13g2_dfrbp_1 _18200_ (.CLK(net5561),
    .RESET_B(net6070),
    .D(_00792_),
    .Q_N(_07823_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][10] ));
 sg13g2_dfrbp_1 _18201_ (.CLK(net5563),
    .RESET_B(net6072),
    .D(_00793_),
    .Q_N(_07824_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][11] ));
 sg13g2_dfrbp_1 _18202_ (.CLK(net5491),
    .RESET_B(net6000),
    .D(_00794_),
    .Q_N(_07825_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][12] ));
 sg13g2_dfrbp_1 _18203_ (.CLK(net5491),
    .RESET_B(net6000),
    .D(_00795_),
    .Q_N(_07826_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][13] ));
 sg13g2_dfrbp_1 _18204_ (.CLK(net5488),
    .RESET_B(net5997),
    .D(_00796_),
    .Q_N(_07827_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][14] ));
 sg13g2_dfrbp_1 _18205_ (.CLK(net5487),
    .RESET_B(net5996),
    .D(_00797_),
    .Q_N(_07828_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][15] ));
 sg13g2_dfrbp_1 _18206_ (.CLK(net5488),
    .RESET_B(net5997),
    .D(_00798_),
    .Q_N(_07829_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][16] ));
 sg13g2_dfrbp_1 _18207_ (.CLK(net5484),
    .RESET_B(net5993),
    .D(_00799_),
    .Q_N(_07830_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][17] ));
 sg13g2_dfrbp_1 _18208_ (.CLK(net5487),
    .RESET_B(net5996),
    .D(_00800_),
    .Q_N(_07831_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][18] ));
 sg13g2_dfrbp_1 _18209_ (.CLK(net5558),
    .RESET_B(net6067),
    .D(_00772_),
    .Q_N(_07832_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_dfrbp_1 _18210_ (.CLK(net5558),
    .RESET_B(net6067),
    .D(_00782_),
    .Q_N(_07833_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_dfrbp_1 _18211_ (.CLK(net5557),
    .RESET_B(net6066),
    .D(_00783_),
    .Q_N(_07834_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_dfrbp_1 _18212_ (.CLK(net5560),
    .RESET_B(net6069),
    .D(_00784_),
    .Q_N(_07835_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_dfrbp_1 _18213_ (.CLK(net5560),
    .RESET_B(net6069),
    .D(_00785_),
    .Q_N(_07836_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_dfrbp_1 _18214_ (.CLK(net5560),
    .RESET_B(net6069),
    .D(_00786_),
    .Q_N(_07837_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_dfrbp_1 _18215_ (.CLK(net5557),
    .RESET_B(net6066),
    .D(_00787_),
    .Q_N(_07838_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_dfrbp_1 _18216_ (.CLK(net5557),
    .RESET_B(net6066),
    .D(_00788_),
    .Q_N(_07839_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_dfrbp_1 _18217_ (.CLK(net5559),
    .RESET_B(net6068),
    .D(_00789_),
    .Q_N(_07840_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_dfrbp_1 _18218_ (.CLK(net5490),
    .RESET_B(net5999),
    .D(_00790_),
    .Q_N(_07841_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_dfrbp_1 _18219_ (.CLK(net5490),
    .RESET_B(net5999),
    .D(_00773_),
    .Q_N(_07842_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_dfrbp_1 _18220_ (.CLK(net5489),
    .RESET_B(net5998),
    .D(_00774_),
    .Q_N(_07843_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_dfrbp_1 _18221_ (.CLK(net5489),
    .RESET_B(net5998),
    .D(_00775_),
    .Q_N(_07844_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_dfrbp_1 _18222_ (.CLK(net5486),
    .RESET_B(net5995),
    .D(_00776_),
    .Q_N(_07845_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_dfrbp_1 _18223_ (.CLK(net5486),
    .RESET_B(net5995),
    .D(_00777_),
    .Q_N(_07846_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_dfrbp_1 _18224_ (.CLK(net5485),
    .RESET_B(net5994),
    .D(_00778_),
    .Q_N(_07847_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_dfrbp_1 _18225_ (.CLK(net5485),
    .RESET_B(net5994),
    .D(_00779_),
    .Q_N(_07848_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[16] ));
 sg13g2_dfrbp_1 _18226_ (.CLK(net5485),
    .RESET_B(net5994),
    .D(_00780_),
    .Q_N(_07849_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_dfrbp_1 _18227_ (.CLK(net5485),
    .RESET_B(net5994),
    .D(_00781_),
    .Q_N(_07850_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.u2.reg_value[18] ));
 sg13g2_dfrbp_1 _18228_ (.CLK(net5558),
    .RESET_B(net6067),
    .D(_00772_),
    .Q_N(_07851_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_dfrbp_1 _18229_ (.CLK(net5558),
    .RESET_B(net6067),
    .D(_00782_),
    .Q_N(_07852_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_dfrbp_1 _18230_ (.CLK(net5560),
    .RESET_B(net6069),
    .D(_00783_),
    .Q_N(_07853_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_dfrbp_1 _18231_ (.CLK(net5560),
    .RESET_B(net6069),
    .D(_00784_),
    .Q_N(_07854_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_dfrbp_1 _18232_ (.CLK(net5562),
    .RESET_B(net6070),
    .D(_00785_),
    .Q_N(_07855_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_dfrbp_1 _18233_ (.CLK(net5562),
    .RESET_B(net6071),
    .D(_00786_),
    .Q_N(_07856_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_dfrbp_1 _18234_ (.CLK(net5562),
    .RESET_B(net6071),
    .D(_00787_),
    .Q_N(_07857_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_dfrbp_1 _18235_ (.CLK(net5560),
    .RESET_B(net6069),
    .D(_00788_),
    .Q_N(_07858_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_dfrbp_1 _18236_ (.CLK(net5557),
    .RESET_B(net6066),
    .D(_00789_),
    .Q_N(_07859_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_dfrbp_1 _18237_ (.CLK(net5559),
    .RESET_B(net6068),
    .D(_00790_),
    .Q_N(_07860_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_dfrbp_1 _18238_ (.CLK(net5490),
    .RESET_B(net5999),
    .D(_00773_),
    .Q_N(_07861_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_dfrbp_1 _18239_ (.CLK(net5490),
    .RESET_B(net5999),
    .D(_00774_),
    .Q_N(_07862_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_dfrbp_1 _18240_ (.CLK(net5489),
    .RESET_B(net5998),
    .D(_00775_),
    .Q_N(_07863_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_dfrbp_1 _18241_ (.CLK(net5489),
    .RESET_B(net5998),
    .D(_00776_),
    .Q_N(_07864_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_dfrbp_1 _18242_ (.CLK(net5485),
    .RESET_B(net5994),
    .D(_00777_),
    .Q_N(_07865_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_dfrbp_1 _18243_ (.CLK(net5485),
    .RESET_B(net5994),
    .D(_00778_),
    .Q_N(_07866_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_dfrbp_1 _18244_ (.CLK(net5487),
    .RESET_B(net5996),
    .D(_00779_),
    .Q_N(_07867_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_dfrbp_1 _18245_ (.CLK(net5487),
    .RESET_B(net5996),
    .D(_00780_),
    .Q_N(_07868_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_dfrbp_1 _18246_ (.CLK(net5485),
    .RESET_B(net5994),
    .D(_00781_),
    .Q_N(_07869_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator2_out[18] ));
 sg13g2_dfrbp_1 _18247_ (.CLK(net5559),
    .RESET_B(net6068),
    .D(_01190_),
    .Q_N(_01190_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[0] ));
 sg13g2_dfrbp_1 _18248_ (.CLK(net5558),
    .RESET_B(net6067),
    .D(_00763_),
    .Q_N(_07870_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_dfrbp_1 _18249_ (.CLK(net5557),
    .RESET_B(net6066),
    .D(_00764_),
    .Q_N(_07871_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_dfrbp_1 _18250_ (.CLK(net5557),
    .RESET_B(net6066),
    .D(_00765_),
    .Q_N(_07872_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_dfrbp_1 _18251_ (.CLK(net5557),
    .RESET_B(net6066),
    .D(_00766_),
    .Q_N(_07873_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[4] ));
 sg13g2_dfrbp_1 _18252_ (.CLK(net5557),
    .RESET_B(net6066),
    .D(_00767_),
    .Q_N(_07874_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_dfrbp_1 _18253_ (.CLK(net5559),
    .RESET_B(net6068),
    .D(_00768_),
    .Q_N(_07875_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_dfrbp_1 _18254_ (.CLK(net5559),
    .RESET_B(net6068),
    .D(_00769_),
    .Q_N(_07876_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_dfrbp_1 _18255_ (.CLK(net5490),
    .RESET_B(net5999),
    .D(_00770_),
    .Q_N(_07877_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_dfrbp_1 _18256_ (.CLK(net5490),
    .RESET_B(net5999),
    .D(_00771_),
    .Q_N(_07878_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_dfrbp_1 _18257_ (.CLK(net5489),
    .RESET_B(net5998),
    .D(_00754_),
    .Q_N(_07879_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_dfrbp_1 _18258_ (.CLK(net5489),
    .RESET_B(net5998),
    .D(_00755_),
    .Q_N(_07880_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_dfrbp_1 _18259_ (.CLK(net5489),
    .RESET_B(net5998),
    .D(_00756_),
    .Q_N(_07881_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_dfrbp_1 _18260_ (.CLK(net5486),
    .RESET_B(net5995),
    .D(_00757_),
    .Q_N(_07882_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_dfrbp_1 _18261_ (.CLK(net5486),
    .RESET_B(net5995),
    .D(_00758_),
    .Q_N(_07883_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_dfrbp_1 _18262_ (.CLK(net5486),
    .RESET_B(net5995),
    .D(_00759_),
    .Q_N(_07884_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_dfrbp_1 _18263_ (.CLK(net5486),
    .RESET_B(net5995),
    .D(_00760_),
    .Q_N(_07885_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_dfrbp_1 _18264_ (.CLK(net5486),
    .RESET_B(net5995),
    .D(_00761_),
    .Q_N(_07886_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_dfrbp_1 _18265_ (.CLK(net5485),
    .RESET_B(net5994),
    .D(_00762_),
    .Q_N(_07887_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.u_top_module.integrator1_out[18] ));
 sg13g2_dfrbp_1 _18266_ (.CLK(net5143),
    .RESET_B(net636),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][0] ),
    .Q_N(_07888_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18267_ (.CLK(net5143),
    .RESET_B(net637),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][1] ),
    .Q_N(_07889_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18268_ (.CLK(net5146),
    .RESET_B(net638),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][2] ),
    .Q_N(_07890_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18269_ (.CLK(net5146),
    .RESET_B(net639),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][3] ),
    .Q_N(_07891_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18270_ (.CLK(net5148),
    .RESET_B(net640),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][4] ),
    .Q_N(_07892_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18271_ (.CLK(net5149),
    .RESET_B(net641),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][5] ),
    .Q_N(_07893_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18272_ (.CLK(net5149),
    .RESET_B(net642),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][6] ),
    .Q_N(_07894_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18273_ (.CLK(net5149),
    .RESET_B(net643),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][7] ),
    .Q_N(_07895_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18274_ (.CLK(net5148),
    .RESET_B(net644),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][8] ),
    .Q_N(_07896_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18275_ (.CLK(net5147),
    .RESET_B(net645),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][9] ),
    .Q_N(_07897_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18276_ (.CLK(net5143),
    .RESET_B(net646),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][10] ),
    .Q_N(_07898_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18277_ (.CLK(net5144),
    .RESET_B(net647),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][11] ),
    .Q_N(_07899_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18278_ (.CLK(net5135),
    .RESET_B(net648),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][12] ),
    .Q_N(_07900_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18279_ (.CLK(net5135),
    .RESET_B(net649),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][13] ),
    .Q_N(_07901_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18280_ (.CLK(net5135),
    .RESET_B(net650),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][14] ),
    .Q_N(_07902_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18281_ (.CLK(net5134),
    .RESET_B(net651),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][15] ),
    .Q_N(_07903_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18282_ (.CLK(net5134),
    .RESET_B(net652),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][16] ),
    .Q_N(_07904_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18283_ (.CLK(net5138),
    .RESET_B(net653),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][17] ),
    .Q_N(_07905_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18284_ (.CLK(net5134),
    .RESET_B(net654),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[0][18] ),
    .Q_N(_07906_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18285_ (.CLK(net5142),
    .RESET_B(net655),
    .D(_00716_),
    .Q_N(_07907_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][0] ));
 sg13g2_dfrbp_1 _18286_ (.CLK(net5142),
    .RESET_B(net656),
    .D(_00726_),
    .Q_N(_07908_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][1] ));
 sg13g2_dfrbp_1 _18287_ (.CLK(net5143),
    .RESET_B(net657),
    .D(_00727_),
    .Q_N(_07909_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][2] ));
 sg13g2_dfrbp_1 _18288_ (.CLK(net5146),
    .RESET_B(net658),
    .D(_00728_),
    .Q_N(_07910_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][3] ));
 sg13g2_dfrbp_1 _18289_ (.CLK(net5148),
    .RESET_B(net659),
    .D(_00729_),
    .Q_N(_07911_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][4] ));
 sg13g2_dfrbp_1 _18290_ (.CLK(net5154),
    .RESET_B(net660),
    .D(_00730_),
    .Q_N(_07912_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][5] ));
 sg13g2_dfrbp_1 _18291_ (.CLK(net5154),
    .RESET_B(net661),
    .D(_00731_),
    .Q_N(_07913_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][6] ));
 sg13g2_dfrbp_1 _18292_ (.CLK(net5154),
    .RESET_B(net662),
    .D(_00732_),
    .Q_N(_07914_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][7] ));
 sg13g2_dfrbp_1 _18293_ (.CLK(net5155),
    .RESET_B(net663),
    .D(_00733_),
    .Q_N(_07915_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][8] ));
 sg13g2_dfrbp_1 _18294_ (.CLK(net5148),
    .RESET_B(net664),
    .D(_00734_),
    .Q_N(_07916_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][9] ));
 sg13g2_dfrbp_1 _18295_ (.CLK(net5147),
    .RESET_B(net665),
    .D(_00717_),
    .Q_N(_07917_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][10] ));
 sg13g2_dfrbp_1 _18296_ (.CLK(net5143),
    .RESET_B(net666),
    .D(_00718_),
    .Q_N(_07918_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][11] ));
 sg13g2_dfrbp_1 _18297_ (.CLK(net5141),
    .RESET_B(net667),
    .D(_00719_),
    .Q_N(_07919_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][12] ));
 sg13g2_dfrbp_1 _18298_ (.CLK(net5141),
    .RESET_B(net668),
    .D(_00720_),
    .Q_N(_07920_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][13] ));
 sg13g2_dfrbp_1 _18299_ (.CLK(net5137),
    .RESET_B(net669),
    .D(_00721_),
    .Q_N(_07921_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][14] ));
 sg13g2_dfrbp_1 _18300_ (.CLK(net5136),
    .RESET_B(net670),
    .D(_00722_),
    .Q_N(_07922_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][15] ));
 sg13g2_dfrbp_1 _18301_ (.CLK(net5136),
    .RESET_B(net671),
    .D(_00723_),
    .Q_N(_07923_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][16] ));
 sg13g2_dfrbp_1 _18302_ (.CLK(net5130),
    .RESET_B(net672),
    .D(_00724_),
    .Q_N(_07924_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][17] ));
 sg13g2_dfrbp_1 _18303_ (.CLK(net5130),
    .RESET_B(net179),
    .D(_00725_),
    .Q_N(_06440_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][18] ));
 sg13g2_dfrbp_1 _18304_ (.CLK(_01610_),
    .RESET_B(net178),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[0] ),
    .Q_N(_06439_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18305_ (.CLK(_01611_),
    .RESET_B(net177),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[1] ),
    .Q_N(_06438_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18306_ (.CLK(_01612_),
    .RESET_B(net176),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[2] ),
    .Q_N(_06437_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18307_ (.CLK(_01613_),
    .RESET_B(net175),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[3] ),
    .Q_N(_06436_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18308_ (.CLK(_01614_),
    .RESET_B(net174),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[4] ),
    .Q_N(_06435_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18309_ (.CLK(_01615_),
    .RESET_B(net173),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[5] ),
    .Q_N(_06434_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18310_ (.CLK(_01616_),
    .RESET_B(net172),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[6] ),
    .Q_N(_06433_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18311_ (.CLK(_01617_),
    .RESET_B(net171),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[7] ),
    .Q_N(_06432_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18312_ (.CLK(_01618_),
    .RESET_B(net170),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[8] ),
    .Q_N(_06431_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18313_ (.CLK(_01619_),
    .RESET_B(net169),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[9] ),
    .Q_N(_06430_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18314_ (.CLK(_01620_),
    .RESET_B(net168),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[10] ),
    .Q_N(_06429_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18315_ (.CLK(_01621_),
    .RESET_B(net167),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[11] ),
    .Q_N(_06428_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _18316_ (.CLK(_01622_),
    .RESET_B(net166),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[12] ),
    .Q_N(_06427_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _18317_ (.CLK(_01623_),
    .RESET_B(net165),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[13] ),
    .Q_N(_06426_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _18318_ (.CLK(_01624_),
    .RESET_B(net164),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[14] ),
    .Q_N(_06425_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _18319_ (.CLK(_01625_),
    .RESET_B(net163),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[15] ),
    .Q_N(_06424_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _18320_ (.CLK(_01626_),
    .RESET_B(net162),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[16] ),
    .Q_N(_06423_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _18321_ (.CLK(_01627_),
    .RESET_B(net161),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[17] ),
    .Q_N(_06422_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _18322_ (.CLK(_01628_),
    .RESET_B(net673),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.temp_delay[18] ),
    .Q_N(_07925_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[1].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _18323_ (.CLK(net5141),
    .RESET_B(net674),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][0] ),
    .Q_N(_07926_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18324_ (.CLK(net5142),
    .RESET_B(net675),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][1] ),
    .Q_N(_07927_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18325_ (.CLK(net5142),
    .RESET_B(net676),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][2] ),
    .Q_N(_07928_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18326_ (.CLK(net5146),
    .RESET_B(net677),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][3] ),
    .Q_N(_07929_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18327_ (.CLK(net5148),
    .RESET_B(net678),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][4] ),
    .Q_N(_07930_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18328_ (.CLK(net5154),
    .RESET_B(net679),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][5] ),
    .Q_N(_07931_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18329_ (.CLK(net5155),
    .RESET_B(net680),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][6] ),
    .Q_N(_07932_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18330_ (.CLK(net5155),
    .RESET_B(net681),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][7] ),
    .Q_N(_07933_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18331_ (.CLK(net5154),
    .RESET_B(net682),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][8] ),
    .Q_N(_07934_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18332_ (.CLK(net5150),
    .RESET_B(net683),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][9] ),
    .Q_N(_07935_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18333_ (.CLK(net5153),
    .RESET_B(net684),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][10] ),
    .Q_N(_07936_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18334_ (.CLK(net5147),
    .RESET_B(net685),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][11] ),
    .Q_N(_07937_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18335_ (.CLK(net5141),
    .RESET_B(net686),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][12] ),
    .Q_N(_07938_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18336_ (.CLK(net5145),
    .RESET_B(net687),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][13] ),
    .Q_N(_07939_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18337_ (.CLK(net5137),
    .RESET_B(net688),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][14] ),
    .Q_N(_07940_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18338_ (.CLK(net5136),
    .RESET_B(net689),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][15] ),
    .Q_N(_07941_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18339_ (.CLK(net5136),
    .RESET_B(net690),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][16] ),
    .Q_N(_07942_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18340_ (.CLK(net5133),
    .RESET_B(net691),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][17] ),
    .Q_N(_07943_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18341_ (.CLK(net5130),
    .RESET_B(net692),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.comb_data[1][18] ),
    .Q_N(_07944_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18342_ (.CLK(net5141),
    .RESET_B(net693),
    .D(_00735_),
    .Q_N(_07945_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18343_ (.CLK(net5141),
    .RESET_B(net694),
    .D(_00745_),
    .Q_N(_07946_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18344_ (.CLK(net5141),
    .RESET_B(net695),
    .D(_00746_),
    .Q_N(_07947_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18345_ (.CLK(net5142),
    .RESET_B(net696),
    .D(_00747_),
    .Q_N(_07948_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18346_ (.CLK(net5147),
    .RESET_B(net697),
    .D(_00748_),
    .Q_N(_07949_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18347_ (.CLK(net5150),
    .RESET_B(net698),
    .D(_00749_),
    .Q_N(_07950_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18348_ (.CLK(net5156),
    .RESET_B(net699),
    .D(_00750_),
    .Q_N(_07951_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18349_ (.CLK(net5156),
    .RESET_B(net700),
    .D(_00751_),
    .Q_N(_07952_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18350_ (.CLK(net5156),
    .RESET_B(net701),
    .D(_00752_),
    .Q_N(_07953_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18351_ (.CLK(net5150),
    .RESET_B(net702),
    .D(_00753_),
    .Q_N(_07954_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18352_ (.CLK(net5150),
    .RESET_B(net703),
    .D(_00736_),
    .Q_N(_07955_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18353_ (.CLK(net5153),
    .RESET_B(net704),
    .D(_00737_),
    .Q_N(_07956_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18354_ (.CLK(net5145),
    .RESET_B(net705),
    .D(_00738_),
    .Q_N(_07957_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18355_ (.CLK(net5145),
    .RESET_B(net706),
    .D(_00739_),
    .Q_N(_07958_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18356_ (.CLK(net5145),
    .RESET_B(net707),
    .D(_00740_),
    .Q_N(_07959_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18357_ (.CLK(net5136),
    .RESET_B(net708),
    .D(_00741_),
    .Q_N(_07960_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18358_ (.CLK(net5133),
    .RESET_B(net709),
    .D(_00742_),
    .Q_N(_07961_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18359_ (.CLK(net5133),
    .RESET_B(net710),
    .D(_00743_),
    .Q_N(_07962_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18360_ (.CLK(net5131),
    .RESET_B(net160),
    .D(_00744_),
    .Q_N(_06421_),
    .Q(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18361_ (.CLK(_01629_),
    .RESET_B(net159),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[0] ),
    .Q_N(_06420_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18362_ (.CLK(_01630_),
    .RESET_B(net158),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[1] ),
    .Q_N(_06419_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18363_ (.CLK(_01631_),
    .RESET_B(net157),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[2] ),
    .Q_N(_06418_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18364_ (.CLK(_01632_),
    .RESET_B(net156),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[3] ),
    .Q_N(_06417_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18365_ (.CLK(_01633_),
    .RESET_B(net155),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[4] ),
    .Q_N(_06416_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18366_ (.CLK(_01634_),
    .RESET_B(net154),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[5] ),
    .Q_N(_06415_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18367_ (.CLK(_01635_),
    .RESET_B(net153),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[6] ),
    .Q_N(_06414_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18368_ (.CLK(_01636_),
    .RESET_B(net152),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[7] ),
    .Q_N(_06413_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18369_ (.CLK(_01637_),
    .RESET_B(net151),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[8] ),
    .Q_N(_06412_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18370_ (.CLK(_01638_),
    .RESET_B(net150),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[9] ),
    .Q_N(_06411_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18371_ (.CLK(_01639_),
    .RESET_B(net149),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[10] ),
    .Q_N(_06410_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18372_ (.CLK(_01640_),
    .RESET_B(net148),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[11] ),
    .Q_N(_06409_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _18373_ (.CLK(_01641_),
    .RESET_B(net147),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[12] ),
    .Q_N(_06408_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _18374_ (.CLK(_01642_),
    .RESET_B(net146),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[13] ),
    .Q_N(_06407_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _18375_ (.CLK(_01643_),
    .RESET_B(net145),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[14] ),
    .Q_N(_06406_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _18376_ (.CLK(_01644_),
    .RESET_B(net144),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[15] ),
    .Q_N(_06405_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _18377_ (.CLK(_01645_),
    .RESET_B(net143),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[16] ),
    .Q_N(_06404_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _18378_ (.CLK(_01646_),
    .RESET_B(net142),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[17] ),
    .Q_N(_06403_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _18379_ (.CLK(_01647_),
    .RESET_B(net711),
    .D(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.temp_delay[18] ),
    .Q_N(_07963_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.genblk1[2].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _18380_ (.CLK(net5436),
    .RESET_B(net5945),
    .D(_00697_),
    .Q_N(_07964_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_dfrbp_1 _18381_ (.CLK(net5430),
    .RESET_B(net5939),
    .D(_00707_),
    .Q_N(_07965_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_dfrbp_1 _18382_ (.CLK(net5476),
    .RESET_B(net5985),
    .D(_00708_),
    .Q_N(_07966_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_dfrbp_1 _18383_ (.CLK(net5477),
    .RESET_B(net5986),
    .D(_00709_),
    .Q_N(_07967_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_dfrbp_1 _18384_ (.CLK(net5477),
    .RESET_B(net5986),
    .D(_00710_),
    .Q_N(_07968_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_dfrbp_1 _18385_ (.CLK(net5477),
    .RESET_B(net5986),
    .D(_00711_),
    .Q_N(_07969_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_dfrbp_1 _18386_ (.CLK(net5477),
    .RESET_B(net5986),
    .D(_00712_),
    .Q_N(_07970_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_dfrbp_1 _18387_ (.CLK(net5430),
    .RESET_B(net5939),
    .D(_00713_),
    .Q_N(_07971_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_dfrbp_1 _18388_ (.CLK(net5429),
    .RESET_B(net5938),
    .D(_00714_),
    .Q_N(_07972_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_dfrbp_1 _18389_ (.CLK(net5433),
    .RESET_B(net5947),
    .D(_00715_),
    .Q_N(_07973_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_dfrbp_1 _18390_ (.CLK(net5438),
    .RESET_B(net5942),
    .D(_00698_),
    .Q_N(_07974_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_dfrbp_1 _18391_ (.CLK(net5433),
    .RESET_B(net5942),
    .D(_00699_),
    .Q_N(_07975_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_dfrbp_1 _18392_ (.CLK(net5433),
    .RESET_B(net5942),
    .D(_00700_),
    .Q_N(_07976_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_dfrbp_1 _18393_ (.CLK(net5423),
    .RESET_B(net5932),
    .D(_00701_),
    .Q_N(_07977_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_dfrbp_1 _18394_ (.CLK(net5423),
    .RESET_B(net5933),
    .D(_00702_),
    .Q_N(_07978_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_dfrbp_1 _18395_ (.CLK(net5424),
    .RESET_B(net5932),
    .D(_00703_),
    .Q_N(_07979_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_dfrbp_1 _18396_ (.CLK(net5424),
    .RESET_B(net5933),
    .D(_00704_),
    .Q_N(_07980_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_dfrbp_1 _18397_ (.CLK(net5424),
    .RESET_B(net5933),
    .D(_00705_),
    .Q_N(_07981_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_dfrbp_1 _18398_ (.CLK(net5421),
    .RESET_B(net5930),
    .D(_00706_),
    .Q_N(_07982_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u3.reg_value[18] ));
 sg13g2_dfrbp_1 _18399_ (.CLK(net5436),
    .RESET_B(net5945),
    .D(_00697_),
    .Q_N(_07983_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][0] ));
 sg13g2_dfrbp_1 _18400_ (.CLK(net5436),
    .RESET_B(net5945),
    .D(_00707_),
    .Q_N(_07984_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][1] ));
 sg13g2_dfrbp_1 _18401_ (.CLK(net5480),
    .RESET_B(net5989),
    .D(_00708_),
    .Q_N(_07985_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][2] ));
 sg13g2_dfrbp_1 _18402_ (.CLK(net5476),
    .RESET_B(net5985),
    .D(_00709_),
    .Q_N(_07986_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][3] ));
 sg13g2_dfrbp_1 _18403_ (.CLK(net5477),
    .RESET_B(net5986),
    .D(_00710_),
    .Q_N(_07987_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][4] ));
 sg13g2_dfrbp_1 _18404_ (.CLK(net5477),
    .RESET_B(net5986),
    .D(_00711_),
    .Q_N(_07988_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][5] ));
 sg13g2_dfrbp_1 _18405_ (.CLK(net5477),
    .RESET_B(net5986),
    .D(_00712_),
    .Q_N(_07989_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][6] ));
 sg13g2_dfrbp_1 _18406_ (.CLK(net5436),
    .RESET_B(net5945),
    .D(_00713_),
    .Q_N(_07990_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][7] ));
 sg13g2_dfrbp_1 _18407_ (.CLK(net5436),
    .RESET_B(net5945),
    .D(_00714_),
    .Q_N(_07991_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][8] ));
 sg13g2_dfrbp_1 _18408_ (.CLK(net5433),
    .RESET_B(net5942),
    .D(_00715_),
    .Q_N(_07992_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][9] ));
 sg13g2_dfrbp_1 _18409_ (.CLK(net5433),
    .RESET_B(net5942),
    .D(_00698_),
    .Q_N(_07993_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][10] ));
 sg13g2_dfrbp_1 _18410_ (.CLK(net5433),
    .RESET_B(net5942),
    .D(_00699_),
    .Q_N(_07994_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][11] ));
 sg13g2_dfrbp_1 _18411_ (.CLK(net5423),
    .RESET_B(net5932),
    .D(_00700_),
    .Q_N(_07995_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][12] ));
 sg13g2_dfrbp_1 _18412_ (.CLK(net5423),
    .RESET_B(net5932),
    .D(_00701_),
    .Q_N(_07996_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][13] ));
 sg13g2_dfrbp_1 _18413_ (.CLK(net5423),
    .RESET_B(net5932),
    .D(_00702_),
    .Q_N(_07997_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][14] ));
 sg13g2_dfrbp_1 _18414_ (.CLK(net5423),
    .RESET_B(net5932),
    .D(_00703_),
    .Q_N(_07998_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][15] ));
 sg13g2_dfrbp_1 _18415_ (.CLK(net5423),
    .RESET_B(net5932),
    .D(_00704_),
    .Q_N(_07999_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][16] ));
 sg13g2_dfrbp_1 _18416_ (.CLK(net5423),
    .RESET_B(net5932),
    .D(_00705_),
    .Q_N(_08000_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][17] ));
 sg13g2_dfrbp_1 _18417_ (.CLK(net5424),
    .RESET_B(net5933),
    .D(_00706_),
    .Q_N(_08001_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][18] ));
 sg13g2_dfrbp_1 _18418_ (.CLK(net5476),
    .RESET_B(net5985),
    .D(_00678_),
    .Q_N(_08002_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_dfrbp_1 _18419_ (.CLK(net5476),
    .RESET_B(net5985),
    .D(_00688_),
    .Q_N(_08003_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_dfrbp_1 _18420_ (.CLK(net5474),
    .RESET_B(net5983),
    .D(_00689_),
    .Q_N(_08004_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_dfrbp_1 _18421_ (.CLK(net5474),
    .RESET_B(net5983),
    .D(_00690_),
    .Q_N(_08005_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_dfrbp_1 _18422_ (.CLK(net5474),
    .RESET_B(net5983),
    .D(_00691_),
    .Q_N(_08006_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_dfrbp_1 _18423_ (.CLK(net5474),
    .RESET_B(net5984),
    .D(_00692_),
    .Q_N(_08007_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_dfrbp_1 _18424_ (.CLK(net5475),
    .RESET_B(net5984),
    .D(_00693_),
    .Q_N(_08008_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_dfrbp_1 _18425_ (.CLK(net5475),
    .RESET_B(net5984),
    .D(_00694_),
    .Q_N(_08009_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_dfrbp_1 _18426_ (.CLK(net5431),
    .RESET_B(net5940),
    .D(_00695_),
    .Q_N(_08010_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_dfrbp_1 _18427_ (.CLK(net5429),
    .RESET_B(net5938),
    .D(_00696_),
    .Q_N(_08011_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_dfrbp_1 _18428_ (.CLK(net5429),
    .RESET_B(net5938),
    .D(_00679_),
    .Q_N(_08012_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_dfrbp_1 _18429_ (.CLK(net5427),
    .RESET_B(net5936),
    .D(_00680_),
    .Q_N(_08013_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_dfrbp_1 _18430_ (.CLK(net5427),
    .RESET_B(net5936),
    .D(_00681_),
    .Q_N(_08014_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_dfrbp_1 _18431_ (.CLK(net5427),
    .RESET_B(net5936),
    .D(_00682_),
    .Q_N(_08015_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_dfrbp_1 _18432_ (.CLK(net5426),
    .RESET_B(net5935),
    .D(_00683_),
    .Q_N(_08016_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_dfrbp_1 _18433_ (.CLK(net5426),
    .RESET_B(net5935),
    .D(_00684_),
    .Q_N(_08017_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_dfrbp_1 _18434_ (.CLK(net5426),
    .RESET_B(net5935),
    .D(_00685_),
    .Q_N(_08018_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[16] ));
 sg13g2_dfrbp_1 _18435_ (.CLK(net5426),
    .RESET_B(net5935),
    .D(_00686_),
    .Q_N(_08019_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_dfrbp_1 _18436_ (.CLK(net5426),
    .RESET_B(net5935),
    .D(_00687_),
    .Q_N(_08020_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.u2.reg_value[18] ));
 sg13g2_dfrbp_1 _18437_ (.CLK(net5430),
    .RESET_B(net5939),
    .D(_00678_),
    .Q_N(_08021_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_dfrbp_1 _18438_ (.CLK(net5476),
    .RESET_B(net5985),
    .D(_00688_),
    .Q_N(_08022_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_dfrbp_1 _18439_ (.CLK(net5476),
    .RESET_B(net5985),
    .D(_00689_),
    .Q_N(_08023_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_dfrbp_1 _18440_ (.CLK(net5478),
    .RESET_B(net5987),
    .D(_00690_),
    .Q_N(_08024_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_dfrbp_1 _18441_ (.CLK(net5474),
    .RESET_B(net5983),
    .D(_00691_),
    .Q_N(_08025_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_dfrbp_1 _18442_ (.CLK(net5474),
    .RESET_B(net5983),
    .D(_00692_),
    .Q_N(_08026_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_dfrbp_1 _18443_ (.CLK(net5476),
    .RESET_B(net5985),
    .D(_00693_),
    .Q_N(_08027_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_dfrbp_1 _18444_ (.CLK(net5430),
    .RESET_B(net5939),
    .D(_00694_),
    .Q_N(_08028_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_dfrbp_1 _18445_ (.CLK(net5430),
    .RESET_B(net5939),
    .D(_00695_),
    .Q_N(_08029_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_dfrbp_1 _18446_ (.CLK(net5429),
    .RESET_B(net5938),
    .D(_00696_),
    .Q_N(_08030_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_dfrbp_1 _18447_ (.CLK(net5429),
    .RESET_B(net5938),
    .D(_00679_),
    .Q_N(_08031_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_dfrbp_1 _18448_ (.CLK(net5427),
    .RESET_B(net5936),
    .D(_00680_),
    .Q_N(_08032_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_dfrbp_1 _18449_ (.CLK(net5427),
    .RESET_B(net5936),
    .D(_00681_),
    .Q_N(_08033_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_dfrbp_1 _18450_ (.CLK(net5426),
    .RESET_B(net5935),
    .D(_00682_),
    .Q_N(_08034_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_dfrbp_1 _18451_ (.CLK(net5426),
    .RESET_B(net5935),
    .D(_00683_),
    .Q_N(_08035_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_dfrbp_1 _18452_ (.CLK(net5427),
    .RESET_B(net5936),
    .D(_00684_),
    .Q_N(_08036_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_dfrbp_1 _18453_ (.CLK(net5421),
    .RESET_B(net5930),
    .D(_00685_),
    .Q_N(_08037_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_dfrbp_1 _18454_ (.CLK(net5422),
    .RESET_B(net5931),
    .D(_00686_),
    .Q_N(_08038_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_dfrbp_1 _18455_ (.CLK(net5426),
    .RESET_B(net5935),
    .D(_00687_),
    .Q_N(_08039_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator2_out[18] ));
 sg13g2_dfrbp_1 _18456_ (.CLK(net5475),
    .RESET_B(net5984),
    .D(_01191_),
    .Q_N(_01191_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[0] ));
 sg13g2_dfrbp_1 _18457_ (.CLK(net5475),
    .RESET_B(net5984),
    .D(_00669_),
    .Q_N(_08040_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_dfrbp_1 _18458_ (.CLK(net5475),
    .RESET_B(net5983),
    .D(_00670_),
    .Q_N(_08041_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_dfrbp_1 _18459_ (.CLK(net5478),
    .RESET_B(net5987),
    .D(_00671_),
    .Q_N(_08042_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_dfrbp_1 _18460_ (.CLK(net5474),
    .RESET_B(net5983),
    .D(_00672_),
    .Q_N(_08043_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[4] ));
 sg13g2_dfrbp_1 _18461_ (.CLK(net5474),
    .RESET_B(net5983),
    .D(_00673_),
    .Q_N(_08044_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_dfrbp_1 _18462_ (.CLK(net5475),
    .RESET_B(net5984),
    .D(_00674_),
    .Q_N(_08045_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_dfrbp_1 _18463_ (.CLK(net5475),
    .RESET_B(net5984),
    .D(_00675_),
    .Q_N(_08046_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_dfrbp_1 _18464_ (.CLK(net5431),
    .RESET_B(net5940),
    .D(_00676_),
    .Q_N(_08047_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_dfrbp_1 _18465_ (.CLK(net5431),
    .RESET_B(net5940),
    .D(_00677_),
    .Q_N(_08048_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_dfrbp_1 _18466_ (.CLK(net5431),
    .RESET_B(net5940),
    .D(_00660_),
    .Q_N(_08049_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_dfrbp_1 _18467_ (.CLK(net5431),
    .RESET_B(net5940),
    .D(_00661_),
    .Q_N(_08050_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_dfrbp_1 _18468_ (.CLK(net5428),
    .RESET_B(net5937),
    .D(_00662_),
    .Q_N(_08051_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_dfrbp_1 _18469_ (.CLK(net5428),
    .RESET_B(net5937),
    .D(_00663_),
    .Q_N(_08052_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_dfrbp_1 _18470_ (.CLK(net5428),
    .RESET_B(net5937),
    .D(_00664_),
    .Q_N(_08053_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_dfrbp_1 _18471_ (.CLK(net5428),
    .RESET_B(net5937),
    .D(_00665_),
    .Q_N(_08054_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_dfrbp_1 _18472_ (.CLK(net5428),
    .RESET_B(net5937),
    .D(_00666_),
    .Q_N(_08055_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_dfrbp_1 _18473_ (.CLK(net5428),
    .RESET_B(net5937),
    .D(_00667_),
    .Q_N(_08056_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_dfrbp_1 _18474_ (.CLK(net5428),
    .RESET_B(net5937),
    .D(_00668_),
    .Q_N(_08057_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.u_top_module.integrator1_out[18] ));
 sg13g2_dfrbp_1 _18475_ (.CLK(net5113),
    .RESET_B(net712),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][0] ),
    .Q_N(_08058_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18476_ (.CLK(net5115),
    .RESET_B(net713),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][1] ),
    .Q_N(_08059_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18477_ (.CLK(net5116),
    .RESET_B(net714),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][2] ),
    .Q_N(_08060_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18478_ (.CLK(net5131),
    .RESET_B(net715),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][3] ),
    .Q_N(_08061_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18479_ (.CLK(net5130),
    .RESET_B(net716),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][4] ),
    .Q_N(_08062_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18480_ (.CLK(net5130),
    .RESET_B(net717),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][5] ),
    .Q_N(_08063_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18481_ (.CLK(net5131),
    .RESET_B(net718),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][6] ),
    .Q_N(_08064_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18482_ (.CLK(net5116),
    .RESET_B(net719),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][7] ),
    .Q_N(_08065_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18483_ (.CLK(net5113),
    .RESET_B(net720),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][8] ),
    .Q_N(_08066_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18484_ (.CLK(net5112),
    .RESET_B(net721),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][9] ),
    .Q_N(_08067_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18485_ (.CLK(net5112),
    .RESET_B(net722),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][10] ),
    .Q_N(_08068_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18486_ (.CLK(net5108),
    .RESET_B(net723),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][11] ),
    .Q_N(_08069_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18487_ (.CLK(net5108),
    .RESET_B(net724),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][12] ),
    .Q_N(_08070_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18488_ (.CLK(net5109),
    .RESET_B(net725),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][13] ),
    .Q_N(_08071_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18489_ (.CLK(net5107),
    .RESET_B(net726),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][14] ),
    .Q_N(_08072_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18490_ (.CLK(net5111),
    .RESET_B(net727),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][15] ),
    .Q_N(_08073_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18491_ (.CLK(net5107),
    .RESET_B(net728),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][16] ),
    .Q_N(_08074_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18492_ (.CLK(net5108),
    .RESET_B(net729),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][17] ),
    .Q_N(_08075_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18493_ (.CLK(net5110),
    .RESET_B(net730),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[0][18] ),
    .Q_N(_08076_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18494_ (.CLK(net5126),
    .RESET_B(net731),
    .D(_00622_),
    .Q_N(_08077_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][0] ));
 sg13g2_dfrbp_1 _18495_ (.CLK(net5126),
    .RESET_B(net732),
    .D(_00632_),
    .Q_N(_08078_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][1] ));
 sg13g2_dfrbp_1 _18496_ (.CLK(net5116),
    .RESET_B(net733),
    .D(_00633_),
    .Q_N(_08079_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][2] ));
 sg13g2_dfrbp_1 _18497_ (.CLK(net5118),
    .RESET_B(net734),
    .D(_00634_),
    .Q_N(_08080_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][3] ));
 sg13g2_dfrbp_1 _18498_ (.CLK(net5132),
    .RESET_B(net735),
    .D(_00635_),
    .Q_N(_08081_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][4] ));
 sg13g2_dfrbp_1 _18499_ (.CLK(net5132),
    .RESET_B(net736),
    .D(_00636_),
    .Q_N(_08082_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][5] ));
 sg13g2_dfrbp_1 _18500_ (.CLK(net5132),
    .RESET_B(net737),
    .D(_00637_),
    .Q_N(_08083_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][6] ));
 sg13g2_dfrbp_1 _18501_ (.CLK(net5116),
    .RESET_B(net738),
    .D(_00638_),
    .Q_N(_08084_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][7] ));
 sg13g2_dfrbp_1 _18502_ (.CLK(net5114),
    .RESET_B(net739),
    .D(_00639_),
    .Q_N(_08085_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][8] ));
 sg13g2_dfrbp_1 _18503_ (.CLK(net5114),
    .RESET_B(net740),
    .D(_00640_),
    .Q_N(_08086_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][9] ));
 sg13g2_dfrbp_1 _18504_ (.CLK(net5120),
    .RESET_B(net741),
    .D(_00623_),
    .Q_N(_08087_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][10] ));
 sg13g2_dfrbp_1 _18505_ (.CLK(net5124),
    .RESET_B(net742),
    .D(_00624_),
    .Q_N(_08088_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][11] ));
 sg13g2_dfrbp_1 _18506_ (.CLK(net5121),
    .RESET_B(net743),
    .D(_00625_),
    .Q_N(_08089_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][12] ));
 sg13g2_dfrbp_1 _18507_ (.CLK(net5121),
    .RESET_B(net744),
    .D(_00626_),
    .Q_N(_08090_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][13] ));
 sg13g2_dfrbp_1 _18508_ (.CLK(net5121),
    .RESET_B(net745),
    .D(_00627_),
    .Q_N(_08091_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][14] ));
 sg13g2_dfrbp_1 _18509_ (.CLK(net5121),
    .RESET_B(net746),
    .D(_00628_),
    .Q_N(_08092_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][15] ));
 sg13g2_dfrbp_1 _18510_ (.CLK(net5119),
    .RESET_B(net747),
    .D(_00629_),
    .Q_N(_08093_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][16] ));
 sg13g2_dfrbp_1 _18511_ (.CLK(net5120),
    .RESET_B(net748),
    .D(_00630_),
    .Q_N(_08094_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][17] ));
 sg13g2_dfrbp_1 _18512_ (.CLK(net5110),
    .RESET_B(net141),
    .D(_00631_),
    .Q_N(_06402_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][18] ));
 sg13g2_dfrbp_1 _18513_ (.CLK(_01648_),
    .RESET_B(net140),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[0] ),
    .Q_N(_06401_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18514_ (.CLK(_01649_),
    .RESET_B(net139),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[1] ),
    .Q_N(_06400_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18515_ (.CLK(_01650_),
    .RESET_B(net138),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[2] ),
    .Q_N(_06399_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18516_ (.CLK(_01651_),
    .RESET_B(net137),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[3] ),
    .Q_N(_06398_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18517_ (.CLK(_01652_),
    .RESET_B(net136),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[4] ),
    .Q_N(_06397_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18518_ (.CLK(_01653_),
    .RESET_B(net135),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[5] ),
    .Q_N(_06396_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18519_ (.CLK(_01654_),
    .RESET_B(net134),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[6] ),
    .Q_N(_06395_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18520_ (.CLK(_01655_),
    .RESET_B(net133),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[7] ),
    .Q_N(_06394_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18521_ (.CLK(_01656_),
    .RESET_B(net132),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[8] ),
    .Q_N(_06393_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18522_ (.CLK(_01657_),
    .RESET_B(net131),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[9] ),
    .Q_N(_06392_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18523_ (.CLK(_01658_),
    .RESET_B(net130),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[10] ),
    .Q_N(_06391_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18524_ (.CLK(_01659_),
    .RESET_B(net129),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[11] ),
    .Q_N(_06390_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _18525_ (.CLK(_01660_),
    .RESET_B(net128),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[12] ),
    .Q_N(_06389_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _18526_ (.CLK(_01661_),
    .RESET_B(net127),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[13] ),
    .Q_N(_06388_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _18527_ (.CLK(_01662_),
    .RESET_B(net126),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[14] ),
    .Q_N(_06387_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _18528_ (.CLK(_01663_),
    .RESET_B(net125),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[15] ),
    .Q_N(_06386_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _18529_ (.CLK(_01664_),
    .RESET_B(net124),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[16] ),
    .Q_N(_06385_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _18530_ (.CLK(_01665_),
    .RESET_B(net123),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[17] ),
    .Q_N(_06384_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _18531_ (.CLK(_01666_),
    .RESET_B(net749),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.temp_delay[18] ),
    .Q_N(_08095_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[1].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _18532_ (.CLK(net5125),
    .RESET_B(net750),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][0] ),
    .Q_N(_08096_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18533_ (.CLK(net5125),
    .RESET_B(net751),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][1] ),
    .Q_N(_08097_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18534_ (.CLK(net5125),
    .RESET_B(net752),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][2] ),
    .Q_N(_08098_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18535_ (.CLK(net5127),
    .RESET_B(net753),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][3] ),
    .Q_N(_08099_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18536_ (.CLK(net5139),
    .RESET_B(net754),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][4] ),
    .Q_N(_08100_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18537_ (.CLK(net5139),
    .RESET_B(net755),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][5] ),
    .Q_N(_08101_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18538_ (.CLK(net5132),
    .RESET_B(net756),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][6] ),
    .Q_N(_08102_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18539_ (.CLK(net5127),
    .RESET_B(net757),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][7] ),
    .Q_N(_08103_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18540_ (.CLK(net5125),
    .RESET_B(net758),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][8] ),
    .Q_N(_08104_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18541_ (.CLK(net5119),
    .RESET_B(net759),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][9] ),
    .Q_N(_08105_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18542_ (.CLK(net5124),
    .RESET_B(net760),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][10] ),
    .Q_N(_08106_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18543_ (.CLK(net5121),
    .RESET_B(net761),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][11] ),
    .Q_N(_08107_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18544_ (.CLK(net5122),
    .RESET_B(net762),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][12] ),
    .Q_N(_08108_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18545_ (.CLK(net5123),
    .RESET_B(net763),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][13] ),
    .Q_N(_08109_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18546_ (.CLK(net5122),
    .RESET_B(net764),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][14] ),
    .Q_N(_08110_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18547_ (.CLK(net5122),
    .RESET_B(net765),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][15] ),
    .Q_N(_08111_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18548_ (.CLK(net5121),
    .RESET_B(net766),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][16] ),
    .Q_N(_08112_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18549_ (.CLK(net5119),
    .RESET_B(net767),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][17] ),
    .Q_N(_08113_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18550_ (.CLK(net5120),
    .RESET_B(net768),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.comb_data[1][18] ),
    .Q_N(_08114_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18551_ (.CLK(net5125),
    .RESET_B(net769),
    .D(_00641_),
    .Q_N(_08115_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18552_ (.CLK(net5128),
    .RESET_B(net770),
    .D(_00651_),
    .Q_N(_08116_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18553_ (.CLK(net5128),
    .RESET_B(net771),
    .D(_00652_),
    .Q_N(_08117_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18554_ (.CLK(net5140),
    .RESET_B(net772),
    .D(_00653_),
    .Q_N(_08118_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18555_ (.CLK(net5140),
    .RESET_B(net773),
    .D(_00654_),
    .Q_N(_08119_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18556_ (.CLK(net5139),
    .RESET_B(net774),
    .D(_00655_),
    .Q_N(_08120_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18557_ (.CLK(net5139),
    .RESET_B(net775),
    .D(_00656_),
    .Q_N(_08121_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18558_ (.CLK(net5139),
    .RESET_B(net776),
    .D(_00657_),
    .Q_N(_08122_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18559_ (.CLK(net5127),
    .RESET_B(net777),
    .D(_00658_),
    .Q_N(_08123_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18560_ (.CLK(net5128),
    .RESET_B(net778),
    .D(_00659_),
    .Q_N(_08124_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18561_ (.CLK(net5128),
    .RESET_B(net779),
    .D(_00642_),
    .Q_N(_08125_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18562_ (.CLK(net5124),
    .RESET_B(net780),
    .D(_00643_),
    .Q_N(_08126_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18563_ (.CLK(net5124),
    .RESET_B(net781),
    .D(_00644_),
    .Q_N(_08127_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18564_ (.CLK(net5124),
    .RESET_B(net782),
    .D(_00645_),
    .Q_N(_08128_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18565_ (.CLK(net5124),
    .RESET_B(net783),
    .D(_00646_),
    .Q_N(_08129_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18566_ (.CLK(net5123),
    .RESET_B(net784),
    .D(_00647_),
    .Q_N(_08130_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18567_ (.CLK(net5121),
    .RESET_B(net785),
    .D(_00648_),
    .Q_N(_08131_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18568_ (.CLK(net5119),
    .RESET_B(net786),
    .D(_00649_),
    .Q_N(_08132_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18569_ (.CLK(net5119),
    .RESET_B(net122),
    .D(_00650_),
    .Q_N(_06383_),
    .Q(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18570_ (.CLK(_01667_),
    .RESET_B(net120),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[0] ),
    .Q_N(_06382_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18571_ (.CLK(_01668_),
    .RESET_B(net119),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[1] ),
    .Q_N(_06381_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18572_ (.CLK(_01669_),
    .RESET_B(net118),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[2] ),
    .Q_N(_06380_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18573_ (.CLK(_01670_),
    .RESET_B(net117),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[3] ),
    .Q_N(_06379_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18574_ (.CLK(_01671_),
    .RESET_B(net116),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[4] ),
    .Q_N(_06378_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18575_ (.CLK(_01672_),
    .RESET_B(net115),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[5] ),
    .Q_N(_06377_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18576_ (.CLK(_01673_),
    .RESET_B(net114),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[6] ),
    .Q_N(_06376_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18577_ (.CLK(_01674_),
    .RESET_B(net113),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[7] ),
    .Q_N(_06375_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18578_ (.CLK(_01675_),
    .RESET_B(net112),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[8] ),
    .Q_N(_06374_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18579_ (.CLK(_01676_),
    .RESET_B(net111),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[9] ),
    .Q_N(_06373_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18580_ (.CLK(_01677_),
    .RESET_B(net110),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[10] ),
    .Q_N(_06372_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18581_ (.CLK(_01678_),
    .RESET_B(net109),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[11] ),
    .Q_N(_06371_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _18582_ (.CLK(_01679_),
    .RESET_B(net108),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[12] ),
    .Q_N(_06370_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _18583_ (.CLK(_01680_),
    .RESET_B(net107),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[13] ),
    .Q_N(_06369_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _18584_ (.CLK(_01681_),
    .RESET_B(net106),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[14] ),
    .Q_N(_06368_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _18585_ (.CLK(_01682_),
    .RESET_B(net105),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[15] ),
    .Q_N(_06367_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _18586_ (.CLK(_01683_),
    .RESET_B(net104),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[16] ),
    .Q_N(_06366_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _18587_ (.CLK(_01684_),
    .RESET_B(net103),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[17] ),
    .Q_N(_06365_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _18588_ (.CLK(_01685_),
    .RESET_B(net787),
    .D(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.temp_delay[18] ),
    .Q_N(_08133_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.genblk1[2].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _18589_ (.CLK(net5270),
    .RESET_B(net5780),
    .D(_00603_),
    .Q_N(_08134_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_dfrbp_1 _18590_ (.CLK(net5270),
    .RESET_B(net5780),
    .D(_00613_),
    .Q_N(_08135_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_dfrbp_1 _18591_ (.CLK(net5270),
    .RESET_B(net5780),
    .D(_00614_),
    .Q_N(_08136_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_dfrbp_1 _18592_ (.CLK(net5270),
    .RESET_B(net5780),
    .D(_00615_),
    .Q_N(_08137_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_dfrbp_1 _18593_ (.CLK(net5270),
    .RESET_B(net5780),
    .D(_00616_),
    .Q_N(_08138_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_dfrbp_1 _18594_ (.CLK(net5268),
    .RESET_B(net5778),
    .D(_00617_),
    .Q_N(_08139_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_dfrbp_1 _18595_ (.CLK(net5269),
    .RESET_B(net5779),
    .D(_00618_),
    .Q_N(_08140_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_dfrbp_1 _18596_ (.CLK(net5268),
    .RESET_B(net5778),
    .D(_00619_),
    .Q_N(_08141_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_dfrbp_1 _18597_ (.CLK(net5268),
    .RESET_B(net5778),
    .D(_00620_),
    .Q_N(_08142_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_dfrbp_1 _18598_ (.CLK(net5259),
    .RESET_B(net5769),
    .D(_00621_),
    .Q_N(_08143_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_dfrbp_1 _18599_ (.CLK(net5260),
    .RESET_B(net5770),
    .D(_00604_),
    .Q_N(_08144_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_dfrbp_1 _18600_ (.CLK(net5261),
    .RESET_B(net5771),
    .D(_00605_),
    .Q_N(_08145_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_dfrbp_1 _18601_ (.CLK(net5259),
    .RESET_B(net5769),
    .D(_00606_),
    .Q_N(_08146_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_dfrbp_1 _18602_ (.CLK(net5259),
    .RESET_B(net5769),
    .D(_00607_),
    .Q_N(_08147_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_dfrbp_1 _18603_ (.CLK(net5257),
    .RESET_B(net5767),
    .D(_00608_),
    .Q_N(_08148_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_dfrbp_1 _18604_ (.CLK(net5257),
    .RESET_B(net5767),
    .D(_00609_),
    .Q_N(_08149_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_dfrbp_1 _18605_ (.CLK(net5257),
    .RESET_B(net5767),
    .D(_00610_),
    .Q_N(_08150_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_dfrbp_1 _18606_ (.CLK(net5255),
    .RESET_B(net5765),
    .D(_00611_),
    .Q_N(_08151_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_dfrbp_1 _18607_ (.CLK(net5255),
    .RESET_B(net5765),
    .D(_00612_),
    .Q_N(_08152_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u3.reg_value[18] ));
 sg13g2_dfrbp_1 _18608_ (.CLK(net5271),
    .RESET_B(net5781),
    .D(_00603_),
    .Q_N(_08153_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][0] ));
 sg13g2_dfrbp_1 _18609_ (.CLK(net5271),
    .RESET_B(net5781),
    .D(_00613_),
    .Q_N(_08154_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][1] ));
 sg13g2_dfrbp_1 _18610_ (.CLK(net5271),
    .RESET_B(net5781),
    .D(_00614_),
    .Q_N(_08155_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][2] ));
 sg13g2_dfrbp_1 _18611_ (.CLK(net5271),
    .RESET_B(net5781),
    .D(_00615_),
    .Q_N(_08156_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][3] ));
 sg13g2_dfrbp_1 _18612_ (.CLK(net5270),
    .RESET_B(net5780),
    .D(_00616_),
    .Q_N(_08157_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][4] ));
 sg13g2_dfrbp_1 _18613_ (.CLK(net5270),
    .RESET_B(net5780),
    .D(_00617_),
    .Q_N(_08158_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][5] ));
 sg13g2_dfrbp_1 _18614_ (.CLK(net5270),
    .RESET_B(net5780),
    .D(_00618_),
    .Q_N(_08159_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][6] ));
 sg13g2_dfrbp_1 _18615_ (.CLK(net5268),
    .RESET_B(net5778),
    .D(_00619_),
    .Q_N(_08160_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][7] ));
 sg13g2_dfrbp_1 _18616_ (.CLK(net5268),
    .RESET_B(net5778),
    .D(_00620_),
    .Q_N(_08161_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][8] ));
 sg13g2_dfrbp_1 _18617_ (.CLK(net5268),
    .RESET_B(net5778),
    .D(_00621_),
    .Q_N(_08162_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][9] ));
 sg13g2_dfrbp_1 _18618_ (.CLK(net5261),
    .RESET_B(net5771),
    .D(_00604_),
    .Q_N(_08163_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][10] ));
 sg13g2_dfrbp_1 _18619_ (.CLK(net5259),
    .RESET_B(net5769),
    .D(_00605_),
    .Q_N(_08164_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][11] ));
 sg13g2_dfrbp_1 _18620_ (.CLK(net5259),
    .RESET_B(net5769),
    .D(_00606_),
    .Q_N(_08165_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][12] ));
 sg13g2_dfrbp_1 _18621_ (.CLK(net5259),
    .RESET_B(net5769),
    .D(_00607_),
    .Q_N(_08166_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][13] ));
 sg13g2_dfrbp_1 _18622_ (.CLK(net5260),
    .RESET_B(net5770),
    .D(_00608_),
    .Q_N(_08167_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][14] ));
 sg13g2_dfrbp_1 _18623_ (.CLK(net5258),
    .RESET_B(net5768),
    .D(_00609_),
    .Q_N(_08168_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][15] ));
 sg13g2_dfrbp_1 _18624_ (.CLK(net5257),
    .RESET_B(net5767),
    .D(_00610_),
    .Q_N(_08169_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][16] ));
 sg13g2_dfrbp_1 _18625_ (.CLK(net5257),
    .RESET_B(net5767),
    .D(_00611_),
    .Q_N(_08170_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][17] ));
 sg13g2_dfrbp_1 _18626_ (.CLK(net5255),
    .RESET_B(net5765),
    .D(_00612_),
    .Q_N(_08171_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][18] ));
 sg13g2_dfrbp_1 _18627_ (.CLK(net5272),
    .RESET_B(net5782),
    .D(_00584_),
    .Q_N(_08172_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_dfrbp_1 _18628_ (.CLK(net5272),
    .RESET_B(net5782),
    .D(_00594_),
    .Q_N(_08173_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_dfrbp_1 _18629_ (.CLK(net5272),
    .RESET_B(net5782),
    .D(_00595_),
    .Q_N(_08174_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_dfrbp_1 _18630_ (.CLK(net5273),
    .RESET_B(net5783),
    .D(_00596_),
    .Q_N(_08175_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_dfrbp_1 _18631_ (.CLK(net5273),
    .RESET_B(net5783),
    .D(_00597_),
    .Q_N(_08176_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_dfrbp_1 _18632_ (.CLK(net5273),
    .RESET_B(net5783),
    .D(_00598_),
    .Q_N(_08177_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_dfrbp_1 _18633_ (.CLK(net5266),
    .RESET_B(net5776),
    .D(_00599_),
    .Q_N(_08178_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_dfrbp_1 _18634_ (.CLK(net5266),
    .RESET_B(net5775),
    .D(_00600_),
    .Q_N(_08179_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_dfrbp_1 _18635_ (.CLK(net5265),
    .RESET_B(net5775),
    .D(_00601_),
    .Q_N(_08180_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_dfrbp_1 _18636_ (.CLK(net5265),
    .RESET_B(net5775),
    .D(_00602_),
    .Q_N(_08181_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_dfrbp_1 _18637_ (.CLK(net5263),
    .RESET_B(net5773),
    .D(_00585_),
    .Q_N(_08182_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_dfrbp_1 _18638_ (.CLK(net5262),
    .RESET_B(net5772),
    .D(_00586_),
    .Q_N(_08183_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_dfrbp_1 _18639_ (.CLK(net5263),
    .RESET_B(net5773),
    .D(_00587_),
    .Q_N(_08184_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_dfrbp_1 _18640_ (.CLK(net5256),
    .RESET_B(net5766),
    .D(_00588_),
    .Q_N(_08185_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_dfrbp_1 _18641_ (.CLK(net5256),
    .RESET_B(net5765),
    .D(_00589_),
    .Q_N(_08186_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_dfrbp_1 _18642_ (.CLK(net5255),
    .RESET_B(net5765),
    .D(_00590_),
    .Q_N(_08187_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_dfrbp_1 _18643_ (.CLK(net5256),
    .RESET_B(net5766),
    .D(_00591_),
    .Q_N(_08188_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[16] ));
 sg13g2_dfrbp_1 _18644_ (.CLK(net5217),
    .RESET_B(net5726),
    .D(_00592_),
    .Q_N(_08189_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_dfrbp_1 _18645_ (.CLK(net5220),
    .RESET_B(net5730),
    .D(_00593_),
    .Q_N(_08190_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.u2.reg_value[18] ));
 sg13g2_dfrbp_1 _18646_ (.CLK(net5272),
    .RESET_B(net5782),
    .D(_00584_),
    .Q_N(_08191_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_dfrbp_1 _18647_ (.CLK(net5272),
    .RESET_B(net5782),
    .D(_00594_),
    .Q_N(_08192_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_dfrbp_1 _18648_ (.CLK(net5272),
    .RESET_B(net5782),
    .D(_00595_),
    .Q_N(_08193_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_dfrbp_1 _18649_ (.CLK(net5272),
    .RESET_B(net5782),
    .D(_00596_),
    .Q_N(_08194_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_dfrbp_1 _18650_ (.CLK(net5272),
    .RESET_B(net5782),
    .D(_00597_),
    .Q_N(_08195_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_dfrbp_1 _18651_ (.CLK(net5268),
    .RESET_B(net5778),
    .D(_00598_),
    .Q_N(_08196_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_dfrbp_1 _18652_ (.CLK(net5268),
    .RESET_B(net5778),
    .D(_00599_),
    .Q_N(_08197_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_dfrbp_1 _18653_ (.CLK(net5265),
    .RESET_B(net5775),
    .D(_00600_),
    .Q_N(_08198_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_dfrbp_1 _18654_ (.CLK(net5265),
    .RESET_B(net5775),
    .D(_00601_),
    .Q_N(_08199_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_dfrbp_1 _18655_ (.CLK(net5265),
    .RESET_B(net5775),
    .D(_00602_),
    .Q_N(_08200_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_dfrbp_1 _18656_ (.CLK(net5259),
    .RESET_B(net5769),
    .D(_00585_),
    .Q_N(_08201_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_dfrbp_1 _18657_ (.CLK(net5259),
    .RESET_B(net5769),
    .D(_00586_),
    .Q_N(_08202_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_dfrbp_1 _18658_ (.CLK(net5257),
    .RESET_B(net5771),
    .D(_00587_),
    .Q_N(_08203_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_dfrbp_1 _18659_ (.CLK(net5261),
    .RESET_B(net5771),
    .D(_00588_),
    .Q_N(_08204_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_dfrbp_1 _18660_ (.CLK(net5261),
    .RESET_B(net5767),
    .D(_00589_),
    .Q_N(_08205_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_dfrbp_1 _18661_ (.CLK(net5255),
    .RESET_B(net5765),
    .D(_00590_),
    .Q_N(_08206_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_dfrbp_1 _18662_ (.CLK(net5256),
    .RESET_B(net5766),
    .D(_00591_),
    .Q_N(_08207_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_dfrbp_1 _18663_ (.CLK(net5255),
    .RESET_B(net5766),
    .D(_00592_),
    .Q_N(_08208_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_dfrbp_1 _18664_ (.CLK(net5217),
    .RESET_B(net5726),
    .D(_00593_),
    .Q_N(_08209_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator2_out[18] ));
 sg13g2_dfrbp_1 _18665_ (.CLK(net5273),
    .RESET_B(net5783),
    .D(_01192_),
    .Q_N(_01192_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[0] ));
 sg13g2_dfrbp_1 _18666_ (.CLK(net5273),
    .RESET_B(net5783),
    .D(_00575_),
    .Q_N(_08210_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_dfrbp_1 _18667_ (.CLK(net5273),
    .RESET_B(net5783),
    .D(_00576_),
    .Q_N(_08211_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_dfrbp_1 _18668_ (.CLK(net5273),
    .RESET_B(net5783),
    .D(_00577_),
    .Q_N(_08212_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_dfrbp_1 _18669_ (.CLK(net5266),
    .RESET_B(net5776),
    .D(_00578_),
    .Q_N(_08213_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[4] ));
 sg13g2_dfrbp_1 _18670_ (.CLK(net5265),
    .RESET_B(net5776),
    .D(_00579_),
    .Q_N(_08214_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_dfrbp_1 _18671_ (.CLK(net5266),
    .RESET_B(net5776),
    .D(_00580_),
    .Q_N(_08215_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_dfrbp_1 _18672_ (.CLK(net5266),
    .RESET_B(net5776),
    .D(_00581_),
    .Q_N(_08216_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_dfrbp_1 _18673_ (.CLK(net5265),
    .RESET_B(net5775),
    .D(_00582_),
    .Q_N(_08217_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_dfrbp_1 _18674_ (.CLK(net5265),
    .RESET_B(net5775),
    .D(_00583_),
    .Q_N(_08218_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_dfrbp_1 _18675_ (.CLK(net5263),
    .RESET_B(net5773),
    .D(_00566_),
    .Q_N(_08219_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_dfrbp_1 _18676_ (.CLK(net5263),
    .RESET_B(net5773),
    .D(_00567_),
    .Q_N(_08220_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_dfrbp_1 _18677_ (.CLK(net5262),
    .RESET_B(net5772),
    .D(_00568_),
    .Q_N(_08221_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_dfrbp_1 _18678_ (.CLK(net5262),
    .RESET_B(net5772),
    .D(_00569_),
    .Q_N(_08222_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_dfrbp_1 _18679_ (.CLK(net5262),
    .RESET_B(net5772),
    .D(_00570_),
    .Q_N(_08223_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_dfrbp_1 _18680_ (.CLK(net5262),
    .RESET_B(net5772),
    .D(_00571_),
    .Q_N(_08224_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_dfrbp_1 _18681_ (.CLK(net5262),
    .RESET_B(net5772),
    .D(_00572_),
    .Q_N(_08225_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_dfrbp_1 _18682_ (.CLK(net5220),
    .RESET_B(net5730),
    .D(_00573_),
    .Q_N(_08226_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_dfrbp_1 _18683_ (.CLK(net5220),
    .RESET_B(net5730),
    .D(_00574_),
    .Q_N(_08227_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.u_top_module.integrator1_out[18] ));
 sg13g2_dfrbp_1 _18684_ (.CLK(net5053),
    .RESET_B(net788),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][0] ),
    .Q_N(_08228_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18685_ (.CLK(net5052),
    .RESET_B(net789),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][1] ),
    .Q_N(_08229_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18686_ (.CLK(net5052),
    .RESET_B(net790),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][2] ),
    .Q_N(_08230_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18687_ (.CLK(net5052),
    .RESET_B(net791),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][3] ),
    .Q_N(_08231_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18688_ (.CLK(net5052),
    .RESET_B(net792),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][4] ),
    .Q_N(_08232_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18689_ (.CLK(net5050),
    .RESET_B(net793),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][5] ),
    .Q_N(_08233_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18690_ (.CLK(net5050),
    .RESET_B(net794),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][6] ),
    .Q_N(_08234_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18691_ (.CLK(net5049),
    .RESET_B(net795),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][7] ),
    .Q_N(_08235_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18692_ (.CLK(net5053),
    .RESET_B(net796),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][8] ),
    .Q_N(_08236_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18693_ (.CLK(net5048),
    .RESET_B(net797),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][9] ),
    .Q_N(_08237_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18694_ (.CLK(net5048),
    .RESET_B(net798),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][10] ),
    .Q_N(_08238_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18695_ (.CLK(net5048),
    .RESET_B(net799),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][11] ),
    .Q_N(_08239_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18696_ (.CLK(net5046),
    .RESET_B(net800),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][12] ),
    .Q_N(_08240_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18697_ (.CLK(net5046),
    .RESET_B(net801),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][13] ),
    .Q_N(_08241_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18698_ (.CLK(net5045),
    .RESET_B(net802),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][14] ),
    .Q_N(_08242_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18699_ (.CLK(net5045),
    .RESET_B(net803),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][15] ),
    .Q_N(_08243_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18700_ (.CLK(net5047),
    .RESET_B(net804),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][16] ),
    .Q_N(_08244_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18701_ (.CLK(net5047),
    .RESET_B(net805),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][17] ),
    .Q_N(_08245_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18702_ (.CLK(net5047),
    .RESET_B(net806),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[0][18] ),
    .Q_N(_08246_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18703_ (.CLK(net5070),
    .RESET_B(net807),
    .D(_00528_),
    .Q_N(_08247_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][0] ));
 sg13g2_dfrbp_1 _18704_ (.CLK(net5070),
    .RESET_B(net808),
    .D(_00538_),
    .Q_N(_08248_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][1] ));
 sg13g2_dfrbp_1 _18705_ (.CLK(net5070),
    .RESET_B(net809),
    .D(_00539_),
    .Q_N(_08249_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][2] ));
 sg13g2_dfrbp_1 _18706_ (.CLK(net5070),
    .RESET_B(net810),
    .D(_00540_),
    .Q_N(_08250_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][3] ));
 sg13g2_dfrbp_1 _18707_ (.CLK(net5068),
    .RESET_B(net811),
    .D(_00541_),
    .Q_N(_08251_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][4] ));
 sg13g2_dfrbp_1 _18708_ (.CLK(net5068),
    .RESET_B(net812),
    .D(_00542_),
    .Q_N(_08252_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][5] ));
 sg13g2_dfrbp_1 _18709_ (.CLK(net5068),
    .RESET_B(net813),
    .D(_00543_),
    .Q_N(_08253_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][6] ));
 sg13g2_dfrbp_1 _18710_ (.CLK(net5051),
    .RESET_B(net814),
    .D(_00544_),
    .Q_N(_08254_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][7] ));
 sg13g2_dfrbp_1 _18711_ (.CLK(net5051),
    .RESET_B(net815),
    .D(_00545_),
    .Q_N(_08255_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][8] ));
 sg13g2_dfrbp_1 _18712_ (.CLK(net5051),
    .RESET_B(net816),
    .D(_00546_),
    .Q_N(_08256_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][9] ));
 sg13g2_dfrbp_1 _18713_ (.CLK(net5050),
    .RESET_B(net817),
    .D(_00529_),
    .Q_N(_08257_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][10] ));
 sg13g2_dfrbp_1 _18714_ (.CLK(net5050),
    .RESET_B(net818),
    .D(_00530_),
    .Q_N(_08258_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][11] ));
 sg13g2_dfrbp_1 _18715_ (.CLK(net5050),
    .RESET_B(net819),
    .D(_00531_),
    .Q_N(_08259_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][12] ));
 sg13g2_dfrbp_1 _18716_ (.CLK(net5043),
    .RESET_B(net820),
    .D(_00532_),
    .Q_N(_08260_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][13] ));
 sg13g2_dfrbp_1 _18717_ (.CLK(net5043),
    .RESET_B(net821),
    .D(_00533_),
    .Q_N(_08261_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][14] ));
 sg13g2_dfrbp_1 _18718_ (.CLK(net5048),
    .RESET_B(net822),
    .D(_00534_),
    .Q_N(_08262_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][15] ));
 sg13g2_dfrbp_1 _18719_ (.CLK(net5048),
    .RESET_B(net823),
    .D(_00535_),
    .Q_N(_08263_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][16] ));
 sg13g2_dfrbp_1 _18720_ (.CLK(net5045),
    .RESET_B(net824),
    .D(_00536_),
    .Q_N(_08264_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][17] ));
 sg13g2_dfrbp_1 _18721_ (.CLK(net5045),
    .RESET_B(net102),
    .D(_00537_),
    .Q_N(_06364_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][18] ));
 sg13g2_dfrbp_1 _18722_ (.CLK(_01686_),
    .RESET_B(net101),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[0] ),
    .Q_N(_06363_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18723_ (.CLK(_01687_),
    .RESET_B(net100),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[1] ),
    .Q_N(_06362_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18724_ (.CLK(_01688_),
    .RESET_B(net99),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[2] ),
    .Q_N(_06361_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18725_ (.CLK(_01689_),
    .RESET_B(net98),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[3] ),
    .Q_N(_06360_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18726_ (.CLK(_01690_),
    .RESET_B(net97),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[4] ),
    .Q_N(_06359_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18727_ (.CLK(_01691_),
    .RESET_B(net96),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[5] ),
    .Q_N(_06358_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18728_ (.CLK(_01692_),
    .RESET_B(net95),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[6] ),
    .Q_N(_06357_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18729_ (.CLK(_01693_),
    .RESET_B(net94),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[7] ),
    .Q_N(_06356_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18730_ (.CLK(_01694_),
    .RESET_B(net93),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[8] ),
    .Q_N(_06355_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18731_ (.CLK(_01695_),
    .RESET_B(net92),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[9] ),
    .Q_N(_06354_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18732_ (.CLK(_01696_),
    .RESET_B(net91),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[10] ),
    .Q_N(_06353_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18733_ (.CLK(_01697_),
    .RESET_B(net90),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[11] ),
    .Q_N(_06352_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _18734_ (.CLK(_01698_),
    .RESET_B(net89),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[12] ),
    .Q_N(_06351_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _18735_ (.CLK(_01699_),
    .RESET_B(net88),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[13] ),
    .Q_N(_06350_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _18736_ (.CLK(_01700_),
    .RESET_B(net86),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[14] ),
    .Q_N(_06349_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _18737_ (.CLK(_01701_),
    .RESET_B(net85),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[15] ),
    .Q_N(_06348_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _18738_ (.CLK(_01702_),
    .RESET_B(net84),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[16] ),
    .Q_N(_06347_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _18739_ (.CLK(_01703_),
    .RESET_B(net83),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[17] ),
    .Q_N(_06346_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _18740_ (.CLK(_01704_),
    .RESET_B(net825),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.temp_delay[18] ),
    .Q_N(_08265_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[1].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _18741_ (.CLK(net5072),
    .RESET_B(net826),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][0] ),
    .Q_N(_08266_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18742_ (.CLK(net5072),
    .RESET_B(net827),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][1] ),
    .Q_N(_08267_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18743_ (.CLK(net5071),
    .RESET_B(net828),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][2] ),
    .Q_N(_08268_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18744_ (.CLK(net5071),
    .RESET_B(net829),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][3] ),
    .Q_N(_08269_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18745_ (.CLK(net5069),
    .RESET_B(net830),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][4] ),
    .Q_N(_08270_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18746_ (.CLK(net5069),
    .RESET_B(net831),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][5] ),
    .Q_N(_08271_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18747_ (.CLK(net5069),
    .RESET_B(net832),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][6] ),
    .Q_N(_08272_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18748_ (.CLK(net5068),
    .RESET_B(net833),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][7] ),
    .Q_N(_08273_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18749_ (.CLK(net5068),
    .RESET_B(net834),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][8] ),
    .Q_N(_08274_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18750_ (.CLK(net5051),
    .RESET_B(net835),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][9] ),
    .Q_N(_08275_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18751_ (.CLK(net5051),
    .RESET_B(net836),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][10] ),
    .Q_N(_08276_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18752_ (.CLK(net5042),
    .RESET_B(net837),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][11] ),
    .Q_N(_08277_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18753_ (.CLK(net5042),
    .RESET_B(net838),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][12] ),
    .Q_N(_08278_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18754_ (.CLK(net5043),
    .RESET_B(net839),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][13] ),
    .Q_N(_08279_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18755_ (.CLK(net5042),
    .RESET_B(net840),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][14] ),
    .Q_N(_08280_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18756_ (.CLK(net5042),
    .RESET_B(net841),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][15] ),
    .Q_N(_08281_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18757_ (.CLK(net5049),
    .RESET_B(net842),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][16] ),
    .Q_N(_08282_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18758_ (.CLK(net5048),
    .RESET_B(net843),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][17] ),
    .Q_N(_08283_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18759_ (.CLK(net5045),
    .RESET_B(net844),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.comb_data[1][18] ),
    .Q_N(_08284_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18760_ (.CLK(net5071),
    .RESET_B(net845),
    .D(_00547_),
    .Q_N(_08285_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18761_ (.CLK(net5079),
    .RESET_B(net846),
    .D(_00557_),
    .Q_N(_08286_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18762_ (.CLK(net5079),
    .RESET_B(net847),
    .D(_00558_),
    .Q_N(_08287_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18763_ (.CLK(net5071),
    .RESET_B(net848),
    .D(_00559_),
    .Q_N(_08288_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18764_ (.CLK(net5074),
    .RESET_B(net849),
    .D(_00560_),
    .Q_N(_08289_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18765_ (.CLK(net5071),
    .RESET_B(net850),
    .D(_00561_),
    .Q_N(_08290_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18766_ (.CLK(net5062),
    .RESET_B(net851),
    .D(_00562_),
    .Q_N(_08291_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18767_ (.CLK(net5062),
    .RESET_B(net852),
    .D(_00563_),
    .Q_N(_08292_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18768_ (.CLK(net5062),
    .RESET_B(net853),
    .D(_00564_),
    .Q_N(_08293_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18769_ (.CLK(net5062),
    .RESET_B(net854),
    .D(_00565_),
    .Q_N(_08294_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18770_ (.CLK(net5062),
    .RESET_B(net855),
    .D(_00548_),
    .Q_N(_08295_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18771_ (.CLK(net5061),
    .RESET_B(net856),
    .D(_00549_),
    .Q_N(_08296_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18772_ (.CLK(net5061),
    .RESET_B(net857),
    .D(_00550_),
    .Q_N(_08297_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18773_ (.CLK(net5061),
    .RESET_B(net858),
    .D(_00551_),
    .Q_N(_08298_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18774_ (.CLK(net5061),
    .RESET_B(net859),
    .D(_00552_),
    .Q_N(_08299_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18775_ (.CLK(net5061),
    .RESET_B(net860),
    .D(_00553_),
    .Q_N(_08300_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18776_ (.CLK(net5061),
    .RESET_B(net861),
    .D(_00554_),
    .Q_N(_08301_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18777_ (.CLK(net5042),
    .RESET_B(net862),
    .D(_00555_),
    .Q_N(_08302_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18778_ (.CLK(net5048),
    .RESET_B(net82),
    .D(_00556_),
    .Q_N(_06345_),
    .Q(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18779_ (.CLK(_01705_),
    .RESET_B(net81),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[0] ),
    .Q_N(_06344_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18780_ (.CLK(_01706_),
    .RESET_B(net80),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[1] ),
    .Q_N(_06343_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18781_ (.CLK(_01707_),
    .RESET_B(net79),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[2] ),
    .Q_N(_06342_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18782_ (.CLK(_01708_),
    .RESET_B(net78),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[3] ),
    .Q_N(_06341_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18783_ (.CLK(_01709_),
    .RESET_B(net77),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[4] ),
    .Q_N(_06340_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18784_ (.CLK(_01710_),
    .RESET_B(net76),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[5] ),
    .Q_N(_06339_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18785_ (.CLK(_01711_),
    .RESET_B(net75),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[6] ),
    .Q_N(_06338_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18786_ (.CLK(_01712_),
    .RESET_B(net74),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[7] ),
    .Q_N(_06337_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18787_ (.CLK(_01713_),
    .RESET_B(net73),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[8] ),
    .Q_N(_06336_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18788_ (.CLK(_01714_),
    .RESET_B(net72),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[9] ),
    .Q_N(_06335_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18789_ (.CLK(_01715_),
    .RESET_B(net71),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[10] ),
    .Q_N(_06334_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18790_ (.CLK(_01716_),
    .RESET_B(net70),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[11] ),
    .Q_N(_06333_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _18791_ (.CLK(_01717_),
    .RESET_B(net69),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[12] ),
    .Q_N(_06332_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _18792_ (.CLK(_01718_),
    .RESET_B(net68),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[13] ),
    .Q_N(_06331_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _18793_ (.CLK(_01719_),
    .RESET_B(net67),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[14] ),
    .Q_N(_06330_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _18794_ (.CLK(_01720_),
    .RESET_B(net66),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[15] ),
    .Q_N(_06329_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _18795_ (.CLK(_01721_),
    .RESET_B(net65),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[16] ),
    .Q_N(_06328_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _18796_ (.CLK(_01722_),
    .RESET_B(net64),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[17] ),
    .Q_N(_06327_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _18797_ (.CLK(_01723_),
    .RESET_B(net863),
    .D(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.temp_delay[18] ),
    .Q_N(_08303_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.genblk1[2].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _18798_ (.CLK(net5196),
    .RESET_B(net5706),
    .D(_00509_),
    .Q_N(_08304_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[0] ));
 sg13g2_dfrbp_1 _18799_ (.CLK(net5196),
    .RESET_B(net5706),
    .D(_00519_),
    .Q_N(_08305_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[1] ));
 sg13g2_dfrbp_1 _18800_ (.CLK(net5196),
    .RESET_B(net5706),
    .D(_00520_),
    .Q_N(_08306_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[2] ));
 sg13g2_dfrbp_1 _18801_ (.CLK(net5196),
    .RESET_B(net5706),
    .D(_00521_),
    .Q_N(_08307_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[3] ));
 sg13g2_dfrbp_1 _18802_ (.CLK(net5197),
    .RESET_B(net5707),
    .D(_00522_),
    .Q_N(_08308_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[4] ));
 sg13g2_dfrbp_1 _18803_ (.CLK(net5197),
    .RESET_B(net5707),
    .D(_00523_),
    .Q_N(_08309_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[5] ));
 sg13g2_dfrbp_1 _18804_ (.CLK(net5225),
    .RESET_B(net5735),
    .D(_00524_),
    .Q_N(_08310_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[6] ));
 sg13g2_dfrbp_1 _18805_ (.CLK(net5224),
    .RESET_B(net5734),
    .D(_00525_),
    .Q_N(_08311_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[7] ));
 sg13g2_dfrbp_1 _18806_ (.CLK(net5223),
    .RESET_B(net5734),
    .D(_00526_),
    .Q_N(_08312_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[8] ));
 sg13g2_dfrbp_1 _18807_ (.CLK(net5223),
    .RESET_B(net5733),
    .D(_00527_),
    .Q_N(_08313_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[9] ));
 sg13g2_dfrbp_1 _18808_ (.CLK(net5227),
    .RESET_B(net5737),
    .D(_00510_),
    .Q_N(_08314_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[10] ));
 sg13g2_dfrbp_1 _18809_ (.CLK(net5227),
    .RESET_B(net5737),
    .D(_00511_),
    .Q_N(_08315_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[11] ));
 sg13g2_dfrbp_1 _18810_ (.CLK(net5227),
    .RESET_B(net5737),
    .D(_00512_),
    .Q_N(_08316_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[12] ));
 sg13g2_dfrbp_1 _18811_ (.CLK(net5227),
    .RESET_B(net5737),
    .D(_00513_),
    .Q_N(_08317_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[13] ));
 sg13g2_dfrbp_1 _18812_ (.CLK(net5228),
    .RESET_B(net5738),
    .D(_00514_),
    .Q_N(_08318_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[14] ));
 sg13g2_dfrbp_1 _18813_ (.CLK(net5227),
    .RESET_B(net5738),
    .D(_00515_),
    .Q_N(_08319_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[15] ));
 sg13g2_dfrbp_1 _18814_ (.CLK(net5228),
    .RESET_B(net5737),
    .D(_00516_),
    .Q_N(_08320_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[16] ));
 sg13g2_dfrbp_1 _18815_ (.CLK(net5228),
    .RESET_B(net5738),
    .D(_00517_),
    .Q_N(_08321_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[17] ));
 sg13g2_dfrbp_1 _18816_ (.CLK(net5228),
    .RESET_B(net5738),
    .D(_00518_),
    .Q_N(_08322_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u3.reg_value[18] ));
 sg13g2_dfrbp_1 _18817_ (.CLK(net5226),
    .RESET_B(net5735),
    .D(_00509_),
    .Q_N(_08323_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][0] ));
 sg13g2_dfrbp_1 _18818_ (.CLK(net5225),
    .RESET_B(net5736),
    .D(_00519_),
    .Q_N(_08324_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][1] ));
 sg13g2_dfrbp_1 _18819_ (.CLK(net5225),
    .RESET_B(net5735),
    .D(_00520_),
    .Q_N(_08325_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][2] ));
 sg13g2_dfrbp_1 _18820_ (.CLK(net5225),
    .RESET_B(net5735),
    .D(_00521_),
    .Q_N(_08326_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][3] ));
 sg13g2_dfrbp_1 _18821_ (.CLK(net5225),
    .RESET_B(net5735),
    .D(_00522_),
    .Q_N(_08327_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][4] ));
 sg13g2_dfrbp_1 _18822_ (.CLK(net5225),
    .RESET_B(net5735),
    .D(_00523_),
    .Q_N(_08328_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][5] ));
 sg13g2_dfrbp_1 _18823_ (.CLK(net5226),
    .RESET_B(net5736),
    .D(_00524_),
    .Q_N(_08329_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][6] ));
 sg13g2_dfrbp_1 _18824_ (.CLK(net5224),
    .RESET_B(net5733),
    .D(_00525_),
    .Q_N(_08330_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][7] ));
 sg13g2_dfrbp_1 _18825_ (.CLK(net5227),
    .RESET_B(net5737),
    .D(_00526_),
    .Q_N(_08331_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][8] ));
 sg13g2_dfrbp_1 _18826_ (.CLK(net5227),
    .RESET_B(net5737),
    .D(_00527_),
    .Q_N(_08332_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][9] ));
 sg13g2_dfrbp_1 _18827_ (.CLK(net5227),
    .RESET_B(net5737),
    .D(_00510_),
    .Q_N(_08333_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][10] ));
 sg13g2_dfrbp_1 _18828_ (.CLK(net5237),
    .RESET_B(net5747),
    .D(_00511_),
    .Q_N(_08334_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][11] ));
 sg13g2_dfrbp_1 _18829_ (.CLK(net5237),
    .RESET_B(net5747),
    .D(_00512_),
    .Q_N(_08335_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][12] ));
 sg13g2_dfrbp_1 _18830_ (.CLK(net5238),
    .RESET_B(net5748),
    .D(_00513_),
    .Q_N(_08336_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][13] ));
 sg13g2_dfrbp_1 _18831_ (.CLK(net5238),
    .RESET_B(net5748),
    .D(_00514_),
    .Q_N(_08337_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][14] ));
 sg13g2_dfrbp_1 _18832_ (.CLK(net5237),
    .RESET_B(net5747),
    .D(_00515_),
    .Q_N(_08338_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][15] ));
 sg13g2_dfrbp_1 _18833_ (.CLK(net5237),
    .RESET_B(net5747),
    .D(_00516_),
    .Q_N(_08339_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][16] ));
 sg13g2_dfrbp_1 _18834_ (.CLK(net5237),
    .RESET_B(net5747),
    .D(_00517_),
    .Q_N(_08340_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][17] ));
 sg13g2_dfrbp_1 _18835_ (.CLK(net5237),
    .RESET_B(net5747),
    .D(_00518_),
    .Q_N(_08341_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][18] ));
 sg13g2_dfrbp_1 _18836_ (.CLK(net5191),
    .RESET_B(net5701),
    .D(_00490_),
    .Q_N(_08342_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[0] ));
 sg13g2_dfrbp_1 _18837_ (.CLK(net5191),
    .RESET_B(net5701),
    .D(_00500_),
    .Q_N(_08343_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[1] ));
 sg13g2_dfrbp_1 _18838_ (.CLK(net5191),
    .RESET_B(net5701),
    .D(_00501_),
    .Q_N(_08344_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[2] ));
 sg13g2_dfrbp_1 _18839_ (.CLK(net5192),
    .RESET_B(net5702),
    .D(_00502_),
    .Q_N(_08345_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[3] ));
 sg13g2_dfrbp_1 _18840_ (.CLK(net5189),
    .RESET_B(net5699),
    .D(_00503_),
    .Q_N(_08346_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[4] ));
 sg13g2_dfrbp_1 _18841_ (.CLK(net5189),
    .RESET_B(net5699),
    .D(_00504_),
    .Q_N(_08347_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[5] ));
 sg13g2_dfrbp_1 _18842_ (.CLK(net5190),
    .RESET_B(net5700),
    .D(_00505_),
    .Q_N(_08348_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[6] ));
 sg13g2_dfrbp_1 _18843_ (.CLK(net5190),
    .RESET_B(net5700),
    .D(_00506_),
    .Q_N(_08349_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[7] ));
 sg13g2_dfrbp_1 _18844_ (.CLK(net5195),
    .RESET_B(net5705),
    .D(_00507_),
    .Q_N(_08350_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[8] ));
 sg13g2_dfrbp_1 _18845_ (.CLK(net5193),
    .RESET_B(net5703),
    .D(_00508_),
    .Q_N(_08351_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[9] ));
 sg13g2_dfrbp_1 _18846_ (.CLK(net5193),
    .RESET_B(net5703),
    .D(_00491_),
    .Q_N(_08352_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[10] ));
 sg13g2_dfrbp_1 _18847_ (.CLK(net5193),
    .RESET_B(net5703),
    .D(_00492_),
    .Q_N(_08353_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[11] ));
 sg13g2_dfrbp_1 _18848_ (.CLK(net5194),
    .RESET_B(net5704),
    .D(_00493_),
    .Q_N(_08354_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[12] ));
 sg13g2_dfrbp_1 _18849_ (.CLK(net5194),
    .RESET_B(net5704),
    .D(_00494_),
    .Q_N(_08355_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[13] ));
 sg13g2_dfrbp_1 _18850_ (.CLK(net5194),
    .RESET_B(net5704),
    .D(_00495_),
    .Q_N(_08356_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[14] ));
 sg13g2_dfrbp_1 _18851_ (.CLK(net5194),
    .RESET_B(net5704),
    .D(_00496_),
    .Q_N(_08357_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[15] ));
 sg13g2_dfrbp_1 _18852_ (.CLK(net5194),
    .RESET_B(net5704),
    .D(_00497_),
    .Q_N(_08358_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[16] ));
 sg13g2_dfrbp_1 _18853_ (.CLK(net5224),
    .RESET_B(net5734),
    .D(_00498_),
    .Q_N(_08359_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[17] ));
 sg13g2_dfrbp_1 _18854_ (.CLK(net5224),
    .RESET_B(net5734),
    .D(_00499_),
    .Q_N(_08360_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.u2.reg_value[18] ));
 sg13g2_dfrbp_1 _18855_ (.CLK(net5192),
    .RESET_B(net5702),
    .D(_00490_),
    .Q_N(_08361_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[0] ));
 sg13g2_dfrbp_1 _18856_ (.CLK(net5192),
    .RESET_B(net5702),
    .D(_00500_),
    .Q_N(_08362_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[1] ));
 sg13g2_dfrbp_1 _18857_ (.CLK(net5192),
    .RESET_B(net5702),
    .D(_00501_),
    .Q_N(_08363_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[2] ));
 sg13g2_dfrbp_1 _18858_ (.CLK(net5192),
    .RESET_B(net5702),
    .D(_00502_),
    .Q_N(_08364_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[3] ));
 sg13g2_dfrbp_1 _18859_ (.CLK(net5196),
    .RESET_B(net5706),
    .D(_00503_),
    .Q_N(_08365_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[4] ));
 sg13g2_dfrbp_1 _18860_ (.CLK(net5196),
    .RESET_B(net5706),
    .D(_00504_),
    .Q_N(_08366_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[5] ));
 sg13g2_dfrbp_1 _18861_ (.CLK(net5193),
    .RESET_B(net5703),
    .D(_00505_),
    .Q_N(_08367_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[6] ));
 sg13g2_dfrbp_1 _18862_ (.CLK(net5193),
    .RESET_B(net5703),
    .D(_00506_),
    .Q_N(_08368_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[7] ));
 sg13g2_dfrbp_1 _18863_ (.CLK(net5195),
    .RESET_B(net5704),
    .D(_00507_),
    .Q_N(_08369_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[8] ));
 sg13g2_dfrbp_1 _18864_ (.CLK(net5194),
    .RESET_B(net5705),
    .D(_00508_),
    .Q_N(_08370_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[9] ));
 sg13g2_dfrbp_1 _18865_ (.CLK(net5224),
    .RESET_B(net5734),
    .D(_00491_),
    .Q_N(_08371_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[10] ));
 sg13g2_dfrbp_1 _18866_ (.CLK(net5224),
    .RESET_B(net5734),
    .D(_00492_),
    .Q_N(_08372_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[11] ));
 sg13g2_dfrbp_1 _18867_ (.CLK(net5224),
    .RESET_B(net5734),
    .D(_00493_),
    .Q_N(_08373_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[12] ));
 sg13g2_dfrbp_1 _18868_ (.CLK(net5223),
    .RESET_B(net5733),
    .D(_00494_),
    .Q_N(_08374_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[13] ));
 sg13g2_dfrbp_1 _18869_ (.CLK(net5223),
    .RESET_B(net5733),
    .D(_00495_),
    .Q_N(_08375_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[14] ));
 sg13g2_dfrbp_1 _18870_ (.CLK(net5223),
    .RESET_B(net5733),
    .D(_00496_),
    .Q_N(_08376_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[15] ));
 sg13g2_dfrbp_1 _18871_ (.CLK(net5223),
    .RESET_B(net5733),
    .D(_00497_),
    .Q_N(_08377_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[16] ));
 sg13g2_dfrbp_1 _18872_ (.CLK(net5223),
    .RESET_B(net5733),
    .D(_00498_),
    .Q_N(_08378_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[17] ));
 sg13g2_dfrbp_1 _18873_ (.CLK(net5223),
    .RESET_B(net5733),
    .D(_00499_),
    .Q_N(_08379_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator2_out[18] ));
 sg13g2_dfrbp_1 _18874_ (.CLK(net5191),
    .RESET_B(net5701),
    .D(_01193_),
    .Q_N(_01193_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[0] ));
 sg13g2_dfrbp_1 _18875_ (.CLK(net5191),
    .RESET_B(net5701),
    .D(_00481_),
    .Q_N(_08380_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[1] ));
 sg13g2_dfrbp_1 _18876_ (.CLK(net5191),
    .RESET_B(net5701),
    .D(_00482_),
    .Q_N(_08381_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[2] ));
 sg13g2_dfrbp_1 _18877_ (.CLK(net5190),
    .RESET_B(net5700),
    .D(_00483_),
    .Q_N(_08382_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[3] ));
 sg13g2_dfrbp_1 _18878_ (.CLK(net5190),
    .RESET_B(net5700),
    .D(_00484_),
    .Q_N(_08383_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[4] ));
 sg13g2_dfrbp_1 _18879_ (.CLK(net5190),
    .RESET_B(net5700),
    .D(_00485_),
    .Q_N(_08384_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[5] ));
 sg13g2_dfrbp_1 _18880_ (.CLK(net5190),
    .RESET_B(net5700),
    .D(_00486_),
    .Q_N(_08385_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[6] ));
 sg13g2_dfrbp_1 _18881_ (.CLK(net5190),
    .RESET_B(net5700),
    .D(_00487_),
    .Q_N(_08386_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[7] ));
 sg13g2_dfrbp_1 _18882_ (.CLK(net5189),
    .RESET_B(net5699),
    .D(_00488_),
    .Q_N(_08387_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[8] ));
 sg13g2_dfrbp_1 _18883_ (.CLK(net5189),
    .RESET_B(net5699),
    .D(_00489_),
    .Q_N(_08388_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[9] ));
 sg13g2_dfrbp_1 _18884_ (.CLK(net5189),
    .RESET_B(net5699),
    .D(_00472_),
    .Q_N(_08389_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[10] ));
 sg13g2_dfrbp_1 _18885_ (.CLK(net5189),
    .RESET_B(net5699),
    .D(_00473_),
    .Q_N(_08390_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[11] ));
 sg13g2_dfrbp_1 _18886_ (.CLK(net5189),
    .RESET_B(net5699),
    .D(_00474_),
    .Q_N(_08391_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[12] ));
 sg13g2_dfrbp_1 _18887_ (.CLK(net5189),
    .RESET_B(net5699),
    .D(_00475_),
    .Q_N(_08392_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[13] ));
 sg13g2_dfrbp_1 _18888_ (.CLK(net5193),
    .RESET_B(net5703),
    .D(_00476_),
    .Q_N(_08393_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[14] ));
 sg13g2_dfrbp_1 _18889_ (.CLK(net5193),
    .RESET_B(net5703),
    .D(_00477_),
    .Q_N(_08394_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[15] ));
 sg13g2_dfrbp_1 _18890_ (.CLK(net5193),
    .RESET_B(net5703),
    .D(_00478_),
    .Q_N(_08395_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[16] ));
 sg13g2_dfrbp_1 _18891_ (.CLK(net5194),
    .RESET_B(net5704),
    .D(_00479_),
    .Q_N(_08396_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[17] ));
 sg13g2_dfrbp_1 _18892_ (.CLK(net5194),
    .RESET_B(net5704),
    .D(_00480_),
    .Q_N(_08397_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.u_top_module.integrator1_out[18] ));
 sg13g2_dfrbp_1 _18893_ (.CLK(net5030),
    .RESET_B(net864),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][0] ),
    .Q_N(_08398_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18894_ (.CLK(net5030),
    .RESET_B(net865),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][1] ),
    .Q_N(_08399_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18895_ (.CLK(net5030),
    .RESET_B(net866),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][2] ),
    .Q_N(_08400_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18896_ (.CLK(net5030),
    .RESET_B(net867),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][3] ),
    .Q_N(_08401_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18897_ (.CLK(net5030),
    .RESET_B(net868),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][4] ),
    .Q_N(_08402_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18898_ (.CLK(net5031),
    .RESET_B(net869),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][5] ),
    .Q_N(_08403_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18899_ (.CLK(net5031),
    .RESET_B(net870),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][6] ),
    .Q_N(_08404_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18900_ (.CLK(net5032),
    .RESET_B(net871),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][7] ),
    .Q_N(_08405_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18901_ (.CLK(net5032),
    .RESET_B(net872),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][8] ),
    .Q_N(_08406_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18902_ (.CLK(net5035),
    .RESET_B(net873),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][9] ),
    .Q_N(_08407_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18903_ (.CLK(net5035),
    .RESET_B(net874),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][10] ),
    .Q_N(_08408_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18904_ (.CLK(net5039),
    .RESET_B(net875),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][11] ),
    .Q_N(_08409_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18905_ (.CLK(net5039),
    .RESET_B(net876),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][12] ),
    .Q_N(_08410_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18906_ (.CLK(net5038),
    .RESET_B(net877),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][13] ),
    .Q_N(_08411_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18907_ (.CLK(net5038),
    .RESET_B(net878),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][14] ),
    .Q_N(_08412_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18908_ (.CLK(net5038),
    .RESET_B(net879),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][15] ),
    .Q_N(_08413_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18909_ (.CLK(net5039),
    .RESET_B(net880),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][16] ),
    .Q_N(_08414_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18910_ (.CLK(net5035),
    .RESET_B(net881),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][17] ),
    .Q_N(_08415_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18911_ (.CLK(net5037),
    .RESET_B(net882),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[0][18] ),
    .Q_N(_08416_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18912_ (.CLK(net5036),
    .RESET_B(net883),
    .D(_00434_),
    .Q_N(_08417_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][0] ));
 sg13g2_dfrbp_1 _18913_ (.CLK(net5032),
    .RESET_B(net884),
    .D(_00444_),
    .Q_N(_08418_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][1] ));
 sg13g2_dfrbp_1 _18914_ (.CLK(net5032),
    .RESET_B(net885),
    .D(_00445_),
    .Q_N(_08419_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][2] ));
 sg13g2_dfrbp_1 _18915_ (.CLK(net5033),
    .RESET_B(net886),
    .D(_00446_),
    .Q_N(_08420_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][3] ));
 sg13g2_dfrbp_1 _18916_ (.CLK(net5032),
    .RESET_B(net887),
    .D(_00447_),
    .Q_N(_08421_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][4] ));
 sg13g2_dfrbp_1 _18917_ (.CLK(net5032),
    .RESET_B(net888),
    .D(_00448_),
    .Q_N(_08422_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][5] ));
 sg13g2_dfrbp_1 _18918_ (.CLK(net5035),
    .RESET_B(net889),
    .D(_00449_),
    .Q_N(_08423_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][6] ));
 sg13g2_dfrbp_1 _18919_ (.CLK(net5035),
    .RESET_B(net890),
    .D(_00450_),
    .Q_N(_08424_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][7] ));
 sg13g2_dfrbp_1 _18920_ (.CLK(net5039),
    .RESET_B(net891),
    .D(_00451_),
    .Q_N(_08425_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][8] ));
 sg13g2_dfrbp_1 _18921_ (.CLK(net5041),
    .RESET_B(net892),
    .D(_00452_),
    .Q_N(_08426_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][9] ));
 sg13g2_dfrbp_1 _18922_ (.CLK(net5057),
    .RESET_B(net893),
    .D(_00435_),
    .Q_N(_08427_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][10] ));
 sg13g2_dfrbp_1 _18923_ (.CLK(net5059),
    .RESET_B(net894),
    .D(_00436_),
    .Q_N(_08428_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][11] ));
 sg13g2_dfrbp_1 _18924_ (.CLK(net5059),
    .RESET_B(net895),
    .D(_00437_),
    .Q_N(_08429_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][12] ));
 sg13g2_dfrbp_1 _18925_ (.CLK(net5064),
    .RESET_B(net896),
    .D(_00438_),
    .Q_N(_08430_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][13] ));
 sg13g2_dfrbp_1 _18926_ (.CLK(net5064),
    .RESET_B(net897),
    .D(_00439_),
    .Q_N(_08431_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][14] ));
 sg13g2_dfrbp_1 _18927_ (.CLK(net5060),
    .RESET_B(net898),
    .D(_00440_),
    .Q_N(_08432_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][15] ));
 sg13g2_dfrbp_1 _18928_ (.CLK(net5058),
    .RESET_B(net899),
    .D(_00441_),
    .Q_N(_08433_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][16] ));
 sg13g2_dfrbp_1 _18929_ (.CLK(net5057),
    .RESET_B(net900),
    .D(_00442_),
    .Q_N(_08434_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][17] ));
 sg13g2_dfrbp_1 _18930_ (.CLK(net5039),
    .RESET_B(net63),
    .D(_00443_),
    .Q_N(_06326_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][18] ));
 sg13g2_dfrbp_1 _18931_ (.CLK(_01724_),
    .RESET_B(net62),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[0] ),
    .Q_N(_06325_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18932_ (.CLK(_01725_),
    .RESET_B(net61),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[1] ),
    .Q_N(_06324_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18933_ (.CLK(_01726_),
    .RESET_B(net60),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[2] ),
    .Q_N(_06323_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18934_ (.CLK(_01727_),
    .RESET_B(net59),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[3] ),
    .Q_N(_06322_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18935_ (.CLK(_01728_),
    .RESET_B(net58),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[4] ),
    .Q_N(_06321_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18936_ (.CLK(_01729_),
    .RESET_B(net57),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[5] ),
    .Q_N(_06320_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18937_ (.CLK(_01730_),
    .RESET_B(net56),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[6] ),
    .Q_N(_06319_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18938_ (.CLK(_01731_),
    .RESET_B(net55),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[7] ),
    .Q_N(_06318_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18939_ (.CLK(_01732_),
    .RESET_B(net54),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[8] ),
    .Q_N(_06317_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18940_ (.CLK(_01733_),
    .RESET_B(net52),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[9] ),
    .Q_N(_06316_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18941_ (.CLK(_01734_),
    .RESET_B(net51),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[10] ),
    .Q_N(_06315_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18942_ (.CLK(_01735_),
    .RESET_B(net50),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[11] ),
    .Q_N(_06314_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _18943_ (.CLK(_01736_),
    .RESET_B(net49),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[12] ),
    .Q_N(_06313_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _18944_ (.CLK(_01737_),
    .RESET_B(net48),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[13] ),
    .Q_N(_06312_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _18945_ (.CLK(_01738_),
    .RESET_B(net47),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[14] ),
    .Q_N(_06311_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _18946_ (.CLK(_01739_),
    .RESET_B(net46),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[15] ),
    .Q_N(_06310_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _18947_ (.CLK(_01740_),
    .RESET_B(net45),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[16] ),
    .Q_N(_06309_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _18948_ (.CLK(_01741_),
    .RESET_B(net44),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[17] ),
    .Q_N(_06308_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _18949_ (.CLK(_01742_),
    .RESET_B(net901),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.temp_delay[18] ),
    .Q_N(_08435_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[1].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _18950_ (.CLK(net5040),
    .RESET_B(net902),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][0] ),
    .Q_N(_08436_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[0] ));
 sg13g2_dfrbp_1 _18951_ (.CLK(net5037),
    .RESET_B(net903),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][1] ),
    .Q_N(_08437_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[1] ));
 sg13g2_dfrbp_1 _18952_ (.CLK(net5036),
    .RESET_B(net904),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][2] ),
    .Q_N(_08438_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[2] ));
 sg13g2_dfrbp_1 _18953_ (.CLK(net5036),
    .RESET_B(net905),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][3] ),
    .Q_N(_08439_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[3] ));
 sg13g2_dfrbp_1 _18954_ (.CLK(net5036),
    .RESET_B(net906),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][4] ),
    .Q_N(_08440_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[4] ));
 sg13g2_dfrbp_1 _18955_ (.CLK(net5036),
    .RESET_B(net907),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][5] ),
    .Q_N(_08441_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[5] ));
 sg13g2_dfrbp_1 _18956_ (.CLK(net5036),
    .RESET_B(net908),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][6] ),
    .Q_N(_08442_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[6] ));
 sg13g2_dfrbp_1 _18957_ (.CLK(net5038),
    .RESET_B(net909),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][7] ),
    .Q_N(_08443_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[7] ));
 sg13g2_dfrbp_1 _18958_ (.CLK(net5038),
    .RESET_B(net910),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][8] ),
    .Q_N(_08444_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[8] ));
 sg13g2_dfrbp_1 _18959_ (.CLK(net5057),
    .RESET_B(net911),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][9] ),
    .Q_N(_08445_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[9] ));
 sg13g2_dfrbp_1 _18960_ (.CLK(net5059),
    .RESET_B(net912),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][10] ),
    .Q_N(_08446_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[10] ));
 sg13g2_dfrbp_1 _18961_ (.CLK(net5059),
    .RESET_B(net913),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][11] ),
    .Q_N(_08447_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[11] ));
 sg13g2_dfrbp_1 _18962_ (.CLK(net5064),
    .RESET_B(net914),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][12] ),
    .Q_N(_08448_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[12] ));
 sg13g2_dfrbp_1 _18963_ (.CLK(net5065),
    .RESET_B(net915),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][13] ),
    .Q_N(_08449_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[13] ));
 sg13g2_dfrbp_1 _18964_ (.CLK(net5065),
    .RESET_B(net916),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][14] ),
    .Q_N(_08450_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[14] ));
 sg13g2_dfrbp_1 _18965_ (.CLK(net5064),
    .RESET_B(net917),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][15] ),
    .Q_N(_08451_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[15] ));
 sg13g2_dfrbp_1 _18966_ (.CLK(net5060),
    .RESET_B(net918),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][16] ),
    .Q_N(_08452_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[16] ));
 sg13g2_dfrbp_1 _18967_ (.CLK(net5059),
    .RESET_B(net919),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][17] ),
    .Q_N(_08453_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[17] ));
 sg13g2_dfrbp_1 _18968_ (.CLK(net5057),
    .RESET_B(net920),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.comb_data[1][18] ),
    .Q_N(_08454_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[18] ));
 sg13g2_dfrbp_1 _18969_ (.CLK(net5058),
    .RESET_B(net921),
    .D(_00453_),
    .Q_N(_08455_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18970_ (.CLK(net5058),
    .RESET_B(net922),
    .D(_00463_),
    .Q_N(_08456_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18971_ (.CLK(net5041),
    .RESET_B(net923),
    .D(_00464_),
    .Q_N(_08457_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18972_ (.CLK(net5040),
    .RESET_B(net924),
    .D(_00465_),
    .Q_N(_08458_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18973_ (.CLK(net5040),
    .RESET_B(net925),
    .D(_00466_),
    .Q_N(_08459_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18974_ (.CLK(net5040),
    .RESET_B(net926),
    .D(_00467_),
    .Q_N(_08460_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18975_ (.CLK(net5058),
    .RESET_B(net927),
    .D(_00468_),
    .Q_N(_08461_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18976_ (.CLK(net5058),
    .RESET_B(net928),
    .D(_00469_),
    .Q_N(_08462_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18977_ (.CLK(net5060),
    .RESET_B(net929),
    .D(_00470_),
    .Q_N(_08463_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18978_ (.CLK(net5060),
    .RESET_B(net930),
    .D(_00471_),
    .Q_N(_08464_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18979_ (.CLK(net5064),
    .RESET_B(net931),
    .D(_00454_),
    .Q_N(_08465_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18980_ (.CLK(net5064),
    .RESET_B(net932),
    .D(_00455_),
    .Q_N(_08466_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18981_ (.CLK(net5067),
    .RESET_B(net933),
    .D(_00456_),
    .Q_N(_08467_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18982_ (.CLK(net5067),
    .RESET_B(net934),
    .D(_00457_),
    .Q_N(_08468_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18983_ (.CLK(net5067),
    .RESET_B(net935),
    .D(_00458_),
    .Q_N(_08469_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18984_ (.CLK(net5067),
    .RESET_B(net936),
    .D(_00459_),
    .Q_N(_08470_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18985_ (.CLK(net5066),
    .RESET_B(net937),
    .D(_00460_),
    .Q_N(_08471_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18986_ (.CLK(net5066),
    .RESET_B(net938),
    .D(_00461_),
    .Q_N(_08472_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18987_ (.CLK(net5060),
    .RESET_B(net43),
    .D(_00462_),
    .Q_N(_06307_),
    .Q(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _18988_ (.CLK(_01743_),
    .RESET_B(net42),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[0] ),
    .Q_N(_06306_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[0] ));
 sg13g2_dfrbp_1 _18989_ (.CLK(_01744_),
    .RESET_B(net41),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[1] ),
    .Q_N(_06305_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[1] ));
 sg13g2_dfrbp_1 _18990_ (.CLK(_01745_),
    .RESET_B(net40),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[2] ),
    .Q_N(_06304_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[2] ));
 sg13g2_dfrbp_1 _18991_ (.CLK(_01746_),
    .RESET_B(net39),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[3] ),
    .Q_N(_06303_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[3] ));
 sg13g2_dfrbp_1 _18992_ (.CLK(_01747_),
    .RESET_B(net38),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[4] ),
    .Q_N(_06302_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[4] ));
 sg13g2_dfrbp_1 _18993_ (.CLK(_01748_),
    .RESET_B(net37),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[5] ),
    .Q_N(_06301_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[5] ));
 sg13g2_dfrbp_1 _18994_ (.CLK(_01749_),
    .RESET_B(net36),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[6] ),
    .Q_N(_06300_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[6] ));
 sg13g2_dfrbp_1 _18995_ (.CLK(_01750_),
    .RESET_B(net35),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[7] ),
    .Q_N(_06299_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[7] ));
 sg13g2_dfrbp_1 _18996_ (.CLK(_01751_),
    .RESET_B(net34),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[8] ),
    .Q_N(_06298_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[8] ));
 sg13g2_dfrbp_1 _18997_ (.CLK(_01752_),
    .RESET_B(net33),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[9] ),
    .Q_N(_06297_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[9] ));
 sg13g2_dfrbp_1 _18998_ (.CLK(_01753_),
    .RESET_B(net32),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[10] ),
    .Q_N(_06296_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[10] ));
 sg13g2_dfrbp_1 _18999_ (.CLK(_01754_),
    .RESET_B(net31),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[11] ),
    .Q_N(_06295_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[11] ));
 sg13g2_dfrbp_1 _19000_ (.CLK(_01755_),
    .RESET_B(net30),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[12] ),
    .Q_N(_06294_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[12] ));
 sg13g2_dfrbp_1 _19001_ (.CLK(_01756_),
    .RESET_B(net29),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[13] ),
    .Q_N(_06293_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[13] ));
 sg13g2_dfrbp_1 _19002_ (.CLK(_01757_),
    .RESET_B(net28),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[14] ),
    .Q_N(_06292_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[14] ));
 sg13g2_dfrbp_1 _19003_ (.CLK(_01758_),
    .RESET_B(net27),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[15] ),
    .Q_N(_06291_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[15] ));
 sg13g2_dfrbp_1 _19004_ (.CLK(_01759_),
    .RESET_B(net26),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[16] ),
    .Q_N(_06290_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[16] ));
 sg13g2_dfrbp_1 _19005_ (.CLK(_01760_),
    .RESET_B(net25),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[17] ),
    .Q_N(_06289_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[17] ));
 sg13g2_dfrbp_1 _19006_ (.CLK(_01761_),
    .RESET_B(net24),
    .D(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.temp_delay[18] ),
    .Q_N(_06288_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.genblk1[2].u_comb.delay_line[18] ));
 sg13g2_dfrbp_1 _19007_ (.CLK(_01762_),
    .RESET_B(net939),
    .D(_01807_),
    .Q_N(_08473_),
    .Q(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.out ));
 sg13g2_dfrbp_1 _19008_ (.CLK(net5461),
    .RESET_B(net5969),
    .D(_00287_),
    .Q_N(_06287_),
    .Q(\u_supermic_top_module.u_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _19009_ (.CLK(_01763_),
    .RESET_B(net5969),
    .D(\u_supermic_top_module.u_i2s_bus.u_mux_shift.data ),
    .Q_N(_08474_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _19010_ (.CLK(net5461),
    .RESET_B(net5969),
    .D(_00266_),
    .Q_N(_06286_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19011_ (.CLK(_01764_),
    .RESET_B(net6011),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_08475_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19012_ (.CLK(net5502),
    .RESET_B(net6011),
    .D(_00277_),
    .Q_N(_06285_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19013_ (.CLK(_01765_),
    .RESET_B(net6015),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_08476_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19014_ (.CLK(net5506),
    .RESET_B(net6015),
    .D(_00280_),
    .Q_N(_06284_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19015_ (.CLK(_01766_),
    .RESET_B(net6015),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_08477_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19016_ (.CLK(net5507),
    .RESET_B(net6016),
    .D(_00281_),
    .Q_N(_06283_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19017_ (.CLK(_01767_),
    .RESET_B(net6017),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_08478_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19018_ (.CLK(net5508),
    .RESET_B(net6017),
    .D(_00282_),
    .Q_N(_06282_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19019_ (.CLK(_01768_),
    .RESET_B(net6017),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_08479_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19020_ (.CLK(net5508),
    .RESET_B(net6017),
    .D(_00283_),
    .Q_N(_06281_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19021_ (.CLK(_01769_),
    .RESET_B(net6037),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_08480_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19022_ (.CLK(net5507),
    .RESET_B(net6016),
    .D(_00284_),
    .Q_N(_06280_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19023_ (.CLK(_01770_),
    .RESET_B(net6016),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_08481_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19024_ (.CLK(net5480),
    .RESET_B(net5989),
    .D(_00285_),
    .Q_N(_06279_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19025_ (.CLK(_01771_),
    .RESET_B(net5988),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_08482_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19026_ (.CLK(net5437),
    .RESET_B(net5946),
    .D(_00286_),
    .Q_N(_06278_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19027_ (.CLK(_01772_),
    .RESET_B(net5944),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_08483_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _19028_ (.CLK(net5455),
    .RESET_B(net5964),
    .D(_00256_),
    .Q_N(_06277_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19029_ (.CLK(_01773_),
    .RESET_B(net5948),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_08484_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19030_ (.CLK(net5440),
    .RESET_B(net5949),
    .D(_00257_),
    .Q_N(_06276_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19031_ (.CLK(_01774_),
    .RESET_B(net5952),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_08485_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19032_ (.CLK(net5443),
    .RESET_B(net5952),
    .D(_00258_),
    .Q_N(_06275_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19033_ (.CLK(_01775_),
    .RESET_B(net5952),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_08486_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19034_ (.CLK(net5407),
    .RESET_B(net5916),
    .D(_00259_),
    .Q_N(_06274_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19035_ (.CLK(_01776_),
    .RESET_B(net5916),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_08487_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19036_ (.CLK(net5407),
    .RESET_B(net5916),
    .D(_00260_),
    .Q_N(_06273_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19037_ (.CLK(_01777_),
    .RESET_B(net5910),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_08488_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19038_ (.CLK(net5401),
    .RESET_B(net5910),
    .D(_00261_),
    .Q_N(_06272_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19039_ (.CLK(_01778_),
    .RESET_B(net5910),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_08489_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19040_ (.CLK(net5400),
    .RESET_B(net5909),
    .D(_00262_),
    .Q_N(_06271_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19041_ (.CLK(_01779_),
    .RESET_B(net5910),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_08490_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19042_ (.CLK(net5400),
    .RESET_B(net5909),
    .D(_00263_),
    .Q_N(_06270_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19043_ (.CLK(_01780_),
    .RESET_B(net5909),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_08491_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19044_ (.CLK(net5366),
    .RESET_B(net5875),
    .D(_00264_),
    .Q_N(_06269_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19045_ (.CLK(_01781_),
    .RESET_B(net5888),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_08492_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19046_ (.CLK(net5368),
    .RESET_B(net5876),
    .D(_00265_),
    .Q_N(_06268_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19047_ (.CLK(_01782_),
    .RESET_B(net5876),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_08493_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19048_ (.CLK(net5363),
    .RESET_B(net5872),
    .D(_00267_),
    .Q_N(_06267_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19049_ (.CLK(_01783_),
    .RESET_B(net5873),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_08494_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19050_ (.CLK(net5346),
    .RESET_B(net5855),
    .D(_00268_),
    .Q_N(_06266_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19051_ (.CLK(_01784_),
    .RESET_B(net5855),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_08495_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19052_ (.CLK(net5346),
    .RESET_B(net5855),
    .D(_00269_),
    .Q_N(_06265_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19053_ (.CLK(_01785_),
    .RESET_B(net5863),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_08496_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19054_ (.CLK(net5355),
    .RESET_B(net5863),
    .D(_00270_),
    .Q_N(_06264_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19055_ (.CLK(_01786_),
    .RESET_B(net5863),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_08497_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19056_ (.CLK(net5355),
    .RESET_B(net5863),
    .D(_00271_),
    .Q_N(_06263_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19057_ (.CLK(_01787_),
    .RESET_B(net5863),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_08498_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19058_ (.CLK(net5346),
    .RESET_B(net5855),
    .D(_00272_),
    .Q_N(_06262_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19059_ (.CLK(_01788_),
    .RESET_B(net5855),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_08499_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19060_ (.CLK(net5303),
    .RESET_B(net5812),
    .D(_00273_),
    .Q_N(_06261_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19061_ (.CLK(_01789_),
    .RESET_B(net5811),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_08500_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19062_ (.CLK(net5302),
    .RESET_B(net5811),
    .D(_00274_),
    .Q_N(_06260_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19063_ (.CLK(_01790_),
    .RESET_B(net5811),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_08501_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19064_ (.CLK(net5297),
    .RESET_B(net5807),
    .D(_00275_),
    .Q_N(_06259_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19065_ (.CLK(_01791_),
    .RESET_B(net5807),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_08502_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19066_ (.CLK(net5298),
    .RESET_B(net5808),
    .D(_00276_),
    .Q_N(_06258_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19067_ (.CLK(_01792_),
    .RESET_B(net5808),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_08503_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19068_ (.CLK(net5307),
    .RESET_B(net5816),
    .D(_00278_),
    .Q_N(_06257_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19069_ (.CLK(_01793_),
    .RESET_B(net5816),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_08504_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19070_ (.CLK(net5217),
    .RESET_B(net5731),
    .D(_00279_),
    .Q_N(_06256_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _19071_ (.CLK(_01794_),
    .RESET_B(net5730),
    .D(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_08505_),
    .Q(\u_supermic_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _19072_ (.CLK(net5307),
    .RESET_B(net5816),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][0] ),
    .Q_N(_08506_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][0] ));
 sg13g2_dfrbp_1 _19073_ (.CLK(net5290),
    .RESET_B(net5800),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][1] ),
    .Q_N(_08507_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][1] ));
 sg13g2_dfrbp_1 _19074_ (.CLK(net5291),
    .RESET_B(net5801),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][2] ),
    .Q_N(_08508_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][2] ));
 sg13g2_dfrbp_1 _19075_ (.CLK(net5291),
    .RESET_B(net5801),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][3] ),
    .Q_N(_08509_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][3] ));
 sg13g2_dfrbp_1 _19076_ (.CLK(net5291),
    .RESET_B(net5801),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][4] ),
    .Q_N(_00316_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][4] ));
 sg13g2_dfrbp_1 _19077_ (.CLK(net5291),
    .RESET_B(net5801),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][5] ),
    .Q_N(_00325_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][5] ));
 sg13g2_dfrbp_1 _19078_ (.CLK(net5291),
    .RESET_B(net5801),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][6] ),
    .Q_N(_08510_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][6] ));
 sg13g2_dfrbp_1 _19079_ (.CLK(net5290),
    .RESET_B(net5800),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][7] ),
    .Q_N(_08511_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][7] ));
 sg13g2_dfrbp_1 _19080_ (.CLK(net5298),
    .RESET_B(net5808),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][8] ),
    .Q_N(_00348_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][8] ));
 sg13g2_dfrbp_1 _19081_ (.CLK(net5297),
    .RESET_B(net5807),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][9] ),
    .Q_N(_00357_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][9] ));
 sg13g2_dfrbp_1 _19082_ (.CLK(net5302),
    .RESET_B(net5811),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][10] ),
    .Q_N(_08512_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][10] ));
 sg13g2_dfrbp_1 _19083_ (.CLK(net5303),
    .RESET_B(net5812),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][11] ),
    .Q_N(_08513_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][11] ));
 sg13g2_dfrbp_1 _19084_ (.CLK(net5348),
    .RESET_B(net5856),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][12] ),
    .Q_N(_00380_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][12] ));
 sg13g2_dfrbp_1 _19085_ (.CLK(net5346),
    .RESET_B(net5856),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][13] ),
    .Q_N(_00389_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][13] ));
 sg13g2_dfrbp_1 _19086_ (.CLK(net5347),
    .RESET_B(net5857),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][14] ),
    .Q_N(_08514_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][14] ));
 sg13g2_dfrbp_1 _19087_ (.CLK(net5346),
    .RESET_B(net5857),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][15] ),
    .Q_N(_08515_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][15] ));
 sg13g2_dfrbp_1 _19088_ (.CLK(net5348),
    .RESET_B(net5856),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][16] ),
    .Q_N(_00412_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][16] ));
 sg13g2_dfrbp_1 _19089_ (.CLK(net5313),
    .RESET_B(net5822),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][17] ),
    .Q_N(_08516_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][17] ));
 sg13g2_dfrbp_1 _19090_ (.CLK(net5306),
    .RESET_B(net5815),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][18] ),
    .Q_N(_08517_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[1][18] ));
 sg13g2_dfrbp_1 _19091_ (.CLK(net5290),
    .RESET_B(net5800),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.u_mux_shift.sum_res ),
    .Q_N(_08518_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][0] ));
 sg13g2_dfrbp_1 _19092_ (.CLK(net5291),
    .RESET_B(net5801),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .Q_N(_08519_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][1] ));
 sg13g2_dfrbp_1 _19093_ (.CLK(net5287),
    .RESET_B(net5797),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .Q_N(_08520_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][2] ));
 sg13g2_dfrbp_1 _19094_ (.CLK(net5287),
    .RESET_B(net5797),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .Q_N(_08521_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][3] ));
 sg13g2_dfrbp_1 _19095_ (.CLK(net5287),
    .RESET_B(net5797),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .Q_N(_00315_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][4] ));
 sg13g2_dfrbp_1 _19096_ (.CLK(net5287),
    .RESET_B(net5797),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .Q_N(_00324_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][5] ));
 sg13g2_dfrbp_1 _19097_ (.CLK(net5281),
    .RESET_B(net5791),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .Q_N(_08522_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][6] ));
 sg13g2_dfrbp_1 _19098_ (.CLK(net5283),
    .RESET_B(net5793),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .Q_N(_08523_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][7] ));
 sg13g2_dfrbp_1 _19099_ (.CLK(net5298),
    .RESET_B(net5808),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .Q_N(_00347_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][8] ));
 sg13g2_dfrbp_1 _19100_ (.CLK(net5298),
    .RESET_B(net5808),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .Q_N(_00356_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][9] ));
 sg13g2_dfrbp_1 _19101_ (.CLK(net5297),
    .RESET_B(net5807),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .Q_N(_08524_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][10] ));
 sg13g2_dfrbp_1 _19102_ (.CLK(net5302),
    .RESET_B(net5811),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .Q_N(_08525_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][11] ));
 sg13g2_dfrbp_1 _19103_ (.CLK(net5348),
    .RESET_B(net5856),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .Q_N(_00379_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][12] ));
 sg13g2_dfrbp_1 _19104_ (.CLK(net5348),
    .RESET_B(net5856),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .Q_N(_00388_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][13] ));
 sg13g2_dfrbp_1 _19105_ (.CLK(net5347),
    .RESET_B(net5855),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .Q_N(_08526_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][14] ));
 sg13g2_dfrbp_1 _19106_ (.CLK(net5348),
    .RESET_B(net5856),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .Q_N(_08527_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][15] ));
 sg13g2_dfrbp_1 _19107_ (.CLK(net5303),
    .RESET_B(net5812),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .Q_N(_00411_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][16] ));
 sg13g2_dfrbp_1 _19108_ (.CLK(net5302),
    .RESET_B(net5811),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .Q_N(_08528_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][17] ));
 sg13g2_dfrbp_1 _19109_ (.CLK(net5298),
    .RESET_B(net5808),
    .D(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .Q_N(_08529_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[0].u_delay_line.buffer[0][18] ));
 sg13g2_dfrbp_1 _19110_ (.CLK(net5400),
    .RESET_B(net5909),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][0] ),
    .Q_N(_08530_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][0] ));
 sg13g2_dfrbp_1 _19111_ (.CLK(net5250),
    .RESET_B(net5760),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][1] ),
    .Q_N(_08531_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][1] ));
 sg13g2_dfrbp_1 _19112_ (.CLK(net5245),
    .RESET_B(net5755),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][2] ),
    .Q_N(_08532_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][2] ));
 sg13g2_dfrbp_1 _19113_ (.CLK(net5244),
    .RESET_B(net5754),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][3] ),
    .Q_N(_08533_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][3] ));
 sg13g2_dfrbp_1 _19114_ (.CLK(net5245),
    .RESET_B(net5755),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][4] ),
    .Q_N(_08534_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][4] ));
 sg13g2_dfrbp_1 _19115_ (.CLK(net5251),
    .RESET_B(net5761),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][5] ),
    .Q_N(_08535_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][5] ));
 sg13g2_dfrbp_1 _19116_ (.CLK(net5246),
    .RESET_B(net5756),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][6] ),
    .Q_N(_08536_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][6] ));
 sg13g2_dfrbp_1 _19117_ (.CLK(net5246),
    .RESET_B(net5756),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][7] ),
    .Q_N(_08537_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][7] ));
 sg13g2_dfrbp_1 _19118_ (.CLK(net5239),
    .RESET_B(net5749),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][8] ),
    .Q_N(_08538_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][8] ));
 sg13g2_dfrbp_1 _19119_ (.CLK(net5248),
    .RESET_B(net5758),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][9] ),
    .Q_N(_08539_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][9] ));
 sg13g2_dfrbp_1 _19120_ (.CLK(net5240),
    .RESET_B(net5750),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][10] ),
    .Q_N(_08540_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][10] ));
 sg13g2_dfrbp_1 _19121_ (.CLK(net5239),
    .RESET_B(net5749),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][11] ),
    .Q_N(_08541_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][11] ));
 sg13g2_dfrbp_1 _19122_ (.CLK(net5285),
    .RESET_B(net5795),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][12] ),
    .Q_N(_08542_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][12] ));
 sg13g2_dfrbp_1 _19123_ (.CLK(net5285),
    .RESET_B(net5795),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][13] ),
    .Q_N(_08543_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][13] ));
 sg13g2_dfrbp_1 _19124_ (.CLK(net5287),
    .RESET_B(net5797),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][14] ),
    .Q_N(_08544_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][14] ));
 sg13g2_dfrbp_1 _19125_ (.CLK(net5249),
    .RESET_B(net5759),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][15] ),
    .Q_N(_08545_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][15] ));
 sg13g2_dfrbp_1 _19126_ (.CLK(net5240),
    .RESET_B(net5750),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][16] ),
    .Q_N(_08546_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][16] ));
 sg13g2_dfrbp_1 _19127_ (.CLK(net5292),
    .RESET_B(net5802),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][17] ),
    .Q_N(_08547_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][17] ));
 sg13g2_dfrbp_1 _19128_ (.CLK(net5250),
    .RESET_B(net5760),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][18] ),
    .Q_N(_08548_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[5][18] ));
 sg13g2_dfrbp_1 _19129_ (.CLK(net5401),
    .RESET_B(net5910),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][0] ),
    .Q_N(_08549_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][0] ));
 sg13g2_dfrbp_1 _19130_ (.CLK(net5250),
    .RESET_B(net5760),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][1] ),
    .Q_N(_08550_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][1] ));
 sg13g2_dfrbp_1 _19131_ (.CLK(net5244),
    .RESET_B(net5754),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][2] ),
    .Q_N(_08551_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][2] ));
 sg13g2_dfrbp_1 _19132_ (.CLK(net5244),
    .RESET_B(net5754),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][3] ),
    .Q_N(_08552_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][3] ));
 sg13g2_dfrbp_1 _19133_ (.CLK(net5244),
    .RESET_B(net5754),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][4] ),
    .Q_N(_08553_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][4] ));
 sg13g2_dfrbp_1 _19134_ (.CLK(net5251),
    .RESET_B(net5761),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][5] ),
    .Q_N(_08554_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][5] ));
 sg13g2_dfrbp_1 _19135_ (.CLK(net5246),
    .RESET_B(net5756),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][6] ),
    .Q_N(_08555_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][6] ));
 sg13g2_dfrbp_1 _19136_ (.CLK(net5246),
    .RESET_B(net5756),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][7] ),
    .Q_N(_08556_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][7] ));
 sg13g2_dfrbp_1 _19137_ (.CLK(net5239),
    .RESET_B(net5749),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][8] ),
    .Q_N(_08557_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][8] ));
 sg13g2_dfrbp_1 _19138_ (.CLK(net5248),
    .RESET_B(net5758),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][9] ),
    .Q_N(_08558_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][9] ));
 sg13g2_dfrbp_1 _19139_ (.CLK(net5240),
    .RESET_B(net5750),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][10] ),
    .Q_N(_08559_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][10] ));
 sg13g2_dfrbp_1 _19140_ (.CLK(net5239),
    .RESET_B(net5749),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][11] ),
    .Q_N(_08560_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][11] ));
 sg13g2_dfrbp_1 _19141_ (.CLK(net5285),
    .RESET_B(net5795),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][12] ),
    .Q_N(_08561_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][12] ));
 sg13g2_dfrbp_1 _19142_ (.CLK(net5285),
    .RESET_B(net5795),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][13] ),
    .Q_N(_08562_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][13] ));
 sg13g2_dfrbp_1 _19143_ (.CLK(net5287),
    .RESET_B(net5797),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][14] ),
    .Q_N(_08563_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][14] ));
 sg13g2_dfrbp_1 _19144_ (.CLK(net5249),
    .RESET_B(net5759),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][15] ),
    .Q_N(_08564_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][15] ));
 sg13g2_dfrbp_1 _19145_ (.CLK(net5241),
    .RESET_B(net5751),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][16] ),
    .Q_N(_08565_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][16] ));
 sg13g2_dfrbp_1 _19146_ (.CLK(net5292),
    .RESET_B(net5802),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][17] ),
    .Q_N(_08566_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][17] ));
 sg13g2_dfrbp_1 _19147_ (.CLK(net5250),
    .RESET_B(net5760),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][18] ),
    .Q_N(_08567_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[4][18] ));
 sg13g2_dfrbp_1 _19148_ (.CLK(net5401),
    .RESET_B(net5909),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][0] ),
    .Q_N(_08568_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][0] ));
 sg13g2_dfrbp_1 _19149_ (.CLK(net5245),
    .RESET_B(net5755),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][1] ),
    .Q_N(_08569_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][1] ));
 sg13g2_dfrbp_1 _19150_ (.CLK(net5244),
    .RESET_B(net5754),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][2] ),
    .Q_N(_08570_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][2] ));
 sg13g2_dfrbp_1 _19151_ (.CLK(net5244),
    .RESET_B(net5754),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][3] ),
    .Q_N(_08571_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][3] ));
 sg13g2_dfrbp_1 _19152_ (.CLK(net5244),
    .RESET_B(net5754),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][4] ),
    .Q_N(_08572_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][4] ));
 sg13g2_dfrbp_1 _19153_ (.CLK(net5251),
    .RESET_B(net5761),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][5] ),
    .Q_N(_08573_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][5] ));
 sg13g2_dfrbp_1 _19154_ (.CLK(net5246),
    .RESET_B(net5756),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][6] ),
    .Q_N(_08574_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][6] ));
 sg13g2_dfrbp_1 _19155_ (.CLK(net5246),
    .RESET_B(net5756),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][7] ),
    .Q_N(_08575_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][7] ));
 sg13g2_dfrbp_1 _19156_ (.CLK(net5239),
    .RESET_B(net5749),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][8] ),
    .Q_N(_08576_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][8] ));
 sg13g2_dfrbp_1 _19157_ (.CLK(net5248),
    .RESET_B(net5758),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][9] ),
    .Q_N(_08577_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][9] ));
 sg13g2_dfrbp_1 _19158_ (.CLK(net5239),
    .RESET_B(net5749),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][10] ),
    .Q_N(_08578_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][10] ));
 sg13g2_dfrbp_1 _19159_ (.CLK(net5239),
    .RESET_B(net5749),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][11] ),
    .Q_N(_08579_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][11] ));
 sg13g2_dfrbp_1 _19160_ (.CLK(net5286),
    .RESET_B(net5796),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][12] ),
    .Q_N(_08580_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][12] ));
 sg13g2_dfrbp_1 _19161_ (.CLK(net5285),
    .RESET_B(net5795),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][13] ),
    .Q_N(_08581_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][13] ));
 sg13g2_dfrbp_1 _19162_ (.CLK(net5287),
    .RESET_B(net5797),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][14] ),
    .Q_N(_08582_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][14] ));
 sg13g2_dfrbp_1 _19163_ (.CLK(net5248),
    .RESET_B(net5758),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][15] ),
    .Q_N(_08583_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][15] ));
 sg13g2_dfrbp_1 _19164_ (.CLK(net5241),
    .RESET_B(net5751),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][16] ),
    .Q_N(_08584_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][16] ));
 sg13g2_dfrbp_1 _19165_ (.CLK(net5292),
    .RESET_B(net5802),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][17] ),
    .Q_N(_08585_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][17] ));
 sg13g2_dfrbp_1 _19166_ (.CLK(net5250),
    .RESET_B(net5760),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][18] ),
    .Q_N(_08586_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[3][18] ));
 sg13g2_dfrbp_1 _19167_ (.CLK(net5400),
    .RESET_B(net5909),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][0] ),
    .Q_N(_08587_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][0] ));
 sg13g2_dfrbp_1 _19168_ (.CLK(net5245),
    .RESET_B(net5755),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][1] ),
    .Q_N(_08588_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][1] ));
 sg13g2_dfrbp_1 _19169_ (.CLK(net5243),
    .RESET_B(net5753),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][2] ),
    .Q_N(_08589_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][2] ));
 sg13g2_dfrbp_1 _19170_ (.CLK(net5243),
    .RESET_B(net5753),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][3] ),
    .Q_N(_08590_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][3] ));
 sg13g2_dfrbp_1 _19171_ (.CLK(net5244),
    .RESET_B(net5754),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][4] ),
    .Q_N(_08591_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][4] ));
 sg13g2_dfrbp_1 _19172_ (.CLK(net5251),
    .RESET_B(net5761),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][5] ),
    .Q_N(_08592_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][5] ));
 sg13g2_dfrbp_1 _19173_ (.CLK(net5246),
    .RESET_B(net5756),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][6] ),
    .Q_N(_08593_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][6] ));
 sg13g2_dfrbp_1 _19174_ (.CLK(net5243),
    .RESET_B(net5753),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][7] ),
    .Q_N(_08594_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][7] ));
 sg13g2_dfrbp_1 _19175_ (.CLK(net5242),
    .RESET_B(net5752),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][8] ),
    .Q_N(_08595_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][8] ));
 sg13g2_dfrbp_1 _19176_ (.CLK(net5248),
    .RESET_B(net5758),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][9] ),
    .Q_N(_08596_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][9] ));
 sg13g2_dfrbp_1 _19177_ (.CLK(net5239),
    .RESET_B(net5749),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][10] ),
    .Q_N(_08597_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][10] ));
 sg13g2_dfrbp_1 _19178_ (.CLK(net5242),
    .RESET_B(net5752),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][11] ),
    .Q_N(_08598_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][11] ));
 sg13g2_dfrbp_1 _19179_ (.CLK(net5286),
    .RESET_B(net5796),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][12] ),
    .Q_N(_08599_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][12] ));
 sg13g2_dfrbp_1 _19180_ (.CLK(net5285),
    .RESET_B(net5795),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][13] ),
    .Q_N(_08600_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][13] ));
 sg13g2_dfrbp_1 _19181_ (.CLK(net5287),
    .RESET_B(net5797),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][14] ),
    .Q_N(_08601_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][14] ));
 sg13g2_dfrbp_1 _19182_ (.CLK(net5248),
    .RESET_B(net5758),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][15] ),
    .Q_N(_08602_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][15] ));
 sg13g2_dfrbp_1 _19183_ (.CLK(net5241),
    .RESET_B(net5751),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][16] ),
    .Q_N(_08603_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][16] ));
 sg13g2_dfrbp_1 _19184_ (.CLK(net5291),
    .RESET_B(net5801),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][17] ),
    .Q_N(_08604_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][17] ));
 sg13g2_dfrbp_1 _19185_ (.CLK(net5250),
    .RESET_B(net5760),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][18] ),
    .Q_N(_08605_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[2][18] ));
 sg13g2_dfrbp_1 _19186_ (.CLK(net5381),
    .RESET_B(net5890),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][0] ),
    .Q_N(_08606_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][0] ));
 sg13g2_dfrbp_1 _19187_ (.CLK(net5243),
    .RESET_B(net5753),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][1] ),
    .Q_N(_08607_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][1] ));
 sg13g2_dfrbp_1 _19188_ (.CLK(net5243),
    .RESET_B(net5753),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][2] ),
    .Q_N(_08608_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][2] ));
 sg13g2_dfrbp_1 _19189_ (.CLK(net5247),
    .RESET_B(net5757),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][3] ),
    .Q_N(_08609_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][3] ));
 sg13g2_dfrbp_1 _19190_ (.CLK(net5247),
    .RESET_B(net5757),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][4] ),
    .Q_N(_08610_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][4] ));
 sg13g2_dfrbp_1 _19191_ (.CLK(net5250),
    .RESET_B(net5760),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][5] ),
    .Q_N(_08611_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][5] ));
 sg13g2_dfrbp_1 _19192_ (.CLK(net5243),
    .RESET_B(net5753),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][6] ),
    .Q_N(_08612_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][6] ));
 sg13g2_dfrbp_1 _19193_ (.CLK(net5243),
    .RESET_B(net5753),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][7] ),
    .Q_N(_08613_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][7] ));
 sg13g2_dfrbp_1 _19194_ (.CLK(net5242),
    .RESET_B(net5752),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][8] ),
    .Q_N(_08614_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][8] ));
 sg13g2_dfrbp_1 _19195_ (.CLK(net5248),
    .RESET_B(net5758),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][9] ),
    .Q_N(_08615_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][9] ));
 sg13g2_dfrbp_1 _19196_ (.CLK(net5242),
    .RESET_B(net5752),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][10] ),
    .Q_N(_08616_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][10] ));
 sg13g2_dfrbp_1 _19197_ (.CLK(net5242),
    .RESET_B(net5752),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][11] ),
    .Q_N(_08617_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][11] ));
 sg13g2_dfrbp_1 _19198_ (.CLK(net5285),
    .RESET_B(net5795),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][12] ),
    .Q_N(_08618_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][12] ));
 sg13g2_dfrbp_1 _19199_ (.CLK(net5285),
    .RESET_B(net5795),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][13] ),
    .Q_N(_08619_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][13] ));
 sg13g2_dfrbp_1 _19200_ (.CLK(net5288),
    .RESET_B(net5798),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][14] ),
    .Q_N(_08620_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][14] ));
 sg13g2_dfrbp_1 _19201_ (.CLK(net5248),
    .RESET_B(net5758),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][15] ),
    .Q_N(_08621_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][15] ));
 sg13g2_dfrbp_1 _19202_ (.CLK(net5242),
    .RESET_B(net5752),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][16] ),
    .Q_N(_08622_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][16] ));
 sg13g2_dfrbp_1 _19203_ (.CLK(net5291),
    .RESET_B(net5801),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][17] ),
    .Q_N(_08623_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][17] ));
 sg13g2_dfrbp_1 _19204_ (.CLK(net5246),
    .RESET_B(net5756),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][18] ),
    .Q_N(_08624_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[1][18] ));
 sg13g2_dfrbp_1 _19205_ (.CLK(net5325),
    .RESET_B(net5835),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ),
    .Q_N(_00293_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][0] ));
 sg13g2_dfrbp_1 _19206_ (.CLK(net5269),
    .RESET_B(net5779),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .Q_N(_00294_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][1] ));
 sg13g2_dfrbp_1 _19207_ (.CLK(net5260),
    .RESET_B(net5770),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .Q_N(_00301_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][2] ));
 sg13g2_dfrbp_1 _19208_ (.CLK(net5235),
    .RESET_B(net5745),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .Q_N(_00308_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][3] ));
 sg13g2_dfrbp_1 _19209_ (.CLK(net5235),
    .RESET_B(net5745),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .Q_N(_00317_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][4] ));
 sg13g2_dfrbp_1 _19210_ (.CLK(net5250),
    .RESET_B(net5760),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .Q_N(_00326_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][5] ));
 sg13g2_dfrbp_1 _19211_ (.CLK(net5235),
    .RESET_B(net5745),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .Q_N(_00333_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][6] ));
 sg13g2_dfrbp_1 _19212_ (.CLK(net5235),
    .RESET_B(net5745),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .Q_N(_00340_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][7] ));
 sg13g2_dfrbp_1 _19213_ (.CLK(net5235),
    .RESET_B(net5745),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .Q_N(_00349_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][8] ));
 sg13g2_dfrbp_1 _19214_ (.CLK(net5240),
    .RESET_B(net5750),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .Q_N(_00358_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][9] ));
 sg13g2_dfrbp_1 _19215_ (.CLK(net5234),
    .RESET_B(net5744),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .Q_N(_00365_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][10] ));
 sg13g2_dfrbp_1 _19216_ (.CLK(net5234),
    .RESET_B(net5744),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .Q_N(_00372_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][11] ));
 sg13g2_dfrbp_1 _19217_ (.CLK(net5249),
    .RESET_B(net5759),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .Q_N(_00381_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][12] ));
 sg13g2_dfrbp_1 _19218_ (.CLK(net5249),
    .RESET_B(net5759),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .Q_N(_00390_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][13] ));
 sg13g2_dfrbp_1 _19219_ (.CLK(net5286),
    .RESET_B(net5796),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .Q_N(_00397_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][14] ));
 sg13g2_dfrbp_1 _19220_ (.CLK(net5241),
    .RESET_B(net5751),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .Q_N(_00404_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][15] ));
 sg13g2_dfrbp_1 _19221_ (.CLK(net5242),
    .RESET_B(net5752),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .Q_N(_00413_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][16] ));
 sg13g2_dfrbp_1 _19222_ (.CLK(net5288),
    .RESET_B(net5798),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .Q_N(_00420_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][17] ));
 sg13g2_dfrbp_1 _19223_ (.CLK(net5243),
    .RESET_B(net5753),
    .D(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .Q_N(_00427_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[1].u_delay_line.buffer[0][18] ));
 sg13g2_dfrbp_1 _19224_ (.CLK(net5400),
    .RESET_B(net5909),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][0] ),
    .Q_N(_08625_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][0] ));
 sg13g2_dfrbp_1 _19225_ (.CLK(net5400),
    .RESET_B(net5909),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][1] ),
    .Q_N(_08626_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][1] ));
 sg13g2_dfrbp_1 _19226_ (.CLK(net5367),
    .RESET_B(net5875),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][2] ),
    .Q_N(_08627_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][2] ));
 sg13g2_dfrbp_1 _19227_ (.CLK(net5366),
    .RESET_B(net5876),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][3] ),
    .Q_N(_08628_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][3] ));
 sg13g2_dfrbp_1 _19228_ (.CLK(net5363),
    .RESET_B(net5872),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][4] ),
    .Q_N(_08629_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][4] ));
 sg13g2_dfrbp_1 _19229_ (.CLK(net5358),
    .RESET_B(net5867),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][5] ),
    .Q_N(_08630_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][5] ));
 sg13g2_dfrbp_1 _19230_ (.CLK(net5361),
    .RESET_B(net5870),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][6] ),
    .Q_N(_08631_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][6] ));
 sg13g2_dfrbp_1 _19231_ (.CLK(net5315),
    .RESET_B(net5824),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][7] ),
    .Q_N(_08632_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][7] ));
 sg13g2_dfrbp_1 _19232_ (.CLK(net5314),
    .RESET_B(net5823),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][8] ),
    .Q_N(_08633_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][8] ));
 sg13g2_dfrbp_1 _19233_ (.CLK(net5312),
    .RESET_B(net5821),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][9] ),
    .Q_N(_08634_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][9] ));
 sg13g2_dfrbp_1 _19234_ (.CLK(net5312),
    .RESET_B(net5821),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][10] ),
    .Q_N(_08635_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][10] ));
 sg13g2_dfrbp_1 _19235_ (.CLK(net5357),
    .RESET_B(net5866),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][11] ),
    .Q_N(_08636_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][11] ));
 sg13g2_dfrbp_1 _19236_ (.CLK(net5311),
    .RESET_B(net5820),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][12] ),
    .Q_N(_08637_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][12] ));
 sg13g2_dfrbp_1 _19237_ (.CLK(net5311),
    .RESET_B(net5820),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][13] ),
    .Q_N(_08638_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][13] ));
 sg13g2_dfrbp_1 _19238_ (.CLK(net5311),
    .RESET_B(net5820),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][14] ),
    .Q_N(_08639_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][14] ));
 sg13g2_dfrbp_1 _19239_ (.CLK(net5357),
    .RESET_B(net5866),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][15] ),
    .Q_N(_08640_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][15] ));
 sg13g2_dfrbp_1 _19240_ (.CLK(net5362),
    .RESET_B(net5871),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][16] ),
    .Q_N(_08641_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][16] ));
 sg13g2_dfrbp_1 _19241_ (.CLK(net5365),
    .RESET_B(net5874),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][17] ),
    .Q_N(_08642_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][17] ));
 sg13g2_dfrbp_1 _19242_ (.CLK(net5364),
    .RESET_B(net5873),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][18] ),
    .Q_N(_08643_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[7][18] ));
 sg13g2_dfrbp_1 _19243_ (.CLK(net5388),
    .RESET_B(net5897),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][0] ),
    .Q_N(_08644_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][0] ));
 sg13g2_dfrbp_1 _19244_ (.CLK(net5388),
    .RESET_B(net5897),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][1] ),
    .Q_N(_08645_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][1] ));
 sg13g2_dfrbp_1 _19245_ (.CLK(net5367),
    .RESET_B(net5875),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][2] ),
    .Q_N(_08646_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][2] ));
 sg13g2_dfrbp_1 _19246_ (.CLK(net5366),
    .RESET_B(net5876),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][3] ),
    .Q_N(_08647_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][3] ));
 sg13g2_dfrbp_1 _19247_ (.CLK(net5363),
    .RESET_B(net5872),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][4] ),
    .Q_N(_08648_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][4] ));
 sg13g2_dfrbp_1 _19248_ (.CLK(net5359),
    .RESET_B(net5867),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][5] ),
    .Q_N(_08649_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][5] ));
 sg13g2_dfrbp_1 _19249_ (.CLK(net5358),
    .RESET_B(net5867),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][6] ),
    .Q_N(_08650_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][6] ));
 sg13g2_dfrbp_1 _19250_ (.CLK(net5314),
    .RESET_B(net5824),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][7] ),
    .Q_N(_08651_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][7] ));
 sg13g2_dfrbp_1 _19251_ (.CLK(net5314),
    .RESET_B(net5823),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][8] ),
    .Q_N(_08652_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][8] ));
 sg13g2_dfrbp_1 _19252_ (.CLK(net5312),
    .RESET_B(net5821),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][9] ),
    .Q_N(_08653_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][9] ));
 sg13g2_dfrbp_1 _19253_ (.CLK(net5312),
    .RESET_B(net5821),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][10] ),
    .Q_N(_08654_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][10] ));
 sg13g2_dfrbp_1 _19254_ (.CLK(net5357),
    .RESET_B(net5866),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][11] ),
    .Q_N(_08655_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][11] ));
 sg13g2_dfrbp_1 _19255_ (.CLK(net5310),
    .RESET_B(net5819),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][12] ),
    .Q_N(_08656_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][12] ));
 sg13g2_dfrbp_1 _19256_ (.CLK(net5310),
    .RESET_B(net5819),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][13] ),
    .Q_N(_08657_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][13] ));
 sg13g2_dfrbp_1 _19257_ (.CLK(net5311),
    .RESET_B(net5820),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][14] ),
    .Q_N(_08658_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][14] ));
 sg13g2_dfrbp_1 _19258_ (.CLK(net5313),
    .RESET_B(net5822),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][15] ),
    .Q_N(_08659_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][15] ));
 sg13g2_dfrbp_1 _19259_ (.CLK(net5362),
    .RESET_B(net5871),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][16] ),
    .Q_N(_08660_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][16] ));
 sg13g2_dfrbp_1 _19260_ (.CLK(net5365),
    .RESET_B(net5874),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][17] ),
    .Q_N(_08661_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][17] ));
 sg13g2_dfrbp_1 _19261_ (.CLK(net5362),
    .RESET_B(net5871),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][18] ),
    .Q_N(_08662_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[6][18] ));
 sg13g2_dfrbp_1 _19262_ (.CLK(net5388),
    .RESET_B(net5898),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][0] ),
    .Q_N(_08663_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][0] ));
 sg13g2_dfrbp_1 _19263_ (.CLK(net5389),
    .RESET_B(net5898),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][1] ),
    .Q_N(_08664_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][1] ));
 sg13g2_dfrbp_1 _19264_ (.CLK(net5367),
    .RESET_B(net5875),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][2] ),
    .Q_N(_08665_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][2] ));
 sg13g2_dfrbp_1 _19265_ (.CLK(net5366),
    .RESET_B(net5876),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][3] ),
    .Q_N(_08666_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][3] ));
 sg13g2_dfrbp_1 _19266_ (.CLK(net5363),
    .RESET_B(net5872),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][4] ),
    .Q_N(_08667_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][4] ));
 sg13g2_dfrbp_1 _19267_ (.CLK(net5358),
    .RESET_B(net5868),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][5] ),
    .Q_N(_08668_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][5] ));
 sg13g2_dfrbp_1 _19268_ (.CLK(net5358),
    .RESET_B(net5867),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][6] ),
    .Q_N(_08669_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][6] ));
 sg13g2_dfrbp_1 _19269_ (.CLK(net5315),
    .RESET_B(net5823),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][7] ),
    .Q_N(_08670_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][7] ));
 sg13g2_dfrbp_1 _19270_ (.CLK(net5314),
    .RESET_B(net5823),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][8] ),
    .Q_N(_08671_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][8] ));
 sg13g2_dfrbp_1 _19271_ (.CLK(net5305),
    .RESET_B(net5814),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][9] ),
    .Q_N(_08672_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][9] ));
 sg13g2_dfrbp_1 _19272_ (.CLK(net5312),
    .RESET_B(net5821),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][10] ),
    .Q_N(_08673_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][10] ));
 sg13g2_dfrbp_1 _19273_ (.CLK(net5357),
    .RESET_B(net5866),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][11] ),
    .Q_N(_08674_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][11] ));
 sg13g2_dfrbp_1 _19274_ (.CLK(net5310),
    .RESET_B(net5819),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][12] ),
    .Q_N(_08675_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][12] ));
 sg13g2_dfrbp_1 _19275_ (.CLK(net5310),
    .RESET_B(net5819),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][13] ),
    .Q_N(_08676_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][13] ));
 sg13g2_dfrbp_1 _19276_ (.CLK(net5311),
    .RESET_B(net5820),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][14] ),
    .Q_N(_08677_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][14] ));
 sg13g2_dfrbp_1 _19277_ (.CLK(net5313),
    .RESET_B(net5822),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][15] ),
    .Q_N(_08678_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][15] ));
 sg13g2_dfrbp_1 _19278_ (.CLK(net5364),
    .RESET_B(net5873),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][16] ),
    .Q_N(_08679_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][16] ));
 sg13g2_dfrbp_1 _19279_ (.CLK(net5365),
    .RESET_B(net5874),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][17] ),
    .Q_N(_08680_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][17] ));
 sg13g2_dfrbp_1 _19280_ (.CLK(net5362),
    .RESET_B(net5871),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][18] ),
    .Q_N(_08681_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[5][18] ));
 sg13g2_dfrbp_1 _19281_ (.CLK(net5388),
    .RESET_B(net5897),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][0] ),
    .Q_N(_08682_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][0] ));
 sg13g2_dfrbp_1 _19282_ (.CLK(net5388),
    .RESET_B(net5897),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][1] ),
    .Q_N(_08683_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][1] ));
 sg13g2_dfrbp_1 _19283_ (.CLK(net5359),
    .RESET_B(net5868),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][2] ),
    .Q_N(_08684_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][2] ));
 sg13g2_dfrbp_1 _19284_ (.CLK(net5366),
    .RESET_B(net5876),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][3] ),
    .Q_N(_08685_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][3] ));
 sg13g2_dfrbp_1 _19285_ (.CLK(net5363),
    .RESET_B(net5872),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][4] ),
    .Q_N(_08686_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][4] ));
 sg13g2_dfrbp_1 _19286_ (.CLK(net5359),
    .RESET_B(net5868),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][5] ),
    .Q_N(_08687_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][5] ));
 sg13g2_dfrbp_1 _19287_ (.CLK(net5357),
    .RESET_B(net5866),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][6] ),
    .Q_N(_08688_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][6] ));
 sg13g2_dfrbp_1 _19288_ (.CLK(net5315),
    .RESET_B(net5823),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][7] ),
    .Q_N(_08689_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][7] ));
 sg13g2_dfrbp_1 _19289_ (.CLK(net5308),
    .RESET_B(net5817),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][8] ),
    .Q_N(_08690_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][8] ));
 sg13g2_dfrbp_1 _19290_ (.CLK(net5305),
    .RESET_B(net5814),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][9] ),
    .Q_N(_08691_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][9] ));
 sg13g2_dfrbp_1 _19291_ (.CLK(net5312),
    .RESET_B(net5821),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][10] ),
    .Q_N(_08692_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][10] ));
 sg13g2_dfrbp_1 _19292_ (.CLK(net5357),
    .RESET_B(net5866),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][11] ),
    .Q_N(_08693_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][11] ));
 sg13g2_dfrbp_1 _19293_ (.CLK(net5310),
    .RESET_B(net5819),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][12] ),
    .Q_N(_08694_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][12] ));
 sg13g2_dfrbp_1 _19294_ (.CLK(net5310),
    .RESET_B(net5819),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][13] ),
    .Q_N(_08695_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][13] ));
 sg13g2_dfrbp_1 _19295_ (.CLK(net5311),
    .RESET_B(net5820),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][14] ),
    .Q_N(_08696_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][14] ));
 sg13g2_dfrbp_1 _19296_ (.CLK(net5313),
    .RESET_B(net5822),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][15] ),
    .Q_N(_08697_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][15] ));
 sg13g2_dfrbp_1 _19297_ (.CLK(net5362),
    .RESET_B(net5871),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][16] ),
    .Q_N(_08698_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][16] ));
 sg13g2_dfrbp_1 _19298_ (.CLK(net5365),
    .RESET_B(net5874),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][17] ),
    .Q_N(_08699_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][17] ));
 sg13g2_dfrbp_1 _19299_ (.CLK(net5362),
    .RESET_B(net5871),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][18] ),
    .Q_N(_08700_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[4][18] ));
 sg13g2_dfrbp_1 _19300_ (.CLK(net5388),
    .RESET_B(net5897),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][0] ),
    .Q_N(_08701_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][0] ));
 sg13g2_dfrbp_1 _19301_ (.CLK(net5389),
    .RESET_B(net5897),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][1] ),
    .Q_N(_08702_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][1] ));
 sg13g2_dfrbp_1 _19302_ (.CLK(net5359),
    .RESET_B(net5868),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][2] ),
    .Q_N(_08703_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][2] ));
 sg13g2_dfrbp_1 _19303_ (.CLK(net5366),
    .RESET_B(net5876),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][3] ),
    .Q_N(_08704_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][3] ));
 sg13g2_dfrbp_1 _19304_ (.CLK(net5363),
    .RESET_B(net5872),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][4] ),
    .Q_N(_08705_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][4] ));
 sg13g2_dfrbp_1 _19305_ (.CLK(net5316),
    .RESET_B(net5825),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][5] ),
    .Q_N(_08706_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][5] ));
 sg13g2_dfrbp_1 _19306_ (.CLK(net5358),
    .RESET_B(net5867),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][6] ),
    .Q_N(_08707_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][6] ));
 sg13g2_dfrbp_1 _19307_ (.CLK(net5314),
    .RESET_B(net5824),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][7] ),
    .Q_N(_08708_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][7] ));
 sg13g2_dfrbp_1 _19308_ (.CLK(net5308),
    .RESET_B(net5817),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][8] ),
    .Q_N(_08709_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][8] ));
 sg13g2_dfrbp_1 _19309_ (.CLK(net5305),
    .RESET_B(net5814),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][9] ),
    .Q_N(_08710_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][9] ));
 sg13g2_dfrbp_1 _19310_ (.CLK(net5312),
    .RESET_B(net5821),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][10] ),
    .Q_N(_08711_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][10] ));
 sg13g2_dfrbp_1 _19311_ (.CLK(net5357),
    .RESET_B(net5866),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][11] ),
    .Q_N(_08712_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][11] ));
 sg13g2_dfrbp_1 _19312_ (.CLK(net5310),
    .RESET_B(net5819),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][12] ),
    .Q_N(_08713_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][12] ));
 sg13g2_dfrbp_1 _19313_ (.CLK(net5306),
    .RESET_B(net5815),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][13] ),
    .Q_N(_08714_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][13] ));
 sg13g2_dfrbp_1 _19314_ (.CLK(net5310),
    .RESET_B(net5819),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][14] ),
    .Q_N(_08715_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][14] ));
 sg13g2_dfrbp_1 _19315_ (.CLK(net5313),
    .RESET_B(net5822),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][15] ),
    .Q_N(_08716_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][15] ));
 sg13g2_dfrbp_1 _19316_ (.CLK(net5362),
    .RESET_B(net5871),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][16] ),
    .Q_N(_08717_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][16] ));
 sg13g2_dfrbp_1 _19317_ (.CLK(net5365),
    .RESET_B(net5874),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][17] ),
    .Q_N(_08718_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][17] ));
 sg13g2_dfrbp_1 _19318_ (.CLK(net5362),
    .RESET_B(net5872),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][18] ),
    .Q_N(_08719_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[3][18] ));
 sg13g2_dfrbp_1 _19319_ (.CLK(net5388),
    .RESET_B(net5897),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][0] ),
    .Q_N(_08720_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][0] ));
 sg13g2_dfrbp_1 _19320_ (.CLK(net5388),
    .RESET_B(net5897),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][1] ),
    .Q_N(_08721_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][1] ));
 sg13g2_dfrbp_1 _19321_ (.CLK(net5359),
    .RESET_B(net5868),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][2] ),
    .Q_N(_08722_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][2] ));
 sg13g2_dfrbp_1 _19322_ (.CLK(net5367),
    .RESET_B(net5875),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][3] ),
    .Q_N(_08723_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][3] ));
 sg13g2_dfrbp_1 _19323_ (.CLK(net5363),
    .RESET_B(net5871),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][4] ),
    .Q_N(_08724_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][4] ));
 sg13g2_dfrbp_1 _19324_ (.CLK(net5316),
    .RESET_B(net5825),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][5] ),
    .Q_N(_08725_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][5] ));
 sg13g2_dfrbp_1 _19325_ (.CLK(net5358),
    .RESET_B(net5867),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][6] ),
    .Q_N(_08726_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][6] ));
 sg13g2_dfrbp_1 _19326_ (.CLK(net5315),
    .RESET_B(net5824),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][7] ),
    .Q_N(_08727_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][7] ));
 sg13g2_dfrbp_1 _19327_ (.CLK(net5308),
    .RESET_B(net5817),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][8] ),
    .Q_N(_08728_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][8] ));
 sg13g2_dfrbp_1 _19328_ (.CLK(net5308),
    .RESET_B(net5817),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][9] ),
    .Q_N(_08729_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][9] ));
 sg13g2_dfrbp_1 _19329_ (.CLK(net5305),
    .RESET_B(net5814),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][10] ),
    .Q_N(_08730_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][10] ));
 sg13g2_dfrbp_1 _19330_ (.CLK(net5357),
    .RESET_B(net5866),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][11] ),
    .Q_N(_08731_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][11] ));
 sg13g2_dfrbp_1 _19331_ (.CLK(net5305),
    .RESET_B(net5814),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][12] ),
    .Q_N(_08732_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][12] ));
 sg13g2_dfrbp_1 _19332_ (.CLK(net5306),
    .RESET_B(net5815),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][13] ),
    .Q_N(_08733_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][13] ));
 sg13g2_dfrbp_1 _19333_ (.CLK(net5306),
    .RESET_B(net5815),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][14] ),
    .Q_N(_08734_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][14] ));
 sg13g2_dfrbp_1 _19334_ (.CLK(net5313),
    .RESET_B(net5822),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][15] ),
    .Q_N(_08735_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][15] ));
 sg13g2_dfrbp_1 _19335_ (.CLK(net5361),
    .RESET_B(net5870),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][16] ),
    .Q_N(_08736_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][16] ));
 sg13g2_dfrbp_1 _19336_ (.CLK(net5365),
    .RESET_B(net5874),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][17] ),
    .Q_N(_08737_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][17] ));
 sg13g2_dfrbp_1 _19337_ (.CLK(net5367),
    .RESET_B(net5875),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][18] ),
    .Q_N(_08738_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[2][18] ));
 sg13g2_dfrbp_1 _19338_ (.CLK(net5394),
    .RESET_B(net5903),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][0] ),
    .Q_N(_08739_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][0] ));
 sg13g2_dfrbp_1 _19339_ (.CLK(net5394),
    .RESET_B(net5903),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][1] ),
    .Q_N(_08740_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][1] ));
 sg13g2_dfrbp_1 _19340_ (.CLK(net5359),
    .RESET_B(net5868),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][2] ),
    .Q_N(_08741_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][2] ));
 sg13g2_dfrbp_1 _19341_ (.CLK(net5367),
    .RESET_B(net5875),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][3] ),
    .Q_N(_08742_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][3] ));
 sg13g2_dfrbp_1 _19342_ (.CLK(net5360),
    .RESET_B(net5869),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][4] ),
    .Q_N(_08743_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][4] ));
 sg13g2_dfrbp_1 _19343_ (.CLK(net5330),
    .RESET_B(net5840),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][5] ),
    .Q_N(_08744_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][5] ));
 sg13g2_dfrbp_1 _19344_ (.CLK(net5358),
    .RESET_B(net5867),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][6] ),
    .Q_N(_08745_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][6] ));
 sg13g2_dfrbp_1 _19345_ (.CLK(net5309),
    .RESET_B(net5818),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][7] ),
    .Q_N(_08746_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][7] ));
 sg13g2_dfrbp_1 _19346_ (.CLK(net5309),
    .RESET_B(net5818),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][8] ),
    .Q_N(_08747_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][8] ));
 sg13g2_dfrbp_1 _19347_ (.CLK(net5309),
    .RESET_B(net5818),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][9] ),
    .Q_N(_08748_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][9] ));
 sg13g2_dfrbp_1 _19348_ (.CLK(net5309),
    .RESET_B(net5818),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][10] ),
    .Q_N(_08749_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][10] ));
 sg13g2_dfrbp_1 _19349_ (.CLK(net5313),
    .RESET_B(net5822),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][11] ),
    .Q_N(_08750_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][11] ));
 sg13g2_dfrbp_1 _19350_ (.CLK(net5305),
    .RESET_B(net5814),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][12] ),
    .Q_N(_08751_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][12] ));
 sg13g2_dfrbp_1 _19351_ (.CLK(net5305),
    .RESET_B(net5814),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][13] ),
    .Q_N(_08752_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][13] ));
 sg13g2_dfrbp_1 _19352_ (.CLK(net5305),
    .RESET_B(net5814),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][14] ),
    .Q_N(_08753_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][14] ));
 sg13g2_dfrbp_1 _19353_ (.CLK(net5314),
    .RESET_B(net5823),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][15] ),
    .Q_N(_08754_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][15] ));
 sg13g2_dfrbp_1 _19354_ (.CLK(net5361),
    .RESET_B(net5870),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][16] ),
    .Q_N(_08755_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][16] ));
 sg13g2_dfrbp_1 _19355_ (.CLK(net5367),
    .RESET_B(net5875),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][17] ),
    .Q_N(_08756_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][17] ));
 sg13g2_dfrbp_1 _19356_ (.CLK(net5360),
    .RESET_B(net5869),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][18] ),
    .Q_N(_08757_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[1][18] ));
 sg13g2_dfrbp_1 _19357_ (.CLK(net5382),
    .RESET_B(net5891),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.u_mux_shift.sum_res ),
    .Q_N(_00291_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][0] ));
 sg13g2_dfrbp_1 _19358_ (.CLK(net5382),
    .RESET_B(net5891),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .Q_N(_00295_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][1] ));
 sg13g2_dfrbp_1 _19359_ (.CLK(net5381),
    .RESET_B(net5890),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .Q_N(_00302_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][2] ));
 sg13g2_dfrbp_1 _19360_ (.CLK(net5382),
    .RESET_B(net5891),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .Q_N(_00309_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][3] ));
 sg13g2_dfrbp_1 _19361_ (.CLK(net5360),
    .RESET_B(net5869),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .Q_N(_00318_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][4] ));
 sg13g2_dfrbp_1 _19362_ (.CLK(net5330),
    .RESET_B(net5840),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .Q_N(_00327_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][5] ));
 sg13g2_dfrbp_1 _19363_ (.CLK(net5316),
    .RESET_B(net5825),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .Q_N(_00334_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][6] ));
 sg13g2_dfrbp_1 _19364_ (.CLK(net5308),
    .RESET_B(net5817),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .Q_N(_00341_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][7] ));
 sg13g2_dfrbp_1 _19365_ (.CLK(net5308),
    .RESET_B(net5817),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .Q_N(_00350_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][8] ));
 sg13g2_dfrbp_1 _19366_ (.CLK(net5308),
    .RESET_B(net5817),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .Q_N(_00359_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][9] ));
 sg13g2_dfrbp_1 _19367_ (.CLK(net5308),
    .RESET_B(net5817),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .Q_N(_00366_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][10] ));
 sg13g2_dfrbp_1 _19368_ (.CLK(net5314),
    .RESET_B(net5823),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .Q_N(_00373_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][11] ));
 sg13g2_dfrbp_1 _19369_ (.CLK(net5307),
    .RESET_B(net5816),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .Q_N(_00382_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][12] ));
 sg13g2_dfrbp_1 _19370_ (.CLK(net5307),
    .RESET_B(net5816),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .Q_N(_00391_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][13] ));
 sg13g2_dfrbp_1 _19371_ (.CLK(net5307),
    .RESET_B(net5816),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .Q_N(_00398_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][14] ));
 sg13g2_dfrbp_1 _19372_ (.CLK(net5314),
    .RESET_B(net5823),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .Q_N(_00405_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][15] ));
 sg13g2_dfrbp_1 _19373_ (.CLK(net5358),
    .RESET_B(net5867),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .Q_N(_00414_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][16] ));
 sg13g2_dfrbp_1 _19374_ (.CLK(net5360),
    .RESET_B(net5869),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .Q_N(_00421_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][17] ));
 sg13g2_dfrbp_1 _19375_ (.CLK(net5359),
    .RESET_B(net5868),
    .D(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .Q_N(_00428_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[2].u_delay_line.buffer[0][18] ));
 sg13g2_dfrbp_1 _19376_ (.CLK(net5405),
    .RESET_B(net5914),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][0] ),
    .Q_N(_08758_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][0] ));
 sg13g2_dfrbp_1 _19377_ (.CLK(net5402),
    .RESET_B(net5911),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][1] ),
    .Q_N(_08759_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][1] ));
 sg13g2_dfrbp_1 _19378_ (.CLK(net5406),
    .RESET_B(net5915),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][2] ),
    .Q_N(_08760_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][2] ));
 sg13g2_dfrbp_1 _19379_ (.CLK(net5410),
    .RESET_B(net5919),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][3] ),
    .Q_N(_08761_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][3] ));
 sg13g2_dfrbp_1 _19380_ (.CLK(net5405),
    .RESET_B(net5914),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][4] ),
    .Q_N(_08762_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][4] ));
 sg13g2_dfrbp_1 _19381_ (.CLK(net5402),
    .RESET_B(net5911),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][5] ),
    .Q_N(_08763_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][5] ));
 sg13g2_dfrbp_1 _19382_ (.CLK(net5392),
    .RESET_B(net5901),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][6] ),
    .Q_N(_08764_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][6] ));
 sg13g2_dfrbp_1 _19383_ (.CLK(net5391),
    .RESET_B(net5900),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][7] ),
    .Q_N(_08765_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][7] ));
 sg13g2_dfrbp_1 _19384_ (.CLK(net5386),
    .RESET_B(net5895),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][8] ),
    .Q_N(_08766_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][8] ));
 sg13g2_dfrbp_1 _19385_ (.CLK(net5386),
    .RESET_B(net5895),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][9] ),
    .Q_N(_08767_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][9] ));
 sg13g2_dfrbp_1 _19386_ (.CLK(net5384),
    .RESET_B(net5893),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][10] ),
    .Q_N(_08768_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][10] ));
 sg13g2_dfrbp_1 _19387_ (.CLK(net5384),
    .RESET_B(net5893),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][11] ),
    .Q_N(_08769_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][11] ));
 sg13g2_dfrbp_1 _19388_ (.CLK(net5383),
    .RESET_B(net5892),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][12] ),
    .Q_N(_08770_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][12] ));
 sg13g2_dfrbp_1 _19389_ (.CLK(net5328),
    .RESET_B(net5838),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][13] ),
    .Q_N(_08771_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][13] ));
 sg13g2_dfrbp_1 _19390_ (.CLK(net5381),
    .RESET_B(net5890),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][14] ),
    .Q_N(_08772_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][14] ));
 sg13g2_dfrbp_1 _19391_ (.CLK(net5381),
    .RESET_B(net5890),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][15] ),
    .Q_N(_08773_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][15] ));
 sg13g2_dfrbp_1 _19392_ (.CLK(net5389),
    .RESET_B(net5898),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][16] ),
    .Q_N(_08774_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][16] ));
 sg13g2_dfrbp_1 _19393_ (.CLK(net5392),
    .RESET_B(net5901),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][17] ),
    .Q_N(_08775_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][17] ));
 sg13g2_dfrbp_1 _19394_ (.CLK(net5390),
    .RESET_B(net5899),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][18] ),
    .Q_N(_08776_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[7][18] ));
 sg13g2_dfrbp_1 _19395_ (.CLK(net5405),
    .RESET_B(net5914),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][0] ),
    .Q_N(_08777_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][0] ));
 sg13g2_dfrbp_1 _19396_ (.CLK(net5402),
    .RESET_B(net5911),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][1] ),
    .Q_N(_08778_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][1] ));
 sg13g2_dfrbp_1 _19397_ (.CLK(net5403),
    .RESET_B(net5912),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][2] ),
    .Q_N(_08779_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][2] ));
 sg13g2_dfrbp_1 _19398_ (.CLK(net5410),
    .RESET_B(net5919),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][3] ),
    .Q_N(_08780_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][3] ));
 sg13g2_dfrbp_1 _19399_ (.CLK(net5405),
    .RESET_B(net5914),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][4] ),
    .Q_N(_08781_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][4] ));
 sg13g2_dfrbp_1 _19400_ (.CLK(net5404),
    .RESET_B(net5913),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][5] ),
    .Q_N(_08782_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][5] ));
 sg13g2_dfrbp_1 _19401_ (.CLK(net5392),
    .RESET_B(net5901),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][6] ),
    .Q_N(_08783_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][6] ));
 sg13g2_dfrbp_1 _19402_ (.CLK(net5391),
    .RESET_B(net5900),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][7] ),
    .Q_N(_08784_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][7] ));
 sg13g2_dfrbp_1 _19403_ (.CLK(net5385),
    .RESET_B(net5894),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][8] ),
    .Q_N(_08785_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][8] ));
 sg13g2_dfrbp_1 _19404_ (.CLK(net5385),
    .RESET_B(net5894),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][9] ),
    .Q_N(_08786_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][9] ));
 sg13g2_dfrbp_1 _19405_ (.CLK(net5383),
    .RESET_B(net5892),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][10] ),
    .Q_N(_08787_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][10] ));
 sg13g2_dfrbp_1 _19406_ (.CLK(net5383),
    .RESET_B(net5893),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][11] ),
    .Q_N(_08788_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][11] ));
 sg13g2_dfrbp_1 _19407_ (.CLK(net5383),
    .RESET_B(net5892),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][12] ),
    .Q_N(_08789_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][12] ));
 sg13g2_dfrbp_1 _19408_ (.CLK(net5328),
    .RESET_B(net5838),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][13] ),
    .Q_N(_08790_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][13] ));
 sg13g2_dfrbp_1 _19409_ (.CLK(net5381),
    .RESET_B(net5890),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][14] ),
    .Q_N(_08791_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][14] ));
 sg13g2_dfrbp_1 _19410_ (.CLK(net5381),
    .RESET_B(net5890),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][15] ),
    .Q_N(_08792_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][15] ));
 sg13g2_dfrbp_1 _19411_ (.CLK(net5389),
    .RESET_B(net5898),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][16] ),
    .Q_N(_08793_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][16] ));
 sg13g2_dfrbp_1 _19412_ (.CLK(net5392),
    .RESET_B(net5901),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][17] ),
    .Q_N(_08794_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][17] ));
 sg13g2_dfrbp_1 _19413_ (.CLK(net5390),
    .RESET_B(net5899),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][18] ),
    .Q_N(_08795_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[6][18] ));
 sg13g2_dfrbp_1 _19414_ (.CLK(net5405),
    .RESET_B(net5914),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][0] ),
    .Q_N(_08796_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][0] ));
 sg13g2_dfrbp_1 _19415_ (.CLK(net5402),
    .RESET_B(net5911),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][1] ),
    .Q_N(_08797_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][1] ));
 sg13g2_dfrbp_1 _19416_ (.CLK(net5403),
    .RESET_B(net5912),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][2] ),
    .Q_N(_08798_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][2] ));
 sg13g2_dfrbp_1 _19417_ (.CLK(net5408),
    .RESET_B(net5917),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][3] ),
    .Q_N(_08799_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][3] ));
 sg13g2_dfrbp_1 _19418_ (.CLK(net5410),
    .RESET_B(net5919),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][4] ),
    .Q_N(_08800_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][4] ));
 sg13g2_dfrbp_1 _19419_ (.CLK(net5404),
    .RESET_B(net5913),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][5] ),
    .Q_N(_08801_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][5] ));
 sg13g2_dfrbp_1 _19420_ (.CLK(net5393),
    .RESET_B(net5902),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][6] ),
    .Q_N(_08802_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][6] ));
 sg13g2_dfrbp_1 _19421_ (.CLK(net5391),
    .RESET_B(net5900),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][7] ),
    .Q_N(_08803_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][7] ));
 sg13g2_dfrbp_1 _19422_ (.CLK(net5385),
    .RESET_B(net5894),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][8] ),
    .Q_N(_08804_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][8] ));
 sg13g2_dfrbp_1 _19423_ (.CLK(net5385),
    .RESET_B(net5894),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][9] ),
    .Q_N(_08805_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][9] ));
 sg13g2_dfrbp_1 _19424_ (.CLK(net5384),
    .RESET_B(net5892),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][10] ),
    .Q_N(_08806_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][10] ));
 sg13g2_dfrbp_1 _19425_ (.CLK(net5383),
    .RESET_B(net5893),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][11] ),
    .Q_N(_08807_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][11] ));
 sg13g2_dfrbp_1 _19426_ (.CLK(net5383),
    .RESET_B(net5892),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][12] ),
    .Q_N(_08808_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][12] ));
 sg13g2_dfrbp_1 _19427_ (.CLK(net5328),
    .RESET_B(net5838),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][13] ),
    .Q_N(_08809_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][13] ));
 sg13g2_dfrbp_1 _19428_ (.CLK(net5329),
    .RESET_B(net5839),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][14] ),
    .Q_N(_08810_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][14] ));
 sg13g2_dfrbp_1 _19429_ (.CLK(net5381),
    .RESET_B(net5890),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][15] ),
    .Q_N(_08811_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][15] ));
 sg13g2_dfrbp_1 _19430_ (.CLK(net5389),
    .RESET_B(net5898),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][16] ),
    .Q_N(_08812_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][16] ));
 sg13g2_dfrbp_1 _19431_ (.CLK(net5392),
    .RESET_B(net5901),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][17] ),
    .Q_N(_08813_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][17] ));
 sg13g2_dfrbp_1 _19432_ (.CLK(net5390),
    .RESET_B(net5899),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][18] ),
    .Q_N(_08814_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[5][18] ));
 sg13g2_dfrbp_1 _19433_ (.CLK(net5405),
    .RESET_B(net5914),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][0] ),
    .Q_N(_08815_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][0] ));
 sg13g2_dfrbp_1 _19434_ (.CLK(net5402),
    .RESET_B(net5911),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][1] ),
    .Q_N(_08816_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][1] ));
 sg13g2_dfrbp_1 _19435_ (.CLK(net5403),
    .RESET_B(net5912),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][2] ),
    .Q_N(_08817_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][2] ));
 sg13g2_dfrbp_1 _19436_ (.CLK(net5410),
    .RESET_B(net5919),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][3] ),
    .Q_N(_08818_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][3] ));
 sg13g2_dfrbp_1 _19437_ (.CLK(net5410),
    .RESET_B(net5919),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][4] ),
    .Q_N(_08819_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][4] ));
 sg13g2_dfrbp_1 _19438_ (.CLK(net5404),
    .RESET_B(net5913),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][5] ),
    .Q_N(_08820_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][5] ));
 sg13g2_dfrbp_1 _19439_ (.CLK(net5393),
    .RESET_B(net5902),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][6] ),
    .Q_N(_08821_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][6] ));
 sg13g2_dfrbp_1 _19440_ (.CLK(net5391),
    .RESET_B(net5900),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][7] ),
    .Q_N(_08822_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][7] ));
 sg13g2_dfrbp_1 _19441_ (.CLK(net5385),
    .RESET_B(net5894),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][8] ),
    .Q_N(_08823_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][8] ));
 sg13g2_dfrbp_1 _19442_ (.CLK(net5385),
    .RESET_B(net5894),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][9] ),
    .Q_N(_08824_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][9] ));
 sg13g2_dfrbp_1 _19443_ (.CLK(net5384),
    .RESET_B(net5892),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][10] ),
    .Q_N(_08825_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][10] ));
 sg13g2_dfrbp_1 _19444_ (.CLK(net5383),
    .RESET_B(net5893),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][11] ),
    .Q_N(_08826_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][11] ));
 sg13g2_dfrbp_1 _19445_ (.CLK(net5383),
    .RESET_B(net5892),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][12] ),
    .Q_N(_08827_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][12] ));
 sg13g2_dfrbp_1 _19446_ (.CLK(net5328),
    .RESET_B(net5838),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][13] ),
    .Q_N(_08828_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][13] ));
 sg13g2_dfrbp_1 _19447_ (.CLK(net5328),
    .RESET_B(net5838),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][14] ),
    .Q_N(_08829_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][14] ));
 sg13g2_dfrbp_1 _19448_ (.CLK(net5381),
    .RESET_B(net5890),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][15] ),
    .Q_N(_08830_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][15] ));
 sg13g2_dfrbp_1 _19449_ (.CLK(net5389),
    .RESET_B(net5898),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][16] ),
    .Q_N(_08831_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][16] ));
 sg13g2_dfrbp_1 _19450_ (.CLK(net5392),
    .RESET_B(net5901),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][17] ),
    .Q_N(_08832_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][17] ));
 sg13g2_dfrbp_1 _19451_ (.CLK(net5390),
    .RESET_B(net5899),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][18] ),
    .Q_N(_08833_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[4][18] ));
 sg13g2_dfrbp_1 _19452_ (.CLK(net5405),
    .RESET_B(net5914),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][0] ),
    .Q_N(_08834_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][0] ));
 sg13g2_dfrbp_1 _19453_ (.CLK(net5402),
    .RESET_B(net5911),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][1] ),
    .Q_N(_08835_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][1] ));
 sg13g2_dfrbp_1 _19454_ (.CLK(net5406),
    .RESET_B(net5915),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][2] ),
    .Q_N(_08836_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][2] ));
 sg13g2_dfrbp_1 _19455_ (.CLK(net5410),
    .RESET_B(net5919),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][3] ),
    .Q_N(_08837_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][3] ));
 sg13g2_dfrbp_1 _19456_ (.CLK(net5410),
    .RESET_B(net5919),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][4] ),
    .Q_N(_08838_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][4] ));
 sg13g2_dfrbp_1 _19457_ (.CLK(net5408),
    .RESET_B(net5917),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][5] ),
    .Q_N(_08839_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][5] ));
 sg13g2_dfrbp_1 _19458_ (.CLK(net5393),
    .RESET_B(net5902),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][6] ),
    .Q_N(_08840_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][6] ));
 sg13g2_dfrbp_1 _19459_ (.CLK(net5391),
    .RESET_B(net5900),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][7] ),
    .Q_N(_08841_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][7] ));
 sg13g2_dfrbp_1 _19460_ (.CLK(net5386),
    .RESET_B(net5895),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][8] ),
    .Q_N(_08842_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][8] ));
 sg13g2_dfrbp_1 _19461_ (.CLK(net5385),
    .RESET_B(net5894),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][9] ),
    .Q_N(_08843_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][9] ));
 sg13g2_dfrbp_1 _19462_ (.CLK(net5384),
    .RESET_B(net5892),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][10] ),
    .Q_N(_08844_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][10] ));
 sg13g2_dfrbp_1 _19463_ (.CLK(net5331),
    .RESET_B(net5841),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][11] ),
    .Q_N(_08845_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][11] ));
 sg13g2_dfrbp_1 _19464_ (.CLK(net5331),
    .RESET_B(net5841),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][12] ),
    .Q_N(_08846_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][12] ));
 sg13g2_dfrbp_1 _19465_ (.CLK(net5328),
    .RESET_B(net5838),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][13] ),
    .Q_N(_08847_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][13] ));
 sg13g2_dfrbp_1 _19466_ (.CLK(net5328),
    .RESET_B(net5838),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][14] ),
    .Q_N(_08848_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][14] ));
 sg13g2_dfrbp_1 _19467_ (.CLK(net5382),
    .RESET_B(net5891),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][15] ),
    .Q_N(_08849_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][15] ));
 sg13g2_dfrbp_1 _19468_ (.CLK(net5392),
    .RESET_B(net5901),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][16] ),
    .Q_N(_08850_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][16] ));
 sg13g2_dfrbp_1 _19469_ (.CLK(net5392),
    .RESET_B(net5901),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][17] ),
    .Q_N(_08851_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][17] ));
 sg13g2_dfrbp_1 _19470_ (.CLK(net5390),
    .RESET_B(net5899),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][18] ),
    .Q_N(_08852_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[3][18] ));
 sg13g2_dfrbp_1 _19471_ (.CLK(net5405),
    .RESET_B(net5914),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][0] ),
    .Q_N(_08853_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][0] ));
 sg13g2_dfrbp_1 _19472_ (.CLK(net5402),
    .RESET_B(net5911),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][1] ),
    .Q_N(_08854_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][1] ));
 sg13g2_dfrbp_1 _19473_ (.CLK(net5410),
    .RESET_B(net5919),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][2] ),
    .Q_N(_08855_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][2] ));
 sg13g2_dfrbp_1 _19474_ (.CLK(net5411),
    .RESET_B(net5920),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][3] ),
    .Q_N(_08856_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][3] ));
 sg13g2_dfrbp_1 _19475_ (.CLK(net5411),
    .RESET_B(net5920),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][4] ),
    .Q_N(_08857_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][4] ));
 sg13g2_dfrbp_1 _19476_ (.CLK(net5408),
    .RESET_B(net5917),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][5] ),
    .Q_N(_08858_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][5] ));
 sg13g2_dfrbp_1 _19477_ (.CLK(net5398),
    .RESET_B(net5907),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][6] ),
    .Q_N(_08859_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][6] ));
 sg13g2_dfrbp_1 _19478_ (.CLK(net5398),
    .RESET_B(net5907),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][7] ),
    .Q_N(_08860_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][7] ));
 sg13g2_dfrbp_1 _19479_ (.CLK(net5397),
    .RESET_B(net5906),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][8] ),
    .Q_N(_08861_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][8] ));
 sg13g2_dfrbp_1 _19480_ (.CLK(net5331),
    .RESET_B(net5841),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][9] ),
    .Q_N(_08862_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][9] ));
 sg13g2_dfrbp_1 _19481_ (.CLK(net5385),
    .RESET_B(net5894),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][10] ),
    .Q_N(_08863_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][10] ));
 sg13g2_dfrbp_1 _19482_ (.CLK(net5331),
    .RESET_B(net5841),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][11] ),
    .Q_N(_08864_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][11] ));
 sg13g2_dfrbp_1 _19483_ (.CLK(net5331),
    .RESET_B(net5841),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][12] ),
    .Q_N(_08865_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][12] ));
 sg13g2_dfrbp_1 _19484_ (.CLK(net5329),
    .RESET_B(net5839),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][13] ),
    .Q_N(_08866_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][13] ));
 sg13g2_dfrbp_1 _19485_ (.CLK(net5329),
    .RESET_B(net5839),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][14] ),
    .Q_N(_08867_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][14] ));
 sg13g2_dfrbp_1 _19486_ (.CLK(net5328),
    .RESET_B(net5838),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][15] ),
    .Q_N(_08868_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][15] ));
 sg13g2_dfrbp_1 _19487_ (.CLK(net5390),
    .RESET_B(net5899),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][16] ),
    .Q_N(_08869_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][16] ));
 sg13g2_dfrbp_1 _19488_ (.CLK(net5390),
    .RESET_B(net5899),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][17] ),
    .Q_N(_08870_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][17] ));
 sg13g2_dfrbp_1 _19489_ (.CLK(net5391),
    .RESET_B(net5900),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][18] ),
    .Q_N(_08871_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[2][18] ));
 sg13g2_dfrbp_1 _19490_ (.CLK(net5402),
    .RESET_B(net5911),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][0] ),
    .Q_N(_08872_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][0] ));
 sg13g2_dfrbp_1 _19491_ (.CLK(net5403),
    .RESET_B(net5912),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][1] ),
    .Q_N(_08873_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][1] ));
 sg13g2_dfrbp_1 _19492_ (.CLK(net5408),
    .RESET_B(net5917),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][2] ),
    .Q_N(_08874_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][2] ));
 sg13g2_dfrbp_1 _19493_ (.CLK(net5408),
    .RESET_B(net5917),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][3] ),
    .Q_N(_08875_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][3] ));
 sg13g2_dfrbp_1 _19494_ (.CLK(net5411),
    .RESET_B(net5920),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][4] ),
    .Q_N(_08876_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][4] ));
 sg13g2_dfrbp_1 _19495_ (.CLK(net5409),
    .RESET_B(net5918),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][5] ),
    .Q_N(_08877_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][5] ));
 sg13g2_dfrbp_1 _19496_ (.CLK(net5398),
    .RESET_B(net5907),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][6] ),
    .Q_N(_08878_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][6] ));
 sg13g2_dfrbp_1 _19497_ (.CLK(net5398),
    .RESET_B(net5907),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][7] ),
    .Q_N(_08879_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][7] ));
 sg13g2_dfrbp_1 _19498_ (.CLK(net5397),
    .RESET_B(net5906),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][8] ),
    .Q_N(_08880_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][8] ));
 sg13g2_dfrbp_1 _19499_ (.CLK(net5337),
    .RESET_B(net5847),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][9] ),
    .Q_N(_08881_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][9] ));
 sg13g2_dfrbp_1 _19500_ (.CLK(net5331),
    .RESET_B(net5841),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][10] ),
    .Q_N(_08882_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][10] ));
 sg13g2_dfrbp_1 _19501_ (.CLK(net5331),
    .RESET_B(net5841),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][11] ),
    .Q_N(_08883_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][11] ));
 sg13g2_dfrbp_1 _19502_ (.CLK(net5332),
    .RESET_B(net5842),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][12] ),
    .Q_N(_08884_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][12] ));
 sg13g2_dfrbp_1 _19503_ (.CLK(net5330),
    .RESET_B(net5840),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][13] ),
    .Q_N(_08885_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][13] ));
 sg13g2_dfrbp_1 _19504_ (.CLK(net5330),
    .RESET_B(net5840),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][14] ),
    .Q_N(_08886_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][14] ));
 sg13g2_dfrbp_1 _19505_ (.CLK(net5329),
    .RESET_B(net5839),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][15] ),
    .Q_N(_08887_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][15] ));
 sg13g2_dfrbp_1 _19506_ (.CLK(net5390),
    .RESET_B(net5899),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][16] ),
    .Q_N(_08888_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][16] ));
 sg13g2_dfrbp_1 _19507_ (.CLK(net5391),
    .RESET_B(net5900),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][17] ),
    .Q_N(_08889_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][17] ));
 sg13g2_dfrbp_1 _19508_ (.CLK(net5387),
    .RESET_B(net5896),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][18] ),
    .Q_N(_08890_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[1][18] ));
 sg13g2_dfrbp_1 _19509_ (.CLK(net5403),
    .RESET_B(net5912),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.u_mux_shift.sum_res ),
    .Q_N(_00292_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][0] ));
 sg13g2_dfrbp_1 _19510_ (.CLK(net5403),
    .RESET_B(net5912),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .Q_N(_00296_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][1] ));
 sg13g2_dfrbp_1 _19511_ (.CLK(net5408),
    .RESET_B(net5917),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .Q_N(_00303_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][2] ));
 sg13g2_dfrbp_1 _19512_ (.CLK(net5409),
    .RESET_B(net5918),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .Q_N(_00310_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][3] ));
 sg13g2_dfrbp_1 _19513_ (.CLK(net5409),
    .RESET_B(net5918),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .Q_N(_00319_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][4] ));
 sg13g2_dfrbp_1 _19514_ (.CLK(net5409),
    .RESET_B(net5918),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .Q_N(_00328_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][5] ));
 sg13g2_dfrbp_1 _19515_ (.CLK(net5399),
    .RESET_B(net5908),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .Q_N(_00335_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][6] ));
 sg13g2_dfrbp_1 _19516_ (.CLK(net5398),
    .RESET_B(net5907),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .Q_N(_00342_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][7] ));
 sg13g2_dfrbp_1 _19517_ (.CLK(net5397),
    .RESET_B(net5906),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .Q_N(_00351_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][8] ));
 sg13g2_dfrbp_1 _19518_ (.CLK(net5337),
    .RESET_B(net5847),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .Q_N(_00360_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][9] ));
 sg13g2_dfrbp_1 _19519_ (.CLK(net5332),
    .RESET_B(net5841),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .Q_N(_00367_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][10] ));
 sg13g2_dfrbp_1 _19520_ (.CLK(net5331),
    .RESET_B(net5842),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .Q_N(_00374_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][11] ));
 sg13g2_dfrbp_1 _19521_ (.CLK(net5332),
    .RESET_B(net5842),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .Q_N(_00383_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][12] ));
 sg13g2_dfrbp_1 _19522_ (.CLK(net5330),
    .RESET_B(net5840),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .Q_N(_00392_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][13] ));
 sg13g2_dfrbp_1 _19523_ (.CLK(net5330),
    .RESET_B(net5840),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .Q_N(_00399_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][14] ));
 sg13g2_dfrbp_1 _19524_ (.CLK(net5330),
    .RESET_B(net5840),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .Q_N(_00406_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][15] ));
 sg13g2_dfrbp_1 _19525_ (.CLK(net5387),
    .RESET_B(net5896),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .Q_N(_00415_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][16] ));
 sg13g2_dfrbp_1 _19526_ (.CLK(net5387),
    .RESET_B(net5896),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .Q_N(_00422_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][17] ));
 sg13g2_dfrbp_1 _19527_ (.CLK(net5387),
    .RESET_B(net5896),
    .D(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .Q_N(_00429_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[3].u_delay_line.buffer[0][18] ));
 sg13g2_dfrbp_1 _19528_ (.CLK(net5465),
    .RESET_B(net5974),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][0] ),
    .Q_N(_08891_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][0] ));
 sg13g2_dfrbp_1 _19529_ (.CLK(net5469),
    .RESET_B(net5978),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][1] ),
    .Q_N(_08892_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][1] ));
 sg13g2_dfrbp_1 _19530_ (.CLK(net5467),
    .RESET_B(net5976),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][2] ),
    .Q_N(_08893_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][2] ));
 sg13g2_dfrbp_1 _19531_ (.CLK(net5513),
    .RESET_B(net6022),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][3] ),
    .Q_N(_08894_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][3] ));
 sg13g2_dfrbp_1 _19532_ (.CLK(net5520),
    .RESET_B(net6029),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][4] ),
    .Q_N(_08895_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][4] ));
 sg13g2_dfrbp_1 _19533_ (.CLK(net5518),
    .RESET_B(net6027),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][5] ),
    .Q_N(_08896_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][5] ));
 sg13g2_dfrbp_1 _19534_ (.CLK(net5539),
    .RESET_B(net6048),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][6] ),
    .Q_N(_08897_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][6] ));
 sg13g2_dfrbp_1 _19535_ (.CLK(net5543),
    .RESET_B(net6052),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][7] ),
    .Q_N(_08898_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][7] ));
 sg13g2_dfrbp_1 _19536_ (.CLK(net5544),
    .RESET_B(net6053),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][8] ),
    .Q_N(_08899_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][8] ));
 sg13g2_dfrbp_1 _19537_ (.CLK(net5547),
    .RESET_B(net6055),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][9] ),
    .Q_N(_08900_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][9] ));
 sg13g2_dfrbp_1 _19538_ (.CLK(net5551),
    .RESET_B(net6060),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][10] ),
    .Q_N(_08901_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][10] ));
 sg13g2_dfrbp_1 _19539_ (.CLK(net5552),
    .RESET_B(net6061),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][11] ),
    .Q_N(_08902_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][11] ));
 sg13g2_dfrbp_1 _19540_ (.CLK(net5549),
    .RESET_B(net6058),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][12] ),
    .Q_N(_08903_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][12] ));
 sg13g2_dfrbp_1 _19541_ (.CLK(net5541),
    .RESET_B(net6050),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][13] ),
    .Q_N(_08904_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][13] ));
 sg13g2_dfrbp_1 _19542_ (.CLK(net5522),
    .RESET_B(net6031),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][14] ),
    .Q_N(_08905_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][14] ));
 sg13g2_dfrbp_1 _19543_ (.CLK(net5450),
    .RESET_B(net5959),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][15] ),
    .Q_N(_08906_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][15] ));
 sg13g2_dfrbp_1 _19544_ (.CLK(net5448),
    .RESET_B(net5957),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][16] ),
    .Q_N(_08907_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][16] ));
 sg13g2_dfrbp_1 _19545_ (.CLK(net5444),
    .RESET_B(net5953),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][17] ),
    .Q_N(_08908_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][17] ));
 sg13g2_dfrbp_1 _19546_ (.CLK(net5446),
    .RESET_B(net5955),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][18] ),
    .Q_N(_08909_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][18] ));
 sg13g2_dfrbp_1 _19547_ (.CLK(net5465),
    .RESET_B(net5974),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][0] ),
    .Q_N(_08910_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][0] ));
 sg13g2_dfrbp_1 _19548_ (.CLK(net5469),
    .RESET_B(net5978),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][1] ),
    .Q_N(_08911_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][1] ));
 sg13g2_dfrbp_1 _19549_ (.CLK(net5467),
    .RESET_B(net5976),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][2] ),
    .Q_N(_08912_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][2] ));
 sg13g2_dfrbp_1 _19550_ (.CLK(net5513),
    .RESET_B(net6022),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][3] ),
    .Q_N(_08913_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][3] ));
 sg13g2_dfrbp_1 _19551_ (.CLK(net5521),
    .RESET_B(net6030),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][4] ),
    .Q_N(_08914_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][4] ));
 sg13g2_dfrbp_1 _19552_ (.CLK(net5518),
    .RESET_B(net6027),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][5] ),
    .Q_N(_08915_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][5] ));
 sg13g2_dfrbp_1 _19553_ (.CLK(net5539),
    .RESET_B(net6048),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][6] ),
    .Q_N(_08916_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][6] ));
 sg13g2_dfrbp_1 _19554_ (.CLK(net5543),
    .RESET_B(net6052),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][7] ),
    .Q_N(_08917_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][7] ));
 sg13g2_dfrbp_1 _19555_ (.CLK(net5544),
    .RESET_B(net6053),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][8] ),
    .Q_N(_08918_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][8] ));
 sg13g2_dfrbp_1 _19556_ (.CLK(net5546),
    .RESET_B(net6057),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][9] ),
    .Q_N(_08919_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][9] ));
 sg13g2_dfrbp_1 _19557_ (.CLK(net5551),
    .RESET_B(net6060),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][10] ),
    .Q_N(_08920_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][10] ));
 sg13g2_dfrbp_1 _19558_ (.CLK(net5552),
    .RESET_B(net6062),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][11] ),
    .Q_N(_08921_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][11] ));
 sg13g2_dfrbp_1 _19559_ (.CLK(net5549),
    .RESET_B(net6058),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][12] ),
    .Q_N(_08922_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][12] ));
 sg13g2_dfrbp_1 _19560_ (.CLK(net5541),
    .RESET_B(net6050),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][13] ),
    .Q_N(_08923_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][13] ));
 sg13g2_dfrbp_1 _19561_ (.CLK(net5523),
    .RESET_B(net6031),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][14] ),
    .Q_N(_08924_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][14] ));
 sg13g2_dfrbp_1 _19562_ (.CLK(net5449),
    .RESET_B(net5958),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][15] ),
    .Q_N(_08925_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][15] ));
 sg13g2_dfrbp_1 _19563_ (.CLK(net5448),
    .RESET_B(net5957),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][16] ),
    .Q_N(_08926_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][16] ));
 sg13g2_dfrbp_1 _19564_ (.CLK(net5444),
    .RESET_B(net5953),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][17] ),
    .Q_N(_08927_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][17] ));
 sg13g2_dfrbp_1 _19565_ (.CLK(net5446),
    .RESET_B(net5955),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][18] ),
    .Q_N(_08928_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[6][18] ));
 sg13g2_dfrbp_1 _19566_ (.CLK(net5465),
    .RESET_B(net5974),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][0] ),
    .Q_N(_08929_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][0] ));
 sg13g2_dfrbp_1 _19567_ (.CLK(net5469),
    .RESET_B(net5979),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][1] ),
    .Q_N(_08930_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][1] ));
 sg13g2_dfrbp_1 _19568_ (.CLK(net5467),
    .RESET_B(net5976),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][2] ),
    .Q_N(_08931_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][2] ));
 sg13g2_dfrbp_1 _19569_ (.CLK(net5514),
    .RESET_B(net6022),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][3] ),
    .Q_N(_08932_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][3] ));
 sg13g2_dfrbp_1 _19570_ (.CLK(net5520),
    .RESET_B(net6029),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][4] ),
    .Q_N(_08933_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][4] ));
 sg13g2_dfrbp_1 _19571_ (.CLK(net5518),
    .RESET_B(net6027),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][5] ),
    .Q_N(_08934_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][5] ));
 sg13g2_dfrbp_1 _19572_ (.CLK(net5539),
    .RESET_B(net6048),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][6] ),
    .Q_N(_08935_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][6] ));
 sg13g2_dfrbp_1 _19573_ (.CLK(net5543),
    .RESET_B(net6052),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][7] ),
    .Q_N(_08936_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][7] ));
 sg13g2_dfrbp_1 _19574_ (.CLK(net5548),
    .RESET_B(net6052),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][8] ),
    .Q_N(_08937_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][8] ));
 sg13g2_dfrbp_1 _19575_ (.CLK(net5546),
    .RESET_B(net6055),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][9] ),
    .Q_N(_08938_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][9] ));
 sg13g2_dfrbp_1 _19576_ (.CLK(net5551),
    .RESET_B(net6060),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][10] ),
    .Q_N(_08939_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][10] ));
 sg13g2_dfrbp_1 _19577_ (.CLK(net5552),
    .RESET_B(net6061),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][11] ),
    .Q_N(_08940_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][11] ));
 sg13g2_dfrbp_1 _19578_ (.CLK(net5549),
    .RESET_B(net6058),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][12] ),
    .Q_N(_08941_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][12] ));
 sg13g2_dfrbp_1 _19579_ (.CLK(net5541),
    .RESET_B(net6050),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][13] ),
    .Q_N(_08942_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][13] ));
 sg13g2_dfrbp_1 _19580_ (.CLK(net5522),
    .RESET_B(net6031),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][14] ),
    .Q_N(_08943_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][14] ));
 sg13g2_dfrbp_1 _19581_ (.CLK(net5450),
    .RESET_B(net5959),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][15] ),
    .Q_N(_08944_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][15] ));
 sg13g2_dfrbp_1 _19582_ (.CLK(net5448),
    .RESET_B(net5957),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][16] ),
    .Q_N(_08945_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][16] ));
 sg13g2_dfrbp_1 _19583_ (.CLK(net5444),
    .RESET_B(net5953),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][17] ),
    .Q_N(_08946_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][17] ));
 sg13g2_dfrbp_1 _19584_ (.CLK(net5446),
    .RESET_B(net5955),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][18] ),
    .Q_N(_08947_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][18] ));
 sg13g2_dfrbp_1 _19585_ (.CLK(net5465),
    .RESET_B(net5974),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][0] ),
    .Q_N(_08948_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][0] ));
 sg13g2_dfrbp_1 _19586_ (.CLK(net5469),
    .RESET_B(net5978),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][1] ),
    .Q_N(_08949_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][1] ));
 sg13g2_dfrbp_1 _19587_ (.CLK(net5467),
    .RESET_B(net5976),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][2] ),
    .Q_N(_08950_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][2] ));
 sg13g2_dfrbp_1 _19588_ (.CLK(net5514),
    .RESET_B(net6023),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][3] ),
    .Q_N(_08951_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][3] ));
 sg13g2_dfrbp_1 _19589_ (.CLK(net5520),
    .RESET_B(net6029),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][4] ),
    .Q_N(_08952_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][4] ));
 sg13g2_dfrbp_1 _19590_ (.CLK(net5518),
    .RESET_B(net6027),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][5] ),
    .Q_N(_08953_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][5] ));
 sg13g2_dfrbp_1 _19591_ (.CLK(net5539),
    .RESET_B(net6048),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][6] ),
    .Q_N(_08954_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][6] ));
 sg13g2_dfrbp_1 _19592_ (.CLK(net5543),
    .RESET_B(net6052),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][7] ),
    .Q_N(_08955_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][7] ));
 sg13g2_dfrbp_1 _19593_ (.CLK(net5544),
    .RESET_B(net6053),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][8] ),
    .Q_N(_08956_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][8] ));
 sg13g2_dfrbp_1 _19594_ (.CLK(net5546),
    .RESET_B(net6055),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][9] ),
    .Q_N(_08957_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][9] ));
 sg13g2_dfrbp_1 _19595_ (.CLK(net5551),
    .RESET_B(net6060),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][10] ),
    .Q_N(_08958_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][10] ));
 sg13g2_dfrbp_1 _19596_ (.CLK(net5552),
    .RESET_B(net6062),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][11] ),
    .Q_N(_08959_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][11] ));
 sg13g2_dfrbp_1 _19597_ (.CLK(net5549),
    .RESET_B(net6058),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][12] ),
    .Q_N(_08960_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][12] ));
 sg13g2_dfrbp_1 _19598_ (.CLK(net5541),
    .RESET_B(net6050),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][13] ),
    .Q_N(_08961_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][13] ));
 sg13g2_dfrbp_1 _19599_ (.CLK(net5522),
    .RESET_B(net6031),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][14] ),
    .Q_N(_08962_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][14] ));
 sg13g2_dfrbp_1 _19600_ (.CLK(net5450),
    .RESET_B(net5959),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][15] ),
    .Q_N(_08963_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][15] ));
 sg13g2_dfrbp_1 _19601_ (.CLK(net5448),
    .RESET_B(net5957),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][16] ),
    .Q_N(_08964_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][16] ));
 sg13g2_dfrbp_1 _19602_ (.CLK(net5444),
    .RESET_B(net5953),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][17] ),
    .Q_N(_08965_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][17] ));
 sg13g2_dfrbp_1 _19603_ (.CLK(net5447),
    .RESET_B(net5956),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][18] ),
    .Q_N(_08966_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[5][18] ));
 sg13g2_dfrbp_1 _19604_ (.CLK(net5465),
    .RESET_B(net5974),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][0] ),
    .Q_N(_08967_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][0] ));
 sg13g2_dfrbp_1 _19605_ (.CLK(net5469),
    .RESET_B(net5978),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][1] ),
    .Q_N(_08968_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][1] ));
 sg13g2_dfrbp_1 _19606_ (.CLK(net5467),
    .RESET_B(net5976),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][2] ),
    .Q_N(_08969_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][2] ));
 sg13g2_dfrbp_1 _19607_ (.CLK(net5514),
    .RESET_B(net6023),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][3] ),
    .Q_N(_08970_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][3] ));
 sg13g2_dfrbp_1 _19608_ (.CLK(net5520),
    .RESET_B(net6029),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][4] ),
    .Q_N(_08971_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][4] ));
 sg13g2_dfrbp_1 _19609_ (.CLK(net5518),
    .RESET_B(net6027),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][5] ),
    .Q_N(_08972_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][5] ));
 sg13g2_dfrbp_1 _19610_ (.CLK(net5539),
    .RESET_B(net6048),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][6] ),
    .Q_N(_08973_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][6] ));
 sg13g2_dfrbp_1 _19611_ (.CLK(net5543),
    .RESET_B(net6052),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][7] ),
    .Q_N(_08974_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][7] ));
 sg13g2_dfrbp_1 _19612_ (.CLK(net5544),
    .RESET_B(net6053),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][8] ),
    .Q_N(_08975_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][8] ));
 sg13g2_dfrbp_1 _19613_ (.CLK(net5548),
    .RESET_B(net6055),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][9] ),
    .Q_N(_08976_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][9] ));
 sg13g2_dfrbp_1 _19614_ (.CLK(net5552),
    .RESET_B(net6061),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][10] ),
    .Q_N(_08977_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][10] ));
 sg13g2_dfrbp_1 _19615_ (.CLK(net5553),
    .RESET_B(net6061),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][11] ),
    .Q_N(_08978_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][11] ));
 sg13g2_dfrbp_1 _19616_ (.CLK(net5549),
    .RESET_B(net6058),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][12] ),
    .Q_N(_08979_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][12] ));
 sg13g2_dfrbp_1 _19617_ (.CLK(net5541),
    .RESET_B(net6050),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][13] ),
    .Q_N(_08980_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][13] ));
 sg13g2_dfrbp_1 _19618_ (.CLK(net5522),
    .RESET_B(net6032),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][14] ),
    .Q_N(_08981_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][14] ));
 sg13g2_dfrbp_1 _19619_ (.CLK(net5450),
    .RESET_B(net5959),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][15] ),
    .Q_N(_08982_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][15] ));
 sg13g2_dfrbp_1 _19620_ (.CLK(net5448),
    .RESET_B(net5957),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][16] ),
    .Q_N(_08983_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][16] ));
 sg13g2_dfrbp_1 _19621_ (.CLK(net5444),
    .RESET_B(net5953),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][17] ),
    .Q_N(_08984_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][17] ));
 sg13g2_dfrbp_1 _19622_ (.CLK(net5446),
    .RESET_B(net5955),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][18] ),
    .Q_N(_08985_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[4][18] ));
 sg13g2_dfrbp_1 _19623_ (.CLK(net5465),
    .RESET_B(net5974),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][0] ),
    .Q_N(_08986_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][0] ));
 sg13g2_dfrbp_1 _19624_ (.CLK(net5469),
    .RESET_B(net5978),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][1] ),
    .Q_N(_08987_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][1] ));
 sg13g2_dfrbp_1 _19625_ (.CLK(net5467),
    .RESET_B(net5976),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][2] ),
    .Q_N(_08988_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][2] ));
 sg13g2_dfrbp_1 _19626_ (.CLK(net5513),
    .RESET_B(net6022),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][3] ),
    .Q_N(_08989_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][3] ));
 sg13g2_dfrbp_1 _19627_ (.CLK(net5520),
    .RESET_B(net6029),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][4] ),
    .Q_N(_08990_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][4] ));
 sg13g2_dfrbp_1 _19628_ (.CLK(net5518),
    .RESET_B(net6027),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][5] ),
    .Q_N(_08991_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][5] ));
 sg13g2_dfrbp_1 _19629_ (.CLK(net5539),
    .RESET_B(net6048),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][6] ),
    .Q_N(_08992_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][6] ));
 sg13g2_dfrbp_1 _19630_ (.CLK(net5545),
    .RESET_B(net6054),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][7] ),
    .Q_N(_08993_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][7] ));
 sg13g2_dfrbp_1 _19631_ (.CLK(net5544),
    .RESET_B(net6053),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][8] ),
    .Q_N(_08994_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][8] ));
 sg13g2_dfrbp_1 _19632_ (.CLK(net5546),
    .RESET_B(net6056),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][9] ),
    .Q_N(_08995_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][9] ));
 sg13g2_dfrbp_1 _19633_ (.CLK(net5552),
    .RESET_B(net6060),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][10] ),
    .Q_N(_08996_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][10] ));
 sg13g2_dfrbp_1 _19634_ (.CLK(net5553),
    .RESET_B(net6061),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][11] ),
    .Q_N(_08997_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][11] ));
 sg13g2_dfrbp_1 _19635_ (.CLK(net5549),
    .RESET_B(net6058),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][12] ),
    .Q_N(_08998_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][12] ));
 sg13g2_dfrbp_1 _19636_ (.CLK(net5542),
    .RESET_B(net6051),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][13] ),
    .Q_N(_08999_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][13] ));
 sg13g2_dfrbp_1 _19637_ (.CLK(net5522),
    .RESET_B(net6031),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][14] ),
    .Q_N(_09000_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][14] ));
 sg13g2_dfrbp_1 _19638_ (.CLK(net5451),
    .RESET_B(net5960),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][15] ),
    .Q_N(_09001_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][15] ));
 sg13g2_dfrbp_1 _19639_ (.CLK(net5448),
    .RESET_B(net5957),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][16] ),
    .Q_N(_09002_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][16] ));
 sg13g2_dfrbp_1 _19640_ (.CLK(net5444),
    .RESET_B(net5953),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][17] ),
    .Q_N(_09003_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][17] ));
 sg13g2_dfrbp_1 _19641_ (.CLK(net5446),
    .RESET_B(net5955),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][18] ),
    .Q_N(_09004_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[3][18] ));
 sg13g2_dfrbp_1 _19642_ (.CLK(net5466),
    .RESET_B(net5975),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][0] ),
    .Q_N(_09005_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][0] ));
 sg13g2_dfrbp_1 _19643_ (.CLK(net5469),
    .RESET_B(net5978),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][1] ),
    .Q_N(_09006_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][1] ));
 sg13g2_dfrbp_1 _19644_ (.CLK(net5467),
    .RESET_B(net5976),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][2] ),
    .Q_N(_09007_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][2] ));
 sg13g2_dfrbp_1 _19645_ (.CLK(net5513),
    .RESET_B(net6022),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][3] ),
    .Q_N(_09008_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][3] ));
 sg13g2_dfrbp_1 _19646_ (.CLK(net5520),
    .RESET_B(net6029),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][4] ),
    .Q_N(_09009_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][4] ));
 sg13g2_dfrbp_1 _19647_ (.CLK(net5519),
    .RESET_B(net6028),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][5] ),
    .Q_N(_09010_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][5] ));
 sg13g2_dfrbp_1 _19648_ (.CLK(net5519),
    .RESET_B(net6028),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][6] ),
    .Q_N(_09011_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][6] ));
 sg13g2_dfrbp_1 _19649_ (.CLK(net5545),
    .RESET_B(net6054),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][7] ),
    .Q_N(_09012_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][7] ));
 sg13g2_dfrbp_1 _19650_ (.CLK(net5544),
    .RESET_B(net6053),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][8] ),
    .Q_N(_09013_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][8] ));
 sg13g2_dfrbp_1 _19651_ (.CLK(net5546),
    .RESET_B(net6055),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][9] ),
    .Q_N(_09014_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][9] ));
 sg13g2_dfrbp_1 _19652_ (.CLK(net5551),
    .RESET_B(net6060),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][10] ),
    .Q_N(_09015_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][10] ));
 sg13g2_dfrbp_1 _19653_ (.CLK(net5553),
    .RESET_B(net6062),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][11] ),
    .Q_N(_09016_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][11] ));
 sg13g2_dfrbp_1 _19654_ (.CLK(net5549),
    .RESET_B(net6058),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][12] ),
    .Q_N(_09017_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][12] ));
 sg13g2_dfrbp_1 _19655_ (.CLK(net5542),
    .RESET_B(net6051),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][13] ),
    .Q_N(_09018_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][13] ));
 sg13g2_dfrbp_1 _19656_ (.CLK(net5522),
    .RESET_B(net6031),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][14] ),
    .Q_N(_09019_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][14] ));
 sg13g2_dfrbp_1 _19657_ (.CLK(net5450),
    .RESET_B(net5959),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][15] ),
    .Q_N(_09020_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][15] ));
 sg13g2_dfrbp_1 _19658_ (.CLK(net5449),
    .RESET_B(net5958),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][16] ),
    .Q_N(_09021_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][16] ));
 sg13g2_dfrbp_1 _19659_ (.CLK(net5445),
    .RESET_B(net5954),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][17] ),
    .Q_N(_09022_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][17] ));
 sg13g2_dfrbp_1 _19660_ (.CLK(net5446),
    .RESET_B(net5955),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][18] ),
    .Q_N(_09023_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[2][18] ));
 sg13g2_dfrbp_1 _19661_ (.CLK(net5465),
    .RESET_B(net5974),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][0] ),
    .Q_N(_09024_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][0] ));
 sg13g2_dfrbp_1 _19662_ (.CLK(net5469),
    .RESET_B(net5978),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][1] ),
    .Q_N(_09025_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][1] ));
 sg13g2_dfrbp_1 _19663_ (.CLK(net5467),
    .RESET_B(net5976),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][2] ),
    .Q_N(_09026_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][2] ));
 sg13g2_dfrbp_1 _19664_ (.CLK(net5513),
    .RESET_B(net6022),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][3] ),
    .Q_N(_09027_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][3] ));
 sg13g2_dfrbp_1 _19665_ (.CLK(net5520),
    .RESET_B(net6029),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][4] ),
    .Q_N(_09028_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][4] ));
 sg13g2_dfrbp_1 _19666_ (.CLK(net5518),
    .RESET_B(net6027),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][5] ),
    .Q_N(_09029_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][5] ));
 sg13g2_dfrbp_1 _19667_ (.CLK(net5539),
    .RESET_B(net6048),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][6] ),
    .Q_N(_09030_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][6] ));
 sg13g2_dfrbp_1 _19668_ (.CLK(net5543),
    .RESET_B(net6052),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][7] ),
    .Q_N(_09031_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][7] ));
 sg13g2_dfrbp_1 _19669_ (.CLK(net5548),
    .RESET_B(net6057),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][8] ),
    .Q_N(_09032_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][8] ));
 sg13g2_dfrbp_1 _19670_ (.CLK(net5546),
    .RESET_B(net6055),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][9] ),
    .Q_N(_09033_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][9] ));
 sg13g2_dfrbp_1 _19671_ (.CLK(net5551),
    .RESET_B(net6060),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][10] ),
    .Q_N(_09034_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][10] ));
 sg13g2_dfrbp_1 _19672_ (.CLK(net5552),
    .RESET_B(net6061),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][11] ),
    .Q_N(_09035_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][11] ));
 sg13g2_dfrbp_1 _19673_ (.CLK(net5549),
    .RESET_B(net6058),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][12] ),
    .Q_N(_09036_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][12] ));
 sg13g2_dfrbp_1 _19674_ (.CLK(net5541),
    .RESET_B(net6050),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][13] ),
    .Q_N(_09037_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][13] ));
 sg13g2_dfrbp_1 _19675_ (.CLK(net5522),
    .RESET_B(net6031),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][14] ),
    .Q_N(_09038_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][14] ));
 sg13g2_dfrbp_1 _19676_ (.CLK(net5450),
    .RESET_B(net5959),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][15] ),
    .Q_N(_09039_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][15] ));
 sg13g2_dfrbp_1 _19677_ (.CLK(net5448),
    .RESET_B(net5957),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][16] ),
    .Q_N(_09040_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][16] ));
 sg13g2_dfrbp_1 _19678_ (.CLK(net5444),
    .RESET_B(net5953),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][17] ),
    .Q_N(_09041_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][17] ));
 sg13g2_dfrbp_1 _19679_ (.CLK(net5446),
    .RESET_B(net5955),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[7][18] ),
    .Q_N(_09042_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[8][18] ));
 sg13g2_dfrbp_1 _19680_ (.CLK(net5466),
    .RESET_B(net5975),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][0] ),
    .Q_N(_09043_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][0] ));
 sg13g2_dfrbp_1 _19681_ (.CLK(net5468),
    .RESET_B(net5977),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][1] ),
    .Q_N(_09044_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][1] ));
 sg13g2_dfrbp_1 _19682_ (.CLK(net5468),
    .RESET_B(net5977),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][2] ),
    .Q_N(_09045_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][2] ));
 sg13g2_dfrbp_1 _19683_ (.CLK(net5513),
    .RESET_B(net6022),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][3] ),
    .Q_N(_09046_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][3] ));
 sg13g2_dfrbp_1 _19684_ (.CLK(net5521),
    .RESET_B(net6030),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][4] ),
    .Q_N(_09047_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][4] ));
 sg13g2_dfrbp_1 _19685_ (.CLK(net5518),
    .RESET_B(net6027),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][5] ),
    .Q_N(_09048_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][5] ));
 sg13g2_dfrbp_1 _19686_ (.CLK(net5519),
    .RESET_B(net6028),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][6] ),
    .Q_N(_09049_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][6] ));
 sg13g2_dfrbp_1 _19687_ (.CLK(net5540),
    .RESET_B(net6049),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][7] ),
    .Q_N(_09050_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][7] ));
 sg13g2_dfrbp_1 _19688_ (.CLK(net5540),
    .RESET_B(net6049),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][8] ),
    .Q_N(_09051_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][8] ));
 sg13g2_dfrbp_1 _19689_ (.CLK(net5543),
    .RESET_B(net6052),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][9] ),
    .Q_N(_09052_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][9] ));
 sg13g2_dfrbp_1 _19690_ (.CLK(net5550),
    .RESET_B(net6059),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][10] ),
    .Q_N(_09053_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][10] ));
 sg13g2_dfrbp_1 _19691_ (.CLK(net5550),
    .RESET_B(net6059),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][11] ),
    .Q_N(_09054_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][11] ));
 sg13g2_dfrbp_1 _19692_ (.CLK(net5542),
    .RESET_B(net6051),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][12] ),
    .Q_N(_09055_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][12] ));
 sg13g2_dfrbp_1 _19693_ (.CLK(net5542),
    .RESET_B(net6051),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][13] ),
    .Q_N(_09056_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][13] ));
 sg13g2_dfrbp_1 _19694_ (.CLK(net5523),
    .RESET_B(net6032),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][14] ),
    .Q_N(_09057_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][14] ));
 sg13g2_dfrbp_1 _19695_ (.CLK(net5449),
    .RESET_B(net5958),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][15] ),
    .Q_N(_09058_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][15] ));
 sg13g2_dfrbp_1 _19696_ (.CLK(net5449),
    .RESET_B(net5958),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][16] ),
    .Q_N(_09059_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][16] ));
 sg13g2_dfrbp_1 _19697_ (.CLK(net5445),
    .RESET_B(net5954),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][17] ),
    .Q_N(_09060_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][17] ));
 sg13g2_dfrbp_1 _19698_ (.CLK(net5447),
    .RESET_B(net5956),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][18] ),
    .Q_N(_09061_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[1][18] ));
 sg13g2_dfrbp_1 _19699_ (.CLK(net5471),
    .RESET_B(net5980),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.u_mux_shift.sum_res ),
    .Q_N(_09062_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][0] ));
 sg13g2_dfrbp_1 _19700_ (.CLK(net5466),
    .RESET_B(net5975),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .Q_N(_00297_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][1] ));
 sg13g2_dfrbp_1 _19701_ (.CLK(net5466),
    .RESET_B(net5975),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .Q_N(_00304_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][2] ));
 sg13g2_dfrbp_1 _19702_ (.CLK(net5513),
    .RESET_B(net6022),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .Q_N(_00311_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][3] ));
 sg13g2_dfrbp_1 _19703_ (.CLK(net5517),
    .RESET_B(net6026),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .Q_N(_00320_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][4] ));
 sg13g2_dfrbp_1 _19704_ (.CLK(net5516),
    .RESET_B(net6025),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .Q_N(_00329_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][5] ));
 sg13g2_dfrbp_1 _19705_ (.CLK(net5519),
    .RESET_B(net6028),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .Q_N(_00336_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][6] ));
 sg13g2_dfrbp_1 _19706_ (.CLK(net5540),
    .RESET_B(net6049),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .Q_N(_00343_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][7] ));
 sg13g2_dfrbp_1 _19707_ (.CLK(net5540),
    .RESET_B(net6049),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .Q_N(_00352_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][8] ));
 sg13g2_dfrbp_1 _19708_ (.CLK(net5544),
    .RESET_B(net6053),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .Q_N(_00361_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][9] ));
 sg13g2_dfrbp_1 _19709_ (.CLK(net5550),
    .RESET_B(net6059),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .Q_N(_00368_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][10] ));
 sg13g2_dfrbp_1 _19710_ (.CLK(net5550),
    .RESET_B(net6059),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .Q_N(_00375_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][11] ));
 sg13g2_dfrbp_1 _19711_ (.CLK(net5541),
    .RESET_B(net6050),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .Q_N(_00384_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][12] ));
 sg13g2_dfrbp_1 _19712_ (.CLK(net5522),
    .RESET_B(net6031),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .Q_N(_00393_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][13] ));
 sg13g2_dfrbp_1 _19713_ (.CLK(net5521),
    .RESET_B(net6030),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .Q_N(_00400_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][14] ));
 sg13g2_dfrbp_1 _19714_ (.CLK(net5452),
    .RESET_B(net5961),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .Q_N(_00407_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][15] ));
 sg13g2_dfrbp_1 _19715_ (.CLK(net5445),
    .RESET_B(net5954),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .Q_N(_00416_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][16] ));
 sg13g2_dfrbp_1 _19716_ (.CLK(net5447),
    .RESET_B(net5956),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .Q_N(_00423_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][17] ));
 sg13g2_dfrbp_1 _19717_ (.CLK(net5442),
    .RESET_B(net5951),
    .D(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .Q_N(_00430_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[0][18] ));
 sg13g2_dfrbp_1 _19718_ (.CLK(net5465),
    .RESET_B(net5974),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][0] ),
    .Q_N(_09063_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][0] ));
 sg13g2_dfrbp_1 _19719_ (.CLK(net5470),
    .RESET_B(net5978),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][1] ),
    .Q_N(_09064_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][1] ));
 sg13g2_dfrbp_1 _19720_ (.CLK(net5468),
    .RESET_B(net5977),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][2] ),
    .Q_N(_09065_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][2] ));
 sg13g2_dfrbp_1 _19721_ (.CLK(net5513),
    .RESET_B(net6023),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][3] ),
    .Q_N(_09066_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][3] ));
 sg13g2_dfrbp_1 _19722_ (.CLK(net5520),
    .RESET_B(net6029),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][4] ),
    .Q_N(_09067_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][4] ));
 sg13g2_dfrbp_1 _19723_ (.CLK(net5519),
    .RESET_B(net6028),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][5] ),
    .Q_N(_09068_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][5] ));
 sg13g2_dfrbp_1 _19724_ (.CLK(net5539),
    .RESET_B(net6048),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][6] ),
    .Q_N(_09069_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][6] ));
 sg13g2_dfrbp_1 _19725_ (.CLK(net5546),
    .RESET_B(net6055),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][7] ),
    .Q_N(_09070_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][7] ));
 sg13g2_dfrbp_1 _19726_ (.CLK(net5543),
    .RESET_B(net6057),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][8] ),
    .Q_N(_09071_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][8] ));
 sg13g2_dfrbp_1 _19727_ (.CLK(net5546),
    .RESET_B(net6055),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][9] ),
    .Q_N(_09072_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][9] ));
 sg13g2_dfrbp_1 _19728_ (.CLK(net5551),
    .RESET_B(net6060),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][10] ),
    .Q_N(_09073_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][10] ));
 sg13g2_dfrbp_1 _19729_ (.CLK(net5551),
    .RESET_B(net6061),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][11] ),
    .Q_N(_09074_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][11] ));
 sg13g2_dfrbp_1 _19730_ (.CLK(net5550),
    .RESET_B(net6059),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][12] ),
    .Q_N(_09075_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][12] ));
 sg13g2_dfrbp_1 _19731_ (.CLK(net5541),
    .RESET_B(net6050),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][13] ),
    .Q_N(_09076_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][13] ));
 sg13g2_dfrbp_1 _19732_ (.CLK(net5542),
    .RESET_B(net6051),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][14] ),
    .Q_N(_09077_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][14] ));
 sg13g2_dfrbp_1 _19733_ (.CLK(net5449),
    .RESET_B(net5958),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][15] ),
    .Q_N(_09078_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][15] ));
 sg13g2_dfrbp_1 _19734_ (.CLK(net5448),
    .RESET_B(net5957),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][16] ),
    .Q_N(_09079_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][16] ));
 sg13g2_dfrbp_1 _19735_ (.CLK(net5444),
    .RESET_B(net5953),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][17] ),
    .Q_N(_09080_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][17] ));
 sg13g2_dfrbp_1 _19736_ (.CLK(net5446),
    .RESET_B(net5955),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[9][18] ),
    .Q_N(_09081_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[4].u_delay_line.buffer[10][18] ));
 sg13g2_dfrbp_1 _19737_ (.CLK(net5441),
    .RESET_B(net5950),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][0] ),
    .Q_N(_09082_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][0] ));
 sg13g2_dfrbp_1 _19738_ (.CLK(net5457),
    .RESET_B(net5966),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][1] ),
    .Q_N(_09083_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][1] ));
 sg13g2_dfrbp_1 _19739_ (.CLK(net5503),
    .RESET_B(net6012),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][2] ),
    .Q_N(_09084_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][2] ));
 sg13g2_dfrbp_1 _19740_ (.CLK(net5509),
    .RESET_B(net6018),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][3] ),
    .Q_N(_09085_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][3] ));
 sg13g2_dfrbp_1 _19741_ (.CLK(net5510),
    .RESET_B(net6019),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][4] ),
    .Q_N(_09086_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][4] ));
 sg13g2_dfrbp_1 _19742_ (.CLK(net5525),
    .RESET_B(net6034),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][5] ),
    .Q_N(_09087_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][5] ));
 sg13g2_dfrbp_1 _19743_ (.CLK(net5526),
    .RESET_B(net6035),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][6] ),
    .Q_N(_09088_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][6] ));
 sg13g2_dfrbp_1 _19744_ (.CLK(net5532),
    .RESET_B(net6041),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][7] ),
    .Q_N(_09089_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][7] ));
 sg13g2_dfrbp_1 _19745_ (.CLK(net5533),
    .RESET_B(net6042),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][8] ),
    .Q_N(_09090_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][8] ));
 sg13g2_dfrbp_1 _19746_ (.CLK(net5599),
    .RESET_B(net6108),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][9] ),
    .Q_N(_09091_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][9] ));
 sg13g2_dfrbp_1 _19747_ (.CLK(net5535),
    .RESET_B(net6044),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][10] ),
    .Q_N(_09092_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][10] ));
 sg13g2_dfrbp_1 _19748_ (.CLK(net5607),
    .RESET_B(net6116),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][11] ),
    .Q_N(_09093_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][11] ));
 sg13g2_dfrbp_1 _19749_ (.CLK(net5547),
    .RESET_B(net6056),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][12] ),
    .Q_N(_09094_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][12] ));
 sg13g2_dfrbp_1 _19750_ (.CLK(net5545),
    .RESET_B(net6054),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][13] ),
    .Q_N(_09095_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][13] ));
 sg13g2_dfrbp_1 _19751_ (.CLK(net5516),
    .RESET_B(net6025),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][14] ),
    .Q_N(_09096_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][14] ));
 sg13g2_dfrbp_1 _19752_ (.CLK(net5462),
    .RESET_B(net5970),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][15] ),
    .Q_N(_09097_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][15] ));
 sg13g2_dfrbp_1 _19753_ (.CLK(net5463),
    .RESET_B(net5971),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][16] ),
    .Q_N(_09098_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][16] ));
 sg13g2_dfrbp_1 _19754_ (.CLK(net5460),
    .RESET_B(net5968),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][17] ),
    .Q_N(_09099_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][17] ));
 sg13g2_dfrbp_1 _19755_ (.CLK(net5455),
    .RESET_B(net5964),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][18] ),
    .Q_N(_09100_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][18] ));
 sg13g2_dfrbp_1 _19756_ (.CLK(net5441),
    .RESET_B(net5950),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][0] ),
    .Q_N(_09101_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][0] ));
 sg13g2_dfrbp_1 _19757_ (.CLK(net5457),
    .RESET_B(net5966),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][1] ),
    .Q_N(_09102_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][1] ));
 sg13g2_dfrbp_1 _19758_ (.CLK(net5503),
    .RESET_B(net6012),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][2] ),
    .Q_N(_09103_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][2] ));
 sg13g2_dfrbp_1 _19759_ (.CLK(net5509),
    .RESET_B(net6018),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][3] ),
    .Q_N(_09104_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][3] ));
 sg13g2_dfrbp_1 _19760_ (.CLK(net5510),
    .RESET_B(net6019),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][4] ),
    .Q_N(_09105_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][4] ));
 sg13g2_dfrbp_1 _19761_ (.CLK(net5525),
    .RESET_B(net6034),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][5] ),
    .Q_N(_09106_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][5] ));
 sg13g2_dfrbp_1 _19762_ (.CLK(net5526),
    .RESET_B(net6035),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][6] ),
    .Q_N(_09107_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][6] ));
 sg13g2_dfrbp_1 _19763_ (.CLK(net5532),
    .RESET_B(net6041),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][7] ),
    .Q_N(_09108_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][7] ));
 sg13g2_dfrbp_1 _19764_ (.CLK(net5534),
    .RESET_B(net6043),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][8] ),
    .Q_N(_09109_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][8] ));
 sg13g2_dfrbp_1 _19765_ (.CLK(net5599),
    .RESET_B(net6108),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][9] ),
    .Q_N(_09110_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][9] ));
 sg13g2_dfrbp_1 _19766_ (.CLK(net5535),
    .RESET_B(net6044),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][10] ),
    .Q_N(_09111_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][10] ));
 sg13g2_dfrbp_1 _19767_ (.CLK(net5607),
    .RESET_B(net6116),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][11] ),
    .Q_N(_09112_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][11] ));
 sg13g2_dfrbp_1 _19768_ (.CLK(net5608),
    .RESET_B(net6117),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][12] ),
    .Q_N(_09113_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][12] ));
 sg13g2_dfrbp_1 _19769_ (.CLK(net5545),
    .RESET_B(net6054),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][13] ),
    .Q_N(_09114_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][13] ));
 sg13g2_dfrbp_1 _19770_ (.CLK(net5516),
    .RESET_B(net6025),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][14] ),
    .Q_N(_09115_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][14] ));
 sg13g2_dfrbp_1 _19771_ (.CLK(net5462),
    .RESET_B(net5970),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][15] ),
    .Q_N(_09116_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][15] ));
 sg13g2_dfrbp_1 _19772_ (.CLK(net5463),
    .RESET_B(net5971),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][16] ),
    .Q_N(_09117_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][16] ));
 sg13g2_dfrbp_1 _19773_ (.CLK(net5460),
    .RESET_B(net5968),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][17] ),
    .Q_N(_09118_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][17] ));
 sg13g2_dfrbp_1 _19774_ (.CLK(net5455),
    .RESET_B(net5964),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][18] ),
    .Q_N(_09119_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[6][18] ));
 sg13g2_dfrbp_1 _19775_ (.CLK(net5442),
    .RESET_B(net5950),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][0] ),
    .Q_N(_09120_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][0] ));
 sg13g2_dfrbp_1 _19776_ (.CLK(net5457),
    .RESET_B(net5966),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][1] ),
    .Q_N(_09121_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][1] ));
 sg13g2_dfrbp_1 _19777_ (.CLK(net5503),
    .RESET_B(net6012),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][2] ),
    .Q_N(_09122_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][2] ));
 sg13g2_dfrbp_1 _19778_ (.CLK(net5509),
    .RESET_B(net6018),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][3] ),
    .Q_N(_09123_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][3] ));
 sg13g2_dfrbp_1 _19779_ (.CLK(net5510),
    .RESET_B(net6019),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][4] ),
    .Q_N(_09124_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][4] ));
 sg13g2_dfrbp_1 _19780_ (.CLK(net5525),
    .RESET_B(net6034),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][5] ),
    .Q_N(_09125_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][5] ));
 sg13g2_dfrbp_1 _19781_ (.CLK(net5526),
    .RESET_B(net6035),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][6] ),
    .Q_N(_09126_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][6] ));
 sg13g2_dfrbp_1 _19782_ (.CLK(net5532),
    .RESET_B(net6041),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][7] ),
    .Q_N(_09127_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][7] ));
 sg13g2_dfrbp_1 _19783_ (.CLK(net5533),
    .RESET_B(net6042),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][8] ),
    .Q_N(_09128_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][8] ));
 sg13g2_dfrbp_1 _19784_ (.CLK(net5599),
    .RESET_B(net6118),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][9] ),
    .Q_N(_09129_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][9] ));
 sg13g2_dfrbp_1 _19785_ (.CLK(net5535),
    .RESET_B(net6044),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][10] ),
    .Q_N(_09130_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][10] ));
 sg13g2_dfrbp_1 _19786_ (.CLK(net5607),
    .RESET_B(net6116),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][11] ),
    .Q_N(_09131_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][11] ));
 sg13g2_dfrbp_1 _19787_ (.CLK(net5547),
    .RESET_B(net6056),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][12] ),
    .Q_N(_09132_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][12] ));
 sg13g2_dfrbp_1 _19788_ (.CLK(net5537),
    .RESET_B(net6046),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][13] ),
    .Q_N(_09133_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][13] ));
 sg13g2_dfrbp_1 _19789_ (.CLK(net5516),
    .RESET_B(net6025),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][14] ),
    .Q_N(_09134_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][14] ));
 sg13g2_dfrbp_1 _19790_ (.CLK(net5463),
    .RESET_B(net5970),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][15] ),
    .Q_N(_09135_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][15] ));
 sg13g2_dfrbp_1 _19791_ (.CLK(net5463),
    .RESET_B(net5971),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][16] ),
    .Q_N(_09136_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][16] ));
 sg13g2_dfrbp_1 _19792_ (.CLK(net5460),
    .RESET_B(net5968),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][17] ),
    .Q_N(_09137_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][17] ));
 sg13g2_dfrbp_1 _19793_ (.CLK(net5455),
    .RESET_B(net5964),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][18] ),
    .Q_N(_09138_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][18] ));
 sg13g2_dfrbp_1 _19794_ (.CLK(net5441),
    .RESET_B(net5950),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][0] ),
    .Q_N(_09139_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][0] ));
 sg13g2_dfrbp_1 _19795_ (.CLK(net5457),
    .RESET_B(net5966),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][1] ),
    .Q_N(_09140_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][1] ));
 sg13g2_dfrbp_1 _19796_ (.CLK(net5503),
    .RESET_B(net6012),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][2] ),
    .Q_N(_09141_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][2] ));
 sg13g2_dfrbp_1 _19797_ (.CLK(net5509),
    .RESET_B(net6018),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][3] ),
    .Q_N(_09142_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][3] ));
 sg13g2_dfrbp_1 _19798_ (.CLK(net5510),
    .RESET_B(net6019),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][4] ),
    .Q_N(_09143_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][4] ));
 sg13g2_dfrbp_1 _19799_ (.CLK(net5525),
    .RESET_B(net6034),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][5] ),
    .Q_N(_09144_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][5] ));
 sg13g2_dfrbp_1 _19800_ (.CLK(net5526),
    .RESET_B(net6035),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][6] ),
    .Q_N(_09145_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][6] ));
 sg13g2_dfrbp_1 _19801_ (.CLK(net5532),
    .RESET_B(net6041),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][7] ),
    .Q_N(_09146_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][7] ));
 sg13g2_dfrbp_1 _19802_ (.CLK(net5534),
    .RESET_B(net6043),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][8] ),
    .Q_N(_09147_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][8] ));
 sg13g2_dfrbp_1 _19803_ (.CLK(net5599),
    .RESET_B(net6108),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][9] ),
    .Q_N(_09148_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][9] ));
 sg13g2_dfrbp_1 _19804_ (.CLK(net5536),
    .RESET_B(net6044),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][10] ),
    .Q_N(_09149_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][10] ));
 sg13g2_dfrbp_1 _19805_ (.CLK(net5607),
    .RESET_B(net6116),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][11] ),
    .Q_N(_09150_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][11] ));
 sg13g2_dfrbp_1 _19806_ (.CLK(net5607),
    .RESET_B(net6116),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][12] ),
    .Q_N(_09151_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][12] ));
 sg13g2_dfrbp_1 _19807_ (.CLK(net5545),
    .RESET_B(net6054),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][13] ),
    .Q_N(_09152_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][13] ));
 sg13g2_dfrbp_1 _19808_ (.CLK(net5516),
    .RESET_B(net6025),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][14] ),
    .Q_N(_09153_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][14] ));
 sg13g2_dfrbp_1 _19809_ (.CLK(net5505),
    .RESET_B(net6014),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][15] ),
    .Q_N(_09154_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][15] ));
 sg13g2_dfrbp_1 _19810_ (.CLK(net5463),
    .RESET_B(net5971),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][16] ),
    .Q_N(_09155_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][16] ));
 sg13g2_dfrbp_1 _19811_ (.CLK(net5460),
    .RESET_B(net5968),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][17] ),
    .Q_N(_09156_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][17] ));
 sg13g2_dfrbp_1 _19812_ (.CLK(net5439),
    .RESET_B(net5948),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][18] ),
    .Q_N(_09157_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[5][18] ));
 sg13g2_dfrbp_1 _19813_ (.CLK(net5441),
    .RESET_B(net5950),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][0] ),
    .Q_N(_09158_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][0] ));
 sg13g2_dfrbp_1 _19814_ (.CLK(net5457),
    .RESET_B(net5966),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][1] ),
    .Q_N(_09159_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][1] ));
 sg13g2_dfrbp_1 _19815_ (.CLK(net5503),
    .RESET_B(net6012),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][2] ),
    .Q_N(_09160_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][2] ));
 sg13g2_dfrbp_1 _19816_ (.CLK(net5509),
    .RESET_B(net6018),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][3] ),
    .Q_N(_09161_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][3] ));
 sg13g2_dfrbp_1 _19817_ (.CLK(net5510),
    .RESET_B(net6019),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][4] ),
    .Q_N(_09162_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][4] ));
 sg13g2_dfrbp_1 _19818_ (.CLK(net5525),
    .RESET_B(net6034),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][5] ),
    .Q_N(_09163_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][5] ));
 sg13g2_dfrbp_1 _19819_ (.CLK(net5526),
    .RESET_B(net6035),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][6] ),
    .Q_N(_09164_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][6] ));
 sg13g2_dfrbp_1 _19820_ (.CLK(net5532),
    .RESET_B(net6041),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][7] ),
    .Q_N(_09165_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][7] ));
 sg13g2_dfrbp_1 _19821_ (.CLK(net5532),
    .RESET_B(net6041),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][8] ),
    .Q_N(_09166_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][8] ));
 sg13g2_dfrbp_1 _19822_ (.CLK(net5599),
    .RESET_B(net6108),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][9] ),
    .Q_N(_09167_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][9] ));
 sg13g2_dfrbp_1 _19823_ (.CLK(net5536),
    .RESET_B(net6045),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][10] ),
    .Q_N(_09168_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][10] ));
 sg13g2_dfrbp_1 _19824_ (.CLK(net5608),
    .RESET_B(net6117),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][11] ),
    .Q_N(_09169_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][11] ));
 sg13g2_dfrbp_1 _19825_ (.CLK(net5608),
    .RESET_B(net6117),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][12] ),
    .Q_N(_09170_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][12] ));
 sg13g2_dfrbp_1 _19826_ (.CLK(net5545),
    .RESET_B(net6054),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][13] ),
    .Q_N(_09171_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][13] ));
 sg13g2_dfrbp_1 _19827_ (.CLK(net5516),
    .RESET_B(net6025),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][14] ),
    .Q_N(_09172_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][14] ));
 sg13g2_dfrbp_1 _19828_ (.CLK(net5462),
    .RESET_B(net5970),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][15] ),
    .Q_N(_09173_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][15] ));
 sg13g2_dfrbp_1 _19829_ (.CLK(net5463),
    .RESET_B(net5971),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][16] ),
    .Q_N(_09174_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][16] ));
 sg13g2_dfrbp_1 _19830_ (.CLK(net5460),
    .RESET_B(net5968),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][17] ),
    .Q_N(_09175_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][17] ));
 sg13g2_dfrbp_1 _19831_ (.CLK(net5439),
    .RESET_B(net5948),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][18] ),
    .Q_N(_09176_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[4][18] ));
 sg13g2_dfrbp_1 _19832_ (.CLK(net5442),
    .RESET_B(net5951),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][0] ),
    .Q_N(_09177_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][0] ));
 sg13g2_dfrbp_1 _19833_ (.CLK(net5458),
    .RESET_B(net5967),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][1] ),
    .Q_N(_09178_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][1] ));
 sg13g2_dfrbp_1 _19834_ (.CLK(net5505),
    .RESET_B(net6014),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][2] ),
    .Q_N(_09179_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][2] ));
 sg13g2_dfrbp_1 _19835_ (.CLK(net5504),
    .RESET_B(net6013),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][3] ),
    .Q_N(_09180_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][3] ));
 sg13g2_dfrbp_1 _19836_ (.CLK(net5510),
    .RESET_B(net6019),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][4] ),
    .Q_N(_09181_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][4] ));
 sg13g2_dfrbp_1 _19837_ (.CLK(net5511),
    .RESET_B(net6020),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][5] ),
    .Q_N(_09182_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][5] ));
 sg13g2_dfrbp_1 _19838_ (.CLK(net5525),
    .RESET_B(net6034),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][6] ),
    .Q_N(_09183_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][6] ));
 sg13g2_dfrbp_1 _19839_ (.CLK(net5534),
    .RESET_B(net6043),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][7] ),
    .Q_N(_09184_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][7] ));
 sg13g2_dfrbp_1 _19840_ (.CLK(net5534),
    .RESET_B(net6043),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][8] ),
    .Q_N(_09185_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][8] ));
 sg13g2_dfrbp_1 _19841_ (.CLK(net5609),
    .RESET_B(net6108),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][9] ),
    .Q_N(_09186_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][9] ));
 sg13g2_dfrbp_1 _19842_ (.CLK(net5535),
    .RESET_B(net6044),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][10] ),
    .Q_N(_09187_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][10] ));
 sg13g2_dfrbp_1 _19843_ (.CLK(net5608),
    .RESET_B(net6117),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][11] ),
    .Q_N(_09188_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][11] ));
 sg13g2_dfrbp_1 _19844_ (.CLK(net5547),
    .RESET_B(net6056),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][12] ),
    .Q_N(_09189_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][12] ));
 sg13g2_dfrbp_1 _19845_ (.CLK(net5545),
    .RESET_B(net6054),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][13] ),
    .Q_N(_09190_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][13] ));
 sg13g2_dfrbp_1 _19846_ (.CLK(net5516),
    .RESET_B(net6025),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][14] ),
    .Q_N(_09191_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][14] ));
 sg13g2_dfrbp_1 _19847_ (.CLK(net5462),
    .RESET_B(net5970),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][15] ),
    .Q_N(_09192_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][15] ));
 sg13g2_dfrbp_1 _19848_ (.CLK(net5458),
    .RESET_B(net5967),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][16] ),
    .Q_N(_09193_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][16] ));
 sg13g2_dfrbp_1 _19849_ (.CLK(net5460),
    .RESET_B(net5968),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][17] ),
    .Q_N(_09194_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][17] ));
 sg13g2_dfrbp_1 _19850_ (.CLK(net5439),
    .RESET_B(net5948),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][18] ),
    .Q_N(_09195_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[3][18] ));
 sg13g2_dfrbp_1 _19851_ (.CLK(net5441),
    .RESET_B(net5950),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][0] ),
    .Q_N(_09196_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][0] ));
 sg13g2_dfrbp_1 _19852_ (.CLK(net5457),
    .RESET_B(net5966),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][1] ),
    .Q_N(_09197_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][1] ));
 sg13g2_dfrbp_1 _19853_ (.CLK(net5505),
    .RESET_B(net6014),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][2] ),
    .Q_N(_09198_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][2] ));
 sg13g2_dfrbp_1 _19854_ (.CLK(net5504),
    .RESET_B(net6013),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][3] ),
    .Q_N(_09199_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][3] ));
 sg13g2_dfrbp_1 _19855_ (.CLK(net5509),
    .RESET_B(net6018),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][4] ),
    .Q_N(_09200_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][4] ));
 sg13g2_dfrbp_1 _19856_ (.CLK(net5507),
    .RESET_B(net6016),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][5] ),
    .Q_N(_09201_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][5] ));
 sg13g2_dfrbp_1 _19857_ (.CLK(net5528),
    .RESET_B(net6037),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][6] ),
    .Q_N(_09202_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][6] ));
 sg13g2_dfrbp_1 _19858_ (.CLK(net5538),
    .RESET_B(net6047),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][7] ),
    .Q_N(_09203_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][7] ));
 sg13g2_dfrbp_1 _19859_ (.CLK(net5534),
    .RESET_B(net6043),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][8] ),
    .Q_N(_09204_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][8] ));
 sg13g2_dfrbp_1 _19860_ (.CLK(net5533),
    .RESET_B(net6042),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][9] ),
    .Q_N(_09205_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][9] ));
 sg13g2_dfrbp_1 _19861_ (.CLK(net5535),
    .RESET_B(net6044),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][10] ),
    .Q_N(_09206_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][10] ));
 sg13g2_dfrbp_1 _19862_ (.CLK(net5607),
    .RESET_B(net6116),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][11] ),
    .Q_N(_09207_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][11] ));
 sg13g2_dfrbp_1 _19863_ (.CLK(net5547),
    .RESET_B(net6056),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][12] ),
    .Q_N(_09208_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][12] ));
 sg13g2_dfrbp_1 _19864_ (.CLK(net5540),
    .RESET_B(net6049),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][13] ),
    .Q_N(_09209_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][13] ));
 sg13g2_dfrbp_1 _19865_ (.CLK(net5504),
    .RESET_B(net6013),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][14] ),
    .Q_N(_09210_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][14] ));
 sg13g2_dfrbp_1 _19866_ (.CLK(net5462),
    .RESET_B(net5970),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][15] ),
    .Q_N(_09211_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][15] ));
 sg13g2_dfrbp_1 _19867_ (.CLK(net5458),
    .RESET_B(net5967),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][16] ),
    .Q_N(_09212_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][16] ));
 sg13g2_dfrbp_1 _19868_ (.CLK(net5456),
    .RESET_B(net5965),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][17] ),
    .Q_N(_09213_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][17] ));
 sg13g2_dfrbp_1 _19869_ (.CLK(net5440),
    .RESET_B(net5948),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][18] ),
    .Q_N(_09214_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[2][18] ));
 sg13g2_dfrbp_1 _19870_ (.CLK(net5441),
    .RESET_B(net5951),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][0] ),
    .Q_N(_09215_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][0] ));
 sg13g2_dfrbp_1 _19871_ (.CLK(net5457),
    .RESET_B(net5966),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][1] ),
    .Q_N(_09216_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][1] ));
 sg13g2_dfrbp_1 _19872_ (.CLK(net5503),
    .RESET_B(net6012),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][2] ),
    .Q_N(_09217_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][2] ));
 sg13g2_dfrbp_1 _19873_ (.CLK(net5509),
    .RESET_B(net6018),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][3] ),
    .Q_N(_09218_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][3] ));
 sg13g2_dfrbp_1 _19874_ (.CLK(net5510),
    .RESET_B(net6019),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][4] ),
    .Q_N(_09219_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][4] ));
 sg13g2_dfrbp_1 _19875_ (.CLK(net5525),
    .RESET_B(net6034),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][5] ),
    .Q_N(_09220_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][5] ));
 sg13g2_dfrbp_1 _19876_ (.CLK(net5526),
    .RESET_B(net6035),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][6] ),
    .Q_N(_09221_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][6] ));
 sg13g2_dfrbp_1 _19877_ (.CLK(net5532),
    .RESET_B(net6041),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][7] ),
    .Q_N(_09222_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][7] ));
 sg13g2_dfrbp_1 _19878_ (.CLK(net5533),
    .RESET_B(net6042),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][8] ),
    .Q_N(_09223_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][8] ));
 sg13g2_dfrbp_1 _19879_ (.CLK(net5599),
    .RESET_B(net6108),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][9] ),
    .Q_N(_09224_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][9] ));
 sg13g2_dfrbp_1 _19880_ (.CLK(net5535),
    .RESET_B(net6044),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][10] ),
    .Q_N(_09225_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][10] ));
 sg13g2_dfrbp_1 _19881_ (.CLK(net5607),
    .RESET_B(net6116),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][11] ),
    .Q_N(_09226_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][11] ));
 sg13g2_dfrbp_1 _19882_ (.CLK(net5547),
    .RESET_B(net6056),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][12] ),
    .Q_N(_09227_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][12] ));
 sg13g2_dfrbp_1 _19883_ (.CLK(net5545),
    .RESET_B(net6054),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][13] ),
    .Q_N(_09228_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][13] ));
 sg13g2_dfrbp_1 _19884_ (.CLK(net5516),
    .RESET_B(net6025),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][14] ),
    .Q_N(_09229_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][14] ));
 sg13g2_dfrbp_1 _19885_ (.CLK(net5462),
    .RESET_B(net5970),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][15] ),
    .Q_N(_09230_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][15] ));
 sg13g2_dfrbp_1 _19886_ (.CLK(net5463),
    .RESET_B(net5971),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][16] ),
    .Q_N(_09231_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][16] ));
 sg13g2_dfrbp_1 _19887_ (.CLK(net5460),
    .RESET_B(net5968),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][17] ),
    .Q_N(_09232_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][17] ));
 sg13g2_dfrbp_1 _19888_ (.CLK(net5455),
    .RESET_B(net5964),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[7][18] ),
    .Q_N(_09233_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[8][18] ));
 sg13g2_dfrbp_1 _19889_ (.CLK(net5441),
    .RESET_B(net5950),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][0] ),
    .Q_N(_09234_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][0] ));
 sg13g2_dfrbp_1 _19890_ (.CLK(net5458),
    .RESET_B(net5967),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][1] ),
    .Q_N(_09235_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][1] ));
 sg13g2_dfrbp_1 _19891_ (.CLK(net5505),
    .RESET_B(net6014),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][2] ),
    .Q_N(_09236_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][2] ));
 sg13g2_dfrbp_1 _19892_ (.CLK(net5504),
    .RESET_B(net6013),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][3] ),
    .Q_N(_09237_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][3] ));
 sg13g2_dfrbp_1 _19893_ (.CLK(net5507),
    .RESET_B(net6016),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][4] ),
    .Q_N(_09238_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][4] ));
 sg13g2_dfrbp_1 _19894_ (.CLK(net5507),
    .RESET_B(net6016),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][5] ),
    .Q_N(_09239_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][5] ));
 sg13g2_dfrbp_1 _19895_ (.CLK(net5528),
    .RESET_B(net6037),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][6] ),
    .Q_N(_09240_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][6] ));
 sg13g2_dfrbp_1 _19896_ (.CLK(net5531),
    .RESET_B(net6040),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][7] ),
    .Q_N(_09241_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][7] ));
 sg13g2_dfrbp_1 _19897_ (.CLK(net5531),
    .RESET_B(net6040),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][8] ),
    .Q_N(_09242_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][8] ));
 sg13g2_dfrbp_1 _19898_ (.CLK(net5537),
    .RESET_B(net6046),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][9] ),
    .Q_N(_09243_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][9] ));
 sg13g2_dfrbp_1 _19899_ (.CLK(net5537),
    .RESET_B(net6046),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][10] ),
    .Q_N(_09244_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][10] ));
 sg13g2_dfrbp_1 _19900_ (.CLK(net5535),
    .RESET_B(net6044),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][11] ),
    .Q_N(_09245_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][11] ));
 sg13g2_dfrbp_1 _19901_ (.CLK(net5537),
    .RESET_B(net6046),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][12] ),
    .Q_N(_09246_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][12] ));
 sg13g2_dfrbp_1 _19902_ (.CLK(net5526),
    .RESET_B(net6035),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][13] ),
    .Q_N(_09247_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][13] ));
 sg13g2_dfrbp_1 _19903_ (.CLK(net5503),
    .RESET_B(net6012),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][14] ),
    .Q_N(_09248_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][14] ));
 sg13g2_dfrbp_1 _19904_ (.CLK(net5462),
    .RESET_B(net5970),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][15] ),
    .Q_N(_09249_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][15] ));
 sg13g2_dfrbp_1 _19905_ (.CLK(net5456),
    .RESET_B(net5965),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][16] ),
    .Q_N(_09250_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][16] ));
 sg13g2_dfrbp_1 _19906_ (.CLK(net5456),
    .RESET_B(net5965),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][17] ),
    .Q_N(_09251_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][17] ));
 sg13g2_dfrbp_1 _19907_ (.CLK(net5439),
    .RESET_B(net5949),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][18] ),
    .Q_N(_09252_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[1][18] ));
 sg13g2_dfrbp_1 _19908_ (.CLK(net5439),
    .RESET_B(net5948),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.u_mux_shift.sum_res ),
    .Q_N(_00290_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][0] ));
 sg13g2_dfrbp_1 _19909_ (.CLK(net5459),
    .RESET_B(net5973),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .Q_N(_00298_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][1] ));
 sg13g2_dfrbp_1 _19910_ (.CLK(net5464),
    .RESET_B(net5972),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .Q_N(_00305_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][2] ));
 sg13g2_dfrbp_1 _19911_ (.CLK(net5502),
    .RESET_B(net6011),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .Q_N(_00312_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][3] ));
 sg13g2_dfrbp_1 _19912_ (.CLK(net5502),
    .RESET_B(net6011),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .Q_N(_00321_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][4] ));
 sg13g2_dfrbp_1 _19913_ (.CLK(net5507),
    .RESET_B(net6016),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .Q_N(_00330_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][5] ));
 sg13g2_dfrbp_1 _19914_ (.CLK(net5507),
    .RESET_B(net6016),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .Q_N(_00337_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][6] ));
 sg13g2_dfrbp_1 _19915_ (.CLK(net5528),
    .RESET_B(net6037),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .Q_N(_00344_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][7] ));
 sg13g2_dfrbp_1 _19916_ (.CLK(net5528),
    .RESET_B(net6037),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .Q_N(_00353_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][8] ));
 sg13g2_dfrbp_1 _19917_ (.CLK(net5531),
    .RESET_B(net6040),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .Q_N(_00362_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][9] ));
 sg13g2_dfrbp_1 _19918_ (.CLK(net5537),
    .RESET_B(net6046),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .Q_N(_00369_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][10] ));
 sg13g2_dfrbp_1 _19919_ (.CLK(net5537),
    .RESET_B(net6046),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .Q_N(_00376_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][11] ));
 sg13g2_dfrbp_1 _19920_ (.CLK(net5527),
    .RESET_B(net6036),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .Q_N(_00385_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][12] ));
 sg13g2_dfrbp_1 _19921_ (.CLK(net5527),
    .RESET_B(net6036),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .Q_N(_00394_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][13] ));
 sg13g2_dfrbp_1 _19922_ (.CLK(net5505),
    .RESET_B(net6014),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .Q_N(_00401_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][14] ));
 sg13g2_dfrbp_1 _19923_ (.CLK(net5463),
    .RESET_B(net5971),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .Q_N(_00408_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][15] ));
 sg13g2_dfrbp_1 _19924_ (.CLK(net5455),
    .RESET_B(net5964),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .Q_N(_00417_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][16] ));
 sg13g2_dfrbp_1 _19925_ (.CLK(net5455),
    .RESET_B(net5964),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .Q_N(_00424_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][17] ));
 sg13g2_dfrbp_1 _19926_ (.CLK(net5440),
    .RESET_B(net5949),
    .D(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .Q_N(_00431_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[0][18] ));
 sg13g2_dfrbp_1 _19927_ (.CLK(net5441),
    .RESET_B(net5950),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][0] ),
    .Q_N(_09253_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][0] ));
 sg13g2_dfrbp_1 _19928_ (.CLK(net5457),
    .RESET_B(net5966),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][1] ),
    .Q_N(_09254_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][1] ));
 sg13g2_dfrbp_1 _19929_ (.CLK(net5503),
    .RESET_B(net6012),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][2] ),
    .Q_N(_09255_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][2] ));
 sg13g2_dfrbp_1 _19930_ (.CLK(net5509),
    .RESET_B(net6018),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][3] ),
    .Q_N(_09256_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][3] ));
 sg13g2_dfrbp_1 _19931_ (.CLK(net5510),
    .RESET_B(net6019),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][4] ),
    .Q_N(_09257_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][4] ));
 sg13g2_dfrbp_1 _19932_ (.CLK(net5525),
    .RESET_B(net6034),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][5] ),
    .Q_N(_09258_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][5] ));
 sg13g2_dfrbp_1 _19933_ (.CLK(net5526),
    .RESET_B(net6035),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][6] ),
    .Q_N(_09259_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][6] ));
 sg13g2_dfrbp_1 _19934_ (.CLK(net5532),
    .RESET_B(net6041),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][7] ),
    .Q_N(_09260_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][7] ));
 sg13g2_dfrbp_1 _19935_ (.CLK(net5533),
    .RESET_B(net6042),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][8] ),
    .Q_N(_09261_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][8] ));
 sg13g2_dfrbp_1 _19936_ (.CLK(net5599),
    .RESET_B(net6108),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][9] ),
    .Q_N(_09262_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][9] ));
 sg13g2_dfrbp_1 _19937_ (.CLK(net5535),
    .RESET_B(net6045),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][10] ),
    .Q_N(_09263_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][10] ));
 sg13g2_dfrbp_1 _19938_ (.CLK(net5607),
    .RESET_B(net6116),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][11] ),
    .Q_N(_09264_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][11] ));
 sg13g2_dfrbp_1 _19939_ (.CLK(net5547),
    .RESET_B(net6056),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][12] ),
    .Q_N(_09265_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][12] ));
 sg13g2_dfrbp_1 _19940_ (.CLK(net5537),
    .RESET_B(net6046),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][13] ),
    .Q_N(_09266_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][13] ));
 sg13g2_dfrbp_1 _19941_ (.CLK(net5512),
    .RESET_B(net6021),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][14] ),
    .Q_N(_09267_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][14] ));
 sg13g2_dfrbp_1 _19942_ (.CLK(net5462),
    .RESET_B(net5971),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][15] ),
    .Q_N(_09268_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][15] ));
 sg13g2_dfrbp_1 _19943_ (.CLK(net5458),
    .RESET_B(net5967),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][16] ),
    .Q_N(_09269_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][16] ));
 sg13g2_dfrbp_1 _19944_ (.CLK(net5460),
    .RESET_B(net5968),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][17] ),
    .Q_N(_09270_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][17] ));
 sg13g2_dfrbp_1 _19945_ (.CLK(net5455),
    .RESET_B(net5964),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[9][18] ),
    .Q_N(_09271_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[5].u_delay_line.buffer[10][18] ));
 sg13g2_dfrbp_1 _19946_ (.CLK(net5567),
    .RESET_B(net6076),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][0] ),
    .Q_N(_09272_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][0] ));
 sg13g2_dfrbp_1 _19947_ (.CLK(net5493),
    .RESET_B(net6002),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][1] ),
    .Q_N(_09273_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][1] ));
 sg13g2_dfrbp_1 _19948_ (.CLK(net5498),
    .RESET_B(net6007),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][2] ),
    .Q_N(_09274_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][2] ));
 sg13g2_dfrbp_1 _19949_ (.CLK(net5496),
    .RESET_B(net6005),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][3] ),
    .Q_N(_09275_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][3] ));
 sg13g2_dfrbp_1 _19950_ (.CLK(net5565),
    .RESET_B(net6074),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][4] ),
    .Q_N(_09276_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][4] ));
 sg13g2_dfrbp_1 _19951_ (.CLK(net5570),
    .RESET_B(net6079),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][5] ),
    .Q_N(_09277_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][5] ));
 sg13g2_dfrbp_1 _19952_ (.CLK(net5573),
    .RESET_B(net6082),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][6] ),
    .Q_N(_09278_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][6] ));
 sg13g2_dfrbp_1 _19953_ (.CLK(net5584),
    .RESET_B(net6093),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][7] ),
    .Q_N(_09279_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][7] ));
 sg13g2_dfrbp_1 _19954_ (.CLK(net5587),
    .RESET_B(net6096),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][8] ),
    .Q_N(_09280_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][8] ));
 sg13g2_dfrbp_1 _19955_ (.CLK(net5582),
    .RESET_B(net6091),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][9] ),
    .Q_N(_09281_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][9] ));
 sg13g2_dfrbp_1 _19956_ (.CLK(net5588),
    .RESET_B(net6097),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][10] ),
    .Q_N(_09282_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][10] ));
 sg13g2_dfrbp_1 _19957_ (.CLK(net5576),
    .RESET_B(net6085),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][11] ),
    .Q_N(_09283_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][11] ));
 sg13g2_dfrbp_1 _19958_ (.CLK(net5600),
    .RESET_B(net6109),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][12] ),
    .Q_N(_09284_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][12] ));
 sg13g2_dfrbp_1 _19959_ (.CLK(net5601),
    .RESET_B(net6110),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][13] ),
    .Q_N(_09285_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][13] ));
 sg13g2_dfrbp_1 _19960_ (.CLK(net5595),
    .RESET_B(net6104),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][14] ),
    .Q_N(_09286_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][14] ));
 sg13g2_dfrbp_1 _19961_ (.CLK(net5529),
    .RESET_B(net6038),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][15] ),
    .Q_N(_09287_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][15] ));
 sg13g2_dfrbp_1 _19962_ (.CLK(net5482),
    .RESET_B(net5991),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][16] ),
    .Q_N(_09288_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][16] ));
 sg13g2_dfrbp_1 _19963_ (.CLK(net5437),
    .RESET_B(net5946),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][17] ),
    .Q_N(_09289_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][17] ));
 sg13g2_dfrbp_1 _19964_ (.CLK(net5434),
    .RESET_B(net5943),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][18] ),
    .Q_N(_09290_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][18] ));
 sg13g2_dfrbp_1 _19965_ (.CLK(net5569),
    .RESET_B(net6078),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][0] ),
    .Q_N(_09291_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][0] ));
 sg13g2_dfrbp_1 _19966_ (.CLK(net5494),
    .RESET_B(net6003),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][1] ),
    .Q_N(_09292_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][1] ));
 sg13g2_dfrbp_1 _19967_ (.CLK(net5499),
    .RESET_B(net6008),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][2] ),
    .Q_N(_09293_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][2] ));
 sg13g2_dfrbp_1 _19968_ (.CLK(net5497),
    .RESET_B(net6006),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][3] ),
    .Q_N(_09294_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][3] ));
 sg13g2_dfrbp_1 _19969_ (.CLK(net5564),
    .RESET_B(net6073),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][4] ),
    .Q_N(_09295_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][4] ));
 sg13g2_dfrbp_1 _19970_ (.CLK(net5570),
    .RESET_B(net6079),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][5] ),
    .Q_N(_09296_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][5] ));
 sg13g2_dfrbp_1 _19971_ (.CLK(net5574),
    .RESET_B(net6083),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][6] ),
    .Q_N(_09297_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][6] ));
 sg13g2_dfrbp_1 _19972_ (.CLK(net5582),
    .RESET_B(net6091),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][7] ),
    .Q_N(_09298_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][7] ));
 sg13g2_dfrbp_1 _19973_ (.CLK(net5583),
    .RESET_B(net6092),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][8] ),
    .Q_N(_09299_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][8] ));
 sg13g2_dfrbp_1 _19974_ (.CLK(net5583),
    .RESET_B(net6092),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][9] ),
    .Q_N(_09300_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][9] ));
 sg13g2_dfrbp_1 _19975_ (.CLK(net5588),
    .RESET_B(net6097),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][10] ),
    .Q_N(_09301_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][10] ));
 sg13g2_dfrbp_1 _19976_ (.CLK(net5575),
    .RESET_B(net6085),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][11] ),
    .Q_N(_09302_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][11] ));
 sg13g2_dfrbp_1 _19977_ (.CLK(net5603),
    .RESET_B(net6112),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][12] ),
    .Q_N(_09303_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][12] ));
 sg13g2_dfrbp_1 _19978_ (.CLK(net5601),
    .RESET_B(net6110),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][13] ),
    .Q_N(_09304_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][13] ));
 sg13g2_dfrbp_1 _19979_ (.CLK(net5595),
    .RESET_B(net6104),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][14] ),
    .Q_N(_09305_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][14] ));
 sg13g2_dfrbp_1 _19980_ (.CLK(net5530),
    .RESET_B(net6039),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][15] ),
    .Q_N(_09306_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][15] ));
 sg13g2_dfrbp_1 _19981_ (.CLK(net5481),
    .RESET_B(net5990),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][16] ),
    .Q_N(_09307_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][16] ));
 sg13g2_dfrbp_1 _19982_ (.CLK(net5479),
    .RESET_B(net5988),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][17] ),
    .Q_N(_09308_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][17] ));
 sg13g2_dfrbp_1 _19983_ (.CLK(net5434),
    .RESET_B(net5943),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][18] ),
    .Q_N(_09309_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[12][18] ));
 sg13g2_dfrbp_1 _19984_ (.CLK(net5567),
    .RESET_B(net6076),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][0] ),
    .Q_N(_09310_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][0] ));
 sg13g2_dfrbp_1 _19985_ (.CLK(net5494),
    .RESET_B(net6003),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][1] ),
    .Q_N(_09311_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][1] ));
 sg13g2_dfrbp_1 _19986_ (.CLK(net5498),
    .RESET_B(net6007),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][2] ),
    .Q_N(_09312_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][2] ));
 sg13g2_dfrbp_1 _19987_ (.CLK(net5496),
    .RESET_B(net6005),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][3] ),
    .Q_N(_09313_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][3] ));
 sg13g2_dfrbp_1 _19988_ (.CLK(net5564),
    .RESET_B(net6073),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][4] ),
    .Q_N(_09314_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][4] ));
 sg13g2_dfrbp_1 _19989_ (.CLK(net5570),
    .RESET_B(net6079),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][5] ),
    .Q_N(_09315_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][5] ));
 sg13g2_dfrbp_1 _19990_ (.CLK(net5573),
    .RESET_B(net6082),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][6] ),
    .Q_N(_09316_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][6] ));
 sg13g2_dfrbp_1 _19991_ (.CLK(net5586),
    .RESET_B(net6095),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][7] ),
    .Q_N(_09317_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][7] ));
 sg13g2_dfrbp_1 _19992_ (.CLK(net5587),
    .RESET_B(net6096),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][8] ),
    .Q_N(_09318_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][8] ));
 sg13g2_dfrbp_1 _19993_ (.CLK(net5582),
    .RESET_B(net6091),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][9] ),
    .Q_N(_09319_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][9] ));
 sg13g2_dfrbp_1 _19994_ (.CLK(net5588),
    .RESET_B(net6097),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][10] ),
    .Q_N(_09320_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][10] ));
 sg13g2_dfrbp_1 _19995_ (.CLK(net5576),
    .RESET_B(net6085),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][11] ),
    .Q_N(_09321_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][11] ));
 sg13g2_dfrbp_1 _19996_ (.CLK(net5600),
    .RESET_B(net6109),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][12] ),
    .Q_N(_09322_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][12] ));
 sg13g2_dfrbp_1 _19997_ (.CLK(net5601),
    .RESET_B(net6110),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][13] ),
    .Q_N(_09323_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][13] ));
 sg13g2_dfrbp_1 _19998_ (.CLK(net5595),
    .RESET_B(net6104),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][14] ),
    .Q_N(_09324_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][14] ));
 sg13g2_dfrbp_1 _19999_ (.CLK(net5529),
    .RESET_B(net6038),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][15] ),
    .Q_N(_09325_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][15] ));
 sg13g2_dfrbp_1 _20000_ (.CLK(net5482),
    .RESET_B(net5991),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][16] ),
    .Q_N(_09326_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][16] ));
 sg13g2_dfrbp_1 _20001_ (.CLK(net5437),
    .RESET_B(net5946),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][17] ),
    .Q_N(_09327_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][17] ));
 sg13g2_dfrbp_1 _20002_ (.CLK(net5434),
    .RESET_B(net5943),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][18] ),
    .Q_N(_09328_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[6][18] ));
 sg13g2_dfrbp_1 _20003_ (.CLK(net5567),
    .RESET_B(net6076),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][0] ),
    .Q_N(_09329_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][0] ));
 sg13g2_dfrbp_1 _20004_ (.CLK(net5493),
    .RESET_B(net6002),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][1] ),
    .Q_N(_09330_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][1] ));
 sg13g2_dfrbp_1 _20005_ (.CLK(net5498),
    .RESET_B(net6007),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][2] ),
    .Q_N(_09331_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][2] ));
 sg13g2_dfrbp_1 _20006_ (.CLK(net5496),
    .RESET_B(net6005),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][3] ),
    .Q_N(_09332_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][3] ));
 sg13g2_dfrbp_1 _20007_ (.CLK(net5564),
    .RESET_B(net6073),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][4] ),
    .Q_N(_09333_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][4] ));
 sg13g2_dfrbp_1 _20008_ (.CLK(net5571),
    .RESET_B(net6080),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][5] ),
    .Q_N(_09334_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][5] ));
 sg13g2_dfrbp_1 _20009_ (.CLK(net5572),
    .RESET_B(net6081),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][6] ),
    .Q_N(_09335_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][6] ));
 sg13g2_dfrbp_1 _20010_ (.CLK(net5584),
    .RESET_B(net6093),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][7] ),
    .Q_N(_09336_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][7] ));
 sg13g2_dfrbp_1 _20011_ (.CLK(net5587),
    .RESET_B(net6096),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][8] ),
    .Q_N(_09337_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][8] ));
 sg13g2_dfrbp_1 _20012_ (.CLK(net5583),
    .RESET_B(net6092),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][9] ),
    .Q_N(_09338_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][9] ));
 sg13g2_dfrbp_1 _20013_ (.CLK(net5575),
    .RESET_B(net6084),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][10] ),
    .Q_N(_09339_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][10] ));
 sg13g2_dfrbp_1 _20014_ (.CLK(net5576),
    .RESET_B(net6086),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][11] ),
    .Q_N(_09340_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][11] ));
 sg13g2_dfrbp_1 _20015_ (.CLK(net5600),
    .RESET_B(net6109),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][12] ),
    .Q_N(_09341_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][12] ));
 sg13g2_dfrbp_1 _20016_ (.CLK(net5600),
    .RESET_B(net6109),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][13] ),
    .Q_N(_09342_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][13] ));
 sg13g2_dfrbp_1 _20017_ (.CLK(net5595),
    .RESET_B(net6104),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][14] ),
    .Q_N(_09343_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][14] ));
 sg13g2_dfrbp_1 _20018_ (.CLK(net5530),
    .RESET_B(net6039),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][15] ),
    .Q_N(_09344_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][15] ));
 sg13g2_dfrbp_1 _20019_ (.CLK(net5482),
    .RESET_B(net5991),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][16] ),
    .Q_N(_09345_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][16] ));
 sg13g2_dfrbp_1 _20020_ (.CLK(net5436),
    .RESET_B(net5945),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][17] ),
    .Q_N(_09346_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][17] ));
 sg13g2_dfrbp_1 _20021_ (.CLK(net5434),
    .RESET_B(net5943),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][18] ),
    .Q_N(_09347_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][18] ));
 sg13g2_dfrbp_1 _20022_ (.CLK(net5567),
    .RESET_B(net6076),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][0] ),
    .Q_N(_09348_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][0] ));
 sg13g2_dfrbp_1 _20023_ (.CLK(net5493),
    .RESET_B(net6002),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][1] ),
    .Q_N(_09349_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][1] ));
 sg13g2_dfrbp_1 _20024_ (.CLK(net5498),
    .RESET_B(net6008),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][2] ),
    .Q_N(_09350_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][2] ));
 sg13g2_dfrbp_1 _20025_ (.CLK(net5496),
    .RESET_B(net6005),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][3] ),
    .Q_N(_09351_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][3] ));
 sg13g2_dfrbp_1 _20026_ (.CLK(net5564),
    .RESET_B(net6073),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][4] ),
    .Q_N(_09352_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][4] ));
 sg13g2_dfrbp_1 _20027_ (.CLK(net5570),
    .RESET_B(net6079),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][5] ),
    .Q_N(_09353_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][5] ));
 sg13g2_dfrbp_1 _20028_ (.CLK(net5573),
    .RESET_B(net6082),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][6] ),
    .Q_N(_09354_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][6] ));
 sg13g2_dfrbp_1 _20029_ (.CLK(net5586),
    .RESET_B(net6095),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][7] ),
    .Q_N(_09355_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][7] ));
 sg13g2_dfrbp_1 _20030_ (.CLK(net5587),
    .RESET_B(net6096),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][8] ),
    .Q_N(_09356_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][8] ));
 sg13g2_dfrbp_1 _20031_ (.CLK(net5587),
    .RESET_B(net6096),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][9] ),
    .Q_N(_09357_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][9] ));
 sg13g2_dfrbp_1 _20032_ (.CLK(net5588),
    .RESET_B(net6098),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][10] ),
    .Q_N(_09358_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][10] ));
 sg13g2_dfrbp_1 _20033_ (.CLK(net5576),
    .RESET_B(net6085),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][11] ),
    .Q_N(_09359_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][11] ));
 sg13g2_dfrbp_1 _20034_ (.CLK(net5577),
    .RESET_B(net6086),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][12] ),
    .Q_N(_09360_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][12] ));
 sg13g2_dfrbp_1 _20035_ (.CLK(net5601),
    .RESET_B(net6110),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][13] ),
    .Q_N(_09361_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][13] ));
 sg13g2_dfrbp_1 _20036_ (.CLK(net5596),
    .RESET_B(net6105),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][14] ),
    .Q_N(_09362_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][14] ));
 sg13g2_dfrbp_1 _20037_ (.CLK(net5529),
    .RESET_B(net6038),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][15] ),
    .Q_N(_09363_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][15] ));
 sg13g2_dfrbp_1 _20038_ (.CLK(net5481),
    .RESET_B(net5990),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][16] ),
    .Q_N(_09364_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][16] ));
 sg13g2_dfrbp_1 _20039_ (.CLK(net5437),
    .RESET_B(net5946),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][17] ),
    .Q_N(_09365_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][17] ));
 sg13g2_dfrbp_1 _20040_ (.CLK(net5435),
    .RESET_B(net5944),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][18] ),
    .Q_N(_09366_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[5][18] ));
 sg13g2_dfrbp_1 _20041_ (.CLK(net5568),
    .RESET_B(net6077),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][0] ),
    .Q_N(_09367_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][0] ));
 sg13g2_dfrbp_1 _20042_ (.CLK(net5494),
    .RESET_B(net6003),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][1] ),
    .Q_N(_09368_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][1] ));
 sg13g2_dfrbp_1 _20043_ (.CLK(net5499),
    .RESET_B(net6007),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][2] ),
    .Q_N(_09369_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][2] ));
 sg13g2_dfrbp_1 _20044_ (.CLK(net5496),
    .RESET_B(net6005),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][3] ),
    .Q_N(_09370_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][3] ));
 sg13g2_dfrbp_1 _20045_ (.CLK(net5564),
    .RESET_B(net6073),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][4] ),
    .Q_N(_09371_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][4] ));
 sg13g2_dfrbp_1 _20046_ (.CLK(net5570),
    .RESET_B(net6079),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][5] ),
    .Q_N(_09372_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][5] ));
 sg13g2_dfrbp_1 _20047_ (.CLK(net5572),
    .RESET_B(net6081),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][6] ),
    .Q_N(_09373_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][6] ));
 sg13g2_dfrbp_1 _20048_ (.CLK(net5585),
    .RESET_B(net6094),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][7] ),
    .Q_N(_09374_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][7] ));
 sg13g2_dfrbp_1 _20049_ (.CLK(net5592),
    .RESET_B(net6101),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][8] ),
    .Q_N(_09375_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][8] ));
 sg13g2_dfrbp_1 _20050_ (.CLK(net5585),
    .RESET_B(net6094),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][9] ),
    .Q_N(_09376_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][9] ));
 sg13g2_dfrbp_1 _20051_ (.CLK(net5589),
    .RESET_B(net6098),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][10] ),
    .Q_N(_09377_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][10] ));
 sg13g2_dfrbp_1 _20052_ (.CLK(net5575),
    .RESET_B(net6084),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][11] ),
    .Q_N(_09378_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][11] ));
 sg13g2_dfrbp_1 _20053_ (.CLK(net5577),
    .RESET_B(net6086),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][12] ),
    .Q_N(_09379_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][12] ));
 sg13g2_dfrbp_1 _20054_ (.CLK(net5597),
    .RESET_B(net6106),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][13] ),
    .Q_N(_09380_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][13] ));
 sg13g2_dfrbp_1 _20055_ (.CLK(net5597),
    .RESET_B(net6106),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][14] ),
    .Q_N(_09381_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][14] ));
 sg13g2_dfrbp_1 _20056_ (.CLK(net5529),
    .RESET_B(net6038),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][15] ),
    .Q_N(_09382_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][15] ));
 sg13g2_dfrbp_1 _20057_ (.CLK(net5481),
    .RESET_B(net5990),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][16] ),
    .Q_N(_09383_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][16] ));
 sg13g2_dfrbp_1 _20058_ (.CLK(net5479),
    .RESET_B(net5988),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][17] ),
    .Q_N(_09384_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][17] ));
 sg13g2_dfrbp_1 _20059_ (.CLK(net5435),
    .RESET_B(net5944),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][18] ),
    .Q_N(_09385_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[4][18] ));
 sg13g2_dfrbp_1 _20060_ (.CLK(net5567),
    .RESET_B(net6076),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][0] ),
    .Q_N(_09386_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][0] ));
 sg13g2_dfrbp_1 _20061_ (.CLK(net5493),
    .RESET_B(net6002),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][1] ),
    .Q_N(_09387_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][1] ));
 sg13g2_dfrbp_1 _20062_ (.CLK(net5499),
    .RESET_B(net6008),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][2] ),
    .Q_N(_09388_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][2] ));
 sg13g2_dfrbp_1 _20063_ (.CLK(net5496),
    .RESET_B(net6005),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][3] ),
    .Q_N(_09389_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][3] ));
 sg13g2_dfrbp_1 _20064_ (.CLK(net5564),
    .RESET_B(net6073),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][4] ),
    .Q_N(_09390_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][4] ));
 sg13g2_dfrbp_1 _20065_ (.CLK(net5570),
    .RESET_B(net6079),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][5] ),
    .Q_N(_09391_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][5] ));
 sg13g2_dfrbp_1 _20066_ (.CLK(net5574),
    .RESET_B(net6083),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][6] ),
    .Q_N(_09392_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][6] ));
 sg13g2_dfrbp_1 _20067_ (.CLK(net5582),
    .RESET_B(net6091),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][7] ),
    .Q_N(_09393_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][7] ));
 sg13g2_dfrbp_1 _20068_ (.CLK(net5582),
    .RESET_B(net6091),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][8] ),
    .Q_N(_09394_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][8] ));
 sg13g2_dfrbp_1 _20069_ (.CLK(net5583),
    .RESET_B(net6092),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][9] ),
    .Q_N(_09395_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][9] ));
 sg13g2_dfrbp_1 _20070_ (.CLK(net5588),
    .RESET_B(net6097),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][10] ),
    .Q_N(_09396_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][10] ));
 sg13g2_dfrbp_1 _20071_ (.CLK(net5575),
    .RESET_B(net6084),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][11] ),
    .Q_N(_09397_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][11] ));
 sg13g2_dfrbp_1 _20072_ (.CLK(net5603),
    .RESET_B(net6112),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][12] ),
    .Q_N(_09398_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][12] ));
 sg13g2_dfrbp_1 _20073_ (.CLK(net5601),
    .RESET_B(net6110),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][13] ),
    .Q_N(_09399_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][13] ));
 sg13g2_dfrbp_1 _20074_ (.CLK(net5595),
    .RESET_B(net6104),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][14] ),
    .Q_N(_09400_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][14] ));
 sg13g2_dfrbp_1 _20075_ (.CLK(net5530),
    .RESET_B(net6039),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][15] ),
    .Q_N(_09401_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][15] ));
 sg13g2_dfrbp_1 _20076_ (.CLK(net5481),
    .RESET_B(net5990),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][16] ),
    .Q_N(_09402_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][16] ));
 sg13g2_dfrbp_1 _20077_ (.CLK(net5479),
    .RESET_B(net5988),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][17] ),
    .Q_N(_09403_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][17] ));
 sg13g2_dfrbp_1 _20078_ (.CLK(net5434),
    .RESET_B(net5943),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][18] ),
    .Q_N(_09404_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[11][18] ));
 sg13g2_dfrbp_1 _20079_ (.CLK(net5567),
    .RESET_B(net6076),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][0] ),
    .Q_N(_09405_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][0] ));
 sg13g2_dfrbp_1 _20080_ (.CLK(net5493),
    .RESET_B(net6002),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][1] ),
    .Q_N(_09406_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][1] ));
 sg13g2_dfrbp_1 _20081_ (.CLK(net5500),
    .RESET_B(net6009),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][2] ),
    .Q_N(_09407_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][2] ));
 sg13g2_dfrbp_1 _20082_ (.CLK(net5501),
    .RESET_B(net6010),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][3] ),
    .Q_N(_09408_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][3] ));
 sg13g2_dfrbp_1 _20083_ (.CLK(net5566),
    .RESET_B(net6075),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][4] ),
    .Q_N(_09409_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][4] ));
 sg13g2_dfrbp_1 _20084_ (.CLK(net5571),
    .RESET_B(net6080),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][5] ),
    .Q_N(_09410_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][5] ));
 sg13g2_dfrbp_1 _20085_ (.CLK(net5572),
    .RESET_B(net6081),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][6] ),
    .Q_N(_09411_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][6] ));
 sg13g2_dfrbp_1 _20086_ (.CLK(net5585),
    .RESET_B(net6094),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][7] ),
    .Q_N(_09412_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][7] ));
 sg13g2_dfrbp_1 _20087_ (.CLK(net5592),
    .RESET_B(net6101),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][8] ),
    .Q_N(_09413_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][8] ));
 sg13g2_dfrbp_1 _20088_ (.CLK(net5585),
    .RESET_B(net6094),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][9] ),
    .Q_N(_09414_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][9] ));
 sg13g2_dfrbp_1 _20089_ (.CLK(net5589),
    .RESET_B(net6097),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][10] ),
    .Q_N(_09415_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][10] ));
 sg13g2_dfrbp_1 _20090_ (.CLK(net5576),
    .RESET_B(net6085),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][11] ),
    .Q_N(_09416_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][11] ));
 sg13g2_dfrbp_1 _20091_ (.CLK(net5577),
    .RESET_B(net6086),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][12] ),
    .Q_N(_09417_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][12] ));
 sg13g2_dfrbp_1 _20092_ (.CLK(net5597),
    .RESET_B(net6106),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][13] ),
    .Q_N(_09418_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][13] ));
 sg13g2_dfrbp_1 _20093_ (.CLK(net5597),
    .RESET_B(net6106),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][14] ),
    .Q_N(_09419_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][14] ));
 sg13g2_dfrbp_1 _20094_ (.CLK(net5529),
    .RESET_B(net6038),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][15] ),
    .Q_N(_09420_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][15] ));
 sg13g2_dfrbp_1 _20095_ (.CLK(net5481),
    .RESET_B(net5990),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][16] ),
    .Q_N(_09421_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][16] ));
 sg13g2_dfrbp_1 _20096_ (.CLK(net5479),
    .RESET_B(net5988),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][17] ),
    .Q_N(_09422_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][17] ));
 sg13g2_dfrbp_1 _20097_ (.CLK(net5434),
    .RESET_B(net5944),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][18] ),
    .Q_N(_09423_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[3][18] ));
 sg13g2_dfrbp_1 _20098_ (.CLK(net5568),
    .RESET_B(net6077),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][0] ),
    .Q_N(_09424_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][0] ));
 sg13g2_dfrbp_1 _20099_ (.CLK(net5493),
    .RESET_B(net6002),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][1] ),
    .Q_N(_09425_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][1] ));
 sg13g2_dfrbp_1 _20100_ (.CLK(net5500),
    .RESET_B(net6009),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][2] ),
    .Q_N(_09426_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][2] ));
 sg13g2_dfrbp_1 _20101_ (.CLK(net5501),
    .RESET_B(net6010),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][3] ),
    .Q_N(_09427_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][3] ));
 sg13g2_dfrbp_1 _20102_ (.CLK(net5566),
    .RESET_B(net6075),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][4] ),
    .Q_N(_09428_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][4] ));
 sg13g2_dfrbp_1 _20103_ (.CLK(net5571),
    .RESET_B(net6080),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][5] ),
    .Q_N(_09429_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][5] ));
 sg13g2_dfrbp_1 _20104_ (.CLK(net5572),
    .RESET_B(net6081),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][6] ),
    .Q_N(_09430_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][6] ));
 sg13g2_dfrbp_1 _20105_ (.CLK(net5585),
    .RESET_B(net6094),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][7] ),
    .Q_N(_09431_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][7] ));
 sg13g2_dfrbp_1 _20106_ (.CLK(net5587),
    .RESET_B(net6096),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][8] ),
    .Q_N(_09432_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][8] ));
 sg13g2_dfrbp_1 _20107_ (.CLK(net5586),
    .RESET_B(net6095),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][9] ),
    .Q_N(_09433_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][9] ));
 sg13g2_dfrbp_1 _20108_ (.CLK(net5589),
    .RESET_B(net6098),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][10] ),
    .Q_N(_09434_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][10] ));
 sg13g2_dfrbp_1 _20109_ (.CLK(net5576),
    .RESET_B(net6085),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][11] ),
    .Q_N(_09435_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][11] ));
 sg13g2_dfrbp_1 _20110_ (.CLK(net5577),
    .RESET_B(net6086),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][12] ),
    .Q_N(_09436_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][12] ));
 sg13g2_dfrbp_1 _20111_ (.CLK(net5595),
    .RESET_B(net6104),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][13] ),
    .Q_N(_09437_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][13] ));
 sg13g2_dfrbp_1 _20112_ (.CLK(net5596),
    .RESET_B(net6105),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][14] ),
    .Q_N(_09438_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][14] ));
 sg13g2_dfrbp_1 _20113_ (.CLK(net5529),
    .RESET_B(net6038),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][15] ),
    .Q_N(_09439_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][15] ));
 sg13g2_dfrbp_1 _20114_ (.CLK(net5481),
    .RESET_B(net5990),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][16] ),
    .Q_N(_09440_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][16] ));
 sg13g2_dfrbp_1 _20115_ (.CLK(net5437),
    .RESET_B(net5946),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][17] ),
    .Q_N(_09441_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][17] ));
 sg13g2_dfrbp_1 _20116_ (.CLK(net5435),
    .RESET_B(net5943),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][18] ),
    .Q_N(_09442_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[2][18] ));
 sg13g2_dfrbp_1 _20117_ (.CLK(net5567),
    .RESET_B(net6076),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][0] ),
    .Q_N(_09443_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][0] ));
 sg13g2_dfrbp_1 _20118_ (.CLK(net5493),
    .RESET_B(net6002),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][1] ),
    .Q_N(_09444_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][1] ));
 sg13g2_dfrbp_1 _20119_ (.CLK(net5498),
    .RESET_B(net6007),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][2] ),
    .Q_N(_09445_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][2] ));
 sg13g2_dfrbp_1 _20120_ (.CLK(net5496),
    .RESET_B(net6005),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][3] ),
    .Q_N(_09446_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][3] ));
 sg13g2_dfrbp_1 _20121_ (.CLK(net5564),
    .RESET_B(net6073),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][4] ),
    .Q_N(_09447_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][4] ));
 sg13g2_dfrbp_1 _20122_ (.CLK(net5570),
    .RESET_B(net6079),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][5] ),
    .Q_N(_09448_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][5] ));
 sg13g2_dfrbp_1 _20123_ (.CLK(net5572),
    .RESET_B(net6081),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][6] ),
    .Q_N(_09449_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][6] ));
 sg13g2_dfrbp_1 _20124_ (.CLK(net5584),
    .RESET_B(net6093),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][7] ),
    .Q_N(_09450_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][7] ));
 sg13g2_dfrbp_1 _20125_ (.CLK(net5587),
    .RESET_B(net6096),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][8] ),
    .Q_N(_09451_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][8] ));
 sg13g2_dfrbp_1 _20126_ (.CLK(net5583),
    .RESET_B(net6092),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][9] ),
    .Q_N(_09452_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][9] ));
 sg13g2_dfrbp_1 _20127_ (.CLK(net5575),
    .RESET_B(net6084),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][10] ),
    .Q_N(_09453_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][10] ));
 sg13g2_dfrbp_1 _20128_ (.CLK(net5575),
    .RESET_B(net6084),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][11] ),
    .Q_N(_09454_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][11] ));
 sg13g2_dfrbp_1 _20129_ (.CLK(net5600),
    .RESET_B(net6109),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][12] ),
    .Q_N(_09455_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][12] ));
 sg13g2_dfrbp_1 _20130_ (.CLK(net5601),
    .RESET_B(net6110),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][13] ),
    .Q_N(_09456_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][13] ));
 sg13g2_dfrbp_1 _20131_ (.CLK(net5595),
    .RESET_B(net6104),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][14] ),
    .Q_N(_09457_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][14] ));
 sg13g2_dfrbp_1 _20132_ (.CLK(net5530),
    .RESET_B(net6039),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][15] ),
    .Q_N(_09458_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][15] ));
 sg13g2_dfrbp_1 _20133_ (.CLK(net5482),
    .RESET_B(net5991),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][16] ),
    .Q_N(_09459_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][16] ));
 sg13g2_dfrbp_1 _20134_ (.CLK(net5436),
    .RESET_B(net5945),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][17] ),
    .Q_N(_09460_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][17] ));
 sg13g2_dfrbp_1 _20135_ (.CLK(net5434),
    .RESET_B(net5943),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[7][18] ),
    .Q_N(_09461_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[8][18] ));
 sg13g2_dfrbp_1 _20136_ (.CLK(net5568),
    .RESET_B(net6077),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][0] ),
    .Q_N(_09462_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][0] ));
 sg13g2_dfrbp_1 _20137_ (.CLK(net5495),
    .RESET_B(net6004),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][1] ),
    .Q_N(_09463_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][1] ));
 sg13g2_dfrbp_1 _20138_ (.CLK(net5498),
    .RESET_B(net6007),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][2] ),
    .Q_N(_09464_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][2] ));
 sg13g2_dfrbp_1 _20139_ (.CLK(net5497),
    .RESET_B(net6006),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][3] ),
    .Q_N(_09465_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][3] ));
 sg13g2_dfrbp_1 _20140_ (.CLK(net5565),
    .RESET_B(net6074),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][4] ),
    .Q_N(_09466_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][4] ));
 sg13g2_dfrbp_1 _20141_ (.CLK(net5571),
    .RESET_B(net6080),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][5] ),
    .Q_N(_09467_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][5] ));
 sg13g2_dfrbp_1 _20142_ (.CLK(net5572),
    .RESET_B(net6081),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][6] ),
    .Q_N(_09468_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][6] ));
 sg13g2_dfrbp_1 _20143_ (.CLK(net5585),
    .RESET_B(net6094),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][7] ),
    .Q_N(_09469_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][7] ));
 sg13g2_dfrbp_1 _20144_ (.CLK(net5585),
    .RESET_B(net6094),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][8] ),
    .Q_N(_09470_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][8] ));
 sg13g2_dfrbp_1 _20145_ (.CLK(net5586),
    .RESET_B(net6095),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][9] ),
    .Q_N(_09471_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][9] ));
 sg13g2_dfrbp_1 _20146_ (.CLK(net5583),
    .RESET_B(net6092),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][10] ),
    .Q_N(_09472_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][10] ));
 sg13g2_dfrbp_1 _20147_ (.CLK(net5576),
    .RESET_B(net6085),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][11] ),
    .Q_N(_09473_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][11] ));
 sg13g2_dfrbp_1 _20148_ (.CLK(net5577),
    .RESET_B(net6086),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][12] ),
    .Q_N(_09474_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][12] ));
 sg13g2_dfrbp_1 _20149_ (.CLK(net5598),
    .RESET_B(net6107),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][13] ),
    .Q_N(_09475_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][13] ));
 sg13g2_dfrbp_1 _20150_ (.CLK(net5596),
    .RESET_B(net6105),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][14] ),
    .Q_N(_09476_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][14] ));
 sg13g2_dfrbp_1 _20151_ (.CLK(net5529),
    .RESET_B(net6038),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][15] ),
    .Q_N(_09477_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][15] ));
 sg13g2_dfrbp_1 _20152_ (.CLK(net5481),
    .RESET_B(net5990),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][16] ),
    .Q_N(_09478_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][16] ));
 sg13g2_dfrbp_1 _20153_ (.CLK(net5480),
    .RESET_B(net5989),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][17] ),
    .Q_N(_09479_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][17] ));
 sg13g2_dfrbp_1 _20154_ (.CLK(net5433),
    .RESET_B(net5942),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][18] ),
    .Q_N(_09480_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[1][18] ));
 sg13g2_dfrbp_1 _20155_ (.CLK(net5568),
    .RESET_B(net6077),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.u_mux_shift.sum_res ),
    .Q_N(_00288_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][0] ));
 sg13g2_dfrbp_1 _20156_ (.CLK(net5495),
    .RESET_B(net6004),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .Q_N(_00299_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][1] ));
 sg13g2_dfrbp_1 _20157_ (.CLK(net5498),
    .RESET_B(net6007),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .Q_N(_00306_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][2] ));
 sg13g2_dfrbp_1 _20158_ (.CLK(net5497),
    .RESET_B(net6006),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .Q_N(_00313_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][3] ));
 sg13g2_dfrbp_1 _20159_ (.CLK(net5565),
    .RESET_B(net6074),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .Q_N(_00322_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][4] ));
 sg13g2_dfrbp_1 _20160_ (.CLK(net5571),
    .RESET_B(net6080),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .Q_N(_00331_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][5] ));
 sg13g2_dfrbp_1 _20161_ (.CLK(net5572),
    .RESET_B(net6081),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .Q_N(_00338_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][6] ));
 sg13g2_dfrbp_1 _20162_ (.CLK(net5585),
    .RESET_B(net6094),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .Q_N(_00345_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][7] ));
 sg13g2_dfrbp_1 _20163_ (.CLK(net5586),
    .RESET_B(net6095),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .Q_N(_00354_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][8] ));
 sg13g2_dfrbp_1 _20164_ (.CLK(net5586),
    .RESET_B(net6095),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .Q_N(_00363_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][9] ));
 sg13g2_dfrbp_1 _20165_ (.CLK(net5582),
    .RESET_B(net6091),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .Q_N(_00370_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][10] ));
 sg13g2_dfrbp_1 _20166_ (.CLK(net5575),
    .RESET_B(net6084),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .Q_N(_00377_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][11] ));
 sg13g2_dfrbp_1 _20167_ (.CLK(net5577),
    .RESET_B(net6086),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .Q_N(_00386_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][12] ));
 sg13g2_dfrbp_1 _20168_ (.CLK(net5598),
    .RESET_B(net6107),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .Q_N(_00395_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][13] ));
 sg13g2_dfrbp_1 _20169_ (.CLK(net5598),
    .RESET_B(net6107),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .Q_N(_00402_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][14] ));
 sg13g2_dfrbp_1 _20170_ (.CLK(net5529),
    .RESET_B(net6038),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .Q_N(_00409_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][15] ));
 sg13g2_dfrbp_1 _20171_ (.CLK(net5481),
    .RESET_B(net5990),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .Q_N(_00418_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][16] ));
 sg13g2_dfrbp_1 _20172_ (.CLK(net5436),
    .RESET_B(net5945),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .Q_N(_00425_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][17] ));
 sg13g2_dfrbp_1 _20173_ (.CLK(net5433),
    .RESET_B(net5942),
    .D(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .Q_N(_00432_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[0][18] ));
 sg13g2_dfrbp_1 _20174_ (.CLK(net5567),
    .RESET_B(net6076),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][0] ),
    .Q_N(_09481_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][0] ));
 sg13g2_dfrbp_1 _20175_ (.CLK(net5493),
    .RESET_B(net6002),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][1] ),
    .Q_N(_09482_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][1] ));
 sg13g2_dfrbp_1 _20176_ (.CLK(net5498),
    .RESET_B(net6007),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][2] ),
    .Q_N(_09483_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][2] ));
 sg13g2_dfrbp_1 _20177_ (.CLK(net5496),
    .RESET_B(net6005),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][3] ),
    .Q_N(_09484_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][3] ));
 sg13g2_dfrbp_1 _20178_ (.CLK(net5564),
    .RESET_B(net6073),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][4] ),
    .Q_N(_09485_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][4] ));
 sg13g2_dfrbp_1 _20179_ (.CLK(net5570),
    .RESET_B(net6079),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][5] ),
    .Q_N(_09486_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][5] ));
 sg13g2_dfrbp_1 _20180_ (.CLK(net5572),
    .RESET_B(net6081),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][6] ),
    .Q_N(_09487_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][6] ));
 sg13g2_dfrbp_1 _20181_ (.CLK(net5582),
    .RESET_B(net6091),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][7] ),
    .Q_N(_09488_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][7] ));
 sg13g2_dfrbp_1 _20182_ (.CLK(net5582),
    .RESET_B(net6091),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][8] ),
    .Q_N(_09489_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][8] ));
 sg13g2_dfrbp_1 _20183_ (.CLK(net5583),
    .RESET_B(net6092),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][9] ),
    .Q_N(_09490_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][9] ));
 sg13g2_dfrbp_1 _20184_ (.CLK(net5575),
    .RESET_B(net6084),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][10] ),
    .Q_N(_09491_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][10] ));
 sg13g2_dfrbp_1 _20185_ (.CLK(net5577),
    .RESET_B(net6084),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][11] ),
    .Q_N(_09492_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][11] ));
 sg13g2_dfrbp_1 _20186_ (.CLK(net5603),
    .RESET_B(net6112),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][12] ),
    .Q_N(_09493_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][12] ));
 sg13g2_dfrbp_1 _20187_ (.CLK(net5600),
    .RESET_B(net6109),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][13] ),
    .Q_N(_09494_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][13] ));
 sg13g2_dfrbp_1 _20188_ (.CLK(net5595),
    .RESET_B(net6104),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][14] ),
    .Q_N(_09495_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][14] ));
 sg13g2_dfrbp_1 _20189_ (.CLK(net5530),
    .RESET_B(net6039),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][15] ),
    .Q_N(_09496_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][15] ));
 sg13g2_dfrbp_1 _20190_ (.CLK(net5482),
    .RESET_B(net5991),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][16] ),
    .Q_N(_09497_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][16] ));
 sg13g2_dfrbp_1 _20191_ (.CLK(net5479),
    .RESET_B(net5988),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][17] ),
    .Q_N(_09498_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][17] ));
 sg13g2_dfrbp_1 _20192_ (.CLK(net5434),
    .RESET_B(net5943),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[9][18] ),
    .Q_N(_09499_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[6].u_delay_line.buffer[10][18] ));
 sg13g2_dfrbp_1 _20193_ (.CLK(net5603),
    .RESET_B(net6112),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][0] ),
    .Q_N(_09500_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][0] ));
 sg13g2_dfrbp_1 _20194_ (.CLK(net5616),
    .RESET_B(net6125),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][1] ),
    .Q_N(_09501_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][1] ));
 sg13g2_dfrbp_1 _20195_ (.CLK(net5614),
    .RESET_B(net6123),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][2] ),
    .Q_N(_09502_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][2] ));
 sg13g2_dfrbp_1 _20196_ (.CLK(net5650),
    .RESET_B(net6159),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][3] ),
    .Q_N(_09503_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][3] ));
 sg13g2_dfrbp_1 _20197_ (.CLK(net5658),
    .RESET_B(net6168),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][4] ),
    .Q_N(_09504_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][4] ));
 sg13g2_dfrbp_1 _20198_ (.CLK(net5644),
    .RESET_B(net6153),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][5] ),
    .Q_N(_09505_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][5] ));
 sg13g2_dfrbp_1 _20199_ (.CLK(net5646),
    .RESET_B(net6155),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][6] ),
    .Q_N(_09506_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][6] ));
 sg13g2_dfrbp_1 _20200_ (.CLK(net5672),
    .RESET_B(net6182),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][7] ),
    .Q_N(_09507_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][7] ));
 sg13g2_dfrbp_1 _20201_ (.CLK(net5670),
    .RESET_B(net6180),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][8] ),
    .Q_N(_09508_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][8] ));
 sg13g2_dfrbp_1 _20202_ (.CLK(net5676),
    .RESET_B(net6186),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][9] ),
    .Q_N(_09509_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][9] ));
 sg13g2_dfrbp_1 _20203_ (.CLK(net5676),
    .RESET_B(net6186),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][10] ),
    .Q_N(_09510_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][10] ));
 sg13g2_dfrbp_1 _20204_ (.CLK(net5681),
    .RESET_B(net6191),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][11] ),
    .Q_N(_09511_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][11] ));
 sg13g2_dfrbp_1 _20205_ (.CLK(net5677),
    .RESET_B(net6187),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][12] ),
    .Q_N(_09512_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][12] ));
 sg13g2_dfrbp_1 _20206_ (.CLK(net5664),
    .RESET_B(net6174),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][13] ),
    .Q_N(_09513_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][13] ));
 sg13g2_dfrbp_1 _20207_ (.CLK(net5656),
    .RESET_B(net6166),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][14] ),
    .Q_N(_09514_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][14] ));
 sg13g2_dfrbp_1 _20208_ (.CLK(net5652),
    .RESET_B(net6162),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][15] ),
    .Q_N(_09515_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][15] ));
 sg13g2_dfrbp_1 _20209_ (.CLK(net5621),
    .RESET_B(net6130),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][16] ),
    .Q_N(_09516_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][16] ));
 sg13g2_dfrbp_1 _20210_ (.CLK(net5605),
    .RESET_B(net6114),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][17] ),
    .Q_N(_09517_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][17] ));
 sg13g2_dfrbp_1 _20211_ (.CLK(net5590),
    .RESET_B(net6098),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][18] ),
    .Q_N(_09518_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][18] ));
 sg13g2_dfrbp_1 _20212_ (.CLK(net5604),
    .RESET_B(net6113),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][0] ),
    .Q_N(_09519_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][0] ));
 sg13g2_dfrbp_1 _20213_ (.CLK(net5616),
    .RESET_B(net6125),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][1] ),
    .Q_N(_09520_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][1] ));
 sg13g2_dfrbp_1 _20214_ (.CLK(net5613),
    .RESET_B(net6122),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][2] ),
    .Q_N(_09521_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][2] ));
 sg13g2_dfrbp_1 _20215_ (.CLK(net5650),
    .RESET_B(net6159),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][3] ),
    .Q_N(_09522_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][3] ));
 sg13g2_dfrbp_1 _20216_ (.CLK(net5659),
    .RESET_B(net6169),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][4] ),
    .Q_N(_09523_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][4] ));
 sg13g2_dfrbp_1 _20217_ (.CLK(net5668),
    .RESET_B(net6178),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][5] ),
    .Q_N(_09524_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][5] ));
 sg13g2_dfrbp_1 _20218_ (.CLK(net5646),
    .RESET_B(net6155),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][6] ),
    .Q_N(_09525_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][6] ));
 sg13g2_dfrbp_1 _20219_ (.CLK(net5672),
    .RESET_B(net6182),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][7] ),
    .Q_N(_09526_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][7] ));
 sg13g2_dfrbp_1 _20220_ (.CLK(net5670),
    .RESET_B(net6180),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][8] ),
    .Q_N(_09527_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][8] ));
 sg13g2_dfrbp_1 _20221_ (.CLK(net5669),
    .RESET_B(net6179),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][9] ),
    .Q_N(_09528_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][9] ));
 sg13g2_dfrbp_1 _20222_ (.CLK(net5675),
    .RESET_B(net6185),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][10] ),
    .Q_N(_09529_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][10] ));
 sg13g2_dfrbp_1 _20223_ (.CLK(net5678),
    .RESET_B(net6188),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][11] ),
    .Q_N(_09530_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][11] ));
 sg13g2_dfrbp_1 _20224_ (.CLK(net5677),
    .RESET_B(net6187),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][12] ),
    .Q_N(_09531_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][12] ));
 sg13g2_dfrbp_1 _20225_ (.CLK(net5664),
    .RESET_B(net6174),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][13] ),
    .Q_N(_09532_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][13] ));
 sg13g2_dfrbp_1 _20226_ (.CLK(net5655),
    .RESET_B(net6165),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][14] ),
    .Q_N(_09533_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][14] ));
 sg13g2_dfrbp_1 _20227_ (.CLK(net5652),
    .RESET_B(net6162),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][15] ),
    .Q_N(_09534_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][15] ));
 sg13g2_dfrbp_1 _20228_ (.CLK(net5621),
    .RESET_B(net6130),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][16] ),
    .Q_N(_09535_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][16] ));
 sg13g2_dfrbp_1 _20229_ (.CLK(net5610),
    .RESET_B(net6119),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][17] ),
    .Q_N(_09536_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][17] ));
 sg13g2_dfrbp_1 _20230_ (.CLK(net5612),
    .RESET_B(net6121),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][18] ),
    .Q_N(_09537_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][18] ));
 sg13g2_dfrbp_1 _20231_ (.CLK(net5603),
    .RESET_B(net6112),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][0] ),
    .Q_N(_09538_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][0] ));
 sg13g2_dfrbp_1 _20232_ (.CLK(net5616),
    .RESET_B(net6125),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][1] ),
    .Q_N(_09539_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][1] ));
 sg13g2_dfrbp_1 _20233_ (.CLK(net5619),
    .RESET_B(net6128),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][2] ),
    .Q_N(_09540_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][2] ));
 sg13g2_dfrbp_1 _20234_ (.CLK(net5650),
    .RESET_B(net6159),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][3] ),
    .Q_N(_09541_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][3] ));
 sg13g2_dfrbp_1 _20235_ (.CLK(net5659),
    .RESET_B(net6169),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][4] ),
    .Q_N(_09542_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][4] ));
 sg13g2_dfrbp_1 _20236_ (.CLK(net5644),
    .RESET_B(net6153),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][5] ),
    .Q_N(_09543_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][5] ));
 sg13g2_dfrbp_1 _20237_ (.CLK(net5647),
    .RESET_B(net6156),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][6] ),
    .Q_N(_09544_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][6] ));
 sg13g2_dfrbp_1 _20238_ (.CLK(net5673),
    .RESET_B(net6183),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][7] ),
    .Q_N(_09545_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][7] ));
 sg13g2_dfrbp_1 _20239_ (.CLK(net5671),
    .RESET_B(net6181),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][8] ),
    .Q_N(_09546_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][8] ));
 sg13g2_dfrbp_1 _20240_ (.CLK(net5680),
    .RESET_B(net6190),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][9] ),
    .Q_N(_09547_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][9] ));
 sg13g2_dfrbp_1 _20241_ (.CLK(net5676),
    .RESET_B(net6186),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][10] ),
    .Q_N(_09548_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][10] ));
 sg13g2_dfrbp_1 _20242_ (.CLK(net5681),
    .RESET_B(net6191),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][11] ),
    .Q_N(_09549_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][11] ));
 sg13g2_dfrbp_1 _20243_ (.CLK(net5684),
    .RESET_B(net6194),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][12] ),
    .Q_N(_09550_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][12] ));
 sg13g2_dfrbp_1 _20244_ (.CLK(net5665),
    .RESET_B(net6175),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][13] ),
    .Q_N(_09551_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][13] ));
 sg13g2_dfrbp_1 _20245_ (.CLK(net5656),
    .RESET_B(net6166),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][14] ),
    .Q_N(_09552_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][14] ));
 sg13g2_dfrbp_1 _20246_ (.CLK(net5652),
    .RESET_B(net6162),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][15] ),
    .Q_N(_09553_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][15] ));
 sg13g2_dfrbp_1 _20247_ (.CLK(net5620),
    .RESET_B(net6129),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][16] ),
    .Q_N(_09554_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][16] ));
 sg13g2_dfrbp_1 _20248_ (.CLK(net5605),
    .RESET_B(net6114),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][17] ),
    .Q_N(_09555_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][17] ));
 sg13g2_dfrbp_1 _20249_ (.CLK(net5590),
    .RESET_B(net6098),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][18] ),
    .Q_N(_09556_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[6][18] ));
 sg13g2_dfrbp_1 _20250_ (.CLK(net5604),
    .RESET_B(net6113),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][0] ),
    .Q_N(_09557_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][0] ));
 sg13g2_dfrbp_1 _20251_ (.CLK(net5620),
    .RESET_B(net6129),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][1] ),
    .Q_N(_09558_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][1] ));
 sg13g2_dfrbp_1 _20252_ (.CLK(net5613),
    .RESET_B(net6122),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][2] ),
    .Q_N(_09559_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][2] ));
 sg13g2_dfrbp_1 _20253_ (.CLK(net5650),
    .RESET_B(net6159),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][3] ),
    .Q_N(_09560_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][3] ));
 sg13g2_dfrbp_1 _20254_ (.CLK(net5658),
    .RESET_B(net6168),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][4] ),
    .Q_N(_09561_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][4] ));
 sg13g2_dfrbp_1 _20255_ (.CLK(net5663),
    .RESET_B(net6173),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][5] ),
    .Q_N(_09562_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][5] ));
 sg13g2_dfrbp_1 _20256_ (.CLK(net5647),
    .RESET_B(net6156),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][6] ),
    .Q_N(_09563_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][6] ));
 sg13g2_dfrbp_1 _20257_ (.CLK(net5673),
    .RESET_B(net6183),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][7] ),
    .Q_N(_09564_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][7] ));
 sg13g2_dfrbp_1 _20258_ (.CLK(net5671),
    .RESET_B(net6181),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][8] ),
    .Q_N(_09565_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][8] ));
 sg13g2_dfrbp_1 _20259_ (.CLK(net5676),
    .RESET_B(net6186),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][9] ),
    .Q_N(_09566_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][9] ));
 sg13g2_dfrbp_1 _20260_ (.CLK(net5680),
    .RESET_B(net6190),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][10] ),
    .Q_N(_09567_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][10] ));
 sg13g2_dfrbp_1 _20261_ (.CLK(net5681),
    .RESET_B(net6191),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][11] ),
    .Q_N(_09568_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][11] ));
 sg13g2_dfrbp_1 _20262_ (.CLK(net5684),
    .RESET_B(net6194),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][12] ),
    .Q_N(_09569_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][12] ));
 sg13g2_dfrbp_1 _20263_ (.CLK(net5665),
    .RESET_B(net6175),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][13] ),
    .Q_N(_09570_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][13] ));
 sg13g2_dfrbp_1 _20264_ (.CLK(net5656),
    .RESET_B(net6166),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][14] ),
    .Q_N(_09571_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][14] ));
 sg13g2_dfrbp_1 _20265_ (.CLK(net5654),
    .RESET_B(net6164),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][15] ),
    .Q_N(_09572_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][15] ));
 sg13g2_dfrbp_1 _20266_ (.CLK(net5620),
    .RESET_B(net6130),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][16] ),
    .Q_N(_09573_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][16] ));
 sg13g2_dfrbp_1 _20267_ (.CLK(net5604),
    .RESET_B(net6113),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][17] ),
    .Q_N(_09574_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][17] ));
 sg13g2_dfrbp_1 _20268_ (.CLK(net5612),
    .RESET_B(net6121),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][18] ),
    .Q_N(_09575_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][18] ));
 sg13g2_dfrbp_1 _20269_ (.CLK(net5601),
    .RESET_B(net6110),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][0] ),
    .Q_N(_09576_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][0] ));
 sg13g2_dfrbp_1 _20270_ (.CLK(net5616),
    .RESET_B(net6125),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][1] ),
    .Q_N(_09577_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][1] ));
 sg13g2_dfrbp_1 _20271_ (.CLK(net5614),
    .RESET_B(net6123),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][2] ),
    .Q_N(_09578_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][2] ));
 sg13g2_dfrbp_1 _20272_ (.CLK(net5630),
    .RESET_B(net6139),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][3] ),
    .Q_N(_09579_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][3] ));
 sg13g2_dfrbp_1 _20273_ (.CLK(net5658),
    .RESET_B(net6168),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][4] ),
    .Q_N(_09580_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][4] ));
 sg13g2_dfrbp_1 _20274_ (.CLK(net5644),
    .RESET_B(net6153),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][5] ),
    .Q_N(_09581_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][5] ));
 sg13g2_dfrbp_1 _20275_ (.CLK(net5647),
    .RESET_B(net6156),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][6] ),
    .Q_N(_09582_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][6] ));
 sg13g2_dfrbp_1 _20276_ (.CLK(net5672),
    .RESET_B(net6182),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][7] ),
    .Q_N(_09583_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][7] ));
 sg13g2_dfrbp_1 _20277_ (.CLK(net5671),
    .RESET_B(net6181),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][8] ),
    .Q_N(_09584_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][8] ));
 sg13g2_dfrbp_1 _20278_ (.CLK(net5680),
    .RESET_B(net6190),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][9] ),
    .Q_N(_09585_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][9] ));
 sg13g2_dfrbp_1 _20279_ (.CLK(net5675),
    .RESET_B(net6185),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][10] ),
    .Q_N(_09586_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][10] ));
 sg13g2_dfrbp_1 _20280_ (.CLK(net5681),
    .RESET_B(net6191),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][11] ),
    .Q_N(_09587_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][11] ));
 sg13g2_dfrbp_1 _20281_ (.CLK(net5684),
    .RESET_B(net6194),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][12] ),
    .Q_N(_09588_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][12] ));
 sg13g2_dfrbp_1 _20282_ (.CLK(net5664),
    .RESET_B(net6174),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][13] ),
    .Q_N(_09589_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][13] ));
 sg13g2_dfrbp_1 _20283_ (.CLK(net5656),
    .RESET_B(net6166),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][14] ),
    .Q_N(_09590_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][14] ));
 sg13g2_dfrbp_1 _20284_ (.CLK(net5652),
    .RESET_B(net6162),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][15] ),
    .Q_N(_09591_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][15] ));
 sg13g2_dfrbp_1 _20285_ (.CLK(net5611),
    .RESET_B(net6120),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][16] ),
    .Q_N(_09592_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][16] ));
 sg13g2_dfrbp_1 _20286_ (.CLK(net5605),
    .RESET_B(net6114),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][17] ),
    .Q_N(_09593_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][17] ));
 sg13g2_dfrbp_1 _20287_ (.CLK(net5590),
    .RESET_B(net6098),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][18] ),
    .Q_N(_09594_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[5][18] ));
 sg13g2_dfrbp_1 _20288_ (.CLK(net5604),
    .RESET_B(net6113),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][0] ),
    .Q_N(_09595_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][0] ));
 sg13g2_dfrbp_1 _20289_ (.CLK(net5617),
    .RESET_B(net6125),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][1] ),
    .Q_N(_09596_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][1] ));
 sg13g2_dfrbp_1 _20290_ (.CLK(net5613),
    .RESET_B(net6122),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][2] ),
    .Q_N(_09597_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][2] ));
 sg13g2_dfrbp_1 _20291_ (.CLK(net5651),
    .RESET_B(net6159),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][3] ),
    .Q_N(_09598_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][3] ));
 sg13g2_dfrbp_1 _20292_ (.CLK(net5659),
    .RESET_B(net6169),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][4] ),
    .Q_N(_09599_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][4] ));
 sg13g2_dfrbp_1 _20293_ (.CLK(net5663),
    .RESET_B(net6173),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][5] ),
    .Q_N(_09600_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][5] ));
 sg13g2_dfrbp_1 _20294_ (.CLK(net5646),
    .RESET_B(net6155),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][6] ),
    .Q_N(_09601_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][6] ));
 sg13g2_dfrbp_1 _20295_ (.CLK(net5672),
    .RESET_B(net6182),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][7] ),
    .Q_N(_09602_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][7] ));
 sg13g2_dfrbp_1 _20296_ (.CLK(net5670),
    .RESET_B(net6180),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][8] ),
    .Q_N(_09603_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][8] ));
 sg13g2_dfrbp_1 _20297_ (.CLK(net5669),
    .RESET_B(net6179),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][9] ),
    .Q_N(_09604_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][9] ));
 sg13g2_dfrbp_1 _20298_ (.CLK(net5675),
    .RESET_B(net6185),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][10] ),
    .Q_N(_09605_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][10] ));
 sg13g2_dfrbp_1 _20299_ (.CLK(net5678),
    .RESET_B(net6188),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][11] ),
    .Q_N(_09606_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][11] ));
 sg13g2_dfrbp_1 _20300_ (.CLK(net5677),
    .RESET_B(net6187),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][12] ),
    .Q_N(_09607_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][12] ));
 sg13g2_dfrbp_1 _20301_ (.CLK(net5664),
    .RESET_B(net6174),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][13] ),
    .Q_N(_09608_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][13] ));
 sg13g2_dfrbp_1 _20302_ (.CLK(net5655),
    .RESET_B(net6165),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][14] ),
    .Q_N(_09609_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][14] ));
 sg13g2_dfrbp_1 _20303_ (.CLK(net5652),
    .RESET_B(net6162),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][15] ),
    .Q_N(_09610_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][15] ));
 sg13g2_dfrbp_1 _20304_ (.CLK(net5620),
    .RESET_B(net6129),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][16] ),
    .Q_N(_09611_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][16] ));
 sg13g2_dfrbp_1 _20305_ (.CLK(net5610),
    .RESET_B(net6119),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][17] ),
    .Q_N(_09612_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][17] ));
 sg13g2_dfrbp_1 _20306_ (.CLK(net5612),
    .RESET_B(net6121),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[12][18] ),
    .Q_N(_09613_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][18] ));
 sg13g2_dfrbp_1 _20307_ (.CLK(net5601),
    .RESET_B(net6110),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][0] ),
    .Q_N(_09614_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][0] ));
 sg13g2_dfrbp_1 _20308_ (.CLK(net5616),
    .RESET_B(net6126),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][1] ),
    .Q_N(_09615_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][1] ));
 sg13g2_dfrbp_1 _20309_ (.CLK(net5619),
    .RESET_B(net6128),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][2] ),
    .Q_N(_09616_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][2] ));
 sg13g2_dfrbp_1 _20310_ (.CLK(net5630),
    .RESET_B(net6139),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][3] ),
    .Q_N(_09617_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][3] ));
 sg13g2_dfrbp_1 _20311_ (.CLK(net5658),
    .RESET_B(net6168),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][4] ),
    .Q_N(_09618_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][4] ));
 sg13g2_dfrbp_1 _20312_ (.CLK(net5645),
    .RESET_B(net6154),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][5] ),
    .Q_N(_09619_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][5] ));
 sg13g2_dfrbp_1 _20313_ (.CLK(net5647),
    .RESET_B(net6156),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][6] ),
    .Q_N(_09620_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][6] ));
 sg13g2_dfrbp_1 _20314_ (.CLK(net5672),
    .RESET_B(net6182),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][7] ),
    .Q_N(_09621_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][7] ));
 sg13g2_dfrbp_1 _20315_ (.CLK(net5671),
    .RESET_B(net6181),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][8] ),
    .Q_N(_09622_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][8] ));
 sg13g2_dfrbp_1 _20316_ (.CLK(net5680),
    .RESET_B(net6190),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][9] ),
    .Q_N(_09623_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][9] ));
 sg13g2_dfrbp_1 _20317_ (.CLK(net5675),
    .RESET_B(net6185),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][10] ),
    .Q_N(_09624_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][10] ));
 sg13g2_dfrbp_1 _20318_ (.CLK(net5678),
    .RESET_B(net6188),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][11] ),
    .Q_N(_09625_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][11] ));
 sg13g2_dfrbp_1 _20319_ (.CLK(net5684),
    .RESET_B(net6194),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][12] ),
    .Q_N(_09626_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][12] ));
 sg13g2_dfrbp_1 _20320_ (.CLK(net5665),
    .RESET_B(net6175),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][13] ),
    .Q_N(_09627_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][13] ));
 sg13g2_dfrbp_1 _20321_ (.CLK(net5656),
    .RESET_B(net6166),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][14] ),
    .Q_N(_09628_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][14] ));
 sg13g2_dfrbp_1 _20322_ (.CLK(net5652),
    .RESET_B(net6162),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][15] ),
    .Q_N(_09629_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][15] ));
 sg13g2_dfrbp_1 _20323_ (.CLK(net5611),
    .RESET_B(net6120),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][16] ),
    .Q_N(_09630_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][16] ));
 sg13g2_dfrbp_1 _20324_ (.CLK(net5610),
    .RESET_B(net6119),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][17] ),
    .Q_N(_09631_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][17] ));
 sg13g2_dfrbp_1 _20325_ (.CLK(net5590),
    .RESET_B(net6098),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][18] ),
    .Q_N(_09632_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[4][18] ));
 sg13g2_dfrbp_1 _20326_ (.CLK(net5604),
    .RESET_B(net6113),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][0] ),
    .Q_N(_09633_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][0] ));
 sg13g2_dfrbp_1 _20327_ (.CLK(net5616),
    .RESET_B(net6125),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][1] ),
    .Q_N(_09634_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][1] ));
 sg13g2_dfrbp_1 _20328_ (.CLK(net5613),
    .RESET_B(net6122),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][2] ),
    .Q_N(_09635_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][2] ));
 sg13g2_dfrbp_1 _20329_ (.CLK(net5650),
    .RESET_B(net6159),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][3] ),
    .Q_N(_09636_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][3] ));
 sg13g2_dfrbp_1 _20330_ (.CLK(net5658),
    .RESET_B(net6168),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][4] ),
    .Q_N(_09637_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][4] ));
 sg13g2_dfrbp_1 _20331_ (.CLK(net5668),
    .RESET_B(net6178),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][5] ),
    .Q_N(_09638_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][5] ));
 sg13g2_dfrbp_1 _20332_ (.CLK(net5646),
    .RESET_B(net6155),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][6] ),
    .Q_N(_09639_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][6] ));
 sg13g2_dfrbp_1 _20333_ (.CLK(net5673),
    .RESET_B(net6183),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][7] ),
    .Q_N(_09640_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][7] ));
 sg13g2_dfrbp_1 _20334_ (.CLK(net5670),
    .RESET_B(net6180),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][8] ),
    .Q_N(_09641_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][8] ));
 sg13g2_dfrbp_1 _20335_ (.CLK(net5669),
    .RESET_B(net6179),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][9] ),
    .Q_N(_09642_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][9] ));
 sg13g2_dfrbp_1 _20336_ (.CLK(net5675),
    .RESET_B(net6185),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][10] ),
    .Q_N(_09643_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][10] ));
 sg13g2_dfrbp_1 _20337_ (.CLK(net5681),
    .RESET_B(net6191),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][11] ),
    .Q_N(_09644_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][11] ));
 sg13g2_dfrbp_1 _20338_ (.CLK(net5677),
    .RESET_B(net6187),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][12] ),
    .Q_N(_09645_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][12] ));
 sg13g2_dfrbp_1 _20339_ (.CLK(net5664),
    .RESET_B(net6174),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][13] ),
    .Q_N(_09646_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][13] ));
 sg13g2_dfrbp_1 _20340_ (.CLK(net5656),
    .RESET_B(net6166),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][14] ),
    .Q_N(_09647_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][14] ));
 sg13g2_dfrbp_1 _20341_ (.CLK(net5653),
    .RESET_B(net6163),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][15] ),
    .Q_N(_09648_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][15] ));
 sg13g2_dfrbp_1 _20342_ (.CLK(net5621),
    .RESET_B(net6130),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][16] ),
    .Q_N(_09649_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][16] ));
 sg13g2_dfrbp_1 _20343_ (.CLK(net5610),
    .RESET_B(net6119),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][17] ),
    .Q_N(_09650_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][17] ));
 sg13g2_dfrbp_1 _20344_ (.CLK(net5612),
    .RESET_B(net6121),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][18] ),
    .Q_N(_09651_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[11][18] ));
 sg13g2_dfrbp_1 _20345_ (.CLK(net5602),
    .RESET_B(net6111),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][0] ),
    .Q_N(_09652_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][0] ));
 sg13g2_dfrbp_1 _20346_ (.CLK(net5616),
    .RESET_B(net6125),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][1] ),
    .Q_N(_09653_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][1] ));
 sg13g2_dfrbp_1 _20347_ (.CLK(net5614),
    .RESET_B(net6123),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][2] ),
    .Q_N(_09654_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][2] ));
 sg13g2_dfrbp_1 _20348_ (.CLK(net5630),
    .RESET_B(net6139),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][3] ),
    .Q_N(_09655_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][3] ));
 sg13g2_dfrbp_1 _20349_ (.CLK(net5658),
    .RESET_B(net6168),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][4] ),
    .Q_N(_09656_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][4] ));
 sg13g2_dfrbp_1 _20350_ (.CLK(net5644),
    .RESET_B(net6153),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][5] ),
    .Q_N(_09657_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][5] ));
 sg13g2_dfrbp_1 _20351_ (.CLK(net5647),
    .RESET_B(net6156),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][6] ),
    .Q_N(_09658_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][6] ));
 sg13g2_dfrbp_1 _20352_ (.CLK(net5672),
    .RESET_B(net6182),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][7] ),
    .Q_N(_09659_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][7] ));
 sg13g2_dfrbp_1 _20353_ (.CLK(net5671),
    .RESET_B(net6181),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][8] ),
    .Q_N(_09660_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][8] ));
 sg13g2_dfrbp_1 _20354_ (.CLK(net5680),
    .RESET_B(net6190),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][9] ),
    .Q_N(_09661_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][9] ));
 sg13g2_dfrbp_1 _20355_ (.CLK(net5679),
    .RESET_B(net6189),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][10] ),
    .Q_N(_09662_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][10] ));
 sg13g2_dfrbp_1 _20356_ (.CLK(net5677),
    .RESET_B(net6187),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][11] ),
    .Q_N(_09663_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][11] ));
 sg13g2_dfrbp_1 _20357_ (.CLK(net5684),
    .RESET_B(net6194),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][12] ),
    .Q_N(_09664_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][12] ));
 sg13g2_dfrbp_1 _20358_ (.CLK(net5661),
    .RESET_B(net6171),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][13] ),
    .Q_N(_09665_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][13] ));
 sg13g2_dfrbp_1 _20359_ (.CLK(net5655),
    .RESET_B(net6165),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][14] ),
    .Q_N(_09666_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][14] ));
 sg13g2_dfrbp_1 _20360_ (.CLK(net5652),
    .RESET_B(net6162),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][15] ),
    .Q_N(_09667_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][15] ));
 sg13g2_dfrbp_1 _20361_ (.CLK(net5611),
    .RESET_B(net6120),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][16] ),
    .Q_N(_09668_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][16] ));
 sg13g2_dfrbp_1 _20362_ (.CLK(net5611),
    .RESET_B(net6120),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][17] ),
    .Q_N(_09669_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][17] ));
 sg13g2_dfrbp_1 _20363_ (.CLK(net5588),
    .RESET_B(net6097),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][18] ),
    .Q_N(_09670_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[3][18] ));
 sg13g2_dfrbp_1 _20364_ (.CLK(net5604),
    .RESET_B(net6113),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][0] ),
    .Q_N(_09671_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][0] ));
 sg13g2_dfrbp_1 _20365_ (.CLK(net5619),
    .RESET_B(net6128),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][1] ),
    .Q_N(_09672_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][1] ));
 sg13g2_dfrbp_1 _20366_ (.CLK(net5614),
    .RESET_B(net6123),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][2] ),
    .Q_N(_09673_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][2] ));
 sg13g2_dfrbp_1 _20367_ (.CLK(net5650),
    .RESET_B(net6160),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][3] ),
    .Q_N(_09674_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][3] ));
 sg13g2_dfrbp_1 _20368_ (.CLK(net5658),
    .RESET_B(net6168),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][4] ),
    .Q_N(_09675_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][4] ));
 sg13g2_dfrbp_1 _20369_ (.CLK(net5668),
    .RESET_B(net6178),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][5] ),
    .Q_N(_09676_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][5] ));
 sg13g2_dfrbp_1 _20370_ (.CLK(net5646),
    .RESET_B(net6155),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][6] ),
    .Q_N(_09677_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][6] ));
 sg13g2_dfrbp_1 _20371_ (.CLK(net5672),
    .RESET_B(net6182),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][7] ),
    .Q_N(_09678_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][7] ));
 sg13g2_dfrbp_1 _20372_ (.CLK(net5670),
    .RESET_B(net6180),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][8] ),
    .Q_N(_09679_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][8] ));
 sg13g2_dfrbp_1 _20373_ (.CLK(net5669),
    .RESET_B(net6179),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][9] ),
    .Q_N(_09680_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][9] ));
 sg13g2_dfrbp_1 _20374_ (.CLK(net5675),
    .RESET_B(net6185),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][10] ),
    .Q_N(_09681_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][10] ));
 sg13g2_dfrbp_1 _20375_ (.CLK(net5678),
    .RESET_B(net6188),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][11] ),
    .Q_N(_09682_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][11] ));
 sg13g2_dfrbp_1 _20376_ (.CLK(net5677),
    .RESET_B(net6187),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][12] ),
    .Q_N(_09683_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][12] ));
 sg13g2_dfrbp_1 _20377_ (.CLK(net5664),
    .RESET_B(net6174),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][13] ),
    .Q_N(_09684_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][13] ));
 sg13g2_dfrbp_1 _20378_ (.CLK(net5655),
    .RESET_B(net6165),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][14] ),
    .Q_N(_09685_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][14] ));
 sg13g2_dfrbp_1 _20379_ (.CLK(net5653),
    .RESET_B(net6163),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][15] ),
    .Q_N(_09686_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][15] ));
 sg13g2_dfrbp_1 _20380_ (.CLK(net5620),
    .RESET_B(net6129),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][16] ),
    .Q_N(_09687_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][16] ));
 sg13g2_dfrbp_1 _20381_ (.CLK(net5610),
    .RESET_B(net6119),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][17] ),
    .Q_N(_09688_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][17] ));
 sg13g2_dfrbp_1 _20382_ (.CLK(net5612),
    .RESET_B(net6121),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[13][18] ),
    .Q_N(_09689_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][18] ));
 sg13g2_dfrbp_1 _20383_ (.CLK(net5602),
    .RESET_B(net6111),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][0] ),
    .Q_N(_09690_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][0] ));
 sg13g2_dfrbp_1 _20384_ (.CLK(net5616),
    .RESET_B(net6125),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][1] ),
    .Q_N(_09691_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][1] ));
 sg13g2_dfrbp_1 _20385_ (.CLK(net5613),
    .RESET_B(net6122),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][2] ),
    .Q_N(_09692_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][2] ));
 sg13g2_dfrbp_1 _20386_ (.CLK(net5630),
    .RESET_B(net6139),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][3] ),
    .Q_N(_09693_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][3] ));
 sg13g2_dfrbp_1 _20387_ (.CLK(net5660),
    .RESET_B(net6170),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][4] ),
    .Q_N(_09694_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][4] ));
 sg13g2_dfrbp_1 _20388_ (.CLK(net5644),
    .RESET_B(net6153),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][5] ),
    .Q_N(_09695_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][5] ));
 sg13g2_dfrbp_1 _20389_ (.CLK(net5647),
    .RESET_B(net6156),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][6] ),
    .Q_N(_09696_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][6] ));
 sg13g2_dfrbp_1 _20390_ (.CLK(net5669),
    .RESET_B(net6179),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][7] ),
    .Q_N(_09697_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][7] ));
 sg13g2_dfrbp_1 _20391_ (.CLK(net5670),
    .RESET_B(net6180),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][8] ),
    .Q_N(_09698_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][8] ));
 sg13g2_dfrbp_1 _20392_ (.CLK(net5669),
    .RESET_B(net6179),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][9] ),
    .Q_N(_09699_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][9] ));
 sg13g2_dfrbp_1 _20393_ (.CLK(net5679),
    .RESET_B(net6189),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][10] ),
    .Q_N(_09700_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][10] ));
 sg13g2_dfrbp_1 _20394_ (.CLK(net5677),
    .RESET_B(net6187),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][11] ),
    .Q_N(_09701_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][11] ));
 sg13g2_dfrbp_1 _20395_ (.CLK(net5667),
    .RESET_B(net6177),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][12] ),
    .Q_N(_09702_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][12] ));
 sg13g2_dfrbp_1 _20396_ (.CLK(net5661),
    .RESET_B(net6171),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][13] ),
    .Q_N(_09703_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][13] ));
 sg13g2_dfrbp_1 _20397_ (.CLK(net5655),
    .RESET_B(net6165),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][14] ),
    .Q_N(_09704_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][14] ));
 sg13g2_dfrbp_1 _20398_ (.CLK(net5653),
    .RESET_B(net6163),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][15] ),
    .Q_N(_09705_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][15] ));
 sg13g2_dfrbp_1 _20399_ (.CLK(net5611),
    .RESET_B(net6120),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][16] ),
    .Q_N(_09706_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][16] ));
 sg13g2_dfrbp_1 _20400_ (.CLK(net5605),
    .RESET_B(net6114),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][17] ),
    .Q_N(_09707_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][17] ));
 sg13g2_dfrbp_1 _20401_ (.CLK(net5588),
    .RESET_B(net6097),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][18] ),
    .Q_N(_09708_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[2][18] ));
 sg13g2_dfrbp_1 _20402_ (.CLK(net5606),
    .RESET_B(net6115),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][0] ),
    .Q_N(_09709_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][0] ));
 sg13g2_dfrbp_1 _20403_ (.CLK(net5620),
    .RESET_B(net6129),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][1] ),
    .Q_N(_09710_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][1] ));
 sg13g2_dfrbp_1 _20404_ (.CLK(net5613),
    .RESET_B(net6122),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][2] ),
    .Q_N(_09711_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][2] ));
 sg13g2_dfrbp_1 _20405_ (.CLK(net5650),
    .RESET_B(net6159),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][3] ),
    .Q_N(_09712_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][3] ));
 sg13g2_dfrbp_1 _20406_ (.CLK(net5658),
    .RESET_B(net6168),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][4] ),
    .Q_N(_09713_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][4] ));
 sg13g2_dfrbp_1 _20407_ (.CLK(net5643),
    .RESET_B(net6152),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][5] ),
    .Q_N(_09714_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][5] ));
 sg13g2_dfrbp_1 _20408_ (.CLK(net5646),
    .RESET_B(net6155),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][6] ),
    .Q_N(_09715_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][6] ));
 sg13g2_dfrbp_1 _20409_ (.CLK(net5673),
    .RESET_B(net6183),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][7] ),
    .Q_N(_09716_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][7] ));
 sg13g2_dfrbp_1 _20410_ (.CLK(net5671),
    .RESET_B(net6181),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][8] ),
    .Q_N(_09717_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][8] ));
 sg13g2_dfrbp_1 _20411_ (.CLK(net5676),
    .RESET_B(net6186),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][9] ),
    .Q_N(_09718_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][9] ));
 sg13g2_dfrbp_1 _20412_ (.CLK(net5675),
    .RESET_B(net6185),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][10] ),
    .Q_N(_09719_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][10] ));
 sg13g2_dfrbp_1 _20413_ (.CLK(net5680),
    .RESET_B(net6190),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][11] ),
    .Q_N(_09720_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][11] ));
 sg13g2_dfrbp_1 _20414_ (.CLK(net5684),
    .RESET_B(net6194),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][12] ),
    .Q_N(_09721_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][12] ));
 sg13g2_dfrbp_1 _20415_ (.CLK(net5661),
    .RESET_B(net6171),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][13] ),
    .Q_N(_09722_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][13] ));
 sg13g2_dfrbp_1 _20416_ (.CLK(net5656),
    .RESET_B(net6166),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][14] ),
    .Q_N(_09723_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][14] ));
 sg13g2_dfrbp_1 _20417_ (.CLK(net5654),
    .RESET_B(net6164),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][15] ),
    .Q_N(_09724_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][15] ));
 sg13g2_dfrbp_1 _20418_ (.CLK(net5621),
    .RESET_B(net6130),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][16] ),
    .Q_N(_09725_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][16] ));
 sg13g2_dfrbp_1 _20419_ (.CLK(net5605),
    .RESET_B(net6114),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][17] ),
    .Q_N(_09726_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][17] ));
 sg13g2_dfrbp_1 _20420_ (.CLK(net5590),
    .RESET_B(net6099),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[7][18] ),
    .Q_N(_09727_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[8][18] ));
 sg13g2_dfrbp_1 _20421_ (.CLK(net5600),
    .RESET_B(net6109),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][0] ),
    .Q_N(_09728_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][0] ));
 sg13g2_dfrbp_1 _20422_ (.CLK(net5617),
    .RESET_B(net6126),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][1] ),
    .Q_N(_09729_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][1] ));
 sg13g2_dfrbp_1 _20423_ (.CLK(net5615),
    .RESET_B(net6124),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][2] ),
    .Q_N(_09730_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][2] ));
 sg13g2_dfrbp_1 _20424_ (.CLK(net5630),
    .RESET_B(net6139),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][3] ),
    .Q_N(_09731_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][3] ));
 sg13g2_dfrbp_1 _20425_ (.CLK(net5660),
    .RESET_B(net6170),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][4] ),
    .Q_N(_09732_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][4] ));
 sg13g2_dfrbp_1 _20426_ (.CLK(net5643),
    .RESET_B(net6152),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][5] ),
    .Q_N(_09733_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][5] ));
 sg13g2_dfrbp_1 _20427_ (.CLK(net5648),
    .RESET_B(net6157),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][6] ),
    .Q_N(_09734_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][6] ));
 sg13g2_dfrbp_1 _20428_ (.CLK(net5668),
    .RESET_B(net6178),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][7] ),
    .Q_N(_09735_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][7] ));
 sg13g2_dfrbp_1 _20429_ (.CLK(net5670),
    .RESET_B(net6180),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][8] ),
    .Q_N(_09736_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][8] ));
 sg13g2_dfrbp_1 _20430_ (.CLK(net5669),
    .RESET_B(net6179),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][9] ),
    .Q_N(_09737_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][9] ));
 sg13g2_dfrbp_1 _20431_ (.CLK(net5667),
    .RESET_B(net6177),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][10] ),
    .Q_N(_09738_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][10] ));
 sg13g2_dfrbp_1 _20432_ (.CLK(net5667),
    .RESET_B(net6177),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][11] ),
    .Q_N(_09739_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][11] ));
 sg13g2_dfrbp_1 _20433_ (.CLK(net5667),
    .RESET_B(net6177),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][12] ),
    .Q_N(_09740_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][12] ));
 sg13g2_dfrbp_1 _20434_ (.CLK(net5661),
    .RESET_B(net6171),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][13] ),
    .Q_N(_09741_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][13] ));
 sg13g2_dfrbp_1 _20435_ (.CLK(net5655),
    .RESET_B(net6165),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][14] ),
    .Q_N(_09742_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][14] ));
 sg13g2_dfrbp_1 _20436_ (.CLK(net5652),
    .RESET_B(net6162),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][15] ),
    .Q_N(_09743_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][15] ));
 sg13g2_dfrbp_1 _20437_ (.CLK(net5620),
    .RESET_B(net6129),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][16] ),
    .Q_N(_09744_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][16] ));
 sg13g2_dfrbp_1 _20438_ (.CLK(net5610),
    .RESET_B(net6119),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][17] ),
    .Q_N(_09745_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][17] ));
 sg13g2_dfrbp_1 _20439_ (.CLK(net5590),
    .RESET_B(net6099),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][18] ),
    .Q_N(_09746_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[1][18] ));
 sg13g2_dfrbp_1 _20440_ (.CLK(net5604),
    .RESET_B(net6113),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][0] ),
    .Q_N(_09747_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][0] ));
 sg13g2_dfrbp_1 _20441_ (.CLK(net5619),
    .RESET_B(net6128),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][1] ),
    .Q_N(_09748_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][1] ));
 sg13g2_dfrbp_1 _20442_ (.CLK(net5619),
    .RESET_B(net6128),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][2] ),
    .Q_N(_09749_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][2] ));
 sg13g2_dfrbp_1 _20443_ (.CLK(net5657),
    .RESET_B(net6161),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][3] ),
    .Q_N(_09750_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][3] ));
 sg13g2_dfrbp_1 _20444_ (.CLK(net5659),
    .RESET_B(net6169),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][4] ),
    .Q_N(_09751_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][4] ));
 sg13g2_dfrbp_1 _20445_ (.CLK(net5668),
    .RESET_B(net6178),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][5] ),
    .Q_N(_09752_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][5] ));
 sg13g2_dfrbp_1 _20446_ (.CLK(net5646),
    .RESET_B(net6155),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][6] ),
    .Q_N(_09753_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][6] ));
 sg13g2_dfrbp_1 _20447_ (.CLK(net5672),
    .RESET_B(net6182),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][7] ),
    .Q_N(_09754_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][7] ));
 sg13g2_dfrbp_1 _20448_ (.CLK(net5670),
    .RESET_B(net6180),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][8] ),
    .Q_N(_09755_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][8] ));
 sg13g2_dfrbp_1 _20449_ (.CLK(net5673),
    .RESET_B(net6183),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][9] ),
    .Q_N(_09756_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][9] ));
 sg13g2_dfrbp_1 _20450_ (.CLK(net5675),
    .RESET_B(net6185),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][10] ),
    .Q_N(_09757_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][10] ));
 sg13g2_dfrbp_1 _20451_ (.CLK(net5678),
    .RESET_B(net6188),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][11] ),
    .Q_N(_09758_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][11] ));
 sg13g2_dfrbp_1 _20452_ (.CLK(net5677),
    .RESET_B(net6187),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][12] ),
    .Q_N(_09759_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][12] ));
 sg13g2_dfrbp_1 _20453_ (.CLK(net5664),
    .RESET_B(net6174),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][13] ),
    .Q_N(_09760_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][13] ));
 sg13g2_dfrbp_1 _20454_ (.CLK(net5655),
    .RESET_B(net6165),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][14] ),
    .Q_N(_09761_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][14] ));
 sg13g2_dfrbp_1 _20455_ (.CLK(net5653),
    .RESET_B(net6163),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][15] ),
    .Q_N(_09762_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][15] ));
 sg13g2_dfrbp_1 _20456_ (.CLK(net5621),
    .RESET_B(net6130),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][16] ),
    .Q_N(_09763_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][16] ));
 sg13g2_dfrbp_1 _20457_ (.CLK(net5611),
    .RESET_B(net6120),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][17] ),
    .Q_N(_09764_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][17] ));
 sg13g2_dfrbp_1 _20458_ (.CLK(net5612),
    .RESET_B(net6121),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[14][18] ),
    .Q_N(_09765_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[15][18] ));
 sg13g2_dfrbp_1 _20459_ (.CLK(net5600),
    .RESET_B(net6109),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.u_mux_shift.sum_res ),
    .Q_N(_00289_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][0] ));
 sg13g2_dfrbp_1 _20460_ (.CLK(net5613),
    .RESET_B(net6122),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .Q_N(_00300_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][1] ));
 sg13g2_dfrbp_1 _20461_ (.CLK(net5615),
    .RESET_B(net6124),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .Q_N(_00307_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][2] ));
 sg13g2_dfrbp_1 _20462_ (.CLK(net5630),
    .RESET_B(net6139),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .Q_N(_00314_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][3] ));
 sg13g2_dfrbp_1 _20463_ (.CLK(net5660),
    .RESET_B(net6170),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .Q_N(_00323_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][4] ));
 sg13g2_dfrbp_1 _20464_ (.CLK(net5643),
    .RESET_B(net6152),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .Q_N(_00332_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][5] ));
 sg13g2_dfrbp_1 _20465_ (.CLK(net5645),
    .RESET_B(net6154),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .Q_N(_00339_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][6] ));
 sg13g2_dfrbp_1 _20466_ (.CLK(net5668),
    .RESET_B(net6178),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .Q_N(_00346_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][7] ));
 sg13g2_dfrbp_1 _20467_ (.CLK(net5668),
    .RESET_B(net6178),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .Q_N(_00355_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][8] ));
 sg13g2_dfrbp_1 _20468_ (.CLK(net5669),
    .RESET_B(net6179),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .Q_N(_00364_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][9] ));
 sg13g2_dfrbp_1 _20469_ (.CLK(net5663),
    .RESET_B(net6173),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .Q_N(_00371_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][10] ));
 sg13g2_dfrbp_1 _20470_ (.CLK(net5667),
    .RESET_B(net6177),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .Q_N(_00378_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][11] ));
 sg13g2_dfrbp_1 _20471_ (.CLK(net5666),
    .RESET_B(net6176),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .Q_N(_00387_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][12] ));
 sg13g2_dfrbp_1 _20472_ (.CLK(net5661),
    .RESET_B(net6171),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .Q_N(_00396_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][13] ));
 sg13g2_dfrbp_1 _20473_ (.CLK(net5655),
    .RESET_B(net6165),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .Q_N(_00403_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][14] ));
 sg13g2_dfrbp_1 _20474_ (.CLK(net5651),
    .RESET_B(net6160),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .Q_N(_00410_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][15] ));
 sg13g2_dfrbp_1 _20475_ (.CLK(net5617),
    .RESET_B(net6126),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .Q_N(_00419_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][16] ));
 sg13g2_dfrbp_1 _20476_ (.CLK(net5610),
    .RESET_B(net6119),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .Q_N(_00426_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][17] ));
 sg13g2_dfrbp_1 _20477_ (.CLK(net5588),
    .RESET_B(net6097),
    .D(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .Q_N(_00433_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[0][18] ));
 sg13g2_dfrbp_1 _20478_ (.CLK(net5604),
    .RESET_B(net6113),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][0] ),
    .Q_N(_09766_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][0] ));
 sg13g2_dfrbp_1 _20479_ (.CLK(net5620),
    .RESET_B(net6129),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][1] ),
    .Q_N(_09767_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][1] ));
 sg13g2_dfrbp_1 _20480_ (.CLK(net5613),
    .RESET_B(net6122),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][2] ),
    .Q_N(_09768_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][2] ));
 sg13g2_dfrbp_1 _20481_ (.CLK(net5650),
    .RESET_B(net6159),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][3] ),
    .Q_N(_09769_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][3] ));
 sg13g2_dfrbp_1 _20482_ (.CLK(net5659),
    .RESET_B(net6169),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][4] ),
    .Q_N(_09770_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][4] ));
 sg13g2_dfrbp_1 _20483_ (.CLK(net5668),
    .RESET_B(net6178),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][5] ),
    .Q_N(_09771_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][5] ));
 sg13g2_dfrbp_1 _20484_ (.CLK(net5646),
    .RESET_B(net6155),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][6] ),
    .Q_N(_09772_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][6] ));
 sg13g2_dfrbp_1 _20485_ (.CLK(net5673),
    .RESET_B(net6183),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][7] ),
    .Q_N(_09773_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][7] ));
 sg13g2_dfrbp_1 _20486_ (.CLK(net5671),
    .RESET_B(net6181),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][8] ),
    .Q_N(_09774_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][8] ));
 sg13g2_dfrbp_1 _20487_ (.CLK(net5680),
    .RESET_B(net6190),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][9] ),
    .Q_N(_09775_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][9] ));
 sg13g2_dfrbp_1 _20488_ (.CLK(net5680),
    .RESET_B(net6190),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][10] ),
    .Q_N(_09776_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][10] ));
 sg13g2_dfrbp_1 _20489_ (.CLK(net5681),
    .RESET_B(net6191),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][11] ),
    .Q_N(_09777_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][11] ));
 sg13g2_dfrbp_1 _20490_ (.CLK(net5684),
    .RESET_B(net6194),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][12] ),
    .Q_N(_09778_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][12] ));
 sg13g2_dfrbp_1 _20491_ (.CLK(net5664),
    .RESET_B(net6174),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][13] ),
    .Q_N(_09779_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][13] ));
 sg13g2_dfrbp_1 _20492_ (.CLK(net5656),
    .RESET_B(net6166),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][14] ),
    .Q_N(_09780_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][14] ));
 sg13g2_dfrbp_1 _20493_ (.CLK(net5654),
    .RESET_B(net6164),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][15] ),
    .Q_N(_09781_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][15] ));
 sg13g2_dfrbp_1 _20494_ (.CLK(net5621),
    .RESET_B(net6129),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][16] ),
    .Q_N(_09782_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][16] ));
 sg13g2_dfrbp_1 _20495_ (.CLK(net5610),
    .RESET_B(net6119),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][17] ),
    .Q_N(_09783_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][17] ));
 sg13g2_dfrbp_1 _20496_ (.CLK(net5612),
    .RESET_B(net6121),
    .D(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[9][18] ),
    .Q_N(_06255_),
    .Q(\u_supermic_top_module.u_delay_module.delay_line_gen[7].u_delay_line.buffer[10][18] ));
 sg13g2_dfrbp_1 _20497_ (.CLK(_01795_),
    .RESET_B(net5777),
    .D(net2),
    .Q_N(_06254_),
    .Q(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[1].u_ddr_to_sdr_dual.ddr_data_falling ));
 sg13g2_dfrbp_1 _20498_ (.CLK(_01796_),
    .RESET_B(net5885),
    .D(net3),
    .Q_N(_06253_),
    .Q(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[2].u_ddr_to_sdr_dual.ddr_data_falling ));
 sg13g2_dfrbp_1 _20499_ (.CLK(_01797_),
    .RESET_B(net6133),
    .D(net4),
    .Q_N(_09784_),
    .Q(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[3].u_ddr_to_sdr_dual.ddr_data_falling ));
 sg13g2_dfrbp_1 _20500_ (.CLK(net5185),
    .RESET_B(net5695),
    .D(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[0].u_ddr_to_sdr_dual.ddr_data_falling ),
    .Q_N(_09785_),
    .Q(\u_supermic_top_module.cic_inst[4].u_cic.i_data ));
 sg13g2_dfrbp_1 _20501_ (.CLK(net5186),
    .RESET_B(net5696),
    .D(net1),
    .Q_N(_09786_),
    .Q(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[0].u_ddr_to_sdr_dual.ddr_data_rising ));
 sg13g2_dfrbp_1 _20502_ (.CLK(net5192),
    .RESET_B(net5702),
    .D(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[0].u_ddr_to_sdr_dual.ddr_data_rising ),
    .Q_N(_09787_),
    .Q(\u_supermic_top_module.cic_inst[0].u_cic.i_data ));
 sg13g2_dfrbp_1 _20503_ (.CLK(net5274),
    .RESET_B(net5784),
    .D(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[1].u_ddr_to_sdr_dual.ddr_data_falling ),
    .Q_N(_09788_),
    .Q(\u_supermic_top_module.cic_inst[5].u_cic.i_data ));
 sg13g2_dfrbp_1 _20504_ (.CLK(net5264),
    .RESET_B(net5774),
    .D(net2),
    .Q_N(_09789_),
    .Q(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[1].u_ddr_to_sdr_dual.ddr_data_rising ));
 sg13g2_dfrbp_1 _20505_ (.CLK(net5264),
    .RESET_B(net5774),
    .D(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[1].u_ddr_to_sdr_dual.ddr_data_rising ),
    .Q_N(_09790_),
    .Q(\u_supermic_top_module.cic_inst[1].u_cic.i_data ));
 sg13g2_dfrbp_1 _20506_ (.CLK(net5376),
    .RESET_B(net5885),
    .D(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[2].u_ddr_to_sdr_dual.ddr_data_falling ),
    .Q_N(_09791_),
    .Q(\u_supermic_top_module.cic_inst[6].u_cic.i_data ));
 sg13g2_dfrbp_1 _20507_ (.CLK(net5422),
    .RESET_B(net5931),
    .D(net3),
    .Q_N(_09792_),
    .Q(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[2].u_ddr_to_sdr_dual.ddr_data_rising ));
 sg13g2_dfrbp_1 _20508_ (.CLK(net5422),
    .RESET_B(net5931),
    .D(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[2].u_ddr_to_sdr_dual.ddr_data_rising ),
    .Q_N(_09793_),
    .Q(\u_supermic_top_module.cic_inst[2].u_cic.i_data ));
 sg13g2_dfrbp_1 _20509_ (.CLK(net5624),
    .RESET_B(net6133),
    .D(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[3].u_ddr_to_sdr_dual.ddr_data_falling ),
    .Q_N(_09794_),
    .Q(\u_supermic_top_module.cic_inst[7].u_cic.i_data ));
 sg13g2_dfrbp_1 _20510_ (.CLK(net5491),
    .RESET_B(net6000),
    .D(net4),
    .Q_N(_09795_),
    .Q(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[3].u_ddr_to_sdr_dual.ddr_data_rising ));
 sg13g2_dfrbp_1 _20511_ (.CLK(net5563),
    .RESET_B(net6072),
    .D(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[3].u_ddr_to_sdr_dual.ddr_data_rising ),
    .Q_N(_06252_),
    .Q(\u_supermic_top_module.cic_inst[3].u_cic.i_data ));
 sg13g2_dfrbp_1 _20512_ (.CLK(_01798_),
    .RESET_B(net5695),
    .D(net1),
    .Q_N(_06251_),
    .Q(\u_supermic_top_module.u_top_ddr_to_sdr.ddr_to_sdr_dual_inst[0].u_ddr_to_sdr_dual.ddr_data_falling ));
 sg13g2_tiehi _16815__20 (.L_HI(net20));
 sg13g2_tiehi _16880__21 (.L_HI(net21));
 sg13g2_tiehi _16945__22 (.L_HI(net22));
 sg13g2_tiehi _17010__23 (.L_HI(net23));
 sg13g2_tiehi _19006__24 (.L_HI(net24));
 sg13g2_tiehi _19005__25 (.L_HI(net25));
 sg13g2_tiehi _19004__26 (.L_HI(net26));
 sg13g2_tiehi _19003__27 (.L_HI(net27));
 sg13g2_tiehi _19002__28 (.L_HI(net28));
 sg13g2_tiehi _19001__29 (.L_HI(net29));
 sg13g2_tiehi _19000__30 (.L_HI(net30));
 sg13g2_tiehi _18999__31 (.L_HI(net31));
 sg13g2_tiehi _18998__32 (.L_HI(net32));
 sg13g2_tiehi _18997__33 (.L_HI(net33));
 sg13g2_tiehi _18996__34 (.L_HI(net34));
 sg13g2_tiehi _18995__35 (.L_HI(net35));
 sg13g2_tiehi _18994__36 (.L_HI(net36));
 sg13g2_tiehi _18993__37 (.L_HI(net37));
 sg13g2_tiehi _18992__38 (.L_HI(net38));
 sg13g2_tiehi _18991__39 (.L_HI(net39));
 sg13g2_tiehi _18990__40 (.L_HI(net40));
 sg13g2_tiehi _18989__41 (.L_HI(net41));
 sg13g2_tiehi _18988__42 (.L_HI(net42));
 sg13g2_tiehi _18987__43 (.L_HI(net43));
 sg13g2_tiehi _18948__44 (.L_HI(net44));
 sg13g2_tiehi _18947__45 (.L_HI(net45));
 sg13g2_tiehi _18946__46 (.L_HI(net46));
 sg13g2_tiehi _18945__47 (.L_HI(net47));
 sg13g2_tiehi _18944__48 (.L_HI(net48));
 sg13g2_tiehi _18943__49 (.L_HI(net49));
 sg13g2_tiehi _18942__50 (.L_HI(net50));
 sg13g2_tiehi _18941__51 (.L_HI(net51));
 sg13g2_tiehi _18940__52 (.L_HI(net52));
 sg13g2_tiehi _17075__53 (.L_HI(net53));
 sg13g2_tiehi _18939__54 (.L_HI(net54));
 sg13g2_tiehi _18938__55 (.L_HI(net55));
 sg13g2_tiehi _18937__56 (.L_HI(net56));
 sg13g2_tiehi _18936__57 (.L_HI(net57));
 sg13g2_tiehi _18935__58 (.L_HI(net58));
 sg13g2_tiehi _18934__59 (.L_HI(net59));
 sg13g2_tiehi _18933__60 (.L_HI(net60));
 sg13g2_tiehi _18932__61 (.L_HI(net61));
 sg13g2_tiehi _18931__62 (.L_HI(net62));
 sg13g2_tiehi _18930__63 (.L_HI(net63));
 sg13g2_tiehi _18796__64 (.L_HI(net64));
 sg13g2_tiehi _18795__65 (.L_HI(net65));
 sg13g2_tiehi _18794__66 (.L_HI(net66));
 sg13g2_tiehi _18793__67 (.L_HI(net67));
 sg13g2_tiehi _18792__68 (.L_HI(net68));
 sg13g2_tiehi _18791__69 (.L_HI(net69));
 sg13g2_tiehi _18790__70 (.L_HI(net70));
 sg13g2_tiehi _18789__71 (.L_HI(net71));
 sg13g2_tiehi _18788__72 (.L_HI(net72));
 sg13g2_tiehi _18787__73 (.L_HI(net73));
 sg13g2_tiehi _18786__74 (.L_HI(net74));
 sg13g2_tiehi _18785__75 (.L_HI(net75));
 sg13g2_tiehi _18784__76 (.L_HI(net76));
 sg13g2_tiehi _18783__77 (.L_HI(net77));
 sg13g2_tiehi _18782__78 (.L_HI(net78));
 sg13g2_tiehi _18781__79 (.L_HI(net79));
 sg13g2_tiehi _18780__80 (.L_HI(net80));
 sg13g2_tiehi _18779__81 (.L_HI(net81));
 sg13g2_tiehi _18778__82 (.L_HI(net82));
 sg13g2_tiehi _18739__83 (.L_HI(net83));
 sg13g2_tiehi _18738__84 (.L_HI(net84));
 sg13g2_tiehi _18737__85 (.L_HI(net85));
 sg13g2_tiehi _18736__86 (.L_HI(net86));
 sg13g2_tiehi _17140__87 (.L_HI(net87));
 sg13g2_tiehi _18735__88 (.L_HI(net88));
 sg13g2_tiehi _18734__89 (.L_HI(net89));
 sg13g2_tiehi _18733__90 (.L_HI(net90));
 sg13g2_tiehi _18732__91 (.L_HI(net91));
 sg13g2_tiehi _18731__92 (.L_HI(net92));
 sg13g2_tiehi _18730__93 (.L_HI(net93));
 sg13g2_tiehi _18729__94 (.L_HI(net94));
 sg13g2_tiehi _18728__95 (.L_HI(net95));
 sg13g2_tiehi _18727__96 (.L_HI(net96));
 sg13g2_tiehi _18726__97 (.L_HI(net97));
 sg13g2_tiehi _18725__98 (.L_HI(net98));
 sg13g2_tiehi _18724__99 (.L_HI(net99));
 sg13g2_tiehi _18723__100 (.L_HI(net100));
 sg13g2_tiehi _18722__101 (.L_HI(net101));
 sg13g2_tiehi _18721__102 (.L_HI(net102));
 sg13g2_tiehi _18587__103 (.L_HI(net103));
 sg13g2_tiehi _18586__104 (.L_HI(net104));
 sg13g2_tiehi _18585__105 (.L_HI(net105));
 sg13g2_tiehi _18584__106 (.L_HI(net106));
 sg13g2_tiehi _18583__107 (.L_HI(net107));
 sg13g2_tiehi _18582__108 (.L_HI(net108));
 sg13g2_tiehi _18581__109 (.L_HI(net109));
 sg13g2_tiehi _18580__110 (.L_HI(net110));
 sg13g2_tiehi _18579__111 (.L_HI(net111));
 sg13g2_tiehi _18578__112 (.L_HI(net112));
 sg13g2_tiehi _18577__113 (.L_HI(net113));
 sg13g2_tiehi _18576__114 (.L_HI(net114));
 sg13g2_tiehi _18575__115 (.L_HI(net115));
 sg13g2_tiehi _18574__116 (.L_HI(net116));
 sg13g2_tiehi _18573__117 (.L_HI(net117));
 sg13g2_tiehi _18572__118 (.L_HI(net118));
 sg13g2_tiehi _18571__119 (.L_HI(net119));
 sg13g2_tiehi _18570__120 (.L_HI(net120));
 sg13g2_tiehi _17205__121 (.L_HI(net121));
 sg13g2_tiehi _18569__122 (.L_HI(net122));
 sg13g2_tiehi _18530__123 (.L_HI(net123));
 sg13g2_tiehi _18529__124 (.L_HI(net124));
 sg13g2_tiehi _18528__125 (.L_HI(net125));
 sg13g2_tiehi _18527__126 (.L_HI(net126));
 sg13g2_tiehi _18526__127 (.L_HI(net127));
 sg13g2_tiehi _18525__128 (.L_HI(net128));
 sg13g2_tiehi _18524__129 (.L_HI(net129));
 sg13g2_tiehi _18523__130 (.L_HI(net130));
 sg13g2_tiehi _18522__131 (.L_HI(net131));
 sg13g2_tiehi _18521__132 (.L_HI(net132));
 sg13g2_tiehi _18520__133 (.L_HI(net133));
 sg13g2_tiehi _18519__134 (.L_HI(net134));
 sg13g2_tiehi _18518__135 (.L_HI(net135));
 sg13g2_tiehi _18517__136 (.L_HI(net136));
 sg13g2_tiehi _18516__137 (.L_HI(net137));
 sg13g2_tiehi _18515__138 (.L_HI(net138));
 sg13g2_tiehi _18514__139 (.L_HI(net139));
 sg13g2_tiehi _18513__140 (.L_HI(net140));
 sg13g2_tiehi _18512__141 (.L_HI(net141));
 sg13g2_tiehi _18378__142 (.L_HI(net142));
 sg13g2_tiehi _18377__143 (.L_HI(net143));
 sg13g2_tiehi _18376__144 (.L_HI(net144));
 sg13g2_tiehi _18375__145 (.L_HI(net145));
 sg13g2_tiehi _18374__146 (.L_HI(net146));
 sg13g2_tiehi _18373__147 (.L_HI(net147));
 sg13g2_tiehi _18372__148 (.L_HI(net148));
 sg13g2_tiehi _18371__149 (.L_HI(net149));
 sg13g2_tiehi _18370__150 (.L_HI(net150));
 sg13g2_tiehi _18369__151 (.L_HI(net151));
 sg13g2_tiehi _18368__152 (.L_HI(net152));
 sg13g2_tiehi _18367__153 (.L_HI(net153));
 sg13g2_tiehi _18366__154 (.L_HI(net154));
 sg13g2_tiehi _18365__155 (.L_HI(net155));
 sg13g2_tiehi _18364__156 (.L_HI(net156));
 sg13g2_tiehi _18363__157 (.L_HI(net157));
 sg13g2_tiehi _18362__158 (.L_HI(net158));
 sg13g2_tiehi _18361__159 (.L_HI(net159));
 sg13g2_tiehi _18360__160 (.L_HI(net160));
 sg13g2_tiehi _18321__161 (.L_HI(net161));
 sg13g2_tiehi _18320__162 (.L_HI(net162));
 sg13g2_tiehi _18319__163 (.L_HI(net163));
 sg13g2_tiehi _18318__164 (.L_HI(net164));
 sg13g2_tiehi _18317__165 (.L_HI(net165));
 sg13g2_tiehi _18316__166 (.L_HI(net166));
 sg13g2_tiehi _18315__167 (.L_HI(net167));
 sg13g2_tiehi _18314__168 (.L_HI(net168));
 sg13g2_tiehi _18313__169 (.L_HI(net169));
 sg13g2_tiehi _18312__170 (.L_HI(net170));
 sg13g2_tiehi _18311__171 (.L_HI(net171));
 sg13g2_tiehi _18310__172 (.L_HI(net172));
 sg13g2_tiehi _18309__173 (.L_HI(net173));
 sg13g2_tiehi _18308__174 (.L_HI(net174));
 sg13g2_tiehi _18307__175 (.L_HI(net175));
 sg13g2_tiehi _18306__176 (.L_HI(net176));
 sg13g2_tiehi _18305__177 (.L_HI(net177));
 sg13g2_tiehi _18304__178 (.L_HI(net178));
 sg13g2_tiehi _18303__179 (.L_HI(net179));
 sg13g2_tiehi _18169__180 (.L_HI(net180));
 sg13g2_tiehi _18168__181 (.L_HI(net181));
 sg13g2_tiehi _18167__182 (.L_HI(net182));
 sg13g2_tiehi _18166__183 (.L_HI(net183));
 sg13g2_tiehi _18165__184 (.L_HI(net184));
 sg13g2_tiehi _17430__185 (.L_HI(net185));
 sg13g2_tiehi _17431__186 (.L_HI(net186));
 sg13g2_tiehi _17432__187 (.L_HI(net187));
 sg13g2_tiehi _17433__188 (.L_HI(net188));
 sg13g2_tiehi _17434__189 (.L_HI(net189));
 sg13g2_tiehi _17435__190 (.L_HI(net190));
 sg13g2_tiehi _17436__191 (.L_HI(net191));
 sg13g2_tiehi _17437__192 (.L_HI(net192));
 sg13g2_tiehi _17438__193 (.L_HI(net193));
 sg13g2_tiehi _17439__194 (.L_HI(net194));
 sg13g2_tiehi _17440__195 (.L_HI(net195));
 sg13g2_tiehi _17441__196 (.L_HI(net196));
 sg13g2_tiehi _17442__197 (.L_HI(net197));
 sg13g2_tiehi _17443__198 (.L_HI(net198));
 sg13g2_tiehi _17444__199 (.L_HI(net199));
 sg13g2_tiehi _17445__200 (.L_HI(net200));
 sg13g2_tiehi _17446__201 (.L_HI(net201));
 sg13g2_tiehi _17447__202 (.L_HI(net202));
 sg13g2_tiehi _17448__203 (.L_HI(net203));
 sg13g2_tiehi _17449__204 (.L_HI(net204));
 sg13g2_tiehi _17450__205 (.L_HI(net205));
 sg13g2_tiehi _17451__206 (.L_HI(net206));
 sg13g2_tiehi _17452__207 (.L_HI(net207));
 sg13g2_tiehi _17453__208 (.L_HI(net208));
 sg13g2_tiehi _17454__209 (.L_HI(net209));
 sg13g2_tiehi _17455__210 (.L_HI(net210));
 sg13g2_tiehi _17456__211 (.L_HI(net211));
 sg13g2_tiehi _17457__212 (.L_HI(net212));
 sg13g2_tiehi _17458__213 (.L_HI(net213));
 sg13g2_tiehi _17459__214 (.L_HI(net214));
 sg13g2_tiehi _17460__215 (.L_HI(net215));
 sg13g2_tiehi _17461__216 (.L_HI(net216));
 sg13g2_tiehi _17462__217 (.L_HI(net217));
 sg13g2_tiehi _17463__218 (.L_HI(net218));
 sg13g2_tiehi _17464__219 (.L_HI(net219));
 sg13g2_tiehi _17465__220 (.L_HI(net220));
 sg13g2_tiehi _18164__221 (.L_HI(net221));
 sg13g2_tiehi _18163__222 (.L_HI(net222));
 sg13g2_tiehi _18162__223 (.L_HI(net223));
 sg13g2_tiehi _18161__224 (.L_HI(net224));
 sg13g2_tiehi _18160__225 (.L_HI(net225));
 sg13g2_tiehi _18159__226 (.L_HI(net226));
 sg13g2_tiehi _18158__227 (.L_HI(net227));
 sg13g2_tiehi _18157__228 (.L_HI(net228));
 sg13g2_tiehi _18156__229 (.L_HI(net229));
 sg13g2_tiehi _18155__230 (.L_HI(net230));
 sg13g2_tiehi _18154__231 (.L_HI(net231));
 sg13g2_tiehi _18153__232 (.L_HI(net232));
 sg13g2_tiehi _18152__233 (.L_HI(net233));
 sg13g2_tiehi _18151__234 (.L_HI(net234));
 sg13g2_tiehi _18112__235 (.L_HI(net235));
 sg13g2_tiehi _18111__236 (.L_HI(net236));
 sg13g2_tiehi _18110__237 (.L_HI(net237));
 sg13g2_tiehi _18109__238 (.L_HI(net238));
 sg13g2_tiehi _18108__239 (.L_HI(net239));
 sg13g2_tiehi _17466__240 (.L_HI(net240));
 sg13g2_tiehi _17486__241 (.L_HI(net241));
 sg13g2_tiehi _17487__242 (.L_HI(net242));
 sg13g2_tiehi _17488__243 (.L_HI(net243));
 sg13g2_tiehi _17489__244 (.L_HI(net244));
 sg13g2_tiehi _17490__245 (.L_HI(net245));
 sg13g2_tiehi _17491__246 (.L_HI(net246));
 sg13g2_tiehi _17492__247 (.L_HI(net247));
 sg13g2_tiehi _17493__248 (.L_HI(net248));
 sg13g2_tiehi _17494__249 (.L_HI(net249));
 sg13g2_tiehi _17495__250 (.L_HI(net250));
 sg13g2_tiehi _17496__251 (.L_HI(net251));
 sg13g2_tiehi _17497__252 (.L_HI(net252));
 sg13g2_tiehi _17498__253 (.L_HI(net253));
 sg13g2_tiehi _17499__254 (.L_HI(net254));
 sg13g2_tiehi _17500__255 (.L_HI(net255));
 sg13g2_tiehi _17501__256 (.L_HI(net256));
 sg13g2_tiehi _17502__257 (.L_HI(net257));
 sg13g2_tiehi _17503__258 (.L_HI(net258));
 sg13g2_tiehi _17504__259 (.L_HI(net259));
 sg13g2_tiehi _17505__260 (.L_HI(net260));
 sg13g2_tiehi _17506__261 (.L_HI(net261));
 sg13g2_tiehi _17507__262 (.L_HI(net262));
 sg13g2_tiehi _17508__263 (.L_HI(net263));
 sg13g2_tiehi _17509__264 (.L_HI(net264));
 sg13g2_tiehi _17510__265 (.L_HI(net265));
 sg13g2_tiehi _17511__266 (.L_HI(net266));
 sg13g2_tiehi _17512__267 (.L_HI(net267));
 sg13g2_tiehi _17513__268 (.L_HI(net268));
 sg13g2_tiehi _17514__269 (.L_HI(net269));
 sg13g2_tiehi _17515__270 (.L_HI(net270));
 sg13g2_tiehi _17516__271 (.L_HI(net271));
 sg13g2_tiehi _17517__272 (.L_HI(net272));
 sg13g2_tiehi _17518__273 (.L_HI(net273));
 sg13g2_tiehi _17519__274 (.L_HI(net274));
 sg13g2_tiehi _17520__275 (.L_HI(net275));
 sg13g2_tiehi _17521__276 (.L_HI(net276));
 sg13g2_tiehi _17522__277 (.L_HI(net277));
 sg13g2_tiehi _18107__278 (.L_HI(net278));
 sg13g2_tiehi _18106__279 (.L_HI(net279));
 sg13g2_tiehi _18105__280 (.L_HI(net280));
 sg13g2_tiehi _18104__281 (.L_HI(net281));
 sg13g2_tiehi _18103__282 (.L_HI(net282));
 sg13g2_tiehi _18102__283 (.L_HI(net283));
 sg13g2_tiehi _18101__284 (.L_HI(net284));
 sg13g2_tiehi _18100__285 (.L_HI(net285));
 sg13g2_tiehi _18099__286 (.L_HI(net286));
 sg13g2_tiehi _18098__287 (.L_HI(net287));
 sg13g2_tiehi _18097__288 (.L_HI(net288));
 sg13g2_tiehi _18096__289 (.L_HI(net289));
 sg13g2_tiehi _18095__290 (.L_HI(net290));
 sg13g2_tiehi _18094__291 (.L_HI(net291));
 sg13g2_tiehi _17960__292 (.L_HI(net292));
 sg13g2_tiehi _17959__293 (.L_HI(net293));
 sg13g2_tiehi _17958__294 (.L_HI(net294));
 sg13g2_tiehi _17957__295 (.L_HI(net295));
 sg13g2_tiehi _17956__296 (.L_HI(net296));
 sg13g2_tiehi _17523__297 (.L_HI(net297));
 sg13g2_tiehi _17543__298 (.L_HI(net298));
 sg13g2_tiehi _17639__299 (.L_HI(net299));
 sg13g2_tiehi _17640__300 (.L_HI(net300));
 sg13g2_tiehi _17641__301 (.L_HI(net301));
 sg13g2_tiehi _17642__302 (.L_HI(net302));
 sg13g2_tiehi _17643__303 (.L_HI(net303));
 sg13g2_tiehi _17644__304 (.L_HI(net304));
 sg13g2_tiehi _17645__305 (.L_HI(net305));
 sg13g2_tiehi _17646__306 (.L_HI(net306));
 sg13g2_tiehi _17647__307 (.L_HI(net307));
 sg13g2_tiehi _17648__308 (.L_HI(net308));
 sg13g2_tiehi _17649__309 (.L_HI(net309));
 sg13g2_tiehi _17650__310 (.L_HI(net310));
 sg13g2_tiehi _17651__311 (.L_HI(net311));
 sg13g2_tiehi _17652__312 (.L_HI(net312));
 sg13g2_tiehi _17653__313 (.L_HI(net313));
 sg13g2_tiehi _17654__314 (.L_HI(net314));
 sg13g2_tiehi _17655__315 (.L_HI(net315));
 sg13g2_tiehi _17656__316 (.L_HI(net316));
 sg13g2_tiehi _17657__317 (.L_HI(net317));
 sg13g2_tiehi _17658__318 (.L_HI(net318));
 sg13g2_tiehi _17659__319 (.L_HI(net319));
 sg13g2_tiehi _17660__320 (.L_HI(net320));
 sg13g2_tiehi _17661__321 (.L_HI(net321));
 sg13g2_tiehi _17662__322 (.L_HI(net322));
 sg13g2_tiehi _17663__323 (.L_HI(net323));
 sg13g2_tiehi _17664__324 (.L_HI(net324));
 sg13g2_tiehi _17665__325 (.L_HI(net325));
 sg13g2_tiehi _17666__326 (.L_HI(net326));
 sg13g2_tiehi _17667__327 (.L_HI(net327));
 sg13g2_tiehi _17668__328 (.L_HI(net328));
 sg13g2_tiehi _17669__329 (.L_HI(net329));
 sg13g2_tiehi _17670__330 (.L_HI(net330));
 sg13g2_tiehi _17671__331 (.L_HI(net331));
 sg13g2_tiehi _17672__332 (.L_HI(net332));
 sg13g2_tiehi _17673__333 (.L_HI(net333));
 sg13g2_tiehi _17674__334 (.L_HI(net334));
 sg13g2_tiehi _17955__335 (.L_HI(net335));
 sg13g2_tiehi _17954__336 (.L_HI(net336));
 sg13g2_tiehi _17953__337 (.L_HI(net337));
 sg13g2_tiehi _17952__338 (.L_HI(net338));
 sg13g2_tiehi _17951__339 (.L_HI(net339));
 sg13g2_tiehi _17950__340 (.L_HI(net340));
 sg13g2_tiehi _17949__341 (.L_HI(net341));
 sg13g2_tiehi _17948__342 (.L_HI(net342));
 sg13g2_tiehi _17947__343 (.L_HI(net343));
 sg13g2_tiehi _17946__344 (.L_HI(net344));
 sg13g2_tiehi _17945__345 (.L_HI(net345));
 sg13g2_tiehi _17944__346 (.L_HI(net346));
 sg13g2_tiehi _17943__347 (.L_HI(net347));
 sg13g2_tiehi _17942__348 (.L_HI(net348));
 sg13g2_tiehi _17903__349 (.L_HI(net349));
 sg13g2_tiehi _17902__350 (.L_HI(net350));
 sg13g2_tiehi _17901__351 (.L_HI(net351));
 sg13g2_tiehi _17900__352 (.L_HI(net352));
 sg13g2_tiehi _17899__353 (.L_HI(net353));
 sg13g2_tiehi _17675__354 (.L_HI(net354));
 sg13g2_tiehi _17695__355 (.L_HI(net355));
 sg13g2_tiehi _17696__356 (.L_HI(net356));
 sg13g2_tiehi _17697__357 (.L_HI(net357));
 sg13g2_tiehi _17698__358 (.L_HI(net358));
 sg13g2_tiehi _17699__359 (.L_HI(net359));
 sg13g2_tiehi _17700__360 (.L_HI(net360));
 sg13g2_tiehi _17701__361 (.L_HI(net361));
 sg13g2_tiehi _17702__362 (.L_HI(net362));
 sg13g2_tiehi _17703__363 (.L_HI(net363));
 sg13g2_tiehi _17704__364 (.L_HI(net364));
 sg13g2_tiehi _17705__365 (.L_HI(net365));
 sg13g2_tiehi _17706__366 (.L_HI(net366));
 sg13g2_tiehi _17707__367 (.L_HI(net367));
 sg13g2_tiehi _17708__368 (.L_HI(net368));
 sg13g2_tiehi _17709__369 (.L_HI(net369));
 sg13g2_tiehi _17710__370 (.L_HI(net370));
 sg13g2_tiehi _17711__371 (.L_HI(net371));
 sg13g2_tiehi _17712__372 (.L_HI(net372));
 sg13g2_tiehi _17713__373 (.L_HI(net373));
 sg13g2_tiehi _17714__374 (.L_HI(net374));
 sg13g2_tiehi _17715__375 (.L_HI(net375));
 sg13g2_tiehi _17716__376 (.L_HI(net376));
 sg13g2_tiehi _17717__377 (.L_HI(net377));
 sg13g2_tiehi _17718__378 (.L_HI(net378));
 sg13g2_tiehi _17719__379 (.L_HI(net379));
 sg13g2_tiehi _17720__380 (.L_HI(net380));
 sg13g2_tiehi _17721__381 (.L_HI(net381));
 sg13g2_tiehi _17722__382 (.L_HI(net382));
 sg13g2_tiehi _17723__383 (.L_HI(net383));
 sg13g2_tiehi _17724__384 (.L_HI(net384));
 sg13g2_tiehi _17725__385 (.L_HI(net385));
 sg13g2_tiehi _17726__386 (.L_HI(net386));
 sg13g2_tiehi _17727__387 (.L_HI(net387));
 sg13g2_tiehi _17728__388 (.L_HI(net388));
 sg13g2_tiehi _17729__389 (.L_HI(net389));
 sg13g2_tiehi _17730__390 (.L_HI(net390));
 sg13g2_tiehi _17731__391 (.L_HI(net391));
 sg13g2_tiehi _17898__392 (.L_HI(net392));
 sg13g2_tiehi _17897__393 (.L_HI(net393));
 sg13g2_tiehi _17896__394 (.L_HI(net394));
 sg13g2_tiehi _17895__395 (.L_HI(net395));
 sg13g2_tiehi _17894__396 (.L_HI(net396));
 sg13g2_tiehi _17893__397 (.L_HI(net397));
 sg13g2_tiehi _17892__398 (.L_HI(net398));
 sg13g2_tiehi _17891__399 (.L_HI(net399));
 sg13g2_tiehi _17890__400 (.L_HI(net400));
 sg13g2_tiehi _17889__401 (.L_HI(net401));
 sg13g2_tiehi _17888__402 (.L_HI(net402));
 sg13g2_tiehi _17887__403 (.L_HI(net403));
 sg13g2_tiehi _17886__404 (.L_HI(net404));
 sg13g2_tiehi _17885__405 (.L_HI(net405));
 sg13g2_tiehi _17751__406 (.L_HI(net406));
 sg13g2_tiehi _17750__407 (.L_HI(net407));
 sg13g2_tiehi _17749__408 (.L_HI(net408));
 sg13g2_tiehi _17748__409 (.L_HI(net409));
 sg13g2_tiehi _17747__410 (.L_HI(net410));
 sg13g2_tiehi _17732__411 (.L_HI(net411));
 sg13g2_tiehi _17752__412 (.L_HI(net412));
 sg13g2_tiehi _17848__413 (.L_HI(net413));
 sg13g2_tiehi _17849__414 (.L_HI(net414));
 sg13g2_tiehi _17850__415 (.L_HI(net415));
 sg13g2_tiehi _17851__416 (.L_HI(net416));
 sg13g2_tiehi _17852__417 (.L_HI(net417));
 sg13g2_tiehi _17853__418 (.L_HI(net418));
 sg13g2_tiehi _17854__419 (.L_HI(net419));
 sg13g2_tiehi _17855__420 (.L_HI(net420));
 sg13g2_tiehi _17856__421 (.L_HI(net421));
 sg13g2_tiehi _17857__422 (.L_HI(net422));
 sg13g2_tiehi _17858__423 (.L_HI(net423));
 sg13g2_tiehi _17859__424 (.L_HI(net424));
 sg13g2_tiehi _17860__425 (.L_HI(net425));
 sg13g2_tiehi _17861__426 (.L_HI(net426));
 sg13g2_tiehi _17862__427 (.L_HI(net427));
 sg13g2_tiehi _17863__428 (.L_HI(net428));
 sg13g2_tiehi _17864__429 (.L_HI(net429));
 sg13g2_tiehi _17865__430 (.L_HI(net430));
 sg13g2_tiehi _17866__431 (.L_HI(net431));
 sg13g2_tiehi _17867__432 (.L_HI(net432));
 sg13g2_tiehi _17868__433 (.L_HI(net433));
 sg13g2_tiehi _17869__434 (.L_HI(net434));
 sg13g2_tiehi _17870__435 (.L_HI(net435));
 sg13g2_tiehi _17871__436 (.L_HI(net436));
 sg13g2_tiehi _17872__437 (.L_HI(net437));
 sg13g2_tiehi _17873__438 (.L_HI(net438));
 sg13g2_tiehi _17874__439 (.L_HI(net439));
 sg13g2_tiehi _17875__440 (.L_HI(net440));
 sg13g2_tiehi _17876__441 (.L_HI(net441));
 sg13g2_tiehi _17877__442 (.L_HI(net442));
 sg13g2_tiehi _17878__443 (.L_HI(net443));
 sg13g2_tiehi _17879__444 (.L_HI(net444));
 sg13g2_tiehi _17880__445 (.L_HI(net445));
 sg13g2_tiehi _17881__446 (.L_HI(net446));
 sg13g2_tiehi _17882__447 (.L_HI(net447));
 sg13g2_tiehi _17883__448 (.L_HI(net448));
 sg13g2_tiehi _17746__449 (.L_HI(net449));
 sg13g2_tiehi _17745__450 (.L_HI(net450));
 sg13g2_tiehi _17744__451 (.L_HI(net451));
 sg13g2_tiehi _17743__452 (.L_HI(net452));
 sg13g2_tiehi _17742__453 (.L_HI(net453));
 sg13g2_tiehi _17741__454 (.L_HI(net454));
 sg13g2_tiehi _17740__455 (.L_HI(net455));
 sg13g2_tiehi _17739__456 (.L_HI(net456));
 sg13g2_tiehi _17738__457 (.L_HI(net457));
 sg13g2_tiehi _17737__458 (.L_HI(net458));
 sg13g2_tiehi _17736__459 (.L_HI(net459));
 sg13g2_tiehi _17735__460 (.L_HI(net460));
 sg13g2_tiehi _17734__461 (.L_HI(net461));
 sg13g2_tiehi _17733__462 (.L_HI(net462));
 sg13g2_tiehi _17694__463 (.L_HI(net463));
 sg13g2_tiehi _17693__464 (.L_HI(net464));
 sg13g2_tiehi _17692__465 (.L_HI(net465));
 sg13g2_tiehi _17691__466 (.L_HI(net466));
 sg13g2_tiehi _17690__467 (.L_HI(net467));
 sg13g2_tiehi _17884__468 (.L_HI(net468));
 sg13g2_tiehi _17904__469 (.L_HI(net469));
 sg13g2_tiehi _17905__470 (.L_HI(net470));
 sg13g2_tiehi _17906__471 (.L_HI(net471));
 sg13g2_tiehi _17907__472 (.L_HI(net472));
 sg13g2_tiehi _17908__473 (.L_HI(net473));
 sg13g2_tiehi _17909__474 (.L_HI(net474));
 sg13g2_tiehi _17910__475 (.L_HI(net475));
 sg13g2_tiehi _17911__476 (.L_HI(net476));
 sg13g2_tiehi _17912__477 (.L_HI(net477));
 sg13g2_tiehi _17913__478 (.L_HI(net478));
 sg13g2_tiehi _17914__479 (.L_HI(net479));
 sg13g2_tiehi _17915__480 (.L_HI(net480));
 sg13g2_tiehi _17916__481 (.L_HI(net481));
 sg13g2_tiehi _17917__482 (.L_HI(net482));
 sg13g2_tiehi _17918__483 (.L_HI(net483));
 sg13g2_tiehi _17919__484 (.L_HI(net484));
 sg13g2_tiehi _17920__485 (.L_HI(net485));
 sg13g2_tiehi _17921__486 (.L_HI(net486));
 sg13g2_tiehi _17922__487 (.L_HI(net487));
 sg13g2_tiehi _17923__488 (.L_HI(net488));
 sg13g2_tiehi _17924__489 (.L_HI(net489));
 sg13g2_tiehi _17925__490 (.L_HI(net490));
 sg13g2_tiehi _17926__491 (.L_HI(net491));
 sg13g2_tiehi _17927__492 (.L_HI(net492));
 sg13g2_tiehi _17928__493 (.L_HI(net493));
 sg13g2_tiehi _17929__494 (.L_HI(net494));
 sg13g2_tiehi _17930__495 (.L_HI(net495));
 sg13g2_tiehi _17931__496 (.L_HI(net496));
 sg13g2_tiehi _17932__497 (.L_HI(net497));
 sg13g2_tiehi _17933__498 (.L_HI(net498));
 sg13g2_tiehi _17934__499 (.L_HI(net499));
 sg13g2_tiehi _17935__500 (.L_HI(net500));
 sg13g2_tiehi _17936__501 (.L_HI(net501));
 sg13g2_tiehi _17937__502 (.L_HI(net502));
 sg13g2_tiehi _17938__503 (.L_HI(net503));
 sg13g2_tiehi _17939__504 (.L_HI(net504));
 sg13g2_tiehi _17940__505 (.L_HI(net505));
 sg13g2_tiehi _17689__506 (.L_HI(net506));
 sg13g2_tiehi _17688__507 (.L_HI(net507));
 sg13g2_tiehi _17687__508 (.L_HI(net508));
 sg13g2_tiehi _17686__509 (.L_HI(net509));
 sg13g2_tiehi _17685__510 (.L_HI(net510));
 sg13g2_tiehi _17684__511 (.L_HI(net511));
 sg13g2_tiehi _17683__512 (.L_HI(net512));
 sg13g2_tiehi _17682__513 (.L_HI(net513));
 sg13g2_tiehi _17681__514 (.L_HI(net514));
 sg13g2_tiehi _17680__515 (.L_HI(net515));
 sg13g2_tiehi _17679__516 (.L_HI(net516));
 sg13g2_tiehi _17678__517 (.L_HI(net517));
 sg13g2_tiehi _17677__518 (.L_HI(net518));
 sg13g2_tiehi _17676__519 (.L_HI(net519));
 sg13g2_tiehi _17542__520 (.L_HI(net520));
 sg13g2_tiehi _17541__521 (.L_HI(net521));
 sg13g2_tiehi _17540__522 (.L_HI(net522));
 sg13g2_tiehi _17539__523 (.L_HI(net523));
 sg13g2_tiehi _17538__524 (.L_HI(net524));
 sg13g2_tiehi _17941__525 (.L_HI(net525));
 sg13g2_tiehi _17961__526 (.L_HI(net526));
 sg13g2_tiehi _18057__527 (.L_HI(net527));
 sg13g2_tiehi _18058__528 (.L_HI(net528));
 sg13g2_tiehi _18059__529 (.L_HI(net529));
 sg13g2_tiehi _18060__530 (.L_HI(net530));
 sg13g2_tiehi _18061__531 (.L_HI(net531));
 sg13g2_tiehi _18062__532 (.L_HI(net532));
 sg13g2_tiehi _18063__533 (.L_HI(net533));
 sg13g2_tiehi _18064__534 (.L_HI(net534));
 sg13g2_tiehi _18065__535 (.L_HI(net535));
 sg13g2_tiehi _18066__536 (.L_HI(net536));
 sg13g2_tiehi _18067__537 (.L_HI(net537));
 sg13g2_tiehi _18068__538 (.L_HI(net538));
 sg13g2_tiehi _18069__539 (.L_HI(net539));
 sg13g2_tiehi _18070__540 (.L_HI(net540));
 sg13g2_tiehi _18071__541 (.L_HI(net541));
 sg13g2_tiehi _18072__542 (.L_HI(net542));
 sg13g2_tiehi _18073__543 (.L_HI(net543));
 sg13g2_tiehi _18074__544 (.L_HI(net544));
 sg13g2_tiehi _18075__545 (.L_HI(net545));
 sg13g2_tiehi _18076__546 (.L_HI(net546));
 sg13g2_tiehi _18077__547 (.L_HI(net547));
 sg13g2_tiehi _18078__548 (.L_HI(net548));
 sg13g2_tiehi _18079__549 (.L_HI(net549));
 sg13g2_tiehi _18080__550 (.L_HI(net550));
 sg13g2_tiehi _18081__551 (.L_HI(net551));
 sg13g2_tiehi _18082__552 (.L_HI(net552));
 sg13g2_tiehi _18083__553 (.L_HI(net553));
 sg13g2_tiehi _18084__554 (.L_HI(net554));
 sg13g2_tiehi _18085__555 (.L_HI(net555));
 sg13g2_tiehi _18086__556 (.L_HI(net556));
 sg13g2_tiehi _18087__557 (.L_HI(net557));
 sg13g2_tiehi _18088__558 (.L_HI(net558));
 sg13g2_tiehi _18089__559 (.L_HI(net559));
 sg13g2_tiehi _18090__560 (.L_HI(net560));
 sg13g2_tiehi _18091__561 (.L_HI(net561));
 sg13g2_tiehi _18092__562 (.L_HI(net562));
 sg13g2_tiehi _17537__563 (.L_HI(net563));
 sg13g2_tiehi _17536__564 (.L_HI(net564));
 sg13g2_tiehi _17535__565 (.L_HI(net565));
 sg13g2_tiehi _17534__566 (.L_HI(net566));
 sg13g2_tiehi _17533__567 (.L_HI(net567));
 sg13g2_tiehi _17532__568 (.L_HI(net568));
 sg13g2_tiehi _17531__569 (.L_HI(net569));
 sg13g2_tiehi _17530__570 (.L_HI(net570));
 sg13g2_tiehi _17529__571 (.L_HI(net571));
 sg13g2_tiehi _17528__572 (.L_HI(net572));
 sg13g2_tiehi _17527__573 (.L_HI(net573));
 sg13g2_tiehi _17526__574 (.L_HI(net574));
 sg13g2_tiehi _17525__575 (.L_HI(net575));
 sg13g2_tiehi _17524__576 (.L_HI(net576));
 sg13g2_tiehi _17485__577 (.L_HI(net577));
 sg13g2_tiehi _17484__578 (.L_HI(net578));
 sg13g2_tiehi _17483__579 (.L_HI(net579));
 sg13g2_tiehi _17482__580 (.L_HI(net580));
 sg13g2_tiehi _17481__581 (.L_HI(net581));
 sg13g2_tiehi _18093__582 (.L_HI(net582));
 sg13g2_tiehi _18113__583 (.L_HI(net583));
 sg13g2_tiehi _18114__584 (.L_HI(net584));
 sg13g2_tiehi _18115__585 (.L_HI(net585));
 sg13g2_tiehi _18116__586 (.L_HI(net586));
 sg13g2_tiehi _18117__587 (.L_HI(net587));
 sg13g2_tiehi _18118__588 (.L_HI(net588));
 sg13g2_tiehi _18119__589 (.L_HI(net589));
 sg13g2_tiehi _18120__590 (.L_HI(net590));
 sg13g2_tiehi _18121__591 (.L_HI(net591));
 sg13g2_tiehi _18122__592 (.L_HI(net592));
 sg13g2_tiehi _18123__593 (.L_HI(net593));
 sg13g2_tiehi _18124__594 (.L_HI(net594));
 sg13g2_tiehi _18125__595 (.L_HI(net595));
 sg13g2_tiehi _18126__596 (.L_HI(net596));
 sg13g2_tiehi _18127__597 (.L_HI(net597));
 sg13g2_tiehi _18128__598 (.L_HI(net598));
 sg13g2_tiehi _18129__599 (.L_HI(net599));
 sg13g2_tiehi _18130__600 (.L_HI(net600));
 sg13g2_tiehi _18131__601 (.L_HI(net601));
 sg13g2_tiehi _18132__602 (.L_HI(net602));
 sg13g2_tiehi _18133__603 (.L_HI(net603));
 sg13g2_tiehi _18134__604 (.L_HI(net604));
 sg13g2_tiehi _18135__605 (.L_HI(net605));
 sg13g2_tiehi _18136__606 (.L_HI(net606));
 sg13g2_tiehi _18137__607 (.L_HI(net607));
 sg13g2_tiehi _18138__608 (.L_HI(net608));
 sg13g2_tiehi _18139__609 (.L_HI(net609));
 sg13g2_tiehi _18140__610 (.L_HI(net610));
 sg13g2_tiehi _18141__611 (.L_HI(net611));
 sg13g2_tiehi _18142__612 (.L_HI(net612));
 sg13g2_tiehi _18143__613 (.L_HI(net613));
 sg13g2_tiehi _18144__614 (.L_HI(net614));
 sg13g2_tiehi _18145__615 (.L_HI(net615));
 sg13g2_tiehi _18146__616 (.L_HI(net616));
 sg13g2_tiehi _18147__617 (.L_HI(net617));
 sg13g2_tiehi _18148__618 (.L_HI(net618));
 sg13g2_tiehi _18149__619 (.L_HI(net619));
 sg13g2_tiehi _17480__620 (.L_HI(net620));
 sg13g2_tiehi _17479__621 (.L_HI(net621));
 sg13g2_tiehi _17478__622 (.L_HI(net622));
 sg13g2_tiehi _17477__623 (.L_HI(net623));
 sg13g2_tiehi _17476__624 (.L_HI(net624));
 sg13g2_tiehi _17475__625 (.L_HI(net625));
 sg13g2_tiehi _17474__626 (.L_HI(net626));
 sg13g2_tiehi _17473__627 (.L_HI(net627));
 sg13g2_tiehi _17472__628 (.L_HI(net628));
 sg13g2_tiehi _17471__629 (.L_HI(net629));
 sg13g2_tiehi _17470__630 (.L_HI(net630));
 sg13g2_tiehi _17469__631 (.L_HI(net631));
 sg13g2_tiehi _17468__632 (.L_HI(net632));
 sg13g2_tiehi _17467__633 (.L_HI(net633));
 sg13g2_tiehi _18150__634 (.L_HI(net634));
 sg13g2_tiehi _18170__635 (.L_HI(net635));
 sg13g2_tiehi _18266__636 (.L_HI(net636));
 sg13g2_tiehi _18267__637 (.L_HI(net637));
 sg13g2_tiehi _18268__638 (.L_HI(net638));
 sg13g2_tiehi _18269__639 (.L_HI(net639));
 sg13g2_tiehi _18270__640 (.L_HI(net640));
 sg13g2_tiehi _18271__641 (.L_HI(net641));
 sg13g2_tiehi _18272__642 (.L_HI(net642));
 sg13g2_tiehi _18273__643 (.L_HI(net643));
 sg13g2_tiehi _18274__644 (.L_HI(net644));
 sg13g2_tiehi _18275__645 (.L_HI(net645));
 sg13g2_tiehi _18276__646 (.L_HI(net646));
 sg13g2_tiehi _18277__647 (.L_HI(net647));
 sg13g2_tiehi _18278__648 (.L_HI(net648));
 sg13g2_tiehi _18279__649 (.L_HI(net649));
 sg13g2_tiehi _18280__650 (.L_HI(net650));
 sg13g2_tiehi _18281__651 (.L_HI(net651));
 sg13g2_tiehi _18282__652 (.L_HI(net652));
 sg13g2_tiehi _18283__653 (.L_HI(net653));
 sg13g2_tiehi _18284__654 (.L_HI(net654));
 sg13g2_tiehi _18285__655 (.L_HI(net655));
 sg13g2_tiehi _18286__656 (.L_HI(net656));
 sg13g2_tiehi _18287__657 (.L_HI(net657));
 sg13g2_tiehi _18288__658 (.L_HI(net658));
 sg13g2_tiehi _18289__659 (.L_HI(net659));
 sg13g2_tiehi _18290__660 (.L_HI(net660));
 sg13g2_tiehi _18291__661 (.L_HI(net661));
 sg13g2_tiehi _18292__662 (.L_HI(net662));
 sg13g2_tiehi _18293__663 (.L_HI(net663));
 sg13g2_tiehi _18294__664 (.L_HI(net664));
 sg13g2_tiehi _18295__665 (.L_HI(net665));
 sg13g2_tiehi _18296__666 (.L_HI(net666));
 sg13g2_tiehi _18297__667 (.L_HI(net667));
 sg13g2_tiehi _18298__668 (.L_HI(net668));
 sg13g2_tiehi _18299__669 (.L_HI(net669));
 sg13g2_tiehi _18300__670 (.L_HI(net670));
 sg13g2_tiehi _18301__671 (.L_HI(net671));
 sg13g2_tiehi _18302__672 (.L_HI(net672));
 sg13g2_tiehi _18322__673 (.L_HI(net673));
 sg13g2_tiehi _18323__674 (.L_HI(net674));
 sg13g2_tiehi _18324__675 (.L_HI(net675));
 sg13g2_tiehi _18325__676 (.L_HI(net676));
 sg13g2_tiehi _18326__677 (.L_HI(net677));
 sg13g2_tiehi _18327__678 (.L_HI(net678));
 sg13g2_tiehi _18328__679 (.L_HI(net679));
 sg13g2_tiehi _18329__680 (.L_HI(net680));
 sg13g2_tiehi _18330__681 (.L_HI(net681));
 sg13g2_tiehi _18331__682 (.L_HI(net682));
 sg13g2_tiehi _18332__683 (.L_HI(net683));
 sg13g2_tiehi _18333__684 (.L_HI(net684));
 sg13g2_tiehi _18334__685 (.L_HI(net685));
 sg13g2_tiehi _18335__686 (.L_HI(net686));
 sg13g2_tiehi _18336__687 (.L_HI(net687));
 sg13g2_tiehi _18337__688 (.L_HI(net688));
 sg13g2_tiehi _18338__689 (.L_HI(net689));
 sg13g2_tiehi _18339__690 (.L_HI(net690));
 sg13g2_tiehi _18340__691 (.L_HI(net691));
 sg13g2_tiehi _18341__692 (.L_HI(net692));
 sg13g2_tiehi _18342__693 (.L_HI(net693));
 sg13g2_tiehi _18343__694 (.L_HI(net694));
 sg13g2_tiehi _18344__695 (.L_HI(net695));
 sg13g2_tiehi _18345__696 (.L_HI(net696));
 sg13g2_tiehi _18346__697 (.L_HI(net697));
 sg13g2_tiehi _18347__698 (.L_HI(net698));
 sg13g2_tiehi _18348__699 (.L_HI(net699));
 sg13g2_tiehi _18349__700 (.L_HI(net700));
 sg13g2_tiehi _18350__701 (.L_HI(net701));
 sg13g2_tiehi _18351__702 (.L_HI(net702));
 sg13g2_tiehi _18352__703 (.L_HI(net703));
 sg13g2_tiehi _18353__704 (.L_HI(net704));
 sg13g2_tiehi _18354__705 (.L_HI(net705));
 sg13g2_tiehi _18355__706 (.L_HI(net706));
 sg13g2_tiehi _18356__707 (.L_HI(net707));
 sg13g2_tiehi _18357__708 (.L_HI(net708));
 sg13g2_tiehi _18358__709 (.L_HI(net709));
 sg13g2_tiehi _18359__710 (.L_HI(net710));
 sg13g2_tiehi _18379__711 (.L_HI(net711));
 sg13g2_tiehi _18475__712 (.L_HI(net712));
 sg13g2_tiehi _18476__713 (.L_HI(net713));
 sg13g2_tiehi _18477__714 (.L_HI(net714));
 sg13g2_tiehi _18478__715 (.L_HI(net715));
 sg13g2_tiehi _18479__716 (.L_HI(net716));
 sg13g2_tiehi _18480__717 (.L_HI(net717));
 sg13g2_tiehi _18481__718 (.L_HI(net718));
 sg13g2_tiehi _18482__719 (.L_HI(net719));
 sg13g2_tiehi _18483__720 (.L_HI(net720));
 sg13g2_tiehi _18484__721 (.L_HI(net721));
 sg13g2_tiehi _18485__722 (.L_HI(net722));
 sg13g2_tiehi _18486__723 (.L_HI(net723));
 sg13g2_tiehi _18487__724 (.L_HI(net724));
 sg13g2_tiehi _18488__725 (.L_HI(net725));
 sg13g2_tiehi _18489__726 (.L_HI(net726));
 sg13g2_tiehi _18490__727 (.L_HI(net727));
 sg13g2_tiehi _18491__728 (.L_HI(net728));
 sg13g2_tiehi _18492__729 (.L_HI(net729));
 sg13g2_tiehi _18493__730 (.L_HI(net730));
 sg13g2_tiehi _18494__731 (.L_HI(net731));
 sg13g2_tiehi _18495__732 (.L_HI(net732));
 sg13g2_tiehi _18496__733 (.L_HI(net733));
 sg13g2_tiehi _18497__734 (.L_HI(net734));
 sg13g2_tiehi _18498__735 (.L_HI(net735));
 sg13g2_tiehi _18499__736 (.L_HI(net736));
 sg13g2_tiehi _18500__737 (.L_HI(net737));
 sg13g2_tiehi _18501__738 (.L_HI(net738));
 sg13g2_tiehi _18502__739 (.L_HI(net739));
 sg13g2_tiehi _18503__740 (.L_HI(net740));
 sg13g2_tiehi _18504__741 (.L_HI(net741));
 sg13g2_tiehi _18505__742 (.L_HI(net742));
 sg13g2_tiehi _18506__743 (.L_HI(net743));
 sg13g2_tiehi _18507__744 (.L_HI(net744));
 sg13g2_tiehi _18508__745 (.L_HI(net745));
 sg13g2_tiehi _18509__746 (.L_HI(net746));
 sg13g2_tiehi _18510__747 (.L_HI(net747));
 sg13g2_tiehi _18511__748 (.L_HI(net748));
 sg13g2_tiehi _18531__749 (.L_HI(net749));
 sg13g2_tiehi _18532__750 (.L_HI(net750));
 sg13g2_tiehi _18533__751 (.L_HI(net751));
 sg13g2_tiehi _18534__752 (.L_HI(net752));
 sg13g2_tiehi _18535__753 (.L_HI(net753));
 sg13g2_tiehi _18536__754 (.L_HI(net754));
 sg13g2_tiehi _18537__755 (.L_HI(net755));
 sg13g2_tiehi _18538__756 (.L_HI(net756));
 sg13g2_tiehi _18539__757 (.L_HI(net757));
 sg13g2_tiehi _18540__758 (.L_HI(net758));
 sg13g2_tiehi _18541__759 (.L_HI(net759));
 sg13g2_tiehi _18542__760 (.L_HI(net760));
 sg13g2_tiehi _18543__761 (.L_HI(net761));
 sg13g2_tiehi _18544__762 (.L_HI(net762));
 sg13g2_tiehi _18545__763 (.L_HI(net763));
 sg13g2_tiehi _18546__764 (.L_HI(net764));
 sg13g2_tiehi _18547__765 (.L_HI(net765));
 sg13g2_tiehi _18548__766 (.L_HI(net766));
 sg13g2_tiehi _18549__767 (.L_HI(net767));
 sg13g2_tiehi _18550__768 (.L_HI(net768));
 sg13g2_tiehi _18551__769 (.L_HI(net769));
 sg13g2_tiehi _18552__770 (.L_HI(net770));
 sg13g2_tiehi _18553__771 (.L_HI(net771));
 sg13g2_tiehi _18554__772 (.L_HI(net772));
 sg13g2_tiehi _18555__773 (.L_HI(net773));
 sg13g2_tiehi _18556__774 (.L_HI(net774));
 sg13g2_tiehi _18557__775 (.L_HI(net775));
 sg13g2_tiehi _18558__776 (.L_HI(net776));
 sg13g2_tiehi _18559__777 (.L_HI(net777));
 sg13g2_tiehi _18560__778 (.L_HI(net778));
 sg13g2_tiehi _18561__779 (.L_HI(net779));
 sg13g2_tiehi _18562__780 (.L_HI(net780));
 sg13g2_tiehi _18563__781 (.L_HI(net781));
 sg13g2_tiehi _18564__782 (.L_HI(net782));
 sg13g2_tiehi _18565__783 (.L_HI(net783));
 sg13g2_tiehi _18566__784 (.L_HI(net784));
 sg13g2_tiehi _18567__785 (.L_HI(net785));
 sg13g2_tiehi _18568__786 (.L_HI(net786));
 sg13g2_tiehi _18588__787 (.L_HI(net787));
 sg13g2_tiehi _18684__788 (.L_HI(net788));
 sg13g2_tiehi _18685__789 (.L_HI(net789));
 sg13g2_tiehi _18686__790 (.L_HI(net790));
 sg13g2_tiehi _18687__791 (.L_HI(net791));
 sg13g2_tiehi _18688__792 (.L_HI(net792));
 sg13g2_tiehi _18689__793 (.L_HI(net793));
 sg13g2_tiehi _18690__794 (.L_HI(net794));
 sg13g2_tiehi _18691__795 (.L_HI(net795));
 sg13g2_tiehi _18692__796 (.L_HI(net796));
 sg13g2_tiehi _18693__797 (.L_HI(net797));
 sg13g2_tiehi _18694__798 (.L_HI(net798));
 sg13g2_tiehi _18695__799 (.L_HI(net799));
 sg13g2_tiehi _18696__800 (.L_HI(net800));
 sg13g2_tiehi _18697__801 (.L_HI(net801));
 sg13g2_tiehi _18698__802 (.L_HI(net802));
 sg13g2_tiehi _18699__803 (.L_HI(net803));
 sg13g2_tiehi _18700__804 (.L_HI(net804));
 sg13g2_tiehi _18701__805 (.L_HI(net805));
 sg13g2_tiehi _18702__806 (.L_HI(net806));
 sg13g2_tiehi _18703__807 (.L_HI(net807));
 sg13g2_tiehi _18704__808 (.L_HI(net808));
 sg13g2_tiehi _18705__809 (.L_HI(net809));
 sg13g2_tiehi _18706__810 (.L_HI(net810));
 sg13g2_tiehi _18707__811 (.L_HI(net811));
 sg13g2_tiehi _18708__812 (.L_HI(net812));
 sg13g2_tiehi _18709__813 (.L_HI(net813));
 sg13g2_tiehi _18710__814 (.L_HI(net814));
 sg13g2_tiehi _18711__815 (.L_HI(net815));
 sg13g2_tiehi _18712__816 (.L_HI(net816));
 sg13g2_tiehi _18713__817 (.L_HI(net817));
 sg13g2_tiehi _18714__818 (.L_HI(net818));
 sg13g2_tiehi _18715__819 (.L_HI(net819));
 sg13g2_tiehi _18716__820 (.L_HI(net820));
 sg13g2_tiehi _18717__821 (.L_HI(net821));
 sg13g2_tiehi _18718__822 (.L_HI(net822));
 sg13g2_tiehi _18719__823 (.L_HI(net823));
 sg13g2_tiehi _18720__824 (.L_HI(net824));
 sg13g2_tiehi _18740__825 (.L_HI(net825));
 sg13g2_tiehi _18741__826 (.L_HI(net826));
 sg13g2_tiehi _18742__827 (.L_HI(net827));
 sg13g2_tiehi _18743__828 (.L_HI(net828));
 sg13g2_tiehi _18744__829 (.L_HI(net829));
 sg13g2_tiehi _18745__830 (.L_HI(net830));
 sg13g2_tiehi _18746__831 (.L_HI(net831));
 sg13g2_tiehi _18747__832 (.L_HI(net832));
 sg13g2_tiehi _18748__833 (.L_HI(net833));
 sg13g2_tiehi _18749__834 (.L_HI(net834));
 sg13g2_tiehi _18750__835 (.L_HI(net835));
 sg13g2_tiehi _18751__836 (.L_HI(net836));
 sg13g2_tiehi _18752__837 (.L_HI(net837));
 sg13g2_tiehi _18753__838 (.L_HI(net838));
 sg13g2_tiehi _18754__839 (.L_HI(net839));
 sg13g2_tiehi _18755__840 (.L_HI(net840));
 sg13g2_tiehi _18756__841 (.L_HI(net841));
 sg13g2_tiehi _18757__842 (.L_HI(net842));
 sg13g2_tiehi _18758__843 (.L_HI(net843));
 sg13g2_tiehi _18759__844 (.L_HI(net844));
 sg13g2_tiehi _18760__845 (.L_HI(net845));
 sg13g2_tiehi _18761__846 (.L_HI(net846));
 sg13g2_tiehi _18762__847 (.L_HI(net847));
 sg13g2_tiehi _18763__848 (.L_HI(net848));
 sg13g2_tiehi _18764__849 (.L_HI(net849));
 sg13g2_tiehi _18765__850 (.L_HI(net850));
 sg13g2_tiehi _18766__851 (.L_HI(net851));
 sg13g2_tiehi _18767__852 (.L_HI(net852));
 sg13g2_tiehi _18768__853 (.L_HI(net853));
 sg13g2_tiehi _18769__854 (.L_HI(net854));
 sg13g2_tiehi _18770__855 (.L_HI(net855));
 sg13g2_tiehi _18771__856 (.L_HI(net856));
 sg13g2_tiehi _18772__857 (.L_HI(net857));
 sg13g2_tiehi _18773__858 (.L_HI(net858));
 sg13g2_tiehi _18774__859 (.L_HI(net859));
 sg13g2_tiehi _18775__860 (.L_HI(net860));
 sg13g2_tiehi _18776__861 (.L_HI(net861));
 sg13g2_tiehi _18777__862 (.L_HI(net862));
 sg13g2_tiehi _18797__863 (.L_HI(net863));
 sg13g2_tiehi _18893__864 (.L_HI(net864));
 sg13g2_tiehi _18894__865 (.L_HI(net865));
 sg13g2_tiehi _18895__866 (.L_HI(net866));
 sg13g2_tiehi _18896__867 (.L_HI(net867));
 sg13g2_tiehi _18897__868 (.L_HI(net868));
 sg13g2_tiehi _18898__869 (.L_HI(net869));
 sg13g2_tiehi _18899__870 (.L_HI(net870));
 sg13g2_tiehi _18900__871 (.L_HI(net871));
 sg13g2_tiehi _18901__872 (.L_HI(net872));
 sg13g2_tiehi _18902__873 (.L_HI(net873));
 sg13g2_tiehi _18903__874 (.L_HI(net874));
 sg13g2_tiehi _18904__875 (.L_HI(net875));
 sg13g2_tiehi _18905__876 (.L_HI(net876));
 sg13g2_tiehi _18906__877 (.L_HI(net877));
 sg13g2_tiehi _18907__878 (.L_HI(net878));
 sg13g2_tiehi _18908__879 (.L_HI(net879));
 sg13g2_tiehi _18909__880 (.L_HI(net880));
 sg13g2_tiehi _18910__881 (.L_HI(net881));
 sg13g2_tiehi _18911__882 (.L_HI(net882));
 sg13g2_tiehi _18912__883 (.L_HI(net883));
 sg13g2_tiehi _18913__884 (.L_HI(net884));
 sg13g2_tiehi _18914__885 (.L_HI(net885));
 sg13g2_tiehi _18915__886 (.L_HI(net886));
 sg13g2_tiehi _18916__887 (.L_HI(net887));
 sg13g2_tiehi _18917__888 (.L_HI(net888));
 sg13g2_tiehi _18918__889 (.L_HI(net889));
 sg13g2_tiehi _18919__890 (.L_HI(net890));
 sg13g2_tiehi _18920__891 (.L_HI(net891));
 sg13g2_tiehi _18921__892 (.L_HI(net892));
 sg13g2_tiehi _18922__893 (.L_HI(net893));
 sg13g2_tiehi _18923__894 (.L_HI(net894));
 sg13g2_tiehi _18924__895 (.L_HI(net895));
 sg13g2_tiehi _18925__896 (.L_HI(net896));
 sg13g2_tiehi _18926__897 (.L_HI(net897));
 sg13g2_tiehi _18927__898 (.L_HI(net898));
 sg13g2_tiehi _18928__899 (.L_HI(net899));
 sg13g2_tiehi _18929__900 (.L_HI(net900));
 sg13g2_tiehi _18949__901 (.L_HI(net901));
 sg13g2_tiehi _18950__902 (.L_HI(net902));
 sg13g2_tiehi _18951__903 (.L_HI(net903));
 sg13g2_tiehi _18952__904 (.L_HI(net904));
 sg13g2_tiehi _18953__905 (.L_HI(net905));
 sg13g2_tiehi _18954__906 (.L_HI(net906));
 sg13g2_tiehi _18955__907 (.L_HI(net907));
 sg13g2_tiehi _18956__908 (.L_HI(net908));
 sg13g2_tiehi _18957__909 (.L_HI(net909));
 sg13g2_tiehi _18958__910 (.L_HI(net910));
 sg13g2_tiehi _18959__911 (.L_HI(net911));
 sg13g2_tiehi _18960__912 (.L_HI(net912));
 sg13g2_tiehi _18961__913 (.L_HI(net913));
 sg13g2_tiehi _18962__914 (.L_HI(net914));
 sg13g2_tiehi _18963__915 (.L_HI(net915));
 sg13g2_tiehi _18964__916 (.L_HI(net916));
 sg13g2_tiehi _18965__917 (.L_HI(net917));
 sg13g2_tiehi _18966__918 (.L_HI(net918));
 sg13g2_tiehi _18967__919 (.L_HI(net919));
 sg13g2_tiehi _18968__920 (.L_HI(net920));
 sg13g2_tiehi _18969__921 (.L_HI(net921));
 sg13g2_tiehi _18970__922 (.L_HI(net922));
 sg13g2_tiehi _18971__923 (.L_HI(net923));
 sg13g2_tiehi _18972__924 (.L_HI(net924));
 sg13g2_tiehi _18973__925 (.L_HI(net925));
 sg13g2_tiehi _18974__926 (.L_HI(net926));
 sg13g2_tiehi _18975__927 (.L_HI(net927));
 sg13g2_tiehi _18976__928 (.L_HI(net928));
 sg13g2_tiehi _18977__929 (.L_HI(net929));
 sg13g2_tiehi _18978__930 (.L_HI(net930));
 sg13g2_tiehi _18979__931 (.L_HI(net931));
 sg13g2_tiehi _18980__932 (.L_HI(net932));
 sg13g2_tiehi _18981__933 (.L_HI(net933));
 sg13g2_tiehi _18982__934 (.L_HI(net934));
 sg13g2_tiehi _18983__935 (.L_HI(net935));
 sg13g2_tiehi _18984__936 (.L_HI(net936));
 sg13g2_tiehi _18985__937 (.L_HI(net937));
 sg13g2_tiehi _18986__938 (.L_HI(net938));
 sg13g2_tiehi _19007__939 (.L_HI(net939));
 sg13g2_tiehi tt_um_supermic_arghunter_940 (.L_HI(net940));
 sg13g2_antennanp ANTENNA_1 (.A(_00628_));
 sg13g2_tielo tt_um_supermic_arghunter_7 (.L_LO(net7));
 sg13g2_tielo tt_um_supermic_arghunter_8 (.L_LO(net8));
 sg13g2_tielo tt_um_supermic_arghunter_9 (.L_LO(net9));
 sg13g2_tielo tt_um_supermic_arghunter_10 (.L_LO(net10));
 sg13g2_tielo tt_um_supermic_arghunter_11 (.L_LO(net11));
 sg13g2_tielo tt_um_supermic_arghunter_12 (.L_LO(net12));
 sg13g2_tielo tt_um_supermic_arghunter_13 (.L_LO(net13));
 sg13g2_tielo tt_um_supermic_arghunter_14 (.L_LO(net14));
 sg13g2_tielo tt_um_supermic_arghunter_15 (.L_LO(net15));
 sg13g2_tielo tt_um_supermic_arghunter_16 (.L_LO(net16));
 sg13g2_tielo tt_um_supermic_arghunter_17 (.L_LO(net17));
 sg13g2_tielo tt_um_supermic_arghunter_18 (.L_LO(net18));
 sg13g2_tiehi _16814__19 (.L_HI(net19));
 sg13g2_buf_2 _21448_ (.A(\u_supermic_top_module.i2s_out ),
    .X(uio_out[0]));
 sg13g2_buf_4 _21449_ (.X(uio_out[1]),
    .A(net5029));
 sg13g2_buf_2 _21450_ (.A(\u_supermic_top_module.i2s_bus_inst[0].c_i2s_bus.out ),
    .X(uo_out[0]));
 sg13g2_buf_2 _21451_ (.A(\u_supermic_top_module.i2s_bus_inst[1].c_i2s_bus.out ),
    .X(uo_out[1]));
 sg13g2_buf_2 _21452_ (.A(\u_supermic_top_module.i2s_bus_inst[2].c_i2s_bus.out ),
    .X(uo_out[2]));
 sg13g2_buf_4 _21453_ (.X(uo_out[3]),
    .A(\u_supermic_top_module.i2s_bus_inst[3].c_i2s_bus.out ));
 sg13g2_buf_2 _21454_ (.A(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.out ),
    .X(uo_out[4]));
 sg13g2_buf_2 _21455_ (.A(\u_supermic_top_module.i2s_bus_inst[5].c_i2s_bus.out ),
    .X(uo_out[5]));
 sg13g2_buf_2 _21456_ (.A(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.out ),
    .X(uo_out[6]));
 sg13g2_buf_2 _21457_ (.A(\u_supermic_top_module.i2s_bus_inst[7].c_i2s_bus.out ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout4646 (.X(net4646),
    .A(_04307_));
 sg13g2_buf_2 fanout4647 (.A(_02776_),
    .X(net4647));
 sg13g2_buf_1 fanout4648 (.A(_02776_),
    .X(net4648));
 sg13g2_buf_4 fanout4649 (.X(net4649),
    .A(net4651));
 sg13g2_buf_4 fanout4650 (.X(net4650),
    .A(_02746_));
 sg13g2_buf_2 fanout4651 (.A(_02746_),
    .X(net4651));
 sg13g2_buf_4 fanout4652 (.X(net4652),
    .A(net4653));
 sg13g2_buf_4 fanout4653 (.X(net4653),
    .A(_02744_));
 sg13g2_buf_4 fanout4654 (.X(net4654),
    .A(net4655));
 sg13g2_buf_4 fanout4655 (.X(net4655),
    .A(_02742_));
 sg13g2_buf_4 fanout4656 (.X(net4656),
    .A(net4657));
 sg13g2_buf_4 fanout4657 (.X(net4657),
    .A(_02738_));
 sg13g2_buf_4 fanout4658 (.X(net4658),
    .A(net4660));
 sg13g2_buf_4 fanout4659 (.X(net4659),
    .A(_02735_));
 sg13g2_buf_2 fanout4660 (.A(_02735_),
    .X(net4660));
 sg13g2_buf_4 fanout4661 (.X(net4661),
    .A(net4662));
 sg13g2_buf_2 fanout4662 (.A(_02734_),
    .X(net4662));
 sg13g2_buf_4 fanout4663 (.X(net4663),
    .A(_02734_));
 sg13g2_buf_4 fanout4664 (.X(net4664),
    .A(net4666));
 sg13g2_buf_4 fanout4665 (.X(net4665),
    .A(_02733_));
 sg13g2_buf_2 fanout4666 (.A(_02733_),
    .X(net4666));
 sg13g2_buf_4 fanout4667 (.X(net4667),
    .A(net4668));
 sg13g2_buf_4 fanout4668 (.X(net4668),
    .A(_02836_));
 sg13g2_buf_2 fanout4669 (.A(net4670),
    .X(net4669));
 sg13g2_buf_4 fanout4670 (.X(net4670),
    .A(_02834_));
 sg13g2_buf_4 fanout4671 (.X(net4671),
    .A(net4673));
 sg13g2_buf_4 fanout4672 (.X(net4672),
    .A(net4673));
 sg13g2_buf_4 fanout4673 (.X(net4673),
    .A(_02833_));
 sg13g2_buf_4 fanout4674 (.X(net4674),
    .A(net4675));
 sg13g2_buf_4 fanout4675 (.X(net4675),
    .A(_02831_));
 sg13g2_buf_2 fanout4676 (.A(net4677),
    .X(net4676));
 sg13g2_buf_4 fanout4677 (.X(net4677),
    .A(_02828_));
 sg13g2_buf_2 fanout4678 (.A(net4679),
    .X(net4678));
 sg13g2_buf_1 fanout4679 (.A(net4680),
    .X(net4679));
 sg13g2_buf_2 fanout4680 (.A(net4683),
    .X(net4680));
 sg13g2_buf_2 fanout4681 (.A(net4682),
    .X(net4681));
 sg13g2_buf_2 fanout4682 (.A(net4683),
    .X(net4682));
 sg13g2_buf_2 fanout4683 (.A(_02826_),
    .X(net4683));
 sg13g2_buf_4 fanout4684 (.X(net4684),
    .A(net4686));
 sg13g2_buf_4 fanout4685 (.X(net4685),
    .A(net4686));
 sg13g2_buf_2 fanout4686 (.A(_02825_),
    .X(net4686));
 sg13g2_buf_4 fanout4687 (.X(net4687),
    .A(net4688));
 sg13g2_buf_4 fanout4688 (.X(net4688),
    .A(_02807_));
 sg13g2_buf_4 fanout4689 (.X(net4689),
    .A(net4690));
 sg13g2_buf_4 fanout4690 (.X(net4690),
    .A(_02805_));
 sg13g2_buf_4 fanout4691 (.X(net4691),
    .A(net4692));
 sg13g2_buf_4 fanout4692 (.X(net4692),
    .A(_02802_));
 sg13g2_buf_4 fanout4693 (.X(net4693),
    .A(net4694));
 sg13g2_buf_4 fanout4694 (.X(net4694),
    .A(_02799_));
 sg13g2_buf_4 fanout4695 (.X(net4695),
    .A(net4696));
 sg13g2_buf_4 fanout4696 (.X(net4696),
    .A(_02796_));
 sg13g2_buf_2 fanout4697 (.A(net4700),
    .X(net4697));
 sg13g2_buf_2 fanout4698 (.A(net4700),
    .X(net4698));
 sg13g2_buf_2 fanout4699 (.A(net4700),
    .X(net4699));
 sg13g2_buf_2 fanout4700 (.A(_02793_),
    .X(net4700));
 sg13g2_buf_4 fanout4701 (.X(net4701),
    .A(net4703));
 sg13g2_buf_2 fanout4702 (.A(net4703),
    .X(net4702));
 sg13g2_buf_2 fanout4703 (.A(net4704),
    .X(net4703));
 sg13g2_buf_2 fanout4704 (.A(_02781_),
    .X(net4704));
 sg13g2_buf_2 fanout4705 (.A(net4706),
    .X(net4705));
 sg13g2_buf_2 fanout4706 (.A(net4707),
    .X(net4706));
 sg13g2_buf_2 fanout4707 (.A(net4708),
    .X(net4707));
 sg13g2_buf_2 fanout4708 (.A(_02777_),
    .X(net4708));
 sg13g2_buf_4 fanout4709 (.X(net4709),
    .A(net4710));
 sg13g2_buf_4 fanout4710 (.X(net4710),
    .A(net4711));
 sg13g2_buf_4 fanout4711 (.X(net4711),
    .A(_02719_));
 sg13g2_buf_4 fanout4712 (.X(net4712),
    .A(net4713));
 sg13g2_buf_4 fanout4713 (.X(net4713),
    .A(net4714));
 sg13g2_buf_4 fanout4714 (.X(net4714),
    .A(_02717_));
 sg13g2_buf_4 fanout4715 (.X(net4715),
    .A(net4717));
 sg13g2_buf_2 fanout4716 (.A(net4717),
    .X(net4716));
 sg13g2_buf_4 fanout4717 (.X(net4717),
    .A(net4718));
 sg13g2_buf_2 fanout4718 (.A(_02716_),
    .X(net4718));
 sg13g2_buf_4 fanout4719 (.X(net4719),
    .A(net4725));
 sg13g2_buf_4 fanout4720 (.X(net4720),
    .A(net4721));
 sg13g2_buf_2 fanout4721 (.A(net4722),
    .X(net4721));
 sg13g2_buf_2 fanout4722 (.A(net4724),
    .X(net4722));
 sg13g2_buf_4 fanout4723 (.X(net4723),
    .A(net4724));
 sg13g2_buf_4 fanout4724 (.X(net4724),
    .A(net4725));
 sg13g2_buf_8 fanout4725 (.A(_02715_),
    .X(net4725));
 sg13g2_buf_2 fanout4726 (.A(_02714_),
    .X(net4726));
 sg13g2_buf_4 fanout4727 (.X(net4727),
    .A(net4733));
 sg13g2_buf_4 fanout4728 (.X(net4728),
    .A(net4729));
 sg13g2_buf_4 fanout4729 (.X(net4729),
    .A(net4730));
 sg13g2_buf_4 fanout4730 (.X(net4730),
    .A(net4733));
 sg13g2_buf_4 fanout4731 (.X(net4731),
    .A(net4732));
 sg13g2_buf_4 fanout4732 (.X(net4732),
    .A(net4733));
 sg13g2_buf_8 fanout4733 (.A(_02703_),
    .X(net4733));
 sg13g2_buf_4 fanout4734 (.X(net4734),
    .A(net4735));
 sg13g2_buf_4 fanout4735 (.X(net4735),
    .A(net4736));
 sg13g2_buf_4 fanout4736 (.X(net4736),
    .A(_02702_));
 sg13g2_buf_4 fanout4737 (.X(net4737),
    .A(net4738));
 sg13g2_buf_4 fanout4738 (.X(net4738),
    .A(net4739));
 sg13g2_buf_4 fanout4739 (.X(net4739),
    .A(_02700_));
 sg13g2_buf_4 fanout4740 (.X(net4740),
    .A(net4741));
 sg13g2_buf_4 fanout4741 (.X(net4741),
    .A(net4742));
 sg13g2_buf_4 fanout4742 (.X(net4742),
    .A(_02698_));
 sg13g2_buf_4 fanout4743 (.X(net4743),
    .A(net4745));
 sg13g2_buf_2 fanout4744 (.A(net4745),
    .X(net4744));
 sg13g2_buf_4 fanout4745 (.X(net4745),
    .A(_02682_));
 sg13g2_buf_4 fanout4746 (.X(net4746),
    .A(net4748));
 sg13g2_buf_2 fanout4747 (.A(net4748),
    .X(net4747));
 sg13g2_buf_4 fanout4748 (.X(net4748),
    .A(_02678_));
 sg13g2_buf_4 fanout4749 (.X(net4749),
    .A(_02668_));
 sg13g2_buf_2 fanout4750 (.A(net4751),
    .X(net4750));
 sg13g2_buf_4 fanout4751 (.X(net4751),
    .A(_02668_));
 sg13g2_buf_4 fanout4752 (.X(net4752),
    .A(_02654_));
 sg13g2_buf_2 fanout4753 (.A(net4754),
    .X(net4753));
 sg13g2_buf_4 fanout4754 (.X(net4754),
    .A(_02654_));
 sg13g2_buf_4 fanout4755 (.X(net4755),
    .A(_02653_));
 sg13g2_buf_2 fanout4756 (.A(net4757),
    .X(net4756));
 sg13g2_buf_4 fanout4757 (.X(net4757),
    .A(_02653_));
 sg13g2_buf_4 fanout4758 (.X(net4758),
    .A(_02602_));
 sg13g2_buf_2 fanout4759 (.A(net4760),
    .X(net4759));
 sg13g2_buf_4 fanout4760 (.X(net4760),
    .A(_02602_));
 sg13g2_buf_4 fanout4761 (.X(net4761),
    .A(_02601_));
 sg13g2_buf_2 fanout4762 (.A(net4763),
    .X(net4762));
 sg13g2_buf_4 fanout4763 (.X(net4763),
    .A(_02601_));
 sg13g2_buf_4 fanout4764 (.X(net4764),
    .A(_02595_));
 sg13g2_buf_2 fanout4765 (.A(net4766),
    .X(net4765));
 sg13g2_buf_4 fanout4766 (.X(net4766),
    .A(_02595_));
 sg13g2_buf_4 fanout4767 (.X(net4767),
    .A(net4773));
 sg13g2_buf_4 fanout4768 (.X(net4768),
    .A(net4773));
 sg13g2_buf_4 fanout4769 (.X(net4769),
    .A(net4773));
 sg13g2_buf_1 fanout4770 (.A(net4773),
    .X(net4770));
 sg13g2_buf_4 fanout4771 (.X(net4771),
    .A(net4772));
 sg13g2_buf_2 fanout4772 (.A(net4773),
    .X(net4772));
 sg13g2_buf_4 fanout4773 (.X(net4773),
    .A(_02559_));
 sg13g2_buf_2 fanout4774 (.A(net4775),
    .X(net4774));
 sg13g2_buf_4 fanout4775 (.X(net4775),
    .A(_02792_));
 sg13g2_buf_4 fanout4776 (.X(net4776),
    .A(net4777));
 sg13g2_buf_2 fanout4777 (.A(net4778),
    .X(net4777));
 sg13g2_buf_2 fanout4778 (.A(net4779),
    .X(net4778));
 sg13g2_buf_4 fanout4779 (.X(net4779),
    .A(_02784_));
 sg13g2_buf_4 fanout4780 (.X(net4780),
    .A(net4781));
 sg13g2_buf_2 fanout4781 (.A(net4782),
    .X(net4781));
 sg13g2_buf_2 fanout4782 (.A(net4783),
    .X(net4782));
 sg13g2_buf_4 fanout4783 (.X(net4783),
    .A(_02780_));
 sg13g2_buf_4 fanout4784 (.X(net4784),
    .A(net4785));
 sg13g2_buf_2 fanout4785 (.A(net4786),
    .X(net4785));
 sg13g2_buf_2 fanout4786 (.A(_02779_),
    .X(net4786));
 sg13g2_buf_2 fanout4787 (.A(net4788),
    .X(net4787));
 sg13g2_buf_2 fanout4788 (.A(net4789),
    .X(net4788));
 sg13g2_buf_2 fanout4789 (.A(net4790),
    .X(net4789));
 sg13g2_buf_2 fanout4790 (.A(_02770_),
    .X(net4790));
 sg13g2_buf_4 fanout4791 (.X(net4791),
    .A(_02690_));
 sg13g2_buf_2 fanout4792 (.A(net4793),
    .X(net4792));
 sg13g2_buf_4 fanout4793 (.X(net4793),
    .A(_02690_));
 sg13g2_buf_4 fanout4794 (.X(net4794),
    .A(_02688_));
 sg13g2_buf_2 fanout4795 (.A(net4796),
    .X(net4795));
 sg13g2_buf_4 fanout4796 (.X(net4796),
    .A(_02688_));
 sg13g2_buf_4 fanout4797 (.X(net4797),
    .A(_02684_));
 sg13g2_buf_2 fanout4798 (.A(net4799),
    .X(net4798));
 sg13g2_buf_4 fanout4799 (.X(net4799),
    .A(_02684_));
 sg13g2_buf_4 fanout4800 (.X(net4800),
    .A(net4802));
 sg13g2_buf_4 fanout4801 (.X(net4801),
    .A(net4802));
 sg13g2_buf_4 fanout4802 (.X(net4802),
    .A(_02667_));
 sg13g2_buf_4 fanout4803 (.X(net4803),
    .A(net4806));
 sg13g2_buf_4 fanout4804 (.X(net4804),
    .A(net4806));
 sg13g2_buf_2 fanout4805 (.A(net4806),
    .X(net4805));
 sg13g2_buf_2 fanout4806 (.A(net4807),
    .X(net4806));
 sg13g2_buf_4 fanout4807 (.X(net4807),
    .A(_02667_));
 sg13g2_buf_4 fanout4808 (.X(net4808),
    .A(net4809));
 sg13g2_buf_4 fanout4809 (.X(net4809),
    .A(net4812));
 sg13g2_buf_4 fanout4810 (.X(net4810),
    .A(net4812));
 sg13g2_buf_2 fanout4811 (.A(net4812),
    .X(net4811));
 sg13g2_buf_2 fanout4812 (.A(_02667_),
    .X(net4812));
 sg13g2_buf_4 fanout4813 (.X(net4813),
    .A(_02651_));
 sg13g2_buf_4 fanout4814 (.X(net4814),
    .A(_02651_));
 sg13g2_buf_4 fanout4815 (.X(net4815),
    .A(net4818));
 sg13g2_buf_4 fanout4816 (.X(net4816),
    .A(net4818));
 sg13g2_buf_4 fanout4817 (.X(net4817),
    .A(net4818));
 sg13g2_buf_4 fanout4818 (.X(net4818),
    .A(_02651_));
 sg13g2_buf_2 fanout4819 (.A(net4821),
    .X(net4819));
 sg13g2_buf_4 fanout4820 (.X(net4820),
    .A(net4821));
 sg13g2_buf_4 fanout4821 (.X(net4821),
    .A(_02616_));
 sg13g2_buf_2 fanout4822 (.A(net4825),
    .X(net4822));
 sg13g2_buf_4 fanout4823 (.X(net4823),
    .A(net4825));
 sg13g2_buf_2 fanout4824 (.A(net4825),
    .X(net4824));
 sg13g2_buf_2 fanout4825 (.A(net4826),
    .X(net4825));
 sg13g2_buf_4 fanout4826 (.X(net4826),
    .A(_02558_));
 sg13g2_buf_4 fanout4827 (.X(net4827),
    .A(net4833));
 sg13g2_buf_2 fanout4828 (.A(net4829),
    .X(net4828));
 sg13g2_buf_2 fanout4829 (.A(net4833),
    .X(net4829));
 sg13g2_buf_2 fanout4830 (.A(net4831),
    .X(net4830));
 sg13g2_buf_1 fanout4831 (.A(net4832),
    .X(net4831));
 sg13g2_buf_2 fanout4832 (.A(net4833),
    .X(net4832));
 sg13g2_buf_2 fanout4833 (.A(_02558_),
    .X(net4833));
 sg13g2_buf_4 fanout4834 (.X(net4834),
    .A(net4836));
 sg13g2_buf_2 fanout4835 (.A(net4836),
    .X(net4835));
 sg13g2_buf_4 fanout4836 (.X(net4836),
    .A(net4837));
 sg13g2_buf_4 fanout4837 (.X(net4837),
    .A(net4842));
 sg13g2_buf_2 fanout4838 (.A(net4839),
    .X(net4838));
 sg13g2_buf_4 fanout4839 (.X(net4839),
    .A(net4842));
 sg13g2_buf_4 fanout4840 (.X(net4840),
    .A(net4842));
 sg13g2_buf_1 fanout4841 (.A(net4842),
    .X(net4841));
 sg13g2_buf_2 fanout4842 (.A(_02558_),
    .X(net4842));
 sg13g2_buf_4 fanout4843 (.X(net4843),
    .A(net4845));
 sg13g2_buf_4 fanout4844 (.X(net4844),
    .A(net4845));
 sg13g2_buf_4 fanout4845 (.X(net4845),
    .A(_02787_));
 sg13g2_buf_4 fanout4846 (.X(net4846),
    .A(net4847));
 sg13g2_buf_4 fanout4847 (.X(net4847),
    .A(net4848));
 sg13g2_buf_4 fanout4848 (.X(net4848),
    .A(_02691_));
 sg13g2_buf_4 fanout4849 (.X(net4849),
    .A(net4851));
 sg13g2_buf_2 fanout4850 (.A(net4851),
    .X(net4850));
 sg13g2_buf_4 fanout4851 (.X(net4851),
    .A(net4852));
 sg13g2_buf_4 fanout4852 (.X(net4852),
    .A(_02535_));
 sg13g2_buf_2 fanout4853 (.A(net4854),
    .X(net4853));
 sg13g2_buf_4 fanout4854 (.X(net4854),
    .A(_02530_));
 sg13g2_buf_2 fanout4855 (.A(net4856),
    .X(net4855));
 sg13g2_buf_4 fanout4856 (.X(net4856),
    .A(_02529_));
 sg13g2_buf_8 fanout4857 (.A(_02528_),
    .X(net4857));
 sg13g2_buf_4 fanout4858 (.X(net4858),
    .A(_02528_));
 sg13g2_buf_2 fanout4859 (.A(net4860),
    .X(net4859));
 sg13g2_buf_1 fanout4860 (.A(net4861),
    .X(net4860));
 sg13g2_buf_4 fanout4861 (.X(net4861),
    .A(_02527_));
 sg13g2_buf_4 fanout4862 (.X(net4862),
    .A(_02526_));
 sg13g2_buf_2 fanout4863 (.A(_02526_),
    .X(net4863));
 sg13g2_buf_2 fanout4864 (.A(net4865),
    .X(net4864));
 sg13g2_buf_2 fanout4865 (.A(net4866),
    .X(net4865));
 sg13g2_buf_4 fanout4866 (.X(net4866),
    .A(_02525_));
 sg13g2_buf_2 fanout4867 (.A(net4868),
    .X(net4867));
 sg13g2_buf_2 fanout4868 (.A(_02524_),
    .X(net4868));
 sg13g2_buf_2 fanout4869 (.A(net4870),
    .X(net4869));
 sg13g2_buf_8 fanout4870 (.A(_02523_),
    .X(net4870));
 sg13g2_buf_4 fanout4871 (.X(net4871),
    .A(net4872));
 sg13g2_buf_2 fanout4872 (.A(net4873),
    .X(net4872));
 sg13g2_buf_4 fanout4873 (.X(net4873),
    .A(net4877));
 sg13g2_buf_4 fanout4874 (.X(net4874),
    .A(net4876));
 sg13g2_buf_2 fanout4875 (.A(net4876),
    .X(net4875));
 sg13g2_buf_4 fanout4876 (.X(net4876),
    .A(net4877));
 sg13g2_buf_4 fanout4877 (.X(net4877),
    .A(_02631_));
 sg13g2_buf_2 fanout4878 (.A(net4886),
    .X(net4878));
 sg13g2_buf_2 fanout4879 (.A(net4886),
    .X(net4879));
 sg13g2_buf_2 fanout4880 (.A(net4881),
    .X(net4880));
 sg13g2_buf_1 fanout4881 (.A(net4882),
    .X(net4881));
 sg13g2_buf_2 fanout4882 (.A(net4883),
    .X(net4882));
 sg13g2_buf_2 fanout4883 (.A(net4886),
    .X(net4883));
 sg13g2_buf_2 fanout4884 (.A(net4886),
    .X(net4884));
 sg13g2_buf_2 fanout4885 (.A(net4886),
    .X(net4885));
 sg13g2_buf_4 fanout4886 (.X(net4886),
    .A(net4909));
 sg13g2_buf_4 fanout4887 (.X(net4887),
    .A(net4889));
 sg13g2_buf_2 fanout4888 (.A(net4889),
    .X(net4888));
 sg13g2_buf_2 fanout4889 (.A(net4890),
    .X(net4889));
 sg13g2_buf_4 fanout4890 (.X(net4890),
    .A(net4891));
 sg13g2_buf_8 fanout4891 (.A(net4909),
    .X(net4891));
 sg13g2_buf_4 fanout4892 (.X(net4892),
    .A(net4894));
 sg13g2_buf_4 fanout4893 (.X(net4893),
    .A(net4894));
 sg13g2_buf_4 fanout4894 (.X(net4894),
    .A(net4900));
 sg13g2_buf_4 fanout4895 (.X(net4895),
    .A(net4900));
 sg13g2_buf_2 fanout4896 (.A(net4900),
    .X(net4896));
 sg13g2_buf_4 fanout4897 (.X(net4897),
    .A(net4898));
 sg13g2_buf_4 fanout4898 (.X(net4898),
    .A(net4899));
 sg13g2_buf_4 fanout4899 (.X(net4899),
    .A(net4900));
 sg13g2_buf_4 fanout4900 (.X(net4900),
    .A(net4908));
 sg13g2_buf_2 fanout4901 (.A(net4902),
    .X(net4901));
 sg13g2_buf_2 fanout4902 (.A(net4905),
    .X(net4902));
 sg13g2_buf_2 fanout4903 (.A(net4904),
    .X(net4903));
 sg13g2_buf_4 fanout4904 (.X(net4904),
    .A(net4905));
 sg13g2_buf_1 fanout4905 (.A(net4906),
    .X(net4905));
 sg13g2_buf_4 fanout4906 (.X(net4906),
    .A(net4908));
 sg13g2_buf_4 fanout4907 (.X(net4907),
    .A(net4908));
 sg13g2_buf_4 fanout4908 (.X(net4908),
    .A(net4909));
 sg13g2_buf_8 fanout4909 (.A(net4923),
    .X(net4909));
 sg13g2_buf_4 fanout4910 (.X(net4910),
    .A(net4912));
 sg13g2_buf_2 fanout4911 (.A(net4912),
    .X(net4911));
 sg13g2_buf_8 fanout4912 (.A(net4913),
    .X(net4912));
 sg13g2_buf_4 fanout4913 (.X(net4913),
    .A(net4917));
 sg13g2_buf_4 fanout4914 (.X(net4914),
    .A(net4917));
 sg13g2_buf_2 fanout4915 (.A(net4917),
    .X(net4915));
 sg13g2_buf_8 fanout4916 (.A(net4917),
    .X(net4916));
 sg13g2_buf_2 fanout4917 (.A(net4923),
    .X(net4917));
 sg13g2_buf_4 fanout4918 (.X(net4918),
    .A(net4919));
 sg13g2_buf_2 fanout4919 (.A(net4923),
    .X(net4919));
 sg13g2_buf_4 fanout4920 (.X(net4920),
    .A(net4922));
 sg13g2_buf_4 fanout4921 (.X(net4921),
    .A(net4922));
 sg13g2_buf_4 fanout4922 (.X(net4922),
    .A(net4923));
 sg13g2_buf_8 fanout4923 (.A(_02522_),
    .X(net4923));
 sg13g2_buf_2 fanout4924 (.A(net4925),
    .X(net4924));
 sg13g2_buf_1 fanout4925 (.A(net4928),
    .X(net4925));
 sg13g2_buf_2 fanout4926 (.A(_02521_),
    .X(net4926));
 sg13g2_buf_8 fanout4927 (.A(net4928),
    .X(net4927));
 sg13g2_buf_8 fanout4928 (.A(_02521_),
    .X(net4928));
 sg13g2_buf_4 fanout4929 (.X(net4929),
    .A(net4933));
 sg13g2_buf_4 fanout4930 (.X(net4930),
    .A(net4933));
 sg13g2_buf_2 fanout4931 (.A(net4932),
    .X(net4931));
 sg13g2_buf_4 fanout4932 (.X(net4932),
    .A(net4933));
 sg13g2_buf_2 fanout4933 (.A(_02521_),
    .X(net4933));
 sg13g2_buf_2 fanout4934 (.A(_02499_),
    .X(net4934));
 sg13g2_buf_2 fanout4935 (.A(_02499_),
    .X(net4935));
 sg13g2_buf_2 fanout4936 (.A(net4937),
    .X(net4936));
 sg13g2_buf_2 fanout4937 (.A(_02455_),
    .X(net4937));
 sg13g2_buf_2 fanout4938 (.A(_02446_),
    .X(net4938));
 sg13g2_buf_1 fanout4939 (.A(_02446_),
    .X(net4939));
 sg13g2_buf_4 fanout4940 (.X(net4940),
    .A(_02434_));
 sg13g2_buf_1 fanout4941 (.A(_02434_),
    .X(net4941));
 sg13g2_buf_2 fanout4942 (.A(_02420_),
    .X(net4942));
 sg13g2_buf_2 fanout4943 (.A(_02420_),
    .X(net4943));
 sg13g2_buf_2 fanout4944 (.A(_02404_),
    .X(net4944));
 sg13g2_buf_1 fanout4945 (.A(_02404_),
    .X(net4945));
 sg13g2_buf_2 fanout4946 (.A(_02383_),
    .X(net4946));
 sg13g2_buf_1 fanout4947 (.A(_02383_),
    .X(net4947));
 sg13g2_buf_2 fanout4948 (.A(_02371_),
    .X(net4948));
 sg13g2_buf_2 fanout4949 (.A(_02371_),
    .X(net4949));
 sg13g2_buf_2 fanout4950 (.A(net4951),
    .X(net4950));
 sg13g2_buf_2 fanout4951 (.A(\u_supermic_top_module.cic_inst[3].u_cic.i_data ),
    .X(net4951));
 sg13g2_buf_4 fanout4952 (.X(net4952),
    .A(net4953));
 sg13g2_buf_2 fanout4953 (.A(\u_supermic_top_module.cic_inst[3].u_cic.i_data ),
    .X(net4953));
 sg13g2_buf_2 fanout4954 (.A(net4956),
    .X(net4954));
 sg13g2_buf_1 fanout4955 (.A(net4956),
    .X(net4955));
 sg13g2_buf_1 fanout4956 (.A(\u_supermic_top_module.cic_inst[7].u_cic.i_data ),
    .X(net4956));
 sg13g2_buf_2 fanout4957 (.A(net4958),
    .X(net4957));
 sg13g2_buf_2 fanout4958 (.A(\u_supermic_top_module.cic_inst[7].u_cic.i_data ),
    .X(net4958));
 sg13g2_buf_2 fanout4959 (.A(\u_supermic_top_module.cic_inst[2].u_cic.i_data ),
    .X(net4959));
 sg13g2_buf_2 fanout4960 (.A(\u_supermic_top_module.cic_inst[2].u_cic.i_data ),
    .X(net4960));
 sg13g2_buf_4 fanout4961 (.X(net4961),
    .A(net4962));
 sg13g2_buf_2 fanout4962 (.A(\u_supermic_top_module.cic_inst[2].u_cic.i_data ),
    .X(net4962));
 sg13g2_buf_2 fanout4963 (.A(net4964),
    .X(net4963));
 sg13g2_buf_4 fanout4964 (.X(net4964),
    .A(\u_supermic_top_module.cic_inst[6].u_cic.i_data ));
 sg13g2_buf_4 fanout4965 (.X(net4965),
    .A(net4966));
 sg13g2_buf_2 fanout4966 (.A(\u_supermic_top_module.cic_inst[6].u_cic.i_data ),
    .X(net4966));
 sg13g2_buf_2 fanout4967 (.A(net4969),
    .X(net4967));
 sg13g2_buf_2 fanout4968 (.A(net4969),
    .X(net4968));
 sg13g2_buf_2 fanout4969 (.A(net4971),
    .X(net4969));
 sg13g2_buf_2 fanout4970 (.A(net4971),
    .X(net4970));
 sg13g2_buf_2 fanout4971 (.A(\u_supermic_top_module.cic_inst[1].u_cic.i_data ),
    .X(net4971));
 sg13g2_buf_4 fanout4972 (.X(net4972),
    .A(\u_supermic_top_module.cic_inst[5].u_cic.i_data ));
 sg13g2_buf_2 fanout4973 (.A(\u_supermic_top_module.cic_inst[5].u_cic.i_data ),
    .X(net4973));
 sg13g2_buf_4 fanout4974 (.X(net4974),
    .A(net4975));
 sg13g2_buf_2 fanout4975 (.A(\u_supermic_top_module.cic_inst[5].u_cic.i_data ),
    .X(net4975));
 sg13g2_buf_4 fanout4976 (.X(net4976),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.i_data ));
 sg13g2_buf_2 fanout4977 (.A(\u_supermic_top_module.cic_inst[0].u_cic.i_data ),
    .X(net4977));
 sg13g2_buf_2 fanout4978 (.A(net4979),
    .X(net4978));
 sg13g2_buf_4 fanout4979 (.X(net4979),
    .A(\u_supermic_top_module.cic_inst[0].u_cic.i_data ));
 sg13g2_buf_2 fanout4980 (.A(net4981),
    .X(net4980));
 sg13g2_buf_4 fanout4981 (.X(net4981),
    .A(net4983));
 sg13g2_buf_4 fanout4982 (.X(net4982),
    .A(net4983));
 sg13g2_buf_2 fanout4983 (.A(\u_supermic_top_module.cic_inst[4].u_cic.i_data ),
    .X(net4983));
 sg13g2_buf_2 fanout4984 (.A(net4985),
    .X(net4984));
 sg13g2_buf_1 fanout4985 (.A(_02333_),
    .X(net4985));
 sg13g2_buf_2 fanout4986 (.A(_02332_),
    .X(net4986));
 sg13g2_buf_1 fanout4987 (.A(_02332_),
    .X(net4987));
 sg13g2_buf_2 fanout4988 (.A(net4994),
    .X(net4988));
 sg13g2_buf_1 fanout4989 (.A(net4994),
    .X(net4989));
 sg13g2_buf_2 fanout4990 (.A(net4991),
    .X(net4990));
 sg13g2_buf_1 fanout4991 (.A(net4994),
    .X(net4991));
 sg13g2_buf_2 fanout4992 (.A(net4994),
    .X(net4992));
 sg13g2_buf_1 fanout4993 (.A(net4994),
    .X(net4993));
 sg13g2_buf_2 fanout4994 (.A(net5),
    .X(net4994));
 sg13g2_buf_2 fanout4995 (.A(uio_in[3]),
    .X(net4995));
 sg13g2_buf_2 fanout4996 (.A(uio_in[3]),
    .X(net4996));
 sg13g2_buf_2 fanout4997 (.A(net4999),
    .X(net4997));
 sg13g2_buf_1 fanout4998 (.A(net4999),
    .X(net4998));
 sg13g2_buf_2 fanout4999 (.A(uio_in[3]),
    .X(net4999));
 sg13g2_buf_2 fanout5000 (.A(net5003),
    .X(net5000));
 sg13g2_buf_2 fanout5001 (.A(net5002),
    .X(net5001));
 sg13g2_buf_2 fanout5002 (.A(net5003),
    .X(net5002));
 sg13g2_buf_1 fanout5003 (.A(uio_in[2]),
    .X(net5003));
 sg13g2_buf_2 fanout5004 (.A(net5005),
    .X(net5004));
 sg13g2_buf_2 fanout5005 (.A(net5006),
    .X(net5005));
 sg13g2_buf_1 fanout5006 (.A(net5007),
    .X(net5006));
 sg13g2_buf_2 fanout5007 (.A(uio_in[1]),
    .X(net5007));
 sg13g2_buf_2 fanout5008 (.A(net5010),
    .X(net5008));
 sg13g2_buf_2 fanout5009 (.A(net5010),
    .X(net5009));
 sg13g2_buf_2 fanout5010 (.A(uio_in[0]),
    .X(net5010));
 sg13g2_buf_2 fanout5011 (.A(net5013),
    .X(net5011));
 sg13g2_buf_2 fanout5012 (.A(net5013),
    .X(net5012));
 sg13g2_buf_2 fanout5013 (.A(net5014),
    .X(net5013));
 sg13g2_buf_2 fanout5014 (.A(net5015),
    .X(net5014));
 sg13g2_buf_2 fanout5015 (.A(net5056),
    .X(net5015));
 sg13g2_buf_2 fanout5016 (.A(net5020),
    .X(net5016));
 sg13g2_buf_1 fanout5017 (.A(net5020),
    .X(net5017));
 sg13g2_buf_2 fanout5018 (.A(net5020),
    .X(net5018));
 sg13g2_buf_2 fanout5019 (.A(net5020),
    .X(net5019));
 sg13g2_buf_2 fanout5020 (.A(net5024),
    .X(net5020));
 sg13g2_buf_2 fanout5021 (.A(net5022),
    .X(net5021));
 sg13g2_buf_2 fanout5022 (.A(net5023),
    .X(net5022));
 sg13g2_buf_2 fanout5023 (.A(net5024),
    .X(net5023));
 sg13g2_buf_2 fanout5024 (.A(net5056),
    .X(net5024));
 sg13g2_buf_2 fanout5025 (.A(net5029),
    .X(net5025));
 sg13g2_buf_2 fanout5026 (.A(net5028),
    .X(net5026));
 sg13g2_buf_2 fanout5027 (.A(net5028),
    .X(net5027));
 sg13g2_buf_1 fanout5028 (.A(net5029),
    .X(net5028));
 sg13g2_buf_2 fanout5029 (.A(net5056),
    .X(net5029));
 sg13g2_buf_2 fanout5030 (.A(net5031),
    .X(net5030));
 sg13g2_buf_1 fanout5031 (.A(net5033),
    .X(net5031));
 sg13g2_buf_2 fanout5032 (.A(net5033),
    .X(net5032));
 sg13g2_buf_1 fanout5033 (.A(net5034),
    .X(net5033));
 sg13g2_buf_2 fanout5034 (.A(net5044),
    .X(net5034));
 sg13g2_buf_2 fanout5035 (.A(net5037),
    .X(net5035));
 sg13g2_buf_2 fanout5036 (.A(net5037),
    .X(net5036));
 sg13g2_buf_2 fanout5037 (.A(net5044),
    .X(net5037));
 sg13g2_buf_2 fanout5038 (.A(net5039),
    .X(net5038));
 sg13g2_buf_2 fanout5039 (.A(net5041),
    .X(net5039));
 sg13g2_buf_2 fanout5040 (.A(net5041),
    .X(net5040));
 sg13g2_buf_2 fanout5041 (.A(net5044),
    .X(net5041));
 sg13g2_buf_2 fanout5042 (.A(net5043),
    .X(net5042));
 sg13g2_buf_1 fanout5043 (.A(net5044),
    .X(net5043));
 sg13g2_buf_4 fanout5044 (.X(net5044),
    .A(net5056));
 sg13g2_buf_2 fanout5045 (.A(net5055),
    .X(net5045));
 sg13g2_buf_1 fanout5046 (.A(net5055),
    .X(net5046));
 sg13g2_buf_2 fanout5047 (.A(net5055),
    .X(net5047));
 sg13g2_buf_2 fanout5048 (.A(net5049),
    .X(net5048));
 sg13g2_buf_2 fanout5049 (.A(net5053),
    .X(net5049));
 sg13g2_buf_2 fanout5050 (.A(net5051),
    .X(net5050));
 sg13g2_buf_2 fanout5051 (.A(net5052),
    .X(net5051));
 sg13g2_buf_2 fanout5052 (.A(net5053),
    .X(net5052));
 sg13g2_buf_2 fanout5053 (.A(net5054),
    .X(net5053));
 sg13g2_buf_2 fanout5054 (.A(net5055),
    .X(net5054));
 sg13g2_buf_2 fanout5055 (.A(net5056),
    .X(net5055));
 sg13g2_buf_8 fanout5056 (.A(ui_in[1]),
    .X(net5056));
 sg13g2_buf_2 fanout5057 (.A(net5058),
    .X(net5057));
 sg13g2_buf_2 fanout5058 (.A(net5063),
    .X(net5058));
 sg13g2_buf_2 fanout5059 (.A(net5060),
    .X(net5059));
 sg13g2_buf_2 fanout5060 (.A(net5063),
    .X(net5060));
 sg13g2_buf_2 fanout5061 (.A(net5063),
    .X(net5061));
 sg13g2_buf_1 fanout5062 (.A(net5063),
    .X(net5062));
 sg13g2_buf_2 fanout5063 (.A(net5104),
    .X(net5063));
 sg13g2_buf_2 fanout5064 (.A(net5066),
    .X(net5064));
 sg13g2_buf_1 fanout5065 (.A(net5066),
    .X(net5065));
 sg13g2_buf_2 fanout5066 (.A(net5067),
    .X(net5066));
 sg13g2_buf_2 fanout5067 (.A(net5104),
    .X(net5067));
 sg13g2_buf_2 fanout5068 (.A(net5070),
    .X(net5068));
 sg13g2_buf_2 fanout5069 (.A(net5070),
    .X(net5069));
 sg13g2_buf_2 fanout5070 (.A(net5075),
    .X(net5070));
 sg13g2_buf_2 fanout5071 (.A(net5074),
    .X(net5071));
 sg13g2_buf_2 fanout5072 (.A(net5074),
    .X(net5072));
 sg13g2_buf_2 fanout5073 (.A(net5074),
    .X(net5073));
 sg13g2_buf_2 fanout5074 (.A(net5075),
    .X(net5074));
 sg13g2_buf_1 fanout5075 (.A(net5083),
    .X(net5075));
 sg13g2_buf_2 fanout5076 (.A(net5083),
    .X(net5076));
 sg13g2_buf_1 fanout5077 (.A(net5083),
    .X(net5077));
 sg13g2_buf_2 fanout5078 (.A(net5079),
    .X(net5078));
 sg13g2_buf_2 fanout5079 (.A(net5083),
    .X(net5079));
 sg13g2_buf_2 fanout5080 (.A(net5082),
    .X(net5080));
 sg13g2_buf_2 fanout5081 (.A(net5082),
    .X(net5081));
 sg13g2_buf_2 fanout5082 (.A(net5083),
    .X(net5082));
 sg13g2_buf_2 fanout5083 (.A(net5104),
    .X(net5083));
 sg13g2_buf_2 fanout5084 (.A(net5087),
    .X(net5084));
 sg13g2_buf_2 fanout5085 (.A(net5087),
    .X(net5085));
 sg13g2_buf_2 fanout5086 (.A(net5087),
    .X(net5086));
 sg13g2_buf_1 fanout5087 (.A(net5092),
    .X(net5087));
 sg13g2_buf_2 fanout5088 (.A(net5089),
    .X(net5088));
 sg13g2_buf_2 fanout5089 (.A(net5091),
    .X(net5089));
 sg13g2_buf_2 fanout5090 (.A(net5091),
    .X(net5090));
 sg13g2_buf_2 fanout5091 (.A(net5092),
    .X(net5091));
 sg13g2_buf_2 fanout5092 (.A(net5104),
    .X(net5092));
 sg13g2_buf_2 fanout5093 (.A(net5103),
    .X(net5093));
 sg13g2_buf_2 fanout5094 (.A(net5095),
    .X(net5094));
 sg13g2_buf_2 fanout5095 (.A(net5096),
    .X(net5095));
 sg13g2_buf_2 fanout5096 (.A(net5103),
    .X(net5096));
 sg13g2_buf_2 fanout5097 (.A(net5100),
    .X(net5097));
 sg13g2_buf_2 fanout5098 (.A(net5100),
    .X(net5098));
 sg13g2_buf_2 fanout5099 (.A(net5100),
    .X(net5099));
 sg13g2_buf_1 fanout5100 (.A(net5101),
    .X(net5100));
 sg13g2_buf_1 fanout5101 (.A(net5102),
    .X(net5101));
 sg13g2_buf_2 fanout5102 (.A(net5103),
    .X(net5102));
 sg13g2_buf_2 fanout5103 (.A(net5104),
    .X(net5103));
 sg13g2_buf_8 fanout5104 (.A(ui_in[1]),
    .X(net5104));
 sg13g2_buf_2 fanout5105 (.A(net5111),
    .X(net5105));
 sg13g2_buf_2 fanout5106 (.A(net5111),
    .X(net5106));
 sg13g2_buf_2 fanout5107 (.A(net5108),
    .X(net5107));
 sg13g2_buf_2 fanout5108 (.A(net5110),
    .X(net5108));
 sg13g2_buf_2 fanout5109 (.A(net5110),
    .X(net5109));
 sg13g2_buf_2 fanout5110 (.A(net5111),
    .X(net5110));
 sg13g2_buf_2 fanout5111 (.A(net5118),
    .X(net5111));
 sg13g2_buf_2 fanout5112 (.A(net5114),
    .X(net5112));
 sg13g2_buf_2 fanout5113 (.A(net5114),
    .X(net5113));
 sg13g2_buf_2 fanout5114 (.A(net5118),
    .X(net5114));
 sg13g2_buf_2 fanout5115 (.A(net5116),
    .X(net5115));
 sg13g2_buf_2 fanout5116 (.A(net5118),
    .X(net5116));
 sg13g2_buf_2 fanout5117 (.A(net5118),
    .X(net5117));
 sg13g2_buf_2 fanout5118 (.A(net5176),
    .X(net5118));
 sg13g2_buf_4 fanout5119 (.X(net5119),
    .A(net5129));
 sg13g2_buf_2 fanout5120 (.A(net5129),
    .X(net5120));
 sg13g2_buf_2 fanout5121 (.A(net5122),
    .X(net5121));
 sg13g2_buf_2 fanout5122 (.A(net5123),
    .X(net5122));
 sg13g2_buf_1 fanout5123 (.A(net5124),
    .X(net5123));
 sg13g2_buf_4 fanout5124 (.X(net5124),
    .A(net5129));
 sg13g2_buf_2 fanout5125 (.A(net5126),
    .X(net5125));
 sg13g2_buf_2 fanout5126 (.A(net5127),
    .X(net5126));
 sg13g2_buf_4 fanout5127 (.X(net5127),
    .A(net5128));
 sg13g2_buf_2 fanout5128 (.A(net5129),
    .X(net5128));
 sg13g2_buf_2 fanout5129 (.A(net5176),
    .X(net5129));
 sg13g2_buf_2 fanout5130 (.A(net5138),
    .X(net5130));
 sg13g2_buf_2 fanout5131 (.A(net5133),
    .X(net5131));
 sg13g2_buf_1 fanout5132 (.A(net5133),
    .X(net5132));
 sg13g2_buf_2 fanout5133 (.A(net5138),
    .X(net5133));
 sg13g2_buf_2 fanout5134 (.A(net5137),
    .X(net5134));
 sg13g2_buf_1 fanout5135 (.A(net5137),
    .X(net5135));
 sg13g2_buf_2 fanout5136 (.A(net5137),
    .X(net5136));
 sg13g2_buf_2 fanout5137 (.A(net5138),
    .X(net5137));
 sg13g2_buf_2 fanout5138 (.A(net5140),
    .X(net5138));
 sg13g2_buf_2 fanout5139 (.A(net5140),
    .X(net5139));
 sg13g2_buf_2 fanout5140 (.A(net5176),
    .X(net5140));
 sg13g2_buf_2 fanout5141 (.A(net5144),
    .X(net5141));
 sg13g2_buf_2 fanout5142 (.A(net5143),
    .X(net5142));
 sg13g2_buf_2 fanout5143 (.A(net5144),
    .X(net5143));
 sg13g2_buf_1 fanout5144 (.A(net5145),
    .X(net5144));
 sg13g2_buf_2 fanout5145 (.A(net5175),
    .X(net5145));
 sg13g2_buf_2 fanout5146 (.A(net5147),
    .X(net5146));
 sg13g2_buf_2 fanout5147 (.A(net5153),
    .X(net5147));
 sg13g2_buf_2 fanout5148 (.A(net5150),
    .X(net5148));
 sg13g2_buf_1 fanout5149 (.A(net5150),
    .X(net5149));
 sg13g2_buf_2 fanout5150 (.A(net5153),
    .X(net5150));
 sg13g2_buf_2 fanout5151 (.A(net5152),
    .X(net5151));
 sg13g2_buf_2 fanout5152 (.A(net5153),
    .X(net5152));
 sg13g2_buf_2 fanout5153 (.A(net5175),
    .X(net5153));
 sg13g2_buf_2 fanout5154 (.A(net5155),
    .X(net5154));
 sg13g2_buf_2 fanout5155 (.A(net5156),
    .X(net5155));
 sg13g2_buf_1 fanout5156 (.A(net5164),
    .X(net5156));
 sg13g2_buf_2 fanout5157 (.A(net5158),
    .X(net5157));
 sg13g2_buf_2 fanout5158 (.A(net5159),
    .X(net5158));
 sg13g2_buf_2 fanout5159 (.A(net5163),
    .X(net5159));
 sg13g2_buf_2 fanout5160 (.A(net5162),
    .X(net5160));
 sg13g2_buf_2 fanout5161 (.A(net5162),
    .X(net5161));
 sg13g2_buf_2 fanout5162 (.A(net5163),
    .X(net5162));
 sg13g2_buf_1 fanout5163 (.A(net5164),
    .X(net5163));
 sg13g2_buf_2 fanout5164 (.A(net5174),
    .X(net5164));
 sg13g2_buf_2 fanout5165 (.A(net5166),
    .X(net5165));
 sg13g2_buf_2 fanout5166 (.A(net5173),
    .X(net5166));
 sg13g2_buf_1 fanout5167 (.A(net5173),
    .X(net5167));
 sg13g2_buf_2 fanout5168 (.A(net5170),
    .X(net5168));
 sg13g2_buf_2 fanout5169 (.A(net5170),
    .X(net5169));
 sg13g2_buf_1 fanout5170 (.A(net5172),
    .X(net5170));
 sg13g2_buf_2 fanout5171 (.A(net5172),
    .X(net5171));
 sg13g2_buf_2 fanout5172 (.A(net5173),
    .X(net5172));
 sg13g2_buf_1 fanout5173 (.A(net5174),
    .X(net5173));
 sg13g2_buf_4 fanout5174 (.X(net5174),
    .A(net5175));
 sg13g2_buf_4 fanout5175 (.X(net5175),
    .A(net5176));
 sg13g2_buf_8 fanout5176 (.A(ui_in[1]),
    .X(net5176));
 sg13g2_buf_2 fanout5177 (.A(net5188),
    .X(net5177));
 sg13g2_buf_2 fanout5178 (.A(net5179),
    .X(net5178));
 sg13g2_buf_1 fanout5179 (.A(net5181),
    .X(net5179));
 sg13g2_buf_2 fanout5180 (.A(net5181),
    .X(net5180));
 sg13g2_buf_1 fanout5181 (.A(net5187),
    .X(net5181));
 sg13g2_buf_2 fanout5182 (.A(net5183),
    .X(net5182));
 sg13g2_buf_2 fanout5183 (.A(net5184),
    .X(net5183));
 sg13g2_buf_2 fanout5184 (.A(net5187),
    .X(net5184));
 sg13g2_buf_2 fanout5185 (.A(net5186),
    .X(net5185));
 sg13g2_buf_2 fanout5186 (.A(net5187),
    .X(net5186));
 sg13g2_buf_2 fanout5187 (.A(net5188),
    .X(net5187));
 sg13g2_buf_1 fanout5188 (.A(net5280),
    .X(net5188));
 sg13g2_buf_2 fanout5189 (.A(net5190),
    .X(net5189));
 sg13g2_buf_2 fanout5190 (.A(net5198),
    .X(net5190));
 sg13g2_buf_2 fanout5191 (.A(net5192),
    .X(net5191));
 sg13g2_buf_2 fanout5192 (.A(net5198),
    .X(net5192));
 sg13g2_buf_2 fanout5193 (.A(net5195),
    .X(net5193));
 sg13g2_buf_2 fanout5194 (.A(net5195),
    .X(net5194));
 sg13g2_buf_1 fanout5195 (.A(net5197),
    .X(net5195));
 sg13g2_buf_2 fanout5196 (.A(net5197),
    .X(net5196));
 sg13g2_buf_1 fanout5197 (.A(net5198),
    .X(net5197));
 sg13g2_buf_2 fanout5198 (.A(net5280),
    .X(net5198));
 sg13g2_buf_2 fanout5199 (.A(net5200),
    .X(net5199));
 sg13g2_buf_2 fanout5200 (.A(net5203),
    .X(net5200));
 sg13g2_buf_2 fanout5201 (.A(net5203),
    .X(net5201));
 sg13g2_buf_1 fanout5202 (.A(net5203),
    .X(net5202));
 sg13g2_buf_2 fanout5203 (.A(net5222),
    .X(net5203));
 sg13g2_buf_2 fanout5204 (.A(net5208),
    .X(net5204));
 sg13g2_buf_2 fanout5205 (.A(net5207),
    .X(net5205));
 sg13g2_buf_1 fanout5206 (.A(net5207),
    .X(net5206));
 sg13g2_buf_2 fanout5207 (.A(net5208),
    .X(net5207));
 sg13g2_buf_1 fanout5208 (.A(net5222),
    .X(net5208));
 sg13g2_buf_2 fanout5209 (.A(net5211),
    .X(net5209));
 sg13g2_buf_1 fanout5210 (.A(net5211),
    .X(net5210));
 sg13g2_buf_2 fanout5211 (.A(net5214),
    .X(net5211));
 sg13g2_buf_2 fanout5212 (.A(net5213),
    .X(net5212));
 sg13g2_buf_2 fanout5213 (.A(net5214),
    .X(net5213));
 sg13g2_buf_2 fanout5214 (.A(net5222),
    .X(net5214));
 sg13g2_buf_2 fanout5215 (.A(net5221),
    .X(net5215));
 sg13g2_buf_2 fanout5216 (.A(net5217),
    .X(net5216));
 sg13g2_buf_2 fanout5217 (.A(net5221),
    .X(net5217));
 sg13g2_buf_2 fanout5218 (.A(net5219),
    .X(net5218));
 sg13g2_buf_2 fanout5219 (.A(net5220),
    .X(net5219));
 sg13g2_buf_2 fanout5220 (.A(net5221),
    .X(net5220));
 sg13g2_buf_2 fanout5221 (.A(net5222),
    .X(net5221));
 sg13g2_buf_2 fanout5222 (.A(net5280),
    .X(net5222));
 sg13g2_buf_2 fanout5223 (.A(net5224),
    .X(net5223));
 sg13g2_buf_2 fanout5224 (.A(net5226),
    .X(net5224));
 sg13g2_buf_2 fanout5225 (.A(net5226),
    .X(net5225));
 sg13g2_buf_1 fanout5226 (.A(net5254),
    .X(net5226));
 sg13g2_buf_2 fanout5227 (.A(net5229),
    .X(net5227));
 sg13g2_buf_1 fanout5228 (.A(net5229),
    .X(net5228));
 sg13g2_buf_2 fanout5229 (.A(net5254),
    .X(net5229));
 sg13g2_buf_2 fanout5230 (.A(net5231),
    .X(net5230));
 sg13g2_buf_1 fanout5231 (.A(net5236),
    .X(net5231));
 sg13g2_buf_2 fanout5232 (.A(net5233),
    .X(net5232));
 sg13g2_buf_2 fanout5233 (.A(net5236),
    .X(net5233));
 sg13g2_buf_2 fanout5234 (.A(net5236),
    .X(net5234));
 sg13g2_buf_1 fanout5235 (.A(net5236),
    .X(net5235));
 sg13g2_buf_2 fanout5236 (.A(net5254),
    .X(net5236));
 sg13g2_buf_2 fanout5237 (.A(net5253),
    .X(net5237));
 sg13g2_buf_2 fanout5238 (.A(net5253),
    .X(net5238));
 sg13g2_buf_2 fanout5239 (.A(net5241),
    .X(net5239));
 sg13g2_buf_1 fanout5240 (.A(net5241),
    .X(net5240));
 sg13g2_buf_1 fanout5241 (.A(net5242),
    .X(net5241));
 sg13g2_buf_2 fanout5242 (.A(net5253),
    .X(net5242));
 sg13g2_buf_2 fanout5243 (.A(net5247),
    .X(net5243));
 sg13g2_buf_2 fanout5244 (.A(net5245),
    .X(net5244));
 sg13g2_buf_1 fanout5245 (.A(net5247),
    .X(net5245));
 sg13g2_buf_2 fanout5246 (.A(net5247),
    .X(net5246));
 sg13g2_buf_2 fanout5247 (.A(net5253),
    .X(net5247));
 sg13g2_buf_2 fanout5248 (.A(net5252),
    .X(net5248));
 sg13g2_buf_1 fanout5249 (.A(net5252),
    .X(net5249));
 sg13g2_buf_2 fanout5250 (.A(net5252),
    .X(net5250));
 sg13g2_buf_1 fanout5251 (.A(net5252),
    .X(net5251));
 sg13g2_buf_2 fanout5252 (.A(net5253),
    .X(net5252));
 sg13g2_buf_2 fanout5253 (.A(net5254),
    .X(net5253));
 sg13g2_buf_2 fanout5254 (.A(net5279),
    .X(net5254));
 sg13g2_buf_2 fanout5255 (.A(net5257),
    .X(net5255));
 sg13g2_buf_1 fanout5256 (.A(net5257),
    .X(net5256));
 sg13g2_buf_2 fanout5257 (.A(net5261),
    .X(net5257));
 sg13g2_buf_2 fanout5258 (.A(net5261),
    .X(net5258));
 sg13g2_buf_2 fanout5259 (.A(net5260),
    .X(net5259));
 sg13g2_buf_2 fanout5260 (.A(net5261),
    .X(net5260));
 sg13g2_buf_2 fanout5261 (.A(net5279),
    .X(net5261));
 sg13g2_buf_2 fanout5262 (.A(net5264),
    .X(net5262));
 sg13g2_buf_1 fanout5263 (.A(net5264),
    .X(net5263));
 sg13g2_buf_1 fanout5264 (.A(net5267),
    .X(net5264));
 sg13g2_buf_2 fanout5265 (.A(net5267),
    .X(net5265));
 sg13g2_buf_1 fanout5266 (.A(net5267),
    .X(net5266));
 sg13g2_buf_2 fanout5267 (.A(net5279),
    .X(net5267));
 sg13g2_buf_2 fanout5268 (.A(net5269),
    .X(net5268));
 sg13g2_buf_2 fanout5269 (.A(net5278),
    .X(net5269));
 sg13g2_buf_2 fanout5270 (.A(net5278),
    .X(net5270));
 sg13g2_buf_1 fanout5271 (.A(net5278),
    .X(net5271));
 sg13g2_buf_2 fanout5272 (.A(net5274),
    .X(net5272));
 sg13g2_buf_2 fanout5273 (.A(net5274),
    .X(net5273));
 sg13g2_buf_1 fanout5274 (.A(net5277),
    .X(net5274));
 sg13g2_buf_2 fanout5275 (.A(net5276),
    .X(net5275));
 sg13g2_buf_2 fanout5276 (.A(net5277),
    .X(net5276));
 sg13g2_buf_1 fanout5277 (.A(net5278),
    .X(net5277));
 sg13g2_buf_2 fanout5278 (.A(net5279),
    .X(net5278));
 sg13g2_buf_2 fanout5279 (.A(net5280),
    .X(net5279));
 sg13g2_buf_4 fanout5280 (.X(net5280),
    .A(net5686));
 sg13g2_buf_2 fanout5281 (.A(net5296),
    .X(net5281));
 sg13g2_buf_1 fanout5282 (.A(net5296),
    .X(net5282));
 sg13g2_buf_2 fanout5283 (.A(net5284),
    .X(net5283));
 sg13g2_buf_2 fanout5284 (.A(net5296),
    .X(net5284));
 sg13g2_buf_2 fanout5285 (.A(net5286),
    .X(net5285));
 sg13g2_buf_1 fanout5286 (.A(net5288),
    .X(net5286));
 sg13g2_buf_2 fanout5287 (.A(net5288),
    .X(net5287));
 sg13g2_buf_1 fanout5288 (.A(net5295),
    .X(net5288));
 sg13g2_buf_2 fanout5289 (.A(net5290),
    .X(net5289));
 sg13g2_buf_1 fanout5290 (.A(net5295),
    .X(net5290));
 sg13g2_buf_2 fanout5291 (.A(net5295),
    .X(net5291));
 sg13g2_buf_2 fanout5292 (.A(net5294),
    .X(net5292));
 sg13g2_buf_1 fanout5293 (.A(net5294),
    .X(net5293));
 sg13g2_buf_1 fanout5294 (.A(net5295),
    .X(net5294));
 sg13g2_buf_2 fanout5295 (.A(net5296),
    .X(net5295));
 sg13g2_buf_2 fanout5296 (.A(net5341),
    .X(net5296));
 sg13g2_buf_2 fanout5297 (.A(net5299),
    .X(net5297));
 sg13g2_buf_2 fanout5298 (.A(net5299),
    .X(net5298));
 sg13g2_buf_2 fanout5299 (.A(net5304),
    .X(net5299));
 sg13g2_buf_2 fanout5300 (.A(net5301),
    .X(net5300));
 sg13g2_buf_1 fanout5301 (.A(net5304),
    .X(net5301));
 sg13g2_buf_2 fanout5302 (.A(net5304),
    .X(net5302));
 sg13g2_buf_2 fanout5303 (.A(net5304),
    .X(net5303));
 sg13g2_buf_1 fanout5304 (.A(net5341),
    .X(net5304));
 sg13g2_buf_2 fanout5305 (.A(net5306),
    .X(net5305));
 sg13g2_buf_1 fanout5306 (.A(net5307),
    .X(net5306));
 sg13g2_buf_2 fanout5307 (.A(net5317),
    .X(net5307));
 sg13g2_buf_2 fanout5308 (.A(net5317),
    .X(net5308));
 sg13g2_buf_1 fanout5309 (.A(net5317),
    .X(net5309));
 sg13g2_buf_2 fanout5310 (.A(net5311),
    .X(net5310));
 sg13g2_buf_2 fanout5311 (.A(net5312),
    .X(net5311));
 sg13g2_buf_2 fanout5312 (.A(net5313),
    .X(net5312));
 sg13g2_buf_2 fanout5313 (.A(net5317),
    .X(net5313));
 sg13g2_buf_2 fanout5314 (.A(net5316),
    .X(net5314));
 sg13g2_buf_1 fanout5315 (.A(net5316),
    .X(net5315));
 sg13g2_buf_1 fanout5316 (.A(net5317),
    .X(net5316));
 sg13g2_buf_2 fanout5317 (.A(net5341),
    .X(net5317));
 sg13g2_buf_2 fanout5318 (.A(net5320),
    .X(net5318));
 sg13g2_buf_2 fanout5319 (.A(net5323),
    .X(net5319));
 sg13g2_buf_1 fanout5320 (.A(net5323),
    .X(net5320));
 sg13g2_buf_2 fanout5321 (.A(net5323),
    .X(net5321));
 sg13g2_buf_2 fanout5322 (.A(net5323),
    .X(net5322));
 sg13g2_buf_2 fanout5323 (.A(net5340),
    .X(net5323));
 sg13g2_buf_2 fanout5324 (.A(net5327),
    .X(net5324));
 sg13g2_buf_2 fanout5325 (.A(net5327),
    .X(net5325));
 sg13g2_buf_2 fanout5326 (.A(net5327),
    .X(net5326));
 sg13g2_buf_1 fanout5327 (.A(net5339),
    .X(net5327));
 sg13g2_buf_2 fanout5328 (.A(net5329),
    .X(net5328));
 sg13g2_buf_1 fanout5329 (.A(net5330),
    .X(net5329));
 sg13g2_buf_2 fanout5330 (.A(net5339),
    .X(net5330));
 sg13g2_buf_2 fanout5331 (.A(net5332),
    .X(net5331));
 sg13g2_buf_2 fanout5332 (.A(net5339),
    .X(net5332));
 sg13g2_buf_2 fanout5333 (.A(net5334),
    .X(net5333));
 sg13g2_buf_2 fanout5334 (.A(net5338),
    .X(net5334));
 sg13g2_buf_2 fanout5335 (.A(net5336),
    .X(net5335));
 sg13g2_buf_2 fanout5336 (.A(net5337),
    .X(net5336));
 sg13g2_buf_2 fanout5337 (.A(net5338),
    .X(net5337));
 sg13g2_buf_2 fanout5338 (.A(net5339),
    .X(net5338));
 sg13g2_buf_2 fanout5339 (.A(net5340),
    .X(net5339));
 sg13g2_buf_2 fanout5340 (.A(net5341),
    .X(net5340));
 sg13g2_buf_2 fanout5341 (.A(net5414),
    .X(net5341));
 sg13g2_buf_2 fanout5342 (.A(net5344),
    .X(net5342));
 sg13g2_buf_1 fanout5343 (.A(net5344),
    .X(net5343));
 sg13g2_buf_2 fanout5344 (.A(net5349),
    .X(net5344));
 sg13g2_buf_2 fanout5345 (.A(net5349),
    .X(net5345));
 sg13g2_buf_2 fanout5346 (.A(net5347),
    .X(net5346));
 sg13g2_buf_2 fanout5347 (.A(net5348),
    .X(net5347));
 sg13g2_buf_2 fanout5348 (.A(net5349),
    .X(net5348));
 sg13g2_buf_1 fanout5349 (.A(net5380),
    .X(net5349));
 sg13g2_buf_2 fanout5350 (.A(net5354),
    .X(net5350));
 sg13g2_buf_2 fanout5351 (.A(net5353),
    .X(net5351));
 sg13g2_buf_1 fanout5352 (.A(net5353),
    .X(net5352));
 sg13g2_buf_2 fanout5353 (.A(net5354),
    .X(net5353));
 sg13g2_buf_2 fanout5354 (.A(net5356),
    .X(net5354));
 sg13g2_buf_2 fanout5355 (.A(net5356),
    .X(net5355));
 sg13g2_buf_2 fanout5356 (.A(net5380),
    .X(net5356));
 sg13g2_buf_2 fanout5357 (.A(net5361),
    .X(net5357));
 sg13g2_buf_2 fanout5358 (.A(net5359),
    .X(net5358));
 sg13g2_buf_2 fanout5359 (.A(net5361),
    .X(net5359));
 sg13g2_buf_1 fanout5360 (.A(net5361),
    .X(net5360));
 sg13g2_buf_2 fanout5361 (.A(net5368),
    .X(net5361));
 sg13g2_buf_2 fanout5362 (.A(net5363),
    .X(net5362));
 sg13g2_buf_2 fanout5363 (.A(net5364),
    .X(net5363));
 sg13g2_buf_1 fanout5364 (.A(net5365),
    .X(net5364));
 sg13g2_buf_2 fanout5365 (.A(net5368),
    .X(net5365));
 sg13g2_buf_2 fanout5366 (.A(net5367),
    .X(net5366));
 sg13g2_buf_2 fanout5367 (.A(net5368),
    .X(net5367));
 sg13g2_buf_2 fanout5368 (.A(net5380),
    .X(net5368));
 sg13g2_buf_2 fanout5369 (.A(net5372),
    .X(net5369));
 sg13g2_buf_1 fanout5370 (.A(net5372),
    .X(net5370));
 sg13g2_buf_2 fanout5371 (.A(net5372),
    .X(net5371));
 sg13g2_buf_1 fanout5372 (.A(net5373),
    .X(net5372));
 sg13g2_buf_2 fanout5373 (.A(net5378),
    .X(net5373));
 sg13g2_buf_2 fanout5374 (.A(net5375),
    .X(net5374));
 sg13g2_buf_2 fanout5375 (.A(net5378),
    .X(net5375));
 sg13g2_buf_2 fanout5376 (.A(net5378),
    .X(net5376));
 sg13g2_buf_1 fanout5377 (.A(net5378),
    .X(net5377));
 sg13g2_buf_2 fanout5378 (.A(net5379),
    .X(net5378));
 sg13g2_buf_2 fanout5379 (.A(net5380),
    .X(net5379));
 sg13g2_buf_2 fanout5380 (.A(net5414),
    .X(net5380));
 sg13g2_buf_2 fanout5381 (.A(net5382),
    .X(net5381));
 sg13g2_buf_2 fanout5382 (.A(net5399),
    .X(net5382));
 sg13g2_buf_2 fanout5383 (.A(net5384),
    .X(net5383));
 sg13g2_buf_1 fanout5384 (.A(net5386),
    .X(net5384));
 sg13g2_buf_2 fanout5385 (.A(net5386),
    .X(net5385));
 sg13g2_buf_1 fanout5386 (.A(net5387),
    .X(net5386));
 sg13g2_buf_2 fanout5387 (.A(net5399),
    .X(net5387));
 sg13g2_buf_2 fanout5388 (.A(net5389),
    .X(net5388));
 sg13g2_buf_2 fanout5389 (.A(net5394),
    .X(net5389));
 sg13g2_buf_2 fanout5390 (.A(net5391),
    .X(net5390));
 sg13g2_buf_2 fanout5391 (.A(net5393),
    .X(net5391));
 sg13g2_buf_2 fanout5392 (.A(net5393),
    .X(net5392));
 sg13g2_buf_1 fanout5393 (.A(net5394),
    .X(net5393));
 sg13g2_buf_1 fanout5394 (.A(net5399),
    .X(net5394));
 sg13g2_buf_2 fanout5395 (.A(net5397),
    .X(net5395));
 sg13g2_buf_1 fanout5396 (.A(net5397),
    .X(net5396));
 sg13g2_buf_2 fanout5397 (.A(net5399),
    .X(net5397));
 sg13g2_buf_2 fanout5398 (.A(net5399),
    .X(net5398));
 sg13g2_buf_2 fanout5399 (.A(net5414),
    .X(net5399));
 sg13g2_buf_2 fanout5400 (.A(net5401),
    .X(net5400));
 sg13g2_buf_2 fanout5401 (.A(net5413),
    .X(net5401));
 sg13g2_buf_2 fanout5402 (.A(net5404),
    .X(net5402));
 sg13g2_buf_2 fanout5403 (.A(net5404),
    .X(net5403));
 sg13g2_buf_1 fanout5404 (.A(net5413),
    .X(net5404));
 sg13g2_buf_2 fanout5405 (.A(net5406),
    .X(net5405));
 sg13g2_buf_2 fanout5406 (.A(net5407),
    .X(net5406));
 sg13g2_buf_2 fanout5407 (.A(net5413),
    .X(net5407));
 sg13g2_buf_2 fanout5408 (.A(net5409),
    .X(net5408));
 sg13g2_buf_2 fanout5409 (.A(net5413),
    .X(net5409));
 sg13g2_buf_2 fanout5410 (.A(net5411),
    .X(net5410));
 sg13g2_buf_2 fanout5411 (.A(net5412),
    .X(net5411));
 sg13g2_buf_1 fanout5412 (.A(net5413),
    .X(net5412));
 sg13g2_buf_4 fanout5413 (.X(net5413),
    .A(net5414));
 sg13g2_buf_2 fanout5414 (.A(net5686),
    .X(net5414));
 sg13g2_buf_2 fanout5415 (.A(net5416),
    .X(net5415));
 sg13g2_buf_2 fanout5416 (.A(net5418),
    .X(net5416));
 sg13g2_buf_2 fanout5417 (.A(net5418),
    .X(net5417));
 sg13g2_buf_2 fanout5418 (.A(net5422),
    .X(net5418));
 sg13g2_buf_2 fanout5419 (.A(net5421),
    .X(net5419));
 sg13g2_buf_1 fanout5420 (.A(net5421),
    .X(net5420));
 sg13g2_buf_2 fanout5421 (.A(net5422),
    .X(net5421));
 sg13g2_buf_2 fanout5422 (.A(net5425),
    .X(net5422));
 sg13g2_buf_2 fanout5423 (.A(net5425),
    .X(net5423));
 sg13g2_buf_1 fanout5424 (.A(net5425),
    .X(net5424));
 sg13g2_buf_1 fanout5425 (.A(net5473),
    .X(net5425));
 sg13g2_buf_2 fanout5426 (.A(net5427),
    .X(net5426));
 sg13g2_buf_2 fanout5427 (.A(net5432),
    .X(net5427));
 sg13g2_buf_2 fanout5428 (.A(net5432),
    .X(net5428));
 sg13g2_buf_2 fanout5429 (.A(net5432),
    .X(net5429));
 sg13g2_buf_1 fanout5430 (.A(net5431),
    .X(net5430));
 sg13g2_buf_2 fanout5431 (.A(net5432),
    .X(net5431));
 sg13g2_buf_1 fanout5432 (.A(net5473),
    .X(net5432));
 sg13g2_buf_2 fanout5433 (.A(net5438),
    .X(net5433));
 sg13g2_buf_2 fanout5434 (.A(net5435),
    .X(net5434));
 sg13g2_buf_2 fanout5435 (.A(net5438),
    .X(net5435));
 sg13g2_buf_4 fanout5436 (.X(net5436),
    .A(net5438));
 sg13g2_buf_2 fanout5437 (.A(net5438),
    .X(net5437));
 sg13g2_buf_2 fanout5438 (.A(net5473),
    .X(net5438));
 sg13g2_buf_2 fanout5439 (.A(net5440),
    .X(net5439));
 sg13g2_buf_2 fanout5440 (.A(net5454),
    .X(net5440));
 sg13g2_buf_2 fanout5441 (.A(net5442),
    .X(net5441));
 sg13g2_buf_1 fanout5442 (.A(net5454),
    .X(net5442));
 sg13g2_buf_2 fanout5443 (.A(net5454),
    .X(net5443));
 sg13g2_buf_2 fanout5444 (.A(net5445),
    .X(net5444));
 sg13g2_buf_1 fanout5445 (.A(net5447),
    .X(net5445));
 sg13g2_buf_2 fanout5446 (.A(net5447),
    .X(net5446));
 sg13g2_buf_2 fanout5447 (.A(net5453),
    .X(net5447));
 sg13g2_buf_2 fanout5448 (.A(net5449),
    .X(net5448));
 sg13g2_buf_2 fanout5449 (.A(net5451),
    .X(net5449));
 sg13g2_buf_2 fanout5450 (.A(net5451),
    .X(net5450));
 sg13g2_buf_1 fanout5451 (.A(net5452),
    .X(net5451));
 sg13g2_buf_2 fanout5452 (.A(net5453),
    .X(net5452));
 sg13g2_buf_2 fanout5453 (.A(net5454),
    .X(net5453));
 sg13g2_buf_2 fanout5454 (.A(net5473),
    .X(net5454));
 sg13g2_buf_2 fanout5455 (.A(net5459),
    .X(net5455));
 sg13g2_buf_2 fanout5456 (.A(net5459),
    .X(net5456));
 sg13g2_buf_2 fanout5457 (.A(net5458),
    .X(net5457));
 sg13g2_buf_2 fanout5458 (.A(net5459),
    .X(net5458));
 sg13g2_buf_1 fanout5459 (.A(net5472),
    .X(net5459));
 sg13g2_buf_2 fanout5460 (.A(net5461),
    .X(net5460));
 sg13g2_buf_2 fanout5461 (.A(net5464),
    .X(net5461));
 sg13g2_buf_2 fanout5462 (.A(net5464),
    .X(net5462));
 sg13g2_buf_2 fanout5463 (.A(net5464),
    .X(net5463));
 sg13g2_buf_1 fanout5464 (.A(net5472),
    .X(net5464));
 sg13g2_buf_2 fanout5465 (.A(net5470),
    .X(net5465));
 sg13g2_buf_2 fanout5466 (.A(net5470),
    .X(net5466));
 sg13g2_buf_2 fanout5467 (.A(net5468),
    .X(net5467));
 sg13g2_buf_1 fanout5468 (.A(net5470),
    .X(net5468));
 sg13g2_buf_2 fanout5469 (.A(net5470),
    .X(net5469));
 sg13g2_buf_2 fanout5470 (.A(net5472),
    .X(net5470));
 sg13g2_buf_2 fanout5471 (.A(net5472),
    .X(net5471));
 sg13g2_buf_2 fanout5472 (.A(net5473),
    .X(net5472));
 sg13g2_buf_4 fanout5473 (.X(net5473),
    .A(net5686));
 sg13g2_buf_2 fanout5474 (.A(net5475),
    .X(net5474));
 sg13g2_buf_2 fanout5475 (.A(net5478),
    .X(net5475));
 sg13g2_buf_2 fanout5476 (.A(net5477),
    .X(net5476));
 sg13g2_buf_2 fanout5477 (.A(net5478),
    .X(net5477));
 sg13g2_buf_2 fanout5478 (.A(net5484),
    .X(net5478));
 sg13g2_buf_2 fanout5479 (.A(net5480),
    .X(net5479));
 sg13g2_buf_2 fanout5480 (.A(net5484),
    .X(net5480));
 sg13g2_buf_2 fanout5481 (.A(net5483),
    .X(net5481));
 sg13g2_buf_1 fanout5482 (.A(net5483),
    .X(net5482));
 sg13g2_buf_1 fanout5483 (.A(net5484),
    .X(net5483));
 sg13g2_buf_2 fanout5484 (.A(net5556),
    .X(net5484));
 sg13g2_buf_2 fanout5485 (.A(net5492),
    .X(net5485));
 sg13g2_buf_2 fanout5486 (.A(net5492),
    .X(net5486));
 sg13g2_buf_2 fanout5487 (.A(net5488),
    .X(net5487));
 sg13g2_buf_2 fanout5488 (.A(net5492),
    .X(net5488));
 sg13g2_buf_2 fanout5489 (.A(net5491),
    .X(net5489));
 sg13g2_buf_2 fanout5490 (.A(net5491),
    .X(net5490));
 sg13g2_buf_2 fanout5491 (.A(net5492),
    .X(net5491));
 sg13g2_buf_2 fanout5492 (.A(net5556),
    .X(net5492));
 sg13g2_buf_2 fanout5493 (.A(net5494),
    .X(net5493));
 sg13g2_buf_1 fanout5494 (.A(net5495),
    .X(net5494));
 sg13g2_buf_1 fanout5495 (.A(net5501),
    .X(net5495));
 sg13g2_buf_2 fanout5496 (.A(net5497),
    .X(net5496));
 sg13g2_buf_1 fanout5497 (.A(net5500),
    .X(net5497));
 sg13g2_buf_2 fanout5498 (.A(net5499),
    .X(net5498));
 sg13g2_buf_1 fanout5499 (.A(net5500),
    .X(net5499));
 sg13g2_buf_2 fanout5500 (.A(net5501),
    .X(net5500));
 sg13g2_buf_1 fanout5501 (.A(net5556),
    .X(net5501));
 sg13g2_buf_2 fanout5502 (.A(net5506),
    .X(net5502));
 sg13g2_buf_2 fanout5503 (.A(net5504),
    .X(net5503));
 sg13g2_buf_2 fanout5504 (.A(net5505),
    .X(net5504));
 sg13g2_buf_2 fanout5505 (.A(net5506),
    .X(net5505));
 sg13g2_buf_2 fanout5506 (.A(net5555),
    .X(net5506));
 sg13g2_buf_2 fanout5507 (.A(net5512),
    .X(net5507));
 sg13g2_buf_1 fanout5508 (.A(net5512),
    .X(net5508));
 sg13g2_buf_2 fanout5509 (.A(net5512),
    .X(net5509));
 sg13g2_buf_2 fanout5510 (.A(net5511),
    .X(net5510));
 sg13g2_buf_1 fanout5511 (.A(net5512),
    .X(net5511));
 sg13g2_buf_2 fanout5512 (.A(net5555),
    .X(net5512));
 sg13g2_buf_2 fanout5513 (.A(net5514),
    .X(net5513));
 sg13g2_buf_1 fanout5514 (.A(net5515),
    .X(net5514));
 sg13g2_buf_1 fanout5515 (.A(net5524),
    .X(net5515));
 sg13g2_buf_2 fanout5516 (.A(net5517),
    .X(net5516));
 sg13g2_buf_1 fanout5517 (.A(net5524),
    .X(net5517));
 sg13g2_buf_2 fanout5518 (.A(net5519),
    .X(net5518));
 sg13g2_buf_2 fanout5519 (.A(net5524),
    .X(net5519));
 sg13g2_buf_2 fanout5520 (.A(net5521),
    .X(net5520));
 sg13g2_buf_1 fanout5521 (.A(net5523),
    .X(net5521));
 sg13g2_buf_2 fanout5522 (.A(net5523),
    .X(net5522));
 sg13g2_buf_1 fanout5523 (.A(net5524),
    .X(net5523));
 sg13g2_buf_1 fanout5524 (.A(net5555),
    .X(net5524));
 sg13g2_buf_2 fanout5525 (.A(net5527),
    .X(net5525));
 sg13g2_buf_2 fanout5526 (.A(net5527),
    .X(net5526));
 sg13g2_buf_1 fanout5527 (.A(net5528),
    .X(net5527));
 sg13g2_buf_2 fanout5528 (.A(net5538),
    .X(net5528));
 sg13g2_buf_2 fanout5529 (.A(net5531),
    .X(net5529));
 sg13g2_buf_1 fanout5530 (.A(net5531),
    .X(net5530));
 sg13g2_buf_1 fanout5531 (.A(net5538),
    .X(net5531));
 sg13g2_buf_2 fanout5532 (.A(net5534),
    .X(net5532));
 sg13g2_buf_1 fanout5533 (.A(net5534),
    .X(net5533));
 sg13g2_buf_2 fanout5534 (.A(net5536),
    .X(net5534));
 sg13g2_buf_2 fanout5535 (.A(net5536),
    .X(net5535));
 sg13g2_buf_1 fanout5536 (.A(net5537),
    .X(net5536));
 sg13g2_buf_2 fanout5537 (.A(net5538),
    .X(net5537));
 sg13g2_buf_2 fanout5538 (.A(net5555),
    .X(net5538));
 sg13g2_buf_2 fanout5539 (.A(net5554),
    .X(net5539));
 sg13g2_buf_2 fanout5540 (.A(net5554),
    .X(net5540));
 sg13g2_buf_2 fanout5541 (.A(net5542),
    .X(net5541));
 sg13g2_buf_2 fanout5542 (.A(net5554),
    .X(net5542));
 sg13g2_buf_2 fanout5543 (.A(net5544),
    .X(net5543));
 sg13g2_buf_2 fanout5544 (.A(net5548),
    .X(net5544));
 sg13g2_buf_2 fanout5545 (.A(net5548),
    .X(net5545));
 sg13g2_buf_2 fanout5546 (.A(net5547),
    .X(net5546));
 sg13g2_buf_2 fanout5547 (.A(net5548),
    .X(net5547));
 sg13g2_buf_2 fanout5548 (.A(net5554),
    .X(net5548));
 sg13g2_buf_2 fanout5549 (.A(net5550),
    .X(net5549));
 sg13g2_buf_2 fanout5550 (.A(net5553),
    .X(net5550));
 sg13g2_buf_2 fanout5551 (.A(net5552),
    .X(net5551));
 sg13g2_buf_2 fanout5552 (.A(net5553),
    .X(net5552));
 sg13g2_buf_1 fanout5553 (.A(net5554),
    .X(net5553));
 sg13g2_buf_2 fanout5554 (.A(net5555),
    .X(net5554));
 sg13g2_buf_2 fanout5555 (.A(net5556),
    .X(net5555));
 sg13g2_buf_2 fanout5556 (.A(net5686),
    .X(net5556));
 sg13g2_buf_2 fanout5557 (.A(net5559),
    .X(net5557));
 sg13g2_buf_2 fanout5558 (.A(net5559),
    .X(net5558));
 sg13g2_buf_2 fanout5559 (.A(net5563),
    .X(net5559));
 sg13g2_buf_2 fanout5560 (.A(net5561),
    .X(net5560));
 sg13g2_buf_2 fanout5561 (.A(net5562),
    .X(net5561));
 sg13g2_buf_2 fanout5562 (.A(net5563),
    .X(net5562));
 sg13g2_buf_2 fanout5563 (.A(net5578),
    .X(net5563));
 sg13g2_buf_2 fanout5564 (.A(net5565),
    .X(net5564));
 sg13g2_buf_1 fanout5565 (.A(net5566),
    .X(net5565));
 sg13g2_buf_2 fanout5566 (.A(net5569),
    .X(net5566));
 sg13g2_buf_2 fanout5567 (.A(net5568),
    .X(net5567));
 sg13g2_buf_1 fanout5568 (.A(net5569),
    .X(net5568));
 sg13g2_buf_1 fanout5569 (.A(net5578),
    .X(net5569));
 sg13g2_buf_2 fanout5570 (.A(net5571),
    .X(net5570));
 sg13g2_buf_2 fanout5571 (.A(net5574),
    .X(net5571));
 sg13g2_buf_2 fanout5572 (.A(net5573),
    .X(net5572));
 sg13g2_buf_1 fanout5573 (.A(net5574),
    .X(net5573));
 sg13g2_buf_1 fanout5574 (.A(net5578),
    .X(net5574));
 sg13g2_buf_2 fanout5575 (.A(net5576),
    .X(net5575));
 sg13g2_buf_2 fanout5576 (.A(net5577),
    .X(net5576));
 sg13g2_buf_2 fanout5577 (.A(net5578),
    .X(net5577));
 sg13g2_buf_2 fanout5578 (.A(net5623),
    .X(net5578));
 sg13g2_buf_2 fanout5579 (.A(net5580),
    .X(net5579));
 sg13g2_buf_2 fanout5580 (.A(net5581),
    .X(net5580));
 sg13g2_buf_2 fanout5581 (.A(net5623),
    .X(net5581));
 sg13g2_buf_2 fanout5582 (.A(net5583),
    .X(net5582));
 sg13g2_buf_2 fanout5583 (.A(net5584),
    .X(net5583));
 sg13g2_buf_1 fanout5584 (.A(net5594),
    .X(net5584));
 sg13g2_buf_2 fanout5585 (.A(net5586),
    .X(net5585));
 sg13g2_buf_2 fanout5586 (.A(net5587),
    .X(net5586));
 sg13g2_buf_2 fanout5587 (.A(net5594),
    .X(net5587));
 sg13g2_buf_2 fanout5588 (.A(net5590),
    .X(net5588));
 sg13g2_buf_1 fanout5589 (.A(net5590),
    .X(net5589));
 sg13g2_buf_2 fanout5590 (.A(net5591),
    .X(net5590));
 sg13g2_buf_1 fanout5591 (.A(net5594),
    .X(net5591));
 sg13g2_buf_2 fanout5592 (.A(net5594),
    .X(net5592));
 sg13g2_buf_2 fanout5593 (.A(net5594),
    .X(net5593));
 sg13g2_buf_2 fanout5594 (.A(net5623),
    .X(net5594));
 sg13g2_buf_2 fanout5595 (.A(net5596),
    .X(net5595));
 sg13g2_buf_1 fanout5596 (.A(net5597),
    .X(net5596));
 sg13g2_buf_1 fanout5597 (.A(net5598),
    .X(net5597));
 sg13g2_buf_2 fanout5598 (.A(net5599),
    .X(net5598));
 sg13g2_buf_2 fanout5599 (.A(net5609),
    .X(net5599));
 sg13g2_buf_2 fanout5600 (.A(net5602),
    .X(net5600));
 sg13g2_buf_2 fanout5601 (.A(net5602),
    .X(net5601));
 sg13g2_buf_1 fanout5602 (.A(net5603),
    .X(net5602));
 sg13g2_buf_2 fanout5603 (.A(net5606),
    .X(net5603));
 sg13g2_buf_2 fanout5604 (.A(net5606),
    .X(net5604));
 sg13g2_buf_1 fanout5605 (.A(net5606),
    .X(net5605));
 sg13g2_buf_1 fanout5606 (.A(net5609),
    .X(net5606));
 sg13g2_buf_2 fanout5607 (.A(net5608),
    .X(net5607));
 sg13g2_buf_1 fanout5608 (.A(net5609),
    .X(net5608));
 sg13g2_buf_2 fanout5609 (.A(net5623),
    .X(net5609));
 sg13g2_buf_2 fanout5610 (.A(net5611),
    .X(net5610));
 sg13g2_buf_2 fanout5611 (.A(net5612),
    .X(net5611));
 sg13g2_buf_2 fanout5612 (.A(net5622),
    .X(net5612));
 sg13g2_buf_2 fanout5613 (.A(net5615),
    .X(net5613));
 sg13g2_buf_1 fanout5614 (.A(net5615),
    .X(net5614));
 sg13g2_buf_1 fanout5615 (.A(net5618),
    .X(net5615));
 sg13g2_buf_2 fanout5616 (.A(net5617),
    .X(net5616));
 sg13g2_buf_1 fanout5617 (.A(net5618),
    .X(net5617));
 sg13g2_buf_1 fanout5618 (.A(net5619),
    .X(net5618));
 sg13g2_buf_2 fanout5619 (.A(net5622),
    .X(net5619));
 sg13g2_buf_2 fanout5620 (.A(net5622),
    .X(net5620));
 sg13g2_buf_2 fanout5621 (.A(net5622),
    .X(net5621));
 sg13g2_buf_1 fanout5622 (.A(net5623),
    .X(net5622));
 sg13g2_buf_4 fanout5623 (.X(net5623),
    .A(net5685));
 sg13g2_buf_2 fanout5624 (.A(net5629),
    .X(net5624));
 sg13g2_buf_2 fanout5625 (.A(net5629),
    .X(net5625));
 sg13g2_buf_2 fanout5626 (.A(net5627),
    .X(net5626));
 sg13g2_buf_2 fanout5627 (.A(net5628),
    .X(net5627));
 sg13g2_buf_2 fanout5628 (.A(net5629),
    .X(net5628));
 sg13g2_buf_2 fanout5629 (.A(net5633),
    .X(net5629));
 sg13g2_buf_2 fanout5630 (.A(net5631),
    .X(net5630));
 sg13g2_buf_2 fanout5631 (.A(net5633),
    .X(net5631));
 sg13g2_buf_2 fanout5632 (.A(net5633),
    .X(net5632));
 sg13g2_buf_2 fanout5633 (.A(net5649),
    .X(net5633));
 sg13g2_buf_2 fanout5634 (.A(net5638),
    .X(net5634));
 sg13g2_buf_2 fanout5635 (.A(net5637),
    .X(net5635));
 sg13g2_buf_2 fanout5636 (.A(net5637),
    .X(net5636));
 sg13g2_buf_2 fanout5637 (.A(net5638),
    .X(net5637));
 sg13g2_buf_2 fanout5638 (.A(net5649),
    .X(net5638));
 sg13g2_buf_2 fanout5639 (.A(net5641),
    .X(net5639));
 sg13g2_buf_1 fanout5640 (.A(net5641),
    .X(net5640));
 sg13g2_buf_1 fanout5641 (.A(net5642),
    .X(net5641));
 sg13g2_buf_1 fanout5642 (.A(net5649),
    .X(net5642));
 sg13g2_buf_2 fanout5643 (.A(net5648),
    .X(net5643));
 sg13g2_buf_2 fanout5644 (.A(net5645),
    .X(net5644));
 sg13g2_buf_1 fanout5645 (.A(net5648),
    .X(net5645));
 sg13g2_buf_2 fanout5646 (.A(net5647),
    .X(net5646));
 sg13g2_buf_2 fanout5647 (.A(net5648),
    .X(net5647));
 sg13g2_buf_2 fanout5648 (.A(net5649),
    .X(net5648));
 sg13g2_buf_4 fanout5649 (.X(net5649),
    .A(net5685));
 sg13g2_buf_2 fanout5650 (.A(net5651),
    .X(net5650));
 sg13g2_buf_2 fanout5651 (.A(net5657),
    .X(net5651));
 sg13g2_buf_2 fanout5652 (.A(net5653),
    .X(net5652));
 sg13g2_buf_1 fanout5653 (.A(net5654),
    .X(net5653));
 sg13g2_buf_1 fanout5654 (.A(net5657),
    .X(net5654));
 sg13g2_buf_2 fanout5655 (.A(net5657),
    .X(net5655));
 sg13g2_buf_2 fanout5656 (.A(net5657),
    .X(net5656));
 sg13g2_buf_2 fanout5657 (.A(net5662),
    .X(net5657));
 sg13g2_buf_2 fanout5658 (.A(net5660),
    .X(net5658));
 sg13g2_buf_1 fanout5659 (.A(net5660),
    .X(net5659));
 sg13g2_buf_1 fanout5660 (.A(net5662),
    .X(net5660));
 sg13g2_buf_2 fanout5661 (.A(net5662),
    .X(net5661));
 sg13g2_buf_1 fanout5662 (.A(net5685),
    .X(net5662));
 sg13g2_buf_2 fanout5663 (.A(net5683),
    .X(net5663));
 sg13g2_buf_2 fanout5664 (.A(net5665),
    .X(net5664));
 sg13g2_buf_1 fanout5665 (.A(net5666),
    .X(net5665));
 sg13g2_buf_1 fanout5666 (.A(net5667),
    .X(net5666));
 sg13g2_buf_2 fanout5667 (.A(net5683),
    .X(net5667));
 sg13g2_buf_2 fanout5668 (.A(net5674),
    .X(net5668));
 sg13g2_buf_2 fanout5669 (.A(net5674),
    .X(net5669));
 sg13g2_buf_2 fanout5670 (.A(net5674),
    .X(net5670));
 sg13g2_buf_2 fanout5671 (.A(net5674),
    .X(net5671));
 sg13g2_buf_2 fanout5672 (.A(net5673),
    .X(net5672));
 sg13g2_buf_2 fanout5673 (.A(net5674),
    .X(net5673));
 sg13g2_buf_2 fanout5674 (.A(net5682),
    .X(net5674));
 sg13g2_buf_2 fanout5675 (.A(net5676),
    .X(net5675));
 sg13g2_buf_2 fanout5676 (.A(net5679),
    .X(net5676));
 sg13g2_buf_2 fanout5677 (.A(net5679),
    .X(net5677));
 sg13g2_buf_1 fanout5678 (.A(net5679),
    .X(net5678));
 sg13g2_buf_1 fanout5679 (.A(net5682),
    .X(net5679));
 sg13g2_buf_2 fanout5680 (.A(net5682),
    .X(net5680));
 sg13g2_buf_1 fanout5681 (.A(net5682),
    .X(net5681));
 sg13g2_buf_2 fanout5682 (.A(net5683),
    .X(net5682));
 sg13g2_buf_2 fanout5683 (.A(net5684),
    .X(net5683));
 sg13g2_buf_2 fanout5684 (.A(net5685),
    .X(net5684));
 sg13g2_buf_2 fanout5685 (.A(net5686),
    .X(net5685));
 sg13g2_buf_8 fanout5686 (.A(ui_in[0]),
    .X(net5686));
 sg13g2_buf_4 fanout5687 (.X(net5687),
    .A(net5698));
 sg13g2_buf_4 fanout5688 (.X(net5688),
    .A(net5689));
 sg13g2_buf_2 fanout5689 (.A(net5691),
    .X(net5689));
 sg13g2_buf_4 fanout5690 (.X(net5690),
    .A(net5691));
 sg13g2_buf_2 fanout5691 (.A(net5697),
    .X(net5691));
 sg13g2_buf_4 fanout5692 (.X(net5692),
    .A(net5693));
 sg13g2_buf_4 fanout5693 (.X(net5693),
    .A(net5694));
 sg13g2_buf_4 fanout5694 (.X(net5694),
    .A(net5697));
 sg13g2_buf_4 fanout5695 (.X(net5695),
    .A(net5696));
 sg13g2_buf_4 fanout5696 (.X(net5696),
    .A(net5697));
 sg13g2_buf_2 fanout5697 (.A(net5698),
    .X(net5697));
 sg13g2_buf_2 fanout5698 (.A(net5790),
    .X(net5698));
 sg13g2_buf_4 fanout5699 (.X(net5699),
    .A(net5700));
 sg13g2_buf_4 fanout5700 (.X(net5700),
    .A(net5708));
 sg13g2_buf_4 fanout5701 (.X(net5701),
    .A(net5702));
 sg13g2_buf_4 fanout5702 (.X(net5702),
    .A(net5708));
 sg13g2_buf_4 fanout5703 (.X(net5703),
    .A(net5705));
 sg13g2_buf_4 fanout5704 (.X(net5704),
    .A(net5705));
 sg13g2_buf_2 fanout5705 (.A(net5707),
    .X(net5705));
 sg13g2_buf_4 fanout5706 (.X(net5706),
    .A(net5707));
 sg13g2_buf_2 fanout5707 (.A(net5708),
    .X(net5707));
 sg13g2_buf_4 fanout5708 (.X(net5708),
    .A(net5790));
 sg13g2_buf_4 fanout5709 (.X(net5709),
    .A(net5710));
 sg13g2_buf_4 fanout5710 (.X(net5710),
    .A(net5713));
 sg13g2_buf_4 fanout5711 (.X(net5711),
    .A(net5713));
 sg13g2_buf_2 fanout5712 (.A(net5713),
    .X(net5712));
 sg13g2_buf_2 fanout5713 (.A(net5732),
    .X(net5713));
 sg13g2_buf_4 fanout5714 (.X(net5714),
    .A(net5718));
 sg13g2_buf_4 fanout5715 (.X(net5715),
    .A(net5717));
 sg13g2_buf_2 fanout5716 (.A(net5717),
    .X(net5716));
 sg13g2_buf_4 fanout5717 (.X(net5717),
    .A(net5718));
 sg13g2_buf_2 fanout5718 (.A(net5732),
    .X(net5718));
 sg13g2_buf_4 fanout5719 (.X(net5719),
    .A(net5720));
 sg13g2_buf_4 fanout5720 (.X(net5720),
    .A(net5724));
 sg13g2_buf_4 fanout5721 (.X(net5721),
    .A(net5723));
 sg13g2_buf_2 fanout5722 (.A(net5723),
    .X(net5722));
 sg13g2_buf_4 fanout5723 (.X(net5723),
    .A(net5724));
 sg13g2_buf_2 fanout5724 (.A(net5732),
    .X(net5724));
 sg13g2_buf_4 fanout5725 (.X(net5725),
    .A(net5731));
 sg13g2_buf_2 fanout5726 (.A(net5731),
    .X(net5726));
 sg13g2_buf_4 fanout5727 (.X(net5727),
    .A(net5731));
 sg13g2_buf_4 fanout5728 (.X(net5728),
    .A(net5729));
 sg13g2_buf_4 fanout5729 (.X(net5729),
    .A(net5730));
 sg13g2_buf_4 fanout5730 (.X(net5730),
    .A(net5731));
 sg13g2_buf_2 fanout5731 (.A(net5732),
    .X(net5731));
 sg13g2_buf_2 fanout5732 (.A(net5790),
    .X(net5732));
 sg13g2_buf_4 fanout5733 (.X(net5733),
    .A(net5734));
 sg13g2_buf_4 fanout5734 (.X(net5734),
    .A(net5736));
 sg13g2_buf_4 fanout5735 (.X(net5735),
    .A(net5736));
 sg13g2_buf_2 fanout5736 (.A(net5764),
    .X(net5736));
 sg13g2_buf_4 fanout5737 (.X(net5737),
    .A(net5739));
 sg13g2_buf_2 fanout5738 (.A(net5739),
    .X(net5738));
 sg13g2_buf_2 fanout5739 (.A(net5764),
    .X(net5739));
 sg13g2_buf_4 fanout5740 (.X(net5740),
    .A(net5741));
 sg13g2_buf_2 fanout5741 (.A(net5746),
    .X(net5741));
 sg13g2_buf_4 fanout5742 (.X(net5742),
    .A(net5743));
 sg13g2_buf_2 fanout5743 (.A(net5746),
    .X(net5743));
 sg13g2_buf_4 fanout5744 (.X(net5744),
    .A(net5746));
 sg13g2_buf_2 fanout5745 (.A(net5746),
    .X(net5745));
 sg13g2_buf_2 fanout5746 (.A(net5764),
    .X(net5746));
 sg13g2_buf_4 fanout5747 (.X(net5747),
    .A(net5763));
 sg13g2_buf_2 fanout5748 (.A(net5763),
    .X(net5748));
 sg13g2_buf_4 fanout5749 (.X(net5749),
    .A(net5751));
 sg13g2_buf_2 fanout5750 (.A(net5751),
    .X(net5750));
 sg13g2_buf_2 fanout5751 (.A(net5752),
    .X(net5751));
 sg13g2_buf_4 fanout5752 (.X(net5752),
    .A(net5763));
 sg13g2_buf_4 fanout5753 (.X(net5753),
    .A(net5757));
 sg13g2_buf_4 fanout5754 (.X(net5754),
    .A(net5755));
 sg13g2_buf_2 fanout5755 (.A(net5757),
    .X(net5755));
 sg13g2_buf_4 fanout5756 (.X(net5756),
    .A(net5757));
 sg13g2_buf_2 fanout5757 (.A(net5763),
    .X(net5757));
 sg13g2_buf_4 fanout5758 (.X(net5758),
    .A(net5762));
 sg13g2_buf_2 fanout5759 (.A(net5762),
    .X(net5759));
 sg13g2_buf_4 fanout5760 (.X(net5760),
    .A(net5762));
 sg13g2_buf_2 fanout5761 (.A(net5762),
    .X(net5761));
 sg13g2_buf_2 fanout5762 (.A(net5763),
    .X(net5762));
 sg13g2_buf_2 fanout5763 (.A(net5764),
    .X(net5763));
 sg13g2_buf_2 fanout5764 (.A(net5789),
    .X(net5764));
 sg13g2_buf_4 fanout5765 (.X(net5765),
    .A(net5767));
 sg13g2_buf_2 fanout5766 (.A(net5767),
    .X(net5766));
 sg13g2_buf_4 fanout5767 (.X(net5767),
    .A(net5771));
 sg13g2_buf_4 fanout5768 (.X(net5768),
    .A(net5771));
 sg13g2_buf_4 fanout5769 (.X(net5769),
    .A(net5770));
 sg13g2_buf_4 fanout5770 (.X(net5770),
    .A(net5771));
 sg13g2_buf_4 fanout5771 (.X(net5771),
    .A(net5789));
 sg13g2_buf_4 fanout5772 (.X(net5772),
    .A(net5774));
 sg13g2_buf_2 fanout5773 (.A(net5774),
    .X(net5773));
 sg13g2_buf_2 fanout5774 (.A(net5777),
    .X(net5774));
 sg13g2_buf_4 fanout5775 (.X(net5775),
    .A(net5777));
 sg13g2_buf_2 fanout5776 (.A(net5777),
    .X(net5776));
 sg13g2_buf_2 fanout5777 (.A(net5789),
    .X(net5777));
 sg13g2_buf_4 fanout5778 (.X(net5778),
    .A(net5779));
 sg13g2_buf_4 fanout5779 (.X(net5779),
    .A(net5788));
 sg13g2_buf_4 fanout5780 (.X(net5780),
    .A(net5788));
 sg13g2_buf_2 fanout5781 (.A(net5788),
    .X(net5781));
 sg13g2_buf_4 fanout5782 (.X(net5782),
    .A(net5784));
 sg13g2_buf_4 fanout5783 (.X(net5783),
    .A(net5784));
 sg13g2_buf_2 fanout5784 (.A(net5787),
    .X(net5784));
 sg13g2_buf_4 fanout5785 (.X(net5785),
    .A(net5786));
 sg13g2_buf_4 fanout5786 (.X(net5786),
    .A(net5787));
 sg13g2_buf_2 fanout5787 (.A(net5788),
    .X(net5787));
 sg13g2_buf_2 fanout5788 (.A(net5789),
    .X(net5788));
 sg13g2_buf_2 fanout5789 (.A(net5790),
    .X(net5789));
 sg13g2_buf_4 fanout5790 (.X(net5790),
    .A(net6196));
 sg13g2_buf_4 fanout5791 (.X(net5791),
    .A(net5806));
 sg13g2_buf_2 fanout5792 (.A(net5806),
    .X(net5792));
 sg13g2_buf_4 fanout5793 (.X(net5793),
    .A(net5794));
 sg13g2_buf_2 fanout5794 (.A(net5806),
    .X(net5794));
 sg13g2_buf_4 fanout5795 (.X(net5795),
    .A(net5796));
 sg13g2_buf_2 fanout5796 (.A(net5798),
    .X(net5796));
 sg13g2_buf_4 fanout5797 (.X(net5797),
    .A(net5798));
 sg13g2_buf_2 fanout5798 (.A(net5805),
    .X(net5798));
 sg13g2_buf_4 fanout5799 (.X(net5799),
    .A(net5800));
 sg13g2_buf_2 fanout5800 (.A(net5805),
    .X(net5800));
 sg13g2_buf_4 fanout5801 (.X(net5801),
    .A(net5805));
 sg13g2_buf_4 fanout5802 (.X(net5802),
    .A(net5804));
 sg13g2_buf_2 fanout5803 (.A(net5804),
    .X(net5803));
 sg13g2_buf_2 fanout5804 (.A(net5805),
    .X(net5804));
 sg13g2_buf_2 fanout5805 (.A(net5806),
    .X(net5805));
 sg13g2_buf_2 fanout5806 (.A(net5827),
    .X(net5806));
 sg13g2_buf_4 fanout5807 (.X(net5807),
    .A(net5809));
 sg13g2_buf_4 fanout5808 (.X(net5808),
    .A(net5809));
 sg13g2_buf_4 fanout5809 (.X(net5809),
    .A(net5827));
 sg13g2_buf_4 fanout5810 (.X(net5810),
    .A(net5813));
 sg13g2_buf_4 fanout5811 (.X(net5811),
    .A(net5813));
 sg13g2_buf_4 fanout5812 (.X(net5812),
    .A(net5813));
 sg13g2_buf_2 fanout5813 (.A(net5827),
    .X(net5813));
 sg13g2_buf_4 fanout5814 (.X(net5814),
    .A(net5815));
 sg13g2_buf_2 fanout5815 (.A(net5816),
    .X(net5815));
 sg13g2_buf_4 fanout5816 (.X(net5816),
    .A(net5826));
 sg13g2_buf_4 fanout5817 (.X(net5817),
    .A(net5826));
 sg13g2_buf_2 fanout5818 (.A(net5826),
    .X(net5818));
 sg13g2_buf_4 fanout5819 (.X(net5819),
    .A(net5820));
 sg13g2_buf_4 fanout5820 (.X(net5820),
    .A(net5821));
 sg13g2_buf_4 fanout5821 (.X(net5821),
    .A(net5822));
 sg13g2_buf_4 fanout5822 (.X(net5822),
    .A(net5826));
 sg13g2_buf_4 fanout5823 (.X(net5823),
    .A(net5825));
 sg13g2_buf_2 fanout5824 (.A(net5825),
    .X(net5824));
 sg13g2_buf_2 fanout5825 (.A(net5826),
    .X(net5825));
 sg13g2_buf_2 fanout5826 (.A(net5827),
    .X(net5826));
 sg13g2_buf_2 fanout5827 (.A(net5923),
    .X(net5827));
 sg13g2_buf_4 fanout5828 (.X(net5828),
    .A(net5830));
 sg13g2_buf_4 fanout5829 (.X(net5829),
    .A(net5833));
 sg13g2_buf_2 fanout5830 (.A(net5833),
    .X(net5830));
 sg13g2_buf_4 fanout5831 (.X(net5831),
    .A(net5833));
 sg13g2_buf_4 fanout5832 (.X(net5832),
    .A(net5833));
 sg13g2_buf_2 fanout5833 (.A(net5850),
    .X(net5833));
 sg13g2_buf_4 fanout5834 (.X(net5834),
    .A(net5837));
 sg13g2_buf_2 fanout5835 (.A(net5837),
    .X(net5835));
 sg13g2_buf_4 fanout5836 (.X(net5836),
    .A(net5837));
 sg13g2_buf_2 fanout5837 (.A(net5849),
    .X(net5837));
 sg13g2_buf_4 fanout5838 (.X(net5838),
    .A(net5839));
 sg13g2_buf_2 fanout5839 (.A(net5840),
    .X(net5839));
 sg13g2_buf_4 fanout5840 (.X(net5840),
    .A(net5849));
 sg13g2_buf_4 fanout5841 (.X(net5841),
    .A(net5842));
 sg13g2_buf_4 fanout5842 (.X(net5842),
    .A(net5849));
 sg13g2_buf_4 fanout5843 (.X(net5843),
    .A(net5844));
 sg13g2_buf_4 fanout5844 (.X(net5844),
    .A(net5848));
 sg13g2_buf_4 fanout5845 (.X(net5845),
    .A(net5846));
 sg13g2_buf_4 fanout5846 (.X(net5846),
    .A(net5847));
 sg13g2_buf_4 fanout5847 (.X(net5847),
    .A(net5848));
 sg13g2_buf_2 fanout5848 (.A(net5849),
    .X(net5848));
 sg13g2_buf_2 fanout5849 (.A(net5850),
    .X(net5849));
 sg13g2_buf_4 fanout5850 (.X(net5850),
    .A(net5923));
 sg13g2_buf_4 fanout5851 (.X(net5851),
    .A(net5853));
 sg13g2_buf_2 fanout5852 (.A(net5853),
    .X(net5852));
 sg13g2_buf_4 fanout5853 (.X(net5853),
    .A(net5857));
 sg13g2_buf_4 fanout5854 (.X(net5854),
    .A(net5857));
 sg13g2_buf_4 fanout5855 (.X(net5855),
    .A(net5856));
 sg13g2_buf_4 fanout5856 (.X(net5856),
    .A(net5857));
 sg13g2_buf_2 fanout5857 (.A(net5865),
    .X(net5857));
 sg13g2_buf_4 fanout5858 (.X(net5858),
    .A(net5862));
 sg13g2_buf_4 fanout5859 (.X(net5859),
    .A(net5861));
 sg13g2_buf_2 fanout5860 (.A(net5861),
    .X(net5860));
 sg13g2_buf_4 fanout5861 (.X(net5861),
    .A(net5862));
 sg13g2_buf_2 fanout5862 (.A(net5865),
    .X(net5862));
 sg13g2_buf_4 fanout5863 (.X(net5863),
    .A(net5865));
 sg13g2_buf_2 fanout5864 (.A(net5865),
    .X(net5864));
 sg13g2_buf_2 fanout5865 (.A(net5889),
    .X(net5865));
 sg13g2_buf_4 fanout5866 (.X(net5866),
    .A(net5870));
 sg13g2_buf_4 fanout5867 (.X(net5867),
    .A(net5868));
 sg13g2_buf_4 fanout5868 (.X(net5868),
    .A(net5870));
 sg13g2_buf_2 fanout5869 (.A(net5870),
    .X(net5869));
 sg13g2_buf_4 fanout5870 (.X(net5870),
    .A(net5877));
 sg13g2_buf_4 fanout5871 (.X(net5871),
    .A(net5872));
 sg13g2_buf_4 fanout5872 (.X(net5872),
    .A(net5873));
 sg13g2_buf_2 fanout5873 (.A(net5874),
    .X(net5873));
 sg13g2_buf_4 fanout5874 (.X(net5874),
    .A(net5877));
 sg13g2_buf_4 fanout5875 (.X(net5875),
    .A(net5877));
 sg13g2_buf_4 fanout5876 (.X(net5876),
    .A(net5877));
 sg13g2_buf_2 fanout5877 (.A(net5889),
    .X(net5877));
 sg13g2_buf_4 fanout5878 (.X(net5878),
    .A(net5881));
 sg13g2_buf_2 fanout5879 (.A(net5881),
    .X(net5879));
 sg13g2_buf_4 fanout5880 (.X(net5880),
    .A(net5881));
 sg13g2_buf_2 fanout5881 (.A(net5882),
    .X(net5881));
 sg13g2_buf_4 fanout5882 (.X(net5882),
    .A(net5887));
 sg13g2_buf_4 fanout5883 (.X(net5883),
    .A(net5884));
 sg13g2_buf_4 fanout5884 (.X(net5884),
    .A(net5887));
 sg13g2_buf_4 fanout5885 (.X(net5885),
    .A(net5887));
 sg13g2_buf_2 fanout5886 (.A(net5887),
    .X(net5886));
 sg13g2_buf_2 fanout5887 (.A(net5889),
    .X(net5887));
 sg13g2_buf_8 fanout5888 (.A(net5889),
    .X(net5888));
 sg13g2_buf_2 fanout5889 (.A(net5923),
    .X(net5889));
 sg13g2_buf_4 fanout5890 (.X(net5890),
    .A(net5891));
 sg13g2_buf_2 fanout5891 (.A(net5908),
    .X(net5891));
 sg13g2_buf_4 fanout5892 (.X(net5892),
    .A(net5893));
 sg13g2_buf_2 fanout5893 (.A(net5895),
    .X(net5893));
 sg13g2_buf_4 fanout5894 (.X(net5894),
    .A(net5895));
 sg13g2_buf_2 fanout5895 (.A(net5896),
    .X(net5895));
 sg13g2_buf_2 fanout5896 (.A(net5908),
    .X(net5896));
 sg13g2_buf_4 fanout5897 (.X(net5897),
    .A(net5898));
 sg13g2_buf_4 fanout5898 (.X(net5898),
    .A(net5903));
 sg13g2_buf_4 fanout5899 (.X(net5899),
    .A(net5900));
 sg13g2_buf_4 fanout5900 (.X(net5900),
    .A(net5902));
 sg13g2_buf_4 fanout5901 (.X(net5901),
    .A(net5902));
 sg13g2_buf_2 fanout5902 (.A(net5903),
    .X(net5902));
 sg13g2_buf_2 fanout5903 (.A(net5908),
    .X(net5903));
 sg13g2_buf_4 fanout5904 (.X(net5904),
    .A(net5906));
 sg13g2_buf_2 fanout5905 (.A(net5906),
    .X(net5905));
 sg13g2_buf_4 fanout5906 (.X(net5906),
    .A(net5908));
 sg13g2_buf_4 fanout5907 (.X(net5907),
    .A(net5908));
 sg13g2_buf_4 fanout5908 (.X(net5908),
    .A(net5923));
 sg13g2_buf_4 fanout5909 (.X(net5909),
    .A(net5910));
 sg13g2_buf_4 fanout5910 (.X(net5910),
    .A(net5922));
 sg13g2_buf_4 fanout5911 (.X(net5911),
    .A(net5913));
 sg13g2_buf_4 fanout5912 (.X(net5912),
    .A(net5913));
 sg13g2_buf_2 fanout5913 (.A(net5922),
    .X(net5913));
 sg13g2_buf_4 fanout5914 (.X(net5914),
    .A(net5915));
 sg13g2_buf_4 fanout5915 (.X(net5915),
    .A(net5916));
 sg13g2_buf_4 fanout5916 (.X(net5916),
    .A(net5922));
 sg13g2_buf_4 fanout5917 (.X(net5917),
    .A(net5918));
 sg13g2_buf_4 fanout5918 (.X(net5918),
    .A(net5922));
 sg13g2_buf_4 fanout5919 (.X(net5919),
    .A(net5920));
 sg13g2_buf_4 fanout5920 (.X(net5920),
    .A(net5921));
 sg13g2_buf_2 fanout5921 (.A(net5922),
    .X(net5921));
 sg13g2_buf_4 fanout5922 (.X(net5922),
    .A(net5923));
 sg13g2_buf_8 fanout5923 (.A(net6196),
    .X(net5923));
 sg13g2_buf_4 fanout5924 (.X(net5924),
    .A(net5925));
 sg13g2_buf_2 fanout5925 (.A(net5927),
    .X(net5925));
 sg13g2_buf_4 fanout5926 (.X(net5926),
    .A(net5927));
 sg13g2_buf_4 fanout5927 (.X(net5927),
    .A(net5931));
 sg13g2_buf_4 fanout5928 (.X(net5928),
    .A(net5930));
 sg13g2_buf_2 fanout5929 (.A(net5930),
    .X(net5929));
 sg13g2_buf_4 fanout5930 (.X(net5930),
    .A(net5931));
 sg13g2_buf_2 fanout5931 (.A(net5934),
    .X(net5931));
 sg13g2_buf_4 fanout5932 (.X(net5932),
    .A(net5934));
 sg13g2_buf_2 fanout5933 (.A(net5934),
    .X(net5933));
 sg13g2_buf_2 fanout5934 (.A(net5982),
    .X(net5934));
 sg13g2_buf_4 fanout5935 (.X(net5935),
    .A(net5936));
 sg13g2_buf_4 fanout5936 (.X(net5936),
    .A(net5941));
 sg13g2_buf_4 fanout5937 (.X(net5937),
    .A(net5941));
 sg13g2_buf_4 fanout5938 (.X(net5938),
    .A(net5941));
 sg13g2_buf_2 fanout5939 (.A(net5940),
    .X(net5939));
 sg13g2_buf_4 fanout5940 (.X(net5940),
    .A(net5941));
 sg13g2_buf_2 fanout5941 (.A(net5982),
    .X(net5941));
 sg13g2_buf_4 fanout5942 (.X(net5942),
    .A(net5947));
 sg13g2_buf_4 fanout5943 (.X(net5943),
    .A(net5944));
 sg13g2_buf_2 fanout5944 (.A(net5947),
    .X(net5944));
 sg13g2_buf_4 fanout5945 (.X(net5945),
    .A(net5947));
 sg13g2_buf_4 fanout5946 (.X(net5946),
    .A(net5947));
 sg13g2_buf_2 fanout5947 (.A(net5982),
    .X(net5947));
 sg13g2_buf_4 fanout5948 (.X(net5948),
    .A(net5949));
 sg13g2_buf_4 fanout5949 (.X(net5949),
    .A(net5963));
 sg13g2_buf_4 fanout5950 (.X(net5950),
    .A(net5951));
 sg13g2_buf_2 fanout5951 (.A(net5963),
    .X(net5951));
 sg13g2_buf_4 fanout5952 (.X(net5952),
    .A(net5963));
 sg13g2_buf_4 fanout5953 (.X(net5953),
    .A(net5954));
 sg13g2_buf_2 fanout5954 (.A(net5956),
    .X(net5954));
 sg13g2_buf_4 fanout5955 (.X(net5955),
    .A(net5956));
 sg13g2_buf_2 fanout5956 (.A(net5962),
    .X(net5956));
 sg13g2_buf_4 fanout5957 (.X(net5957),
    .A(net5958));
 sg13g2_buf_4 fanout5958 (.X(net5958),
    .A(net5960));
 sg13g2_buf_4 fanout5959 (.X(net5959),
    .A(net5960));
 sg13g2_buf_2 fanout5960 (.A(net5961),
    .X(net5960));
 sg13g2_buf_4 fanout5961 (.X(net5961),
    .A(net5962));
 sg13g2_buf_4 fanout5962 (.X(net5962),
    .A(net5963));
 sg13g2_buf_2 fanout5963 (.A(net5981),
    .X(net5963));
 sg13g2_buf_4 fanout5964 (.X(net5964),
    .A(net5965));
 sg13g2_buf_4 fanout5965 (.X(net5965),
    .A(net5973));
 sg13g2_buf_4 fanout5966 (.X(net5966),
    .A(net5967));
 sg13g2_buf_2 fanout5967 (.A(net5973),
    .X(net5967));
 sg13g2_buf_4 fanout5968 (.X(net5968),
    .A(net5969));
 sg13g2_buf_4 fanout5969 (.X(net5969),
    .A(net5972));
 sg13g2_buf_4 fanout5970 (.X(net5970),
    .A(net5972));
 sg13g2_buf_4 fanout5971 (.X(net5971),
    .A(net5972));
 sg13g2_buf_2 fanout5972 (.A(net5973),
    .X(net5972));
 sg13g2_buf_2 fanout5973 (.A(net5981),
    .X(net5973));
 sg13g2_buf_4 fanout5974 (.X(net5974),
    .A(net5979));
 sg13g2_buf_4 fanout5975 (.X(net5975),
    .A(net5979));
 sg13g2_buf_4 fanout5976 (.X(net5976),
    .A(net5977));
 sg13g2_buf_2 fanout5977 (.A(net5979),
    .X(net5977));
 sg13g2_buf_4 fanout5978 (.X(net5978),
    .A(net5979));
 sg13g2_buf_2 fanout5979 (.A(net5981),
    .X(net5979));
 sg13g2_buf_4 fanout5980 (.X(net5980),
    .A(net5981));
 sg13g2_buf_2 fanout5981 (.A(net5982),
    .X(net5981));
 sg13g2_buf_2 fanout5982 (.A(net6196),
    .X(net5982));
 sg13g2_buf_4 fanout5983 (.X(net5983),
    .A(net5984));
 sg13g2_buf_4 fanout5984 (.X(net5984),
    .A(net5987));
 sg13g2_buf_4 fanout5985 (.X(net5985),
    .A(net5986));
 sg13g2_buf_4 fanout5986 (.X(net5986),
    .A(net5987));
 sg13g2_buf_2 fanout5987 (.A(net5993),
    .X(net5987));
 sg13g2_buf_4 fanout5988 (.X(net5988),
    .A(net5989));
 sg13g2_buf_4 fanout5989 (.X(net5989),
    .A(net5993));
 sg13g2_buf_4 fanout5990 (.X(net5990),
    .A(net5992));
 sg13g2_buf_2 fanout5991 (.A(net5992),
    .X(net5991));
 sg13g2_buf_2 fanout5992 (.A(net5993),
    .X(net5992));
 sg13g2_buf_2 fanout5993 (.A(net6065),
    .X(net5993));
 sg13g2_buf_4 fanout5994 (.X(net5994),
    .A(net6001));
 sg13g2_buf_4 fanout5995 (.X(net5995),
    .A(net6001));
 sg13g2_buf_4 fanout5996 (.X(net5996),
    .A(net5997));
 sg13g2_buf_2 fanout5997 (.A(net6001),
    .X(net5997));
 sg13g2_buf_4 fanout5998 (.X(net5998),
    .A(net6000));
 sg13g2_buf_4 fanout5999 (.X(net5999),
    .A(net6000));
 sg13g2_buf_4 fanout6000 (.X(net6000),
    .A(net6001));
 sg13g2_buf_2 fanout6001 (.A(net6065),
    .X(net6001));
 sg13g2_buf_4 fanout6002 (.X(net6002),
    .A(net6003));
 sg13g2_buf_2 fanout6003 (.A(net6004),
    .X(net6003));
 sg13g2_buf_2 fanout6004 (.A(net6010),
    .X(net6004));
 sg13g2_buf_4 fanout6005 (.X(net6005),
    .A(net6006));
 sg13g2_buf_2 fanout6006 (.A(net6009),
    .X(net6006));
 sg13g2_buf_4 fanout6007 (.X(net6007),
    .A(net6008));
 sg13g2_buf_2 fanout6008 (.A(net6009),
    .X(net6008));
 sg13g2_buf_2 fanout6009 (.A(net6010),
    .X(net6009));
 sg13g2_buf_2 fanout6010 (.A(net6065),
    .X(net6010));
 sg13g2_buf_4 fanout6011 (.X(net6011),
    .A(net6015));
 sg13g2_buf_4 fanout6012 (.X(net6012),
    .A(net6013));
 sg13g2_buf_2 fanout6013 (.A(net6014),
    .X(net6013));
 sg13g2_buf_4 fanout6014 (.X(net6014),
    .A(net6015));
 sg13g2_buf_2 fanout6015 (.A(net6064),
    .X(net6015));
 sg13g2_buf_4 fanout6016 (.X(net6016),
    .A(net6021));
 sg13g2_buf_2 fanout6017 (.A(net6021),
    .X(net6017));
 sg13g2_buf_4 fanout6018 (.X(net6018),
    .A(net6021));
 sg13g2_buf_4 fanout6019 (.X(net6019),
    .A(net6020));
 sg13g2_buf_2 fanout6020 (.A(net6021),
    .X(net6020));
 sg13g2_buf_2 fanout6021 (.A(net6064),
    .X(net6021));
 sg13g2_buf_4 fanout6022 (.X(net6022),
    .A(net6023));
 sg13g2_buf_2 fanout6023 (.A(net6024),
    .X(net6023));
 sg13g2_buf_2 fanout6024 (.A(net6033),
    .X(net6024));
 sg13g2_buf_4 fanout6025 (.X(net6025),
    .A(net6026));
 sg13g2_buf_2 fanout6026 (.A(net6033),
    .X(net6026));
 sg13g2_buf_4 fanout6027 (.X(net6027),
    .A(net6028));
 sg13g2_buf_4 fanout6028 (.X(net6028),
    .A(net6033));
 sg13g2_buf_4 fanout6029 (.X(net6029),
    .A(net6030));
 sg13g2_buf_2 fanout6030 (.A(net6032),
    .X(net6030));
 sg13g2_buf_4 fanout6031 (.X(net6031),
    .A(net6032));
 sg13g2_buf_2 fanout6032 (.A(net6033),
    .X(net6032));
 sg13g2_buf_2 fanout6033 (.A(net6064),
    .X(net6033));
 sg13g2_buf_4 fanout6034 (.X(net6034),
    .A(net6036));
 sg13g2_buf_4 fanout6035 (.X(net6035),
    .A(net6036));
 sg13g2_buf_2 fanout6036 (.A(net6037),
    .X(net6036));
 sg13g2_buf_4 fanout6037 (.X(net6037),
    .A(net6047));
 sg13g2_buf_4 fanout6038 (.X(net6038),
    .A(net6040));
 sg13g2_buf_2 fanout6039 (.A(net6040),
    .X(net6039));
 sg13g2_buf_2 fanout6040 (.A(net6047),
    .X(net6040));
 sg13g2_buf_4 fanout6041 (.X(net6041),
    .A(net6043));
 sg13g2_buf_2 fanout6042 (.A(net6043),
    .X(net6042));
 sg13g2_buf_4 fanout6043 (.X(net6043),
    .A(net6045));
 sg13g2_buf_4 fanout6044 (.X(net6044),
    .A(net6045));
 sg13g2_buf_2 fanout6045 (.A(net6046),
    .X(net6045));
 sg13g2_buf_4 fanout6046 (.X(net6046),
    .A(net6047));
 sg13g2_buf_2 fanout6047 (.A(net6064),
    .X(net6047));
 sg13g2_buf_4 fanout6048 (.X(net6048),
    .A(net6063));
 sg13g2_buf_2 fanout6049 (.A(net6063),
    .X(net6049));
 sg13g2_buf_4 fanout6050 (.X(net6050),
    .A(net6051));
 sg13g2_buf_4 fanout6051 (.X(net6051),
    .A(net6063));
 sg13g2_buf_4 fanout6052 (.X(net6052),
    .A(net6053));
 sg13g2_buf_4 fanout6053 (.X(net6053),
    .A(net6057));
 sg13g2_buf_4 fanout6054 (.X(net6054),
    .A(net6057));
 sg13g2_buf_4 fanout6055 (.X(net6055),
    .A(net6056));
 sg13g2_buf_4 fanout6056 (.X(net6056),
    .A(net6057));
 sg13g2_buf_4 fanout6057 (.X(net6057),
    .A(net6063));
 sg13g2_buf_4 fanout6058 (.X(net6058),
    .A(net6059));
 sg13g2_buf_4 fanout6059 (.X(net6059),
    .A(net6062));
 sg13g2_buf_4 fanout6060 (.X(net6060),
    .A(net6061));
 sg13g2_buf_4 fanout6061 (.X(net6061),
    .A(net6062));
 sg13g2_buf_2 fanout6062 (.A(net6063),
    .X(net6062));
 sg13g2_buf_2 fanout6063 (.A(net6064),
    .X(net6063));
 sg13g2_buf_2 fanout6064 (.A(net6065),
    .X(net6064));
 sg13g2_buf_2 fanout6065 (.A(net6196),
    .X(net6065));
 sg13g2_buf_4 fanout6066 (.X(net6066),
    .A(net6068));
 sg13g2_buf_4 fanout6067 (.X(net6067),
    .A(net6068));
 sg13g2_buf_4 fanout6068 (.X(net6068),
    .A(net6072));
 sg13g2_buf_4 fanout6069 (.X(net6069),
    .A(net6070));
 sg13g2_buf_4 fanout6070 (.X(net6070),
    .A(net6071));
 sg13g2_buf_4 fanout6071 (.X(net6071),
    .A(net6072));
 sg13g2_buf_2 fanout6072 (.A(net6087),
    .X(net6072));
 sg13g2_buf_4 fanout6073 (.X(net6073),
    .A(net6074));
 sg13g2_buf_2 fanout6074 (.A(net6075),
    .X(net6074));
 sg13g2_buf_4 fanout6075 (.X(net6075),
    .A(net6078));
 sg13g2_buf_4 fanout6076 (.X(net6076),
    .A(net6077));
 sg13g2_buf_2 fanout6077 (.A(net6078),
    .X(net6077));
 sg13g2_buf_2 fanout6078 (.A(net6087),
    .X(net6078));
 sg13g2_buf_4 fanout6079 (.X(net6079),
    .A(net6080));
 sg13g2_buf_4 fanout6080 (.X(net6080),
    .A(net6083));
 sg13g2_buf_4 fanout6081 (.X(net6081),
    .A(net6082));
 sg13g2_buf_2 fanout6082 (.A(net6083),
    .X(net6082));
 sg13g2_buf_2 fanout6083 (.A(net6087),
    .X(net6083));
 sg13g2_buf_4 fanout6084 (.X(net6084),
    .A(net6085));
 sg13g2_buf_4 fanout6085 (.X(net6085),
    .A(net6086));
 sg13g2_buf_4 fanout6086 (.X(net6086),
    .A(net6087));
 sg13g2_buf_2 fanout6087 (.A(net6132),
    .X(net6087));
 sg13g2_buf_4 fanout6088 (.X(net6088),
    .A(net6089));
 sg13g2_buf_4 fanout6089 (.X(net6089),
    .A(net6090));
 sg13g2_buf_4 fanout6090 (.X(net6090),
    .A(net6132));
 sg13g2_buf_4 fanout6091 (.X(net6091),
    .A(net6092));
 sg13g2_buf_4 fanout6092 (.X(net6092),
    .A(net6093));
 sg13g2_buf_2 fanout6093 (.A(net6103),
    .X(net6093));
 sg13g2_buf_4 fanout6094 (.X(net6094),
    .A(net6095));
 sg13g2_buf_4 fanout6095 (.X(net6095),
    .A(net6096));
 sg13g2_buf_4 fanout6096 (.X(net6096),
    .A(net6103));
 sg13g2_buf_4 fanout6097 (.X(net6097),
    .A(net6098));
 sg13g2_buf_4 fanout6098 (.X(net6098),
    .A(net6100));
 sg13g2_buf_2 fanout6099 (.A(net6100),
    .X(net6099));
 sg13g2_buf_2 fanout6100 (.A(net6103),
    .X(net6100));
 sg13g2_buf_4 fanout6101 (.X(net6101),
    .A(net6103));
 sg13g2_buf_2 fanout6102 (.A(net6103),
    .X(net6102));
 sg13g2_buf_2 fanout6103 (.A(net6132),
    .X(net6103));
 sg13g2_buf_4 fanout6104 (.X(net6104),
    .A(net6105));
 sg13g2_buf_2 fanout6105 (.A(net6106),
    .X(net6105));
 sg13g2_buf_2 fanout6106 (.A(net6107),
    .X(net6106));
 sg13g2_buf_2 fanout6107 (.A(net6108),
    .X(net6107));
 sg13g2_buf_4 fanout6108 (.X(net6108),
    .A(net6118));
 sg13g2_buf_4 fanout6109 (.X(net6109),
    .A(net6111));
 sg13g2_buf_4 fanout6110 (.X(net6110),
    .A(net6111));
 sg13g2_buf_2 fanout6111 (.A(net6112),
    .X(net6111));
 sg13g2_buf_4 fanout6112 (.X(net6112),
    .A(net6115));
 sg13g2_buf_4 fanout6113 (.X(net6113),
    .A(net6115));
 sg13g2_buf_2 fanout6114 (.A(net6115),
    .X(net6114));
 sg13g2_buf_2 fanout6115 (.A(net6118),
    .X(net6115));
 sg13g2_buf_4 fanout6116 (.X(net6116),
    .A(net6117));
 sg13g2_buf_2 fanout6117 (.A(net6118),
    .X(net6117));
 sg13g2_buf_2 fanout6118 (.A(net6132),
    .X(net6118));
 sg13g2_buf_4 fanout6119 (.X(net6119),
    .A(net6120));
 sg13g2_buf_4 fanout6120 (.X(net6120),
    .A(net6121));
 sg13g2_buf_4 fanout6121 (.X(net6121),
    .A(net6131));
 sg13g2_buf_4 fanout6122 (.X(net6122),
    .A(net6124));
 sg13g2_buf_2 fanout6123 (.A(net6124),
    .X(net6123));
 sg13g2_buf_2 fanout6124 (.A(net6127),
    .X(net6124));
 sg13g2_buf_4 fanout6125 (.X(net6125),
    .A(net6126));
 sg13g2_buf_2 fanout6126 (.A(net6127),
    .X(net6126));
 sg13g2_buf_2 fanout6127 (.A(net6128),
    .X(net6127));
 sg13g2_buf_4 fanout6128 (.X(net6128),
    .A(net6131));
 sg13g2_buf_4 fanout6129 (.X(net6129),
    .A(net6131));
 sg13g2_buf_4 fanout6130 (.X(net6130),
    .A(net6131));
 sg13g2_buf_2 fanout6131 (.A(net6132),
    .X(net6131));
 sg13g2_buf_4 fanout6132 (.X(net6132),
    .A(net6195));
 sg13g2_buf_4 fanout6133 (.X(net6133),
    .A(net6138));
 sg13g2_buf_4 fanout6134 (.X(net6134),
    .A(net6138));
 sg13g2_buf_4 fanout6135 (.X(net6135),
    .A(net6136));
 sg13g2_buf_4 fanout6136 (.X(net6136),
    .A(net6137));
 sg13g2_buf_4 fanout6137 (.X(net6137),
    .A(net6138));
 sg13g2_buf_4 fanout6138 (.X(net6138),
    .A(net6142));
 sg13g2_buf_4 fanout6139 (.X(net6139),
    .A(net6140));
 sg13g2_buf_2 fanout6140 (.A(net6142),
    .X(net6140));
 sg13g2_buf_4 fanout6141 (.X(net6141),
    .A(net6142));
 sg13g2_buf_2 fanout6142 (.A(net6158),
    .X(net6142));
 sg13g2_buf_4 fanout6143 (.X(net6143),
    .A(net6147));
 sg13g2_buf_4 fanout6144 (.X(net6144),
    .A(net6146));
 sg13g2_buf_4 fanout6145 (.X(net6145),
    .A(net6146));
 sg13g2_buf_2 fanout6146 (.A(net6147),
    .X(net6146));
 sg13g2_buf_2 fanout6147 (.A(net6158),
    .X(net6147));
 sg13g2_buf_4 fanout6148 (.X(net6148),
    .A(net6150));
 sg13g2_buf_2 fanout6149 (.A(net6150),
    .X(net6149));
 sg13g2_buf_2 fanout6150 (.A(net6151),
    .X(net6150));
 sg13g2_buf_2 fanout6151 (.A(net6158),
    .X(net6151));
 sg13g2_buf_4 fanout6152 (.X(net6152),
    .A(net6157));
 sg13g2_buf_4 fanout6153 (.X(net6153),
    .A(net6154));
 sg13g2_buf_2 fanout6154 (.A(net6157),
    .X(net6154));
 sg13g2_buf_4 fanout6155 (.X(net6155),
    .A(net6156));
 sg13g2_buf_4 fanout6156 (.X(net6156),
    .A(net6157));
 sg13g2_buf_2 fanout6157 (.A(net6158),
    .X(net6157));
 sg13g2_buf_2 fanout6158 (.A(net6195),
    .X(net6158));
 sg13g2_buf_4 fanout6159 (.X(net6159),
    .A(net6160));
 sg13g2_buf_2 fanout6160 (.A(net6161),
    .X(net6160));
 sg13g2_buf_2 fanout6161 (.A(net6167),
    .X(net6161));
 sg13g2_buf_4 fanout6162 (.X(net6162),
    .A(net6163));
 sg13g2_buf_2 fanout6163 (.A(net6164),
    .X(net6163));
 sg13g2_buf_2 fanout6164 (.A(net6167),
    .X(net6164));
 sg13g2_buf_4 fanout6165 (.X(net6165),
    .A(net6167));
 sg13g2_buf_4 fanout6166 (.X(net6166),
    .A(net6167));
 sg13g2_buf_2 fanout6167 (.A(net6172),
    .X(net6167));
 sg13g2_buf_4 fanout6168 (.X(net6168),
    .A(net6170));
 sg13g2_buf_2 fanout6169 (.A(net6170),
    .X(net6169));
 sg13g2_buf_2 fanout6170 (.A(net6172),
    .X(net6170));
 sg13g2_buf_4 fanout6171 (.X(net6171),
    .A(net6172));
 sg13g2_buf_2 fanout6172 (.A(net6195),
    .X(net6172));
 sg13g2_buf_4 fanout6173 (.X(net6173),
    .A(net6193));
 sg13g2_buf_4 fanout6174 (.X(net6174),
    .A(net6175));
 sg13g2_buf_2 fanout6175 (.A(net6176),
    .X(net6175));
 sg13g2_buf_2 fanout6176 (.A(net6177),
    .X(net6176));
 sg13g2_buf_2 fanout6177 (.A(net6193),
    .X(net6177));
 sg13g2_buf_4 fanout6178 (.X(net6178),
    .A(net6184));
 sg13g2_buf_4 fanout6179 (.X(net6179),
    .A(net6184));
 sg13g2_buf_4 fanout6180 (.X(net6180),
    .A(net6184));
 sg13g2_buf_4 fanout6181 (.X(net6181),
    .A(net6184));
 sg13g2_buf_4 fanout6182 (.X(net6182),
    .A(net6183));
 sg13g2_buf_4 fanout6183 (.X(net6183),
    .A(net6184));
 sg13g2_buf_2 fanout6184 (.A(net6192),
    .X(net6184));
 sg13g2_buf_4 fanout6185 (.X(net6185),
    .A(net6186));
 sg13g2_buf_4 fanout6186 (.X(net6186),
    .A(net6189));
 sg13g2_buf_4 fanout6187 (.X(net6187),
    .A(net6189));
 sg13g2_buf_2 fanout6188 (.A(net6189),
    .X(net6188));
 sg13g2_buf_2 fanout6189 (.A(net6192),
    .X(net6189));
 sg13g2_buf_4 fanout6190 (.X(net6190),
    .A(net6192));
 sg13g2_buf_4 fanout6191 (.X(net6191),
    .A(net6192));
 sg13g2_buf_2 fanout6192 (.A(net6193),
    .X(net6192));
 sg13g2_buf_2 fanout6193 (.A(net6194),
    .X(net6193));
 sg13g2_buf_4 fanout6194 (.X(net6194),
    .A(net6195));
 sg13g2_buf_2 fanout6195 (.A(net6196),
    .X(net6195));
 sg13g2_buf_8 fanout6196 (.A(rst_n),
    .X(net6196));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ui_in[2]));
 sg13g2_buf_2 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_8 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_16 input4 (.X(net4),
    .A(ui_in[5]));
 sg13g2_buf_8 input5 (.A(uio_in[4]),
    .X(net5));
 sg13g2_tielo tt_um_supermic_arghunter_6 (.L_LO(net6));
 sg13g2_antennanp ANTENNA_2 (.A(rst_n));
 sg13g2_antennanp ANTENNA_3 (.A(rst_n));
 sg13g2_antennanp ANTENNA_4 (.A(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_antennanp ANTENNA_5 (.A(\u_supermic_top_module.i2s_bus_inst[6].c_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_antennanp ANTENNA_6 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_7 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_8 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_9 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_10 (.A(uio_in[1]));
 sg13g2_antennanp ANTENNA_11 (.A(uio_in[1]));
 sg13g2_antennanp ANTENNA_12 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_13 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_14 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_15 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_16 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_17 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_18 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_19 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_20 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_21 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_22 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_23 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_24 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_25 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_26 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_27 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_28 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_29 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_30 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_31 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_32 (.A(net4870));
 sg13g2_antennanp ANTENNA_33 (.A(net4870));
 sg13g2_antennanp ANTENNA_34 (.A(net4870));
 sg13g2_antennanp ANTENNA_35 (.A(net4870));
 sg13g2_antennanp ANTENNA_36 (.A(net4870));
 sg13g2_antennanp ANTENNA_37 (.A(net4870));
 sg13g2_antennanp ANTENNA_38 (.A(net4870));
 sg13g2_antennanp ANTENNA_39 (.A(net4870));
 sg13g2_antennanp ANTENNA_40 (.A(net4870));
 sg13g2_antennanp ANTENNA_41 (.A(net4870));
 sg13g2_antennanp ANTENNA_42 (.A(net4870));
 sg13g2_antennanp ANTENNA_43 (.A(net4870));
 sg13g2_antennanp ANTENNA_44 (.A(net4870));
 sg13g2_antennanp ANTENNA_45 (.A(net4870));
 sg13g2_antennanp ANTENNA_46 (.A(net4870));
 sg13g2_antennanp ANTENNA_47 (.A(net4870));
 sg13g2_antennanp ANTENNA_48 (.A(net4870));
 sg13g2_antennanp ANTENNA_49 (.A(net4870));
 sg13g2_antennanp ANTENNA_50 (.A(net4870));
 sg13g2_antennanp ANTENNA_51 (.A(net4870));
 sg13g2_antennanp ANTENNA_52 (.A(net4870));
 sg13g2_antennanp ANTENNA_53 (.A(net4870));
 sg13g2_antennanp ANTENNA_54 (.A(net4870));
 sg13g2_antennanp ANTENNA_55 (.A(net4870));
 sg13g2_antennanp ANTENNA_56 (.A(net4870));
 sg13g2_antennanp ANTENNA_57 (.A(net4870));
 sg13g2_antennanp ANTENNA_58 (.A(net4870));
 sg13g2_antennanp ANTENNA_59 (.A(net4870));
 sg13g2_antennanp ANTENNA_60 (.A(net4870));
 sg13g2_antennanp ANTENNA_61 (.A(net4870));
 sg13g2_antennanp ANTENNA_62 (.A(net4870));
 sg13g2_antennanp ANTENNA_63 (.A(net4870));
 sg13g2_antennanp ANTENNA_64 (.A(net4870));
 sg13g2_antennanp ANTENNA_65 (.A(net4870));
 sg13g2_antennanp ANTENNA_66 (.A(net5175));
 sg13g2_antennanp ANTENNA_67 (.A(net5175));
 sg13g2_antennanp ANTENNA_68 (.A(net5175));
 sg13g2_antennanp ANTENNA_69 (.A(net5175));
 sg13g2_antennanp ANTENNA_70 (.A(net5280));
 sg13g2_antennanp ANTENNA_71 (.A(net5280));
 sg13g2_antennanp ANTENNA_72 (.A(net5280));
 sg13g2_antennanp ANTENNA_73 (.A(net5280));
 sg13g2_antennanp ANTENNA_74 (.A(net5280));
 sg13g2_antennanp ANTENNA_75 (.A(net5280));
 sg13g2_antennanp ANTENNA_76 (.A(net5280));
 sg13g2_antennanp ANTENNA_77 (.A(net5280));
 sg13g2_antennanp ANTENNA_78 (.A(net4));
 sg13g2_antennanp ANTENNA_79 (.A(net4));
 sg13g2_antennanp ANTENNA_80 (.A(net4));
 sg13g2_antennanp ANTENNA_81 (.A(net4));
 sg13g2_antennanp ANTENNA_82 (.A(net4));
 sg13g2_antennanp ANTENNA_83 (.A(net4));
 sg13g2_antennanp ANTENNA_84 (.A(net4));
 sg13g2_antennanp ANTENNA_85 (.A(net4));
 sg13g2_antennanp ANTENNA_86 (.A(_00627_));
 sg13g2_antennanp ANTENNA_87 (.A(rst_n));
 sg13g2_antennanp ANTENNA_88 (.A(rst_n));
 sg13g2_antennanp ANTENNA_89 (.A(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_antennanp ANTENNA_90 (.A(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_antennanp ANTENNA_91 (.A(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_antennanp ANTENNA_92 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_93 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_94 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_95 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_96 (.A(uio_in[1]));
 sg13g2_antennanp ANTENNA_97 (.A(uio_in[1]));
 sg13g2_antennanp ANTENNA_98 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_99 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_100 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_101 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_102 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_103 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_104 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_105 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_106 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_107 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_108 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_109 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_110 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_111 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_112 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_113 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_114 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_115 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_116 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_117 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_118 (.A(net5175));
 sg13g2_antennanp ANTENNA_119 (.A(net5175));
 sg13g2_antennanp ANTENNA_120 (.A(net5175));
 sg13g2_antennanp ANTENNA_121 (.A(net5175));
 sg13g2_antennanp ANTENNA_122 (.A(net5280));
 sg13g2_antennanp ANTENNA_123 (.A(net5280));
 sg13g2_antennanp ANTENNA_124 (.A(net5280));
 sg13g2_antennanp ANTENNA_125 (.A(net5280));
 sg13g2_antennanp ANTENNA_126 (.A(net5280));
 sg13g2_antennanp ANTENNA_127 (.A(net5280));
 sg13g2_antennanp ANTENNA_128 (.A(net5280));
 sg13g2_antennanp ANTENNA_129 (.A(net5280));
 sg13g2_antennanp ANTENNA_130 (.A(net5280));
 sg13g2_antennanp ANTENNA_131 (.A(net5280));
 sg13g2_antennanp ANTENNA_132 (.A(net5280));
 sg13g2_antennanp ANTENNA_133 (.A(net5280));
 sg13g2_antennanp ANTENNA_134 (.A(net1));
 sg13g2_antennanp ANTENNA_135 (.A(net1));
 sg13g2_antennanp ANTENNA_136 (.A(net1));
 sg13g2_antennanp ANTENNA_137 (.A(net1));
 sg13g2_antennanp ANTENNA_138 (.A(net4));
 sg13g2_antennanp ANTENNA_139 (.A(net4));
 sg13g2_antennanp ANTENNA_140 (.A(net4));
 sg13g2_antennanp ANTENNA_141 (.A(net4));
 sg13g2_antennanp ANTENNA_142 (.A(net4));
 sg13g2_antennanp ANTENNA_143 (.A(rst_n));
 sg13g2_antennanp ANTENNA_144 (.A(rst_n));
 sg13g2_antennanp ANTENNA_145 (.A(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_antennanp ANTENNA_146 (.A(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_antennanp ANTENNA_147 (.A(\u_supermic_top_module.i2s_bus_inst[4].c_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_antennanp ANTENNA_148 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_149 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_150 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_151 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_152 (.A(uio_in[1]));
 sg13g2_antennanp ANTENNA_153 (.A(uio_in[1]));
 sg13g2_antennanp ANTENNA_154 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_155 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_156 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_157 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_158 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_159 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_160 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_161 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_162 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_163 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_164 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_165 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_166 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_167 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_168 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_169 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_170 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_171 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_172 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_173 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_174 (.A(net5175));
 sg13g2_antennanp ANTENNA_175 (.A(net5175));
 sg13g2_antennanp ANTENNA_176 (.A(net5175));
 sg13g2_antennanp ANTENNA_177 (.A(net5175));
 sg13g2_antennanp ANTENNA_178 (.A(net1));
 sg13g2_antennanp ANTENNA_179 (.A(net1));
 sg13g2_antennanp ANTENNA_180 (.A(net1));
 sg13g2_antennanp ANTENNA_181 (.A(net1));
 sg13g2_antennanp ANTENNA_182 (.A(net4));
 sg13g2_antennanp ANTENNA_183 (.A(net4));
 sg13g2_antennanp ANTENNA_184 (.A(net4));
 sg13g2_antennanp ANTENNA_185 (.A(net4));
 sg13g2_antennanp ANTENNA_186 (.A(net4));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_4 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_635 ();
 sg13g2_decap_8 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_649 ();
 sg13g2_decap_8 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_663 ();
 sg13g2_fill_2 FILLER_0_670 ();
 sg13g2_fill_1 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_680 ();
 sg13g2_fill_2 FILLER_0_687 ();
 sg13g2_fill_2 FILLER_0_705 ();
 sg13g2_fill_2 FILLER_0_722 ();
 sg13g2_decap_8 FILLER_0_732 ();
 sg13g2_decap_8 FILLER_0_739 ();
 sg13g2_decap_4 FILLER_0_746 ();
 sg13g2_fill_2 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_778 ();
 sg13g2_decap_8 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_fill_2 FILLER_0_799 ();
 sg13g2_decap_4 FILLER_0_814 ();
 sg13g2_decap_8 FILLER_0_844 ();
 sg13g2_decap_8 FILLER_0_851 ();
 sg13g2_decap_4 FILLER_0_858 ();
 sg13g2_fill_1 FILLER_0_862 ();
 sg13g2_fill_2 FILLER_0_889 ();
 sg13g2_fill_1 FILLER_0_891 ();
 sg13g2_decap_4 FILLER_0_918 ();
 sg13g2_fill_2 FILLER_0_922 ();
 sg13g2_decap_8 FILLER_0_937 ();
 sg13g2_decap_8 FILLER_0_944 ();
 sg13g2_decap_8 FILLER_0_951 ();
 sg13g2_decap_8 FILLER_0_958 ();
 sg13g2_decap_8 FILLER_0_965 ();
 sg13g2_decap_8 FILLER_0_972 ();
 sg13g2_decap_8 FILLER_0_979 ();
 sg13g2_fill_2 FILLER_0_986 ();
 sg13g2_decap_8 FILLER_0_993 ();
 sg13g2_decap_8 FILLER_0_1000 ();
 sg13g2_decap_8 FILLER_0_1007 ();
 sg13g2_decap_8 FILLER_0_1014 ();
 sg13g2_decap_8 FILLER_0_1021 ();
 sg13g2_decap_8 FILLER_0_1028 ();
 sg13g2_decap_8 FILLER_0_1035 ();
 sg13g2_decap_8 FILLER_0_1042 ();
 sg13g2_decap_8 FILLER_0_1049 ();
 sg13g2_decap_8 FILLER_0_1056 ();
 sg13g2_decap_8 FILLER_0_1063 ();
 sg13g2_decap_8 FILLER_0_1070 ();
 sg13g2_decap_8 FILLER_0_1077 ();
 sg13g2_decap_8 FILLER_0_1084 ();
 sg13g2_decap_8 FILLER_0_1091 ();
 sg13g2_decap_8 FILLER_0_1098 ();
 sg13g2_decap_8 FILLER_0_1105 ();
 sg13g2_decap_8 FILLER_0_1112 ();
 sg13g2_decap_8 FILLER_0_1119 ();
 sg13g2_decap_8 FILLER_0_1126 ();
 sg13g2_decap_8 FILLER_0_1133 ();
 sg13g2_decap_8 FILLER_0_1140 ();
 sg13g2_decap_8 FILLER_0_1147 ();
 sg13g2_decap_8 FILLER_0_1154 ();
 sg13g2_decap_8 FILLER_0_1161 ();
 sg13g2_decap_8 FILLER_0_1168 ();
 sg13g2_decap_8 FILLER_0_1175 ();
 sg13g2_decap_8 FILLER_0_1182 ();
 sg13g2_decap_8 FILLER_0_1189 ();
 sg13g2_decap_8 FILLER_0_1196 ();
 sg13g2_decap_8 FILLER_0_1203 ();
 sg13g2_decap_8 FILLER_0_1210 ();
 sg13g2_decap_8 FILLER_0_1217 ();
 sg13g2_fill_2 FILLER_0_1251 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_fill_2 FILLER_0_1281 ();
 sg13g2_decap_8 FILLER_0_1291 ();
 sg13g2_decap_8 FILLER_0_1298 ();
 sg13g2_decap_8 FILLER_0_1305 ();
 sg13g2_decap_8 FILLER_0_1312 ();
 sg13g2_decap_8 FILLER_0_1319 ();
 sg13g2_decap_8 FILLER_0_1326 ();
 sg13g2_decap_8 FILLER_0_1333 ();
 sg13g2_fill_2 FILLER_0_1353 ();
 sg13g2_decap_8 FILLER_0_1360 ();
 sg13g2_fill_2 FILLER_0_1367 ();
 sg13g2_decap_8 FILLER_0_1399 ();
 sg13g2_decap_8 FILLER_0_1406 ();
 sg13g2_decap_4 FILLER_0_1413 ();
 sg13g2_fill_1 FILLER_0_1417 ();
 sg13g2_fill_2 FILLER_0_1427 ();
 sg13g2_decap_8 FILLER_0_1437 ();
 sg13g2_decap_8 FILLER_0_1444 ();
 sg13g2_decap_4 FILLER_0_1451 ();
 sg13g2_fill_2 FILLER_0_1455 ();
 sg13g2_fill_1 FILLER_0_1483 ();
 sg13g2_decap_8 FILLER_0_1502 ();
 sg13g2_decap_8 FILLER_0_1509 ();
 sg13g2_decap_8 FILLER_0_1516 ();
 sg13g2_decap_8 FILLER_0_1523 ();
 sg13g2_decap_8 FILLER_0_1530 ();
 sg13g2_decap_8 FILLER_0_1537 ();
 sg13g2_fill_1 FILLER_0_1544 ();
 sg13g2_decap_8 FILLER_0_1560 ();
 sg13g2_decap_8 FILLER_0_1567 ();
 sg13g2_decap_8 FILLER_0_1574 ();
 sg13g2_decap_8 FILLER_0_1581 ();
 sg13g2_decap_8 FILLER_0_1588 ();
 sg13g2_decap_8 FILLER_0_1608 ();
 sg13g2_fill_1 FILLER_0_1615 ();
 sg13g2_decap_8 FILLER_0_1642 ();
 sg13g2_decap_8 FILLER_0_1649 ();
 sg13g2_decap_8 FILLER_0_1656 ();
 sg13g2_decap_4 FILLER_0_1663 ();
 sg13g2_fill_2 FILLER_0_1667 ();
 sg13g2_fill_2 FILLER_0_1673 ();
 sg13g2_fill_1 FILLER_0_1675 ();
 sg13g2_decap_8 FILLER_0_1689 ();
 sg13g2_decap_8 FILLER_0_1696 ();
 sg13g2_decap_8 FILLER_0_1717 ();
 sg13g2_decap_8 FILLER_0_1724 ();
 sg13g2_decap_8 FILLER_0_1731 ();
 sg13g2_decap_8 FILLER_0_1738 ();
 sg13g2_decap_8 FILLER_0_1745 ();
 sg13g2_decap_4 FILLER_0_1752 ();
 sg13g2_fill_1 FILLER_0_1756 ();
 sg13g2_decap_8 FILLER_0_1790 ();
 sg13g2_decap_8 FILLER_0_1797 ();
 sg13g2_decap_8 FILLER_0_1804 ();
 sg13g2_decap_8 FILLER_0_1811 ();
 sg13g2_decap_4 FILLER_0_1818 ();
 sg13g2_decap_8 FILLER_0_1871 ();
 sg13g2_fill_1 FILLER_0_1878 ();
 sg13g2_fill_2 FILLER_0_1887 ();
 sg13g2_fill_1 FILLER_0_1909 ();
 sg13g2_decap_8 FILLER_0_1936 ();
 sg13g2_decap_8 FILLER_0_1943 ();
 sg13g2_decap_8 FILLER_0_1950 ();
 sg13g2_decap_8 FILLER_0_1957 ();
 sg13g2_decap_8 FILLER_0_1964 ();
 sg13g2_decap_8 FILLER_0_1971 ();
 sg13g2_decap_8 FILLER_0_1978 ();
 sg13g2_decap_8 FILLER_0_1985 ();
 sg13g2_decap_8 FILLER_0_1992 ();
 sg13g2_decap_8 FILLER_0_1999 ();
 sg13g2_decap_8 FILLER_0_2006 ();
 sg13g2_fill_2 FILLER_0_2013 ();
 sg13g2_decap_8 FILLER_0_2031 ();
 sg13g2_fill_1 FILLER_0_2038 ();
 sg13g2_decap_8 FILLER_0_2047 ();
 sg13g2_decap_8 FILLER_0_2054 ();
 sg13g2_decap_8 FILLER_0_2061 ();
 sg13g2_decap_8 FILLER_0_2068 ();
 sg13g2_decap_4 FILLER_0_2075 ();
 sg13g2_fill_1 FILLER_0_2079 ();
 sg13g2_fill_1 FILLER_0_2088 ();
 sg13g2_decap_8 FILLER_0_2112 ();
 sg13g2_decap_8 FILLER_0_2119 ();
 sg13g2_decap_8 FILLER_0_2126 ();
 sg13g2_decap_4 FILLER_0_2133 ();
 sg13g2_decap_8 FILLER_0_2179 ();
 sg13g2_decap_8 FILLER_0_2186 ();
 sg13g2_decap_8 FILLER_0_2193 ();
 sg13g2_decap_8 FILLER_0_2200 ();
 sg13g2_decap_8 FILLER_0_2221 ();
 sg13g2_decap_8 FILLER_0_2228 ();
 sg13g2_decap_8 FILLER_0_2235 ();
 sg13g2_decap_8 FILLER_0_2242 ();
 sg13g2_fill_1 FILLER_0_2249 ();
 sg13g2_decap_8 FILLER_0_2281 ();
 sg13g2_decap_8 FILLER_0_2288 ();
 sg13g2_decap_8 FILLER_0_2295 ();
 sg13g2_decap_8 FILLER_0_2302 ();
 sg13g2_fill_1 FILLER_0_2309 ();
 sg13g2_decap_8 FILLER_0_2349 ();
 sg13g2_decap_4 FILLER_0_2356 ();
 sg13g2_fill_2 FILLER_0_2360 ();
 sg13g2_fill_2 FILLER_0_2375 ();
 sg13g2_decap_8 FILLER_0_2385 ();
 sg13g2_decap_8 FILLER_0_2392 ();
 sg13g2_decap_8 FILLER_0_2399 ();
 sg13g2_decap_4 FILLER_0_2406 ();
 sg13g2_fill_2 FILLER_0_2410 ();
 sg13g2_fill_1 FILLER_0_2430 ();
 sg13g2_decap_8 FILLER_0_2449 ();
 sg13g2_decap_8 FILLER_0_2456 ();
 sg13g2_decap_8 FILLER_0_2463 ();
 sg13g2_fill_2 FILLER_0_2470 ();
 sg13g2_decap_8 FILLER_0_2484 ();
 sg13g2_decap_8 FILLER_0_2491 ();
 sg13g2_decap_8 FILLER_0_2498 ();
 sg13g2_decap_8 FILLER_0_2505 ();
 sg13g2_decap_8 FILLER_0_2512 ();
 sg13g2_decap_8 FILLER_0_2519 ();
 sg13g2_decap_8 FILLER_0_2526 ();
 sg13g2_decap_8 FILLER_0_2533 ();
 sg13g2_decap_8 FILLER_0_2540 ();
 sg13g2_decap_8 FILLER_0_2547 ();
 sg13g2_decap_8 FILLER_0_2554 ();
 sg13g2_decap_8 FILLER_0_2561 ();
 sg13g2_decap_8 FILLER_0_2568 ();
 sg13g2_decap_8 FILLER_0_2575 ();
 sg13g2_decap_8 FILLER_0_2582 ();
 sg13g2_decap_8 FILLER_0_2589 ();
 sg13g2_decap_8 FILLER_0_2596 ();
 sg13g2_decap_8 FILLER_0_2603 ();
 sg13g2_decap_8 FILLER_0_2610 ();
 sg13g2_decap_8 FILLER_0_2617 ();
 sg13g2_decap_8 FILLER_0_2624 ();
 sg13g2_decap_8 FILLER_0_2631 ();
 sg13g2_decap_8 FILLER_0_2638 ();
 sg13g2_decap_8 FILLER_0_2645 ();
 sg13g2_decap_8 FILLER_0_2652 ();
 sg13g2_decap_8 FILLER_0_2659 ();
 sg13g2_decap_8 FILLER_0_2666 ();
 sg13g2_decap_8 FILLER_0_2673 ();
 sg13g2_decap_8 FILLER_0_2680 ();
 sg13g2_decap_8 FILLER_0_2687 ();
 sg13g2_decap_8 FILLER_0_2694 ();
 sg13g2_decap_8 FILLER_0_2701 ();
 sg13g2_decap_8 FILLER_0_2708 ();
 sg13g2_decap_8 FILLER_0_2715 ();
 sg13g2_decap_8 FILLER_0_2722 ();
 sg13g2_decap_8 FILLER_0_2729 ();
 sg13g2_decap_8 FILLER_0_2736 ();
 sg13g2_decap_8 FILLER_0_2743 ();
 sg13g2_decap_8 FILLER_0_2750 ();
 sg13g2_decap_8 FILLER_0_2757 ();
 sg13g2_decap_8 FILLER_0_2764 ();
 sg13g2_decap_8 FILLER_0_2771 ();
 sg13g2_decap_8 FILLER_0_2778 ();
 sg13g2_decap_8 FILLER_0_2785 ();
 sg13g2_decap_8 FILLER_0_2792 ();
 sg13g2_decap_8 FILLER_0_2799 ();
 sg13g2_decap_8 FILLER_0_2806 ();
 sg13g2_decap_8 FILLER_0_2813 ();
 sg13g2_decap_8 FILLER_0_2820 ();
 sg13g2_decap_8 FILLER_0_2827 ();
 sg13g2_decap_8 FILLER_0_2834 ();
 sg13g2_decap_8 FILLER_0_2841 ();
 sg13g2_decap_8 FILLER_0_2848 ();
 sg13g2_decap_8 FILLER_0_2855 ();
 sg13g2_decap_8 FILLER_0_2862 ();
 sg13g2_decap_8 FILLER_0_2869 ();
 sg13g2_decap_8 FILLER_0_2876 ();
 sg13g2_decap_8 FILLER_0_2883 ();
 sg13g2_decap_8 FILLER_0_2890 ();
 sg13g2_decap_8 FILLER_0_2897 ();
 sg13g2_decap_8 FILLER_0_2904 ();
 sg13g2_decap_8 FILLER_0_2911 ();
 sg13g2_decap_8 FILLER_0_2918 ();
 sg13g2_decap_8 FILLER_0_2925 ();
 sg13g2_decap_8 FILLER_0_2932 ();
 sg13g2_decap_8 FILLER_0_2939 ();
 sg13g2_decap_8 FILLER_0_2946 ();
 sg13g2_decap_8 FILLER_0_2953 ();
 sg13g2_decap_8 FILLER_0_2960 ();
 sg13g2_decap_8 FILLER_0_2967 ();
 sg13g2_decap_8 FILLER_0_2974 ();
 sg13g2_decap_8 FILLER_0_2981 ();
 sg13g2_decap_8 FILLER_0_2988 ();
 sg13g2_decap_8 FILLER_0_2995 ();
 sg13g2_decap_8 FILLER_0_3002 ();
 sg13g2_decap_8 FILLER_0_3009 ();
 sg13g2_decap_8 FILLER_0_3016 ();
 sg13g2_decap_8 FILLER_0_3023 ();
 sg13g2_decap_8 FILLER_0_3030 ();
 sg13g2_decap_8 FILLER_0_3037 ();
 sg13g2_decap_8 FILLER_0_3044 ();
 sg13g2_decap_8 FILLER_0_3051 ();
 sg13g2_decap_8 FILLER_0_3058 ();
 sg13g2_decap_8 FILLER_0_3065 ();
 sg13g2_decap_8 FILLER_0_3072 ();
 sg13g2_decap_8 FILLER_0_3079 ();
 sg13g2_decap_8 FILLER_0_3086 ();
 sg13g2_decap_8 FILLER_0_3093 ();
 sg13g2_decap_8 FILLER_0_3100 ();
 sg13g2_decap_8 FILLER_0_3107 ();
 sg13g2_decap_8 FILLER_0_3114 ();
 sg13g2_decap_8 FILLER_0_3121 ();
 sg13g2_decap_8 FILLER_0_3128 ();
 sg13g2_decap_8 FILLER_0_3135 ();
 sg13g2_decap_8 FILLER_0_3142 ();
 sg13g2_decap_8 FILLER_0_3149 ();
 sg13g2_decap_8 FILLER_0_3156 ();
 sg13g2_decap_8 FILLER_0_3163 ();
 sg13g2_decap_8 FILLER_0_3170 ();
 sg13g2_decap_8 FILLER_0_3177 ();
 sg13g2_decap_8 FILLER_0_3184 ();
 sg13g2_decap_8 FILLER_0_3191 ();
 sg13g2_decap_8 FILLER_0_3198 ();
 sg13g2_decap_8 FILLER_0_3205 ();
 sg13g2_decap_8 FILLER_0_3212 ();
 sg13g2_decap_8 FILLER_0_3219 ();
 sg13g2_decap_8 FILLER_0_3226 ();
 sg13g2_decap_8 FILLER_0_3233 ();
 sg13g2_decap_8 FILLER_0_3240 ();
 sg13g2_decap_8 FILLER_0_3247 ();
 sg13g2_decap_8 FILLER_0_3254 ();
 sg13g2_decap_8 FILLER_0_3261 ();
 sg13g2_decap_8 FILLER_0_3268 ();
 sg13g2_decap_8 FILLER_0_3275 ();
 sg13g2_decap_8 FILLER_0_3282 ();
 sg13g2_decap_8 FILLER_0_3289 ();
 sg13g2_decap_8 FILLER_0_3296 ();
 sg13g2_decap_8 FILLER_0_3303 ();
 sg13g2_decap_8 FILLER_0_3310 ();
 sg13g2_decap_8 FILLER_0_3317 ();
 sg13g2_decap_8 FILLER_0_3324 ();
 sg13g2_decap_8 FILLER_0_3331 ();
 sg13g2_decap_8 FILLER_0_3338 ();
 sg13g2_decap_8 FILLER_0_3345 ();
 sg13g2_decap_8 FILLER_0_3352 ();
 sg13g2_decap_8 FILLER_0_3359 ();
 sg13g2_decap_8 FILLER_0_3366 ();
 sg13g2_decap_8 FILLER_0_3373 ();
 sg13g2_decap_8 FILLER_0_3380 ();
 sg13g2_decap_8 FILLER_0_3387 ();
 sg13g2_decap_8 FILLER_0_3394 ();
 sg13g2_decap_8 FILLER_0_3401 ();
 sg13g2_decap_8 FILLER_0_3408 ();
 sg13g2_decap_8 FILLER_0_3415 ();
 sg13g2_decap_8 FILLER_0_3422 ();
 sg13g2_decap_8 FILLER_0_3429 ();
 sg13g2_decap_8 FILLER_0_3436 ();
 sg13g2_decap_8 FILLER_0_3443 ();
 sg13g2_decap_8 FILLER_0_3450 ();
 sg13g2_decap_8 FILLER_0_3457 ();
 sg13g2_decap_8 FILLER_0_3464 ();
 sg13g2_decap_8 FILLER_0_3471 ();
 sg13g2_decap_8 FILLER_0_3478 ();
 sg13g2_decap_8 FILLER_0_3485 ();
 sg13g2_decap_8 FILLER_0_3492 ();
 sg13g2_decap_8 FILLER_0_3499 ();
 sg13g2_decap_8 FILLER_0_3506 ();
 sg13g2_decap_8 FILLER_0_3513 ();
 sg13g2_decap_8 FILLER_0_3520 ();
 sg13g2_decap_8 FILLER_0_3527 ();
 sg13g2_decap_8 FILLER_0_3534 ();
 sg13g2_decap_8 FILLER_0_3541 ();
 sg13g2_decap_8 FILLER_0_3548 ();
 sg13g2_decap_8 FILLER_0_3555 ();
 sg13g2_decap_8 FILLER_0_3562 ();
 sg13g2_decap_8 FILLER_0_3569 ();
 sg13g2_decap_4 FILLER_0_3576 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_641 ();
 sg13g2_fill_2 FILLER_1_648 ();
 sg13g2_decap_8 FILLER_1_741 ();
 sg13g2_decap_8 FILLER_1_748 ();
 sg13g2_decap_8 FILLER_1_781 ();
 sg13g2_decap_8 FILLER_1_788 ();
 sg13g2_fill_2 FILLER_1_795 ();
 sg13g2_fill_2 FILLER_1_823 ();
 sg13g2_decap_8 FILLER_1_856 ();
 sg13g2_decap_4 FILLER_1_863 ();
 sg13g2_decap_8 FILLER_1_893 ();
 sg13g2_decap_4 FILLER_1_900 ();
 sg13g2_fill_1 FILLER_1_904 ();
 sg13g2_fill_1 FILLER_1_934 ();
 sg13g2_fill_2 FILLER_1_987 ();
 sg13g2_fill_2 FILLER_1_994 ();
 sg13g2_fill_1 FILLER_1_996 ();
 sg13g2_decap_8 FILLER_1_1014 ();
 sg13g2_fill_2 FILLER_1_1021 ();
 sg13g2_decap_8 FILLER_1_1049 ();
 sg13g2_decap_8 FILLER_1_1056 ();
 sg13g2_decap_8 FILLER_1_1063 ();
 sg13g2_decap_8 FILLER_1_1070 ();
 sg13g2_decap_8 FILLER_1_1077 ();
 sg13g2_decap_8 FILLER_1_1084 ();
 sg13g2_decap_8 FILLER_1_1091 ();
 sg13g2_decap_8 FILLER_1_1098 ();
 sg13g2_decap_8 FILLER_1_1105 ();
 sg13g2_decap_8 FILLER_1_1112 ();
 sg13g2_decap_8 FILLER_1_1119 ();
 sg13g2_decap_8 FILLER_1_1126 ();
 sg13g2_decap_8 FILLER_1_1133 ();
 sg13g2_decap_8 FILLER_1_1140 ();
 sg13g2_decap_8 FILLER_1_1147 ();
 sg13g2_decap_8 FILLER_1_1154 ();
 sg13g2_decap_8 FILLER_1_1161 ();
 sg13g2_fill_1 FILLER_1_1168 ();
 sg13g2_decap_8 FILLER_1_1177 ();
 sg13g2_decap_8 FILLER_1_1184 ();
 sg13g2_decap_8 FILLER_1_1191 ();
 sg13g2_decap_8 FILLER_1_1198 ();
 sg13g2_decap_8 FILLER_1_1205 ();
 sg13g2_decap_4 FILLER_1_1212 ();
 sg13g2_fill_2 FILLER_1_1216 ();
 sg13g2_fill_1 FILLER_1_1296 ();
 sg13g2_decap_4 FILLER_1_1302 ();
 sg13g2_fill_1 FILLER_1_1306 ();
 sg13g2_decap_8 FILLER_1_1310 ();
 sg13g2_decap_8 FILLER_1_1317 ();
 sg13g2_decap_8 FILLER_1_1324 ();
 sg13g2_decap_4 FILLER_1_1331 ();
 sg13g2_fill_1 FILLER_1_1335 ();
 sg13g2_fill_2 FILLER_1_1372 ();
 sg13g2_fill_1 FILLER_1_1374 ();
 sg13g2_decap_8 FILLER_1_1401 ();
 sg13g2_decap_4 FILLER_1_1408 ();
 sg13g2_decap_8 FILLER_1_1451 ();
 sg13g2_fill_2 FILLER_1_1458 ();
 sg13g2_fill_1 FILLER_1_1460 ();
 sg13g2_decap_8 FILLER_1_1509 ();
 sg13g2_decap_8 FILLER_1_1516 ();
 sg13g2_decap_8 FILLER_1_1523 ();
 sg13g2_decap_4 FILLER_1_1530 ();
 sg13g2_fill_2 FILLER_1_1534 ();
 sg13g2_decap_8 FILLER_1_1570 ();
 sg13g2_decap_8 FILLER_1_1577 ();
 sg13g2_decap_4 FILLER_1_1584 ();
 sg13g2_fill_2 FILLER_1_1614 ();
 sg13g2_decap_8 FILLER_1_1650 ();
 sg13g2_decap_8 FILLER_1_1657 ();
 sg13g2_decap_8 FILLER_1_1727 ();
 sg13g2_decap_8 FILLER_1_1734 ();
 sg13g2_decap_8 FILLER_1_1741 ();
 sg13g2_decap_8 FILLER_1_1795 ();
 sg13g2_decap_8 FILLER_1_1802 ();
 sg13g2_fill_2 FILLER_1_1809 ();
 sg13g2_fill_2 FILLER_1_1840 ();
 sg13g2_fill_2 FILLER_1_1868 ();
 sg13g2_fill_2 FILLER_1_1882 ();
 sg13g2_fill_1 FILLER_1_1884 ();
 sg13g2_decap_8 FILLER_1_1937 ();
 sg13g2_decap_8 FILLER_1_1944 ();
 sg13g2_decap_8 FILLER_1_1951 ();
 sg13g2_decap_8 FILLER_1_1958 ();
 sg13g2_decap_8 FILLER_1_1965 ();
 sg13g2_decap_8 FILLER_1_1972 ();
 sg13g2_decap_8 FILLER_1_1979 ();
 sg13g2_decap_8 FILLER_1_1986 ();
 sg13g2_decap_4 FILLER_1_1993 ();
 sg13g2_fill_2 FILLER_1_1997 ();
 sg13g2_decap_4 FILLER_1_2049 ();
 sg13g2_fill_2 FILLER_1_2073 ();
 sg13g2_fill_2 FILLER_1_2088 ();
 sg13g2_decap_8 FILLER_1_2116 ();
 sg13g2_decap_8 FILLER_1_2123 ();
 sg13g2_fill_1 FILLER_1_2130 ();
 sg13g2_fill_2 FILLER_1_2165 ();
 sg13g2_fill_1 FILLER_1_2184 ();
 sg13g2_decap_8 FILLER_1_2190 ();
 sg13g2_fill_1 FILLER_1_2197 ();
 sg13g2_fill_1 FILLER_1_2206 ();
 sg13g2_decap_8 FILLER_1_2233 ();
 sg13g2_fill_2 FILLER_1_2240 ();
 sg13g2_decap_8 FILLER_1_2294 ();
 sg13g2_decap_4 FILLER_1_2301 ();
 sg13g2_fill_2 FILLER_1_2347 ();
 sg13g2_fill_1 FILLER_1_2349 ();
 sg13g2_decap_4 FILLER_1_2401 ();
 sg13g2_fill_2 FILLER_1_2405 ();
 sg13g2_decap_4 FILLER_1_2449 ();
 sg13g2_decap_8 FILLER_1_2491 ();
 sg13g2_decap_8 FILLER_1_2498 ();
 sg13g2_decap_8 FILLER_1_2505 ();
 sg13g2_decap_8 FILLER_1_2512 ();
 sg13g2_decap_8 FILLER_1_2519 ();
 sg13g2_decap_8 FILLER_1_2526 ();
 sg13g2_decap_8 FILLER_1_2533 ();
 sg13g2_decap_8 FILLER_1_2540 ();
 sg13g2_decap_8 FILLER_1_2547 ();
 sg13g2_decap_8 FILLER_1_2554 ();
 sg13g2_decap_8 FILLER_1_2561 ();
 sg13g2_decap_8 FILLER_1_2568 ();
 sg13g2_decap_8 FILLER_1_2575 ();
 sg13g2_decap_8 FILLER_1_2582 ();
 sg13g2_decap_8 FILLER_1_2589 ();
 sg13g2_decap_8 FILLER_1_2596 ();
 sg13g2_decap_8 FILLER_1_2603 ();
 sg13g2_decap_8 FILLER_1_2610 ();
 sg13g2_decap_8 FILLER_1_2617 ();
 sg13g2_decap_8 FILLER_1_2624 ();
 sg13g2_decap_8 FILLER_1_2631 ();
 sg13g2_decap_8 FILLER_1_2638 ();
 sg13g2_decap_8 FILLER_1_2645 ();
 sg13g2_decap_8 FILLER_1_2652 ();
 sg13g2_decap_8 FILLER_1_2659 ();
 sg13g2_decap_8 FILLER_1_2666 ();
 sg13g2_decap_8 FILLER_1_2673 ();
 sg13g2_decap_8 FILLER_1_2680 ();
 sg13g2_decap_8 FILLER_1_2687 ();
 sg13g2_decap_8 FILLER_1_2694 ();
 sg13g2_decap_8 FILLER_1_2701 ();
 sg13g2_decap_8 FILLER_1_2708 ();
 sg13g2_decap_8 FILLER_1_2715 ();
 sg13g2_decap_8 FILLER_1_2722 ();
 sg13g2_decap_8 FILLER_1_2729 ();
 sg13g2_decap_8 FILLER_1_2736 ();
 sg13g2_decap_8 FILLER_1_2743 ();
 sg13g2_decap_8 FILLER_1_2750 ();
 sg13g2_decap_8 FILLER_1_2757 ();
 sg13g2_decap_8 FILLER_1_2764 ();
 sg13g2_decap_8 FILLER_1_2771 ();
 sg13g2_decap_8 FILLER_1_2778 ();
 sg13g2_decap_8 FILLER_1_2785 ();
 sg13g2_decap_8 FILLER_1_2792 ();
 sg13g2_decap_8 FILLER_1_2799 ();
 sg13g2_decap_8 FILLER_1_2806 ();
 sg13g2_decap_8 FILLER_1_2813 ();
 sg13g2_decap_8 FILLER_1_2820 ();
 sg13g2_decap_8 FILLER_1_2827 ();
 sg13g2_decap_8 FILLER_1_2834 ();
 sg13g2_decap_8 FILLER_1_2841 ();
 sg13g2_decap_8 FILLER_1_2848 ();
 sg13g2_decap_8 FILLER_1_2855 ();
 sg13g2_decap_8 FILLER_1_2862 ();
 sg13g2_decap_8 FILLER_1_2869 ();
 sg13g2_decap_8 FILLER_1_2876 ();
 sg13g2_decap_8 FILLER_1_2883 ();
 sg13g2_decap_8 FILLER_1_2890 ();
 sg13g2_decap_8 FILLER_1_2897 ();
 sg13g2_decap_8 FILLER_1_2904 ();
 sg13g2_decap_8 FILLER_1_2911 ();
 sg13g2_decap_8 FILLER_1_2918 ();
 sg13g2_decap_8 FILLER_1_2925 ();
 sg13g2_decap_8 FILLER_1_2932 ();
 sg13g2_decap_8 FILLER_1_2939 ();
 sg13g2_decap_8 FILLER_1_2946 ();
 sg13g2_decap_8 FILLER_1_2953 ();
 sg13g2_decap_8 FILLER_1_2960 ();
 sg13g2_decap_8 FILLER_1_2967 ();
 sg13g2_decap_8 FILLER_1_2974 ();
 sg13g2_decap_8 FILLER_1_2981 ();
 sg13g2_decap_8 FILLER_1_2988 ();
 sg13g2_decap_8 FILLER_1_2995 ();
 sg13g2_decap_8 FILLER_1_3002 ();
 sg13g2_decap_8 FILLER_1_3009 ();
 sg13g2_decap_8 FILLER_1_3016 ();
 sg13g2_decap_8 FILLER_1_3023 ();
 sg13g2_decap_8 FILLER_1_3030 ();
 sg13g2_decap_8 FILLER_1_3037 ();
 sg13g2_decap_8 FILLER_1_3044 ();
 sg13g2_decap_8 FILLER_1_3051 ();
 sg13g2_decap_8 FILLER_1_3058 ();
 sg13g2_decap_8 FILLER_1_3065 ();
 sg13g2_decap_8 FILLER_1_3072 ();
 sg13g2_decap_8 FILLER_1_3079 ();
 sg13g2_decap_8 FILLER_1_3086 ();
 sg13g2_decap_8 FILLER_1_3093 ();
 sg13g2_decap_8 FILLER_1_3100 ();
 sg13g2_decap_8 FILLER_1_3107 ();
 sg13g2_decap_8 FILLER_1_3114 ();
 sg13g2_decap_8 FILLER_1_3121 ();
 sg13g2_decap_8 FILLER_1_3128 ();
 sg13g2_decap_8 FILLER_1_3135 ();
 sg13g2_decap_8 FILLER_1_3142 ();
 sg13g2_decap_8 FILLER_1_3149 ();
 sg13g2_decap_8 FILLER_1_3156 ();
 sg13g2_decap_8 FILLER_1_3163 ();
 sg13g2_decap_8 FILLER_1_3170 ();
 sg13g2_decap_8 FILLER_1_3177 ();
 sg13g2_decap_8 FILLER_1_3184 ();
 sg13g2_decap_8 FILLER_1_3191 ();
 sg13g2_decap_8 FILLER_1_3198 ();
 sg13g2_decap_8 FILLER_1_3205 ();
 sg13g2_decap_8 FILLER_1_3212 ();
 sg13g2_decap_8 FILLER_1_3219 ();
 sg13g2_decap_8 FILLER_1_3226 ();
 sg13g2_decap_8 FILLER_1_3233 ();
 sg13g2_decap_8 FILLER_1_3240 ();
 sg13g2_decap_8 FILLER_1_3247 ();
 sg13g2_decap_8 FILLER_1_3254 ();
 sg13g2_decap_8 FILLER_1_3261 ();
 sg13g2_decap_8 FILLER_1_3268 ();
 sg13g2_decap_8 FILLER_1_3275 ();
 sg13g2_decap_8 FILLER_1_3282 ();
 sg13g2_decap_8 FILLER_1_3289 ();
 sg13g2_decap_8 FILLER_1_3296 ();
 sg13g2_decap_8 FILLER_1_3303 ();
 sg13g2_decap_8 FILLER_1_3310 ();
 sg13g2_decap_8 FILLER_1_3317 ();
 sg13g2_decap_8 FILLER_1_3324 ();
 sg13g2_decap_8 FILLER_1_3331 ();
 sg13g2_decap_8 FILLER_1_3338 ();
 sg13g2_decap_8 FILLER_1_3345 ();
 sg13g2_decap_8 FILLER_1_3352 ();
 sg13g2_decap_8 FILLER_1_3359 ();
 sg13g2_decap_8 FILLER_1_3366 ();
 sg13g2_decap_8 FILLER_1_3373 ();
 sg13g2_decap_8 FILLER_1_3380 ();
 sg13g2_decap_8 FILLER_1_3387 ();
 sg13g2_decap_8 FILLER_1_3394 ();
 sg13g2_decap_8 FILLER_1_3401 ();
 sg13g2_decap_8 FILLER_1_3408 ();
 sg13g2_decap_8 FILLER_1_3415 ();
 sg13g2_decap_8 FILLER_1_3422 ();
 sg13g2_decap_8 FILLER_1_3429 ();
 sg13g2_decap_8 FILLER_1_3436 ();
 sg13g2_decap_8 FILLER_1_3443 ();
 sg13g2_decap_8 FILLER_1_3450 ();
 sg13g2_decap_8 FILLER_1_3457 ();
 sg13g2_decap_8 FILLER_1_3464 ();
 sg13g2_decap_8 FILLER_1_3471 ();
 sg13g2_decap_8 FILLER_1_3478 ();
 sg13g2_decap_8 FILLER_1_3485 ();
 sg13g2_decap_8 FILLER_1_3492 ();
 sg13g2_decap_8 FILLER_1_3499 ();
 sg13g2_decap_8 FILLER_1_3506 ();
 sg13g2_decap_8 FILLER_1_3513 ();
 sg13g2_decap_8 FILLER_1_3520 ();
 sg13g2_decap_8 FILLER_1_3527 ();
 sg13g2_decap_8 FILLER_1_3534 ();
 sg13g2_decap_8 FILLER_1_3541 ();
 sg13g2_decap_8 FILLER_1_3548 ();
 sg13g2_decap_8 FILLER_1_3555 ();
 sg13g2_decap_8 FILLER_1_3562 ();
 sg13g2_decap_8 FILLER_1_3569 ();
 sg13g2_decap_4 FILLER_1_3576 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_4 FILLER_2_581 ();
 sg13g2_fill_2 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_649 ();
 sg13g2_decap_4 FILLER_2_656 ();
 sg13g2_fill_2 FILLER_2_660 ();
 sg13g2_fill_1 FILLER_2_701 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_fill_2 FILLER_2_756 ();
 sg13g2_fill_2 FILLER_2_789 ();
 sg13g2_decap_8 FILLER_2_863 ();
 sg13g2_decap_8 FILLER_2_870 ();
 sg13g2_decap_8 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_2_884 ();
 sg13g2_decap_8 FILLER_2_891 ();
 sg13g2_decap_4 FILLER_2_898 ();
 sg13g2_fill_1 FILLER_2_902 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_fill_2 FILLER_2_914 ();
 sg13g2_fill_2 FILLER_2_938 ();
 sg13g2_fill_1 FILLER_2_940 ();
 sg13g2_fill_1 FILLER_2_993 ();
 sg13g2_fill_1 FILLER_2_1025 ();
 sg13g2_decap_8 FILLER_2_1060 ();
 sg13g2_decap_8 FILLER_2_1067 ();
 sg13g2_decap_8 FILLER_2_1074 ();
 sg13g2_decap_8 FILLER_2_1081 ();
 sg13g2_decap_8 FILLER_2_1088 ();
 sg13g2_decap_8 FILLER_2_1095 ();
 sg13g2_decap_8 FILLER_2_1102 ();
 sg13g2_decap_8 FILLER_2_1109 ();
 sg13g2_decap_8 FILLER_2_1116 ();
 sg13g2_decap_8 FILLER_2_1123 ();
 sg13g2_decap_8 FILLER_2_1130 ();
 sg13g2_decap_8 FILLER_2_1137 ();
 sg13g2_decap_4 FILLER_2_1144 ();
 sg13g2_fill_1 FILLER_2_1148 ();
 sg13g2_decap_8 FILLER_2_1190 ();
 sg13g2_decap_8 FILLER_2_1197 ();
 sg13g2_decap_4 FILLER_2_1204 ();
 sg13g2_fill_2 FILLER_2_1208 ();
 sg13g2_decap_4 FILLER_2_1312 ();
 sg13g2_fill_1 FILLER_2_1321 ();
 sg13g2_fill_1 FILLER_2_1332 ();
 sg13g2_fill_2 FILLER_2_1346 ();
 sg13g2_fill_1 FILLER_2_1348 ();
 sg13g2_fill_2 FILLER_2_1378 ();
 sg13g2_fill_2 FILLER_2_1419 ();
 sg13g2_fill_1 FILLER_2_1462 ();
 sg13g2_decap_8 FILLER_2_1515 ();
 sg13g2_decap_4 FILLER_2_1522 ();
 sg13g2_fill_2 FILLER_2_1526 ();
 sg13g2_fill_1 FILLER_2_1575 ();
 sg13g2_fill_2 FILLER_2_1659 ();
 sg13g2_decap_4 FILLER_2_1737 ();
 sg13g2_fill_2 FILLER_2_1801 ();
 sg13g2_fill_1 FILLER_2_1803 ();
 sg13g2_fill_2 FILLER_2_1862 ();
 sg13g2_decap_8 FILLER_2_1874 ();
 sg13g2_fill_2 FILLER_2_1897 ();
 sg13g2_decap_8 FILLER_2_1933 ();
 sg13g2_decap_8 FILLER_2_1940 ();
 sg13g2_decap_8 FILLER_2_1947 ();
 sg13g2_decap_8 FILLER_2_1954 ();
 sg13g2_decap_8 FILLER_2_1961 ();
 sg13g2_decap_8 FILLER_2_1968 ();
 sg13g2_decap_8 FILLER_2_1975 ();
 sg13g2_decap_8 FILLER_2_1982 ();
 sg13g2_decap_8 FILLER_2_1989 ();
 sg13g2_fill_1 FILLER_2_1996 ();
 sg13g2_fill_2 FILLER_2_2124 ();
 sg13g2_fill_2 FILLER_2_2173 ();
 sg13g2_decap_4 FILLER_2_2232 ();
 sg13g2_fill_1 FILLER_2_2236 ();
 sg13g2_fill_1 FILLER_2_2245 ();
 sg13g2_fill_1 FILLER_2_2280 ();
 sg13g2_fill_2 FILLER_2_2356 ();
 sg13g2_fill_1 FILLER_2_2358 ();
 sg13g2_decap_8 FILLER_2_2499 ();
 sg13g2_decap_8 FILLER_2_2506 ();
 sg13g2_decap_8 FILLER_2_2513 ();
 sg13g2_decap_8 FILLER_2_2520 ();
 sg13g2_decap_8 FILLER_2_2527 ();
 sg13g2_decap_8 FILLER_2_2534 ();
 sg13g2_decap_8 FILLER_2_2541 ();
 sg13g2_decap_8 FILLER_2_2548 ();
 sg13g2_decap_8 FILLER_2_2555 ();
 sg13g2_decap_8 FILLER_2_2562 ();
 sg13g2_decap_8 FILLER_2_2569 ();
 sg13g2_decap_8 FILLER_2_2576 ();
 sg13g2_decap_8 FILLER_2_2583 ();
 sg13g2_decap_8 FILLER_2_2590 ();
 sg13g2_decap_8 FILLER_2_2597 ();
 sg13g2_decap_8 FILLER_2_2604 ();
 sg13g2_decap_8 FILLER_2_2611 ();
 sg13g2_decap_8 FILLER_2_2618 ();
 sg13g2_decap_8 FILLER_2_2625 ();
 sg13g2_decap_8 FILLER_2_2632 ();
 sg13g2_decap_8 FILLER_2_2639 ();
 sg13g2_decap_8 FILLER_2_2646 ();
 sg13g2_decap_8 FILLER_2_2653 ();
 sg13g2_decap_8 FILLER_2_2660 ();
 sg13g2_decap_8 FILLER_2_2667 ();
 sg13g2_decap_8 FILLER_2_2674 ();
 sg13g2_decap_8 FILLER_2_2681 ();
 sg13g2_decap_8 FILLER_2_2688 ();
 sg13g2_decap_8 FILLER_2_2695 ();
 sg13g2_decap_8 FILLER_2_2702 ();
 sg13g2_decap_8 FILLER_2_2709 ();
 sg13g2_decap_8 FILLER_2_2716 ();
 sg13g2_decap_8 FILLER_2_2723 ();
 sg13g2_decap_8 FILLER_2_2730 ();
 sg13g2_decap_8 FILLER_2_2737 ();
 sg13g2_decap_8 FILLER_2_2744 ();
 sg13g2_decap_8 FILLER_2_2751 ();
 sg13g2_decap_8 FILLER_2_2758 ();
 sg13g2_decap_8 FILLER_2_2765 ();
 sg13g2_decap_8 FILLER_2_2772 ();
 sg13g2_decap_8 FILLER_2_2779 ();
 sg13g2_decap_8 FILLER_2_2786 ();
 sg13g2_decap_8 FILLER_2_2793 ();
 sg13g2_decap_8 FILLER_2_2800 ();
 sg13g2_decap_8 FILLER_2_2807 ();
 sg13g2_decap_8 FILLER_2_2814 ();
 sg13g2_decap_8 FILLER_2_2821 ();
 sg13g2_decap_8 FILLER_2_2828 ();
 sg13g2_decap_8 FILLER_2_2835 ();
 sg13g2_decap_8 FILLER_2_2842 ();
 sg13g2_decap_8 FILLER_2_2849 ();
 sg13g2_decap_8 FILLER_2_2856 ();
 sg13g2_decap_8 FILLER_2_2863 ();
 sg13g2_decap_8 FILLER_2_2870 ();
 sg13g2_decap_8 FILLER_2_2877 ();
 sg13g2_decap_8 FILLER_2_2884 ();
 sg13g2_decap_8 FILLER_2_2891 ();
 sg13g2_decap_8 FILLER_2_2898 ();
 sg13g2_decap_8 FILLER_2_2905 ();
 sg13g2_decap_8 FILLER_2_2912 ();
 sg13g2_decap_8 FILLER_2_2919 ();
 sg13g2_decap_8 FILLER_2_2926 ();
 sg13g2_decap_8 FILLER_2_2933 ();
 sg13g2_decap_8 FILLER_2_2940 ();
 sg13g2_decap_8 FILLER_2_2947 ();
 sg13g2_decap_8 FILLER_2_2954 ();
 sg13g2_decap_8 FILLER_2_2961 ();
 sg13g2_decap_8 FILLER_2_2968 ();
 sg13g2_decap_8 FILLER_2_2975 ();
 sg13g2_decap_8 FILLER_2_2982 ();
 sg13g2_decap_8 FILLER_2_2989 ();
 sg13g2_decap_8 FILLER_2_2996 ();
 sg13g2_decap_8 FILLER_2_3003 ();
 sg13g2_decap_8 FILLER_2_3010 ();
 sg13g2_decap_8 FILLER_2_3017 ();
 sg13g2_decap_8 FILLER_2_3024 ();
 sg13g2_decap_8 FILLER_2_3031 ();
 sg13g2_decap_8 FILLER_2_3038 ();
 sg13g2_decap_8 FILLER_2_3045 ();
 sg13g2_decap_8 FILLER_2_3052 ();
 sg13g2_decap_8 FILLER_2_3059 ();
 sg13g2_decap_8 FILLER_2_3066 ();
 sg13g2_decap_8 FILLER_2_3073 ();
 sg13g2_decap_8 FILLER_2_3080 ();
 sg13g2_decap_8 FILLER_2_3087 ();
 sg13g2_decap_8 FILLER_2_3094 ();
 sg13g2_decap_8 FILLER_2_3101 ();
 sg13g2_decap_8 FILLER_2_3108 ();
 sg13g2_decap_8 FILLER_2_3115 ();
 sg13g2_decap_8 FILLER_2_3122 ();
 sg13g2_decap_8 FILLER_2_3129 ();
 sg13g2_decap_8 FILLER_2_3136 ();
 sg13g2_decap_8 FILLER_2_3143 ();
 sg13g2_decap_8 FILLER_2_3150 ();
 sg13g2_decap_8 FILLER_2_3157 ();
 sg13g2_decap_8 FILLER_2_3164 ();
 sg13g2_decap_8 FILLER_2_3171 ();
 sg13g2_decap_8 FILLER_2_3178 ();
 sg13g2_decap_8 FILLER_2_3185 ();
 sg13g2_decap_8 FILLER_2_3192 ();
 sg13g2_decap_8 FILLER_2_3199 ();
 sg13g2_decap_8 FILLER_2_3206 ();
 sg13g2_decap_8 FILLER_2_3213 ();
 sg13g2_decap_8 FILLER_2_3220 ();
 sg13g2_decap_8 FILLER_2_3227 ();
 sg13g2_decap_8 FILLER_2_3234 ();
 sg13g2_decap_8 FILLER_2_3241 ();
 sg13g2_decap_8 FILLER_2_3248 ();
 sg13g2_decap_8 FILLER_2_3255 ();
 sg13g2_decap_8 FILLER_2_3262 ();
 sg13g2_decap_8 FILLER_2_3269 ();
 sg13g2_decap_8 FILLER_2_3276 ();
 sg13g2_decap_8 FILLER_2_3283 ();
 sg13g2_decap_8 FILLER_2_3290 ();
 sg13g2_decap_8 FILLER_2_3297 ();
 sg13g2_decap_8 FILLER_2_3304 ();
 sg13g2_decap_8 FILLER_2_3311 ();
 sg13g2_decap_8 FILLER_2_3318 ();
 sg13g2_decap_8 FILLER_2_3325 ();
 sg13g2_decap_8 FILLER_2_3332 ();
 sg13g2_decap_8 FILLER_2_3339 ();
 sg13g2_decap_8 FILLER_2_3346 ();
 sg13g2_decap_8 FILLER_2_3353 ();
 sg13g2_decap_8 FILLER_2_3360 ();
 sg13g2_decap_8 FILLER_2_3367 ();
 sg13g2_decap_8 FILLER_2_3374 ();
 sg13g2_decap_8 FILLER_2_3381 ();
 sg13g2_decap_8 FILLER_2_3388 ();
 sg13g2_decap_8 FILLER_2_3395 ();
 sg13g2_decap_8 FILLER_2_3402 ();
 sg13g2_decap_8 FILLER_2_3409 ();
 sg13g2_decap_8 FILLER_2_3416 ();
 sg13g2_decap_8 FILLER_2_3423 ();
 sg13g2_decap_8 FILLER_2_3430 ();
 sg13g2_decap_8 FILLER_2_3437 ();
 sg13g2_decap_8 FILLER_2_3444 ();
 sg13g2_decap_8 FILLER_2_3451 ();
 sg13g2_decap_8 FILLER_2_3458 ();
 sg13g2_decap_8 FILLER_2_3465 ();
 sg13g2_decap_8 FILLER_2_3472 ();
 sg13g2_decap_8 FILLER_2_3479 ();
 sg13g2_decap_8 FILLER_2_3486 ();
 sg13g2_decap_8 FILLER_2_3493 ();
 sg13g2_decap_8 FILLER_2_3500 ();
 sg13g2_decap_8 FILLER_2_3507 ();
 sg13g2_decap_8 FILLER_2_3514 ();
 sg13g2_decap_8 FILLER_2_3521 ();
 sg13g2_decap_8 FILLER_2_3528 ();
 sg13g2_decap_8 FILLER_2_3535 ();
 sg13g2_decap_8 FILLER_2_3542 ();
 sg13g2_decap_8 FILLER_2_3549 ();
 sg13g2_decap_8 FILLER_2_3556 ();
 sg13g2_decap_8 FILLER_2_3563 ();
 sg13g2_decap_8 FILLER_2_3570 ();
 sg13g2_fill_2 FILLER_2_3577 ();
 sg13g2_fill_1 FILLER_2_3579 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_4 FILLER_3_574 ();
 sg13g2_fill_2 FILLER_3_578 ();
 sg13g2_decap_8 FILLER_3_690 ();
 sg13g2_decap_8 FILLER_3_697 ();
 sg13g2_decap_8 FILLER_3_704 ();
 sg13g2_fill_2 FILLER_3_711 ();
 sg13g2_fill_1 FILLER_3_713 ();
 sg13g2_fill_2 FILLER_3_752 ();
 sg13g2_decap_8 FILLER_3_818 ();
 sg13g2_decap_8 FILLER_3_875 ();
 sg13g2_decap_8 FILLER_3_882 ();
 sg13g2_decap_8 FILLER_3_889 ();
 sg13g2_decap_8 FILLER_3_896 ();
 sg13g2_decap_8 FILLER_3_903 ();
 sg13g2_decap_8 FILLER_3_910 ();
 sg13g2_decap_4 FILLER_3_917 ();
 sg13g2_fill_2 FILLER_3_921 ();
 sg13g2_decap_8 FILLER_3_928 ();
 sg13g2_decap_8 FILLER_3_935 ();
 sg13g2_decap_4 FILLER_3_942 ();
 sg13g2_decap_4 FILLER_3_950 ();
 sg13g2_fill_2 FILLER_3_954 ();
 sg13g2_decap_4 FILLER_3_963 ();
 sg13g2_fill_2 FILLER_3_970 ();
 sg13g2_fill_2 FILLER_3_976 ();
 sg13g2_fill_2 FILLER_3_982 ();
 sg13g2_decap_8 FILLER_3_1012 ();
 sg13g2_fill_1 FILLER_3_1019 ();
 sg13g2_fill_1 FILLER_3_1058 ();
 sg13g2_decap_8 FILLER_3_1099 ();
 sg13g2_decap_8 FILLER_3_1106 ();
 sg13g2_decap_8 FILLER_3_1113 ();
 sg13g2_decap_8 FILLER_3_1120 ();
 sg13g2_decap_8 FILLER_3_1127 ();
 sg13g2_decap_4 FILLER_3_1134 ();
 sg13g2_fill_2 FILLER_3_1138 ();
 sg13g2_fill_1 FILLER_3_1161 ();
 sg13g2_decap_8 FILLER_3_1198 ();
 sg13g2_decap_8 FILLER_3_1205 ();
 sg13g2_fill_2 FILLER_3_1212 ();
 sg13g2_fill_1 FILLER_3_1214 ();
 sg13g2_decap_4 FILLER_3_1269 ();
 sg13g2_fill_1 FILLER_3_1273 ();
 sg13g2_fill_2 FILLER_3_1360 ();
 sg13g2_decap_8 FILLER_3_1396 ();
 sg13g2_fill_2 FILLER_3_1403 ();
 sg13g2_fill_1 FILLER_3_1405 ();
 sg13g2_decap_4 FILLER_3_1437 ();
 sg13g2_decap_8 FILLER_3_1454 ();
 sg13g2_decap_8 FILLER_3_1520 ();
 sg13g2_fill_1 FILLER_3_1527 ();
 sg13g2_decap_8 FILLER_3_1572 ();
 sg13g2_decap_8 FILLER_3_1579 ();
 sg13g2_fill_1 FILLER_3_1586 ();
 sg13g2_fill_2 FILLER_3_1595 ();
 sg13g2_fill_1 FILLER_3_1618 ();
 sg13g2_fill_1 FILLER_3_1624 ();
 sg13g2_decap_8 FILLER_3_1652 ();
 sg13g2_decap_4 FILLER_3_1659 ();
 sg13g2_fill_1 FILLER_3_1663 ();
 sg13g2_fill_1 FILLER_3_1687 ();
 sg13g2_fill_2 FILLER_3_1693 ();
 sg13g2_decap_4 FILLER_3_1719 ();
 sg13g2_decap_8 FILLER_3_1739 ();
 sg13g2_fill_1 FILLER_3_1746 ();
 sg13g2_decap_8 FILLER_3_1802 ();
 sg13g2_decap_8 FILLER_3_1809 ();
 sg13g2_fill_2 FILLER_3_1816 ();
 sg13g2_fill_1 FILLER_3_1834 ();
 sg13g2_fill_2 FILLER_3_1874 ();
 sg13g2_fill_1 FILLER_3_1876 ();
 sg13g2_decap_8 FILLER_3_1923 ();
 sg13g2_decap_4 FILLER_3_1930 ();
 sg13g2_fill_2 FILLER_3_1934 ();
 sg13g2_decap_8 FILLER_3_1941 ();
 sg13g2_decap_8 FILLER_3_1948 ();
 sg13g2_decap_8 FILLER_3_1955 ();
 sg13g2_decap_8 FILLER_3_1962 ();
 sg13g2_decap_8 FILLER_3_1969 ();
 sg13g2_decap_4 FILLER_3_1976 ();
 sg13g2_fill_2 FILLER_3_1980 ();
 sg13g2_fill_2 FILLER_3_2077 ();
 sg13g2_fill_1 FILLER_3_2079 ();
 sg13g2_fill_2 FILLER_3_2130 ();
 sg13g2_fill_1 FILLER_3_2132 ();
 sg13g2_fill_1 FILLER_3_2174 ();
 sg13g2_decap_8 FILLER_3_2191 ();
 sg13g2_fill_2 FILLER_3_2198 ();
 sg13g2_decap_8 FILLER_3_2224 ();
 sg13g2_decap_8 FILLER_3_2240 ();
 sg13g2_fill_2 FILLER_3_2247 ();
 sg13g2_fill_1 FILLER_3_2249 ();
 sg13g2_fill_1 FILLER_3_2263 ();
 sg13g2_fill_1 FILLER_3_2286 ();
 sg13g2_decap_8 FILLER_3_2295 ();
 sg13g2_decap_4 FILLER_3_2302 ();
 sg13g2_fill_1 FILLER_3_2306 ();
 sg13g2_fill_2 FILLER_3_2353 ();
 sg13g2_fill_1 FILLER_3_2355 ();
 sg13g2_decap_8 FILLER_3_2401 ();
 sg13g2_decap_4 FILLER_3_2449 ();
 sg13g2_fill_1 FILLER_3_2453 ();
 sg13g2_decap_8 FILLER_3_2498 ();
 sg13g2_decap_8 FILLER_3_2505 ();
 sg13g2_decap_8 FILLER_3_2512 ();
 sg13g2_decap_8 FILLER_3_2519 ();
 sg13g2_decap_8 FILLER_3_2526 ();
 sg13g2_decap_8 FILLER_3_2533 ();
 sg13g2_decap_8 FILLER_3_2540 ();
 sg13g2_decap_8 FILLER_3_2547 ();
 sg13g2_decap_8 FILLER_3_2554 ();
 sg13g2_decap_8 FILLER_3_2561 ();
 sg13g2_decap_8 FILLER_3_2568 ();
 sg13g2_decap_8 FILLER_3_2575 ();
 sg13g2_decap_8 FILLER_3_2582 ();
 sg13g2_decap_8 FILLER_3_2589 ();
 sg13g2_decap_8 FILLER_3_2596 ();
 sg13g2_decap_8 FILLER_3_2603 ();
 sg13g2_decap_8 FILLER_3_2610 ();
 sg13g2_decap_8 FILLER_3_2617 ();
 sg13g2_decap_8 FILLER_3_2624 ();
 sg13g2_decap_8 FILLER_3_2631 ();
 sg13g2_decap_8 FILLER_3_2638 ();
 sg13g2_decap_8 FILLER_3_2645 ();
 sg13g2_decap_8 FILLER_3_2652 ();
 sg13g2_decap_8 FILLER_3_2659 ();
 sg13g2_decap_8 FILLER_3_2666 ();
 sg13g2_decap_8 FILLER_3_2673 ();
 sg13g2_decap_8 FILLER_3_2680 ();
 sg13g2_decap_8 FILLER_3_2687 ();
 sg13g2_decap_8 FILLER_3_2694 ();
 sg13g2_decap_8 FILLER_3_2701 ();
 sg13g2_decap_8 FILLER_3_2708 ();
 sg13g2_decap_8 FILLER_3_2715 ();
 sg13g2_decap_8 FILLER_3_2722 ();
 sg13g2_decap_8 FILLER_3_2729 ();
 sg13g2_decap_8 FILLER_3_2736 ();
 sg13g2_decap_8 FILLER_3_2743 ();
 sg13g2_decap_8 FILLER_3_2750 ();
 sg13g2_decap_8 FILLER_3_2757 ();
 sg13g2_decap_8 FILLER_3_2764 ();
 sg13g2_decap_8 FILLER_3_2771 ();
 sg13g2_decap_8 FILLER_3_2778 ();
 sg13g2_decap_8 FILLER_3_2785 ();
 sg13g2_decap_8 FILLER_3_2792 ();
 sg13g2_decap_8 FILLER_3_2799 ();
 sg13g2_decap_8 FILLER_3_2806 ();
 sg13g2_decap_8 FILLER_3_2813 ();
 sg13g2_decap_8 FILLER_3_2820 ();
 sg13g2_decap_8 FILLER_3_2827 ();
 sg13g2_decap_8 FILLER_3_2834 ();
 sg13g2_decap_8 FILLER_3_2841 ();
 sg13g2_decap_8 FILLER_3_2848 ();
 sg13g2_decap_8 FILLER_3_2855 ();
 sg13g2_decap_8 FILLER_3_2862 ();
 sg13g2_decap_8 FILLER_3_2869 ();
 sg13g2_decap_8 FILLER_3_2876 ();
 sg13g2_decap_8 FILLER_3_2883 ();
 sg13g2_decap_8 FILLER_3_2890 ();
 sg13g2_decap_8 FILLER_3_2897 ();
 sg13g2_decap_8 FILLER_3_2904 ();
 sg13g2_decap_8 FILLER_3_2911 ();
 sg13g2_decap_8 FILLER_3_2918 ();
 sg13g2_decap_8 FILLER_3_2925 ();
 sg13g2_decap_8 FILLER_3_2932 ();
 sg13g2_decap_8 FILLER_3_2939 ();
 sg13g2_decap_8 FILLER_3_2946 ();
 sg13g2_decap_8 FILLER_3_2953 ();
 sg13g2_decap_8 FILLER_3_2960 ();
 sg13g2_decap_8 FILLER_3_2967 ();
 sg13g2_decap_8 FILLER_3_2974 ();
 sg13g2_decap_8 FILLER_3_2981 ();
 sg13g2_decap_8 FILLER_3_2988 ();
 sg13g2_decap_8 FILLER_3_2995 ();
 sg13g2_decap_8 FILLER_3_3002 ();
 sg13g2_decap_8 FILLER_3_3009 ();
 sg13g2_decap_8 FILLER_3_3016 ();
 sg13g2_decap_8 FILLER_3_3023 ();
 sg13g2_decap_8 FILLER_3_3030 ();
 sg13g2_decap_8 FILLER_3_3037 ();
 sg13g2_decap_8 FILLER_3_3044 ();
 sg13g2_decap_8 FILLER_3_3051 ();
 sg13g2_decap_8 FILLER_3_3058 ();
 sg13g2_decap_8 FILLER_3_3065 ();
 sg13g2_decap_8 FILLER_3_3072 ();
 sg13g2_decap_8 FILLER_3_3079 ();
 sg13g2_decap_8 FILLER_3_3086 ();
 sg13g2_decap_8 FILLER_3_3093 ();
 sg13g2_decap_8 FILLER_3_3100 ();
 sg13g2_decap_8 FILLER_3_3107 ();
 sg13g2_decap_8 FILLER_3_3114 ();
 sg13g2_decap_8 FILLER_3_3121 ();
 sg13g2_decap_8 FILLER_3_3128 ();
 sg13g2_decap_8 FILLER_3_3135 ();
 sg13g2_decap_8 FILLER_3_3142 ();
 sg13g2_decap_8 FILLER_3_3149 ();
 sg13g2_decap_8 FILLER_3_3156 ();
 sg13g2_decap_8 FILLER_3_3163 ();
 sg13g2_decap_8 FILLER_3_3170 ();
 sg13g2_decap_8 FILLER_3_3177 ();
 sg13g2_decap_8 FILLER_3_3184 ();
 sg13g2_decap_8 FILLER_3_3191 ();
 sg13g2_decap_8 FILLER_3_3198 ();
 sg13g2_decap_8 FILLER_3_3205 ();
 sg13g2_decap_8 FILLER_3_3212 ();
 sg13g2_decap_8 FILLER_3_3219 ();
 sg13g2_decap_8 FILLER_3_3226 ();
 sg13g2_decap_8 FILLER_3_3233 ();
 sg13g2_decap_8 FILLER_3_3240 ();
 sg13g2_decap_8 FILLER_3_3247 ();
 sg13g2_decap_8 FILLER_3_3254 ();
 sg13g2_decap_8 FILLER_3_3261 ();
 sg13g2_decap_8 FILLER_3_3268 ();
 sg13g2_decap_8 FILLER_3_3275 ();
 sg13g2_decap_8 FILLER_3_3282 ();
 sg13g2_decap_8 FILLER_3_3289 ();
 sg13g2_decap_8 FILLER_3_3296 ();
 sg13g2_decap_8 FILLER_3_3303 ();
 sg13g2_decap_8 FILLER_3_3310 ();
 sg13g2_decap_8 FILLER_3_3317 ();
 sg13g2_decap_8 FILLER_3_3324 ();
 sg13g2_decap_8 FILLER_3_3331 ();
 sg13g2_decap_8 FILLER_3_3338 ();
 sg13g2_decap_8 FILLER_3_3345 ();
 sg13g2_decap_8 FILLER_3_3352 ();
 sg13g2_decap_8 FILLER_3_3359 ();
 sg13g2_decap_8 FILLER_3_3366 ();
 sg13g2_decap_8 FILLER_3_3373 ();
 sg13g2_decap_8 FILLER_3_3380 ();
 sg13g2_decap_8 FILLER_3_3387 ();
 sg13g2_decap_8 FILLER_3_3394 ();
 sg13g2_decap_8 FILLER_3_3401 ();
 sg13g2_decap_8 FILLER_3_3408 ();
 sg13g2_decap_8 FILLER_3_3415 ();
 sg13g2_decap_8 FILLER_3_3422 ();
 sg13g2_decap_8 FILLER_3_3429 ();
 sg13g2_decap_8 FILLER_3_3436 ();
 sg13g2_decap_8 FILLER_3_3443 ();
 sg13g2_decap_8 FILLER_3_3450 ();
 sg13g2_decap_8 FILLER_3_3457 ();
 sg13g2_decap_8 FILLER_3_3464 ();
 sg13g2_decap_8 FILLER_3_3471 ();
 sg13g2_decap_8 FILLER_3_3478 ();
 sg13g2_decap_8 FILLER_3_3485 ();
 sg13g2_decap_8 FILLER_3_3492 ();
 sg13g2_decap_8 FILLER_3_3499 ();
 sg13g2_decap_8 FILLER_3_3506 ();
 sg13g2_decap_8 FILLER_3_3513 ();
 sg13g2_decap_8 FILLER_3_3520 ();
 sg13g2_decap_8 FILLER_3_3527 ();
 sg13g2_decap_8 FILLER_3_3534 ();
 sg13g2_decap_8 FILLER_3_3541 ();
 sg13g2_decap_8 FILLER_3_3548 ();
 sg13g2_decap_8 FILLER_3_3555 ();
 sg13g2_decap_8 FILLER_3_3562 ();
 sg13g2_decap_8 FILLER_3_3569 ();
 sg13g2_decap_4 FILLER_3_3576 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_4 FILLER_4_574 ();
 sg13g2_fill_2 FILLER_4_578 ();
 sg13g2_fill_2 FILLER_4_627 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_4 FILLER_4_714 ();
 sg13g2_fill_1 FILLER_4_718 ();
 sg13g2_decap_8 FILLER_4_744 ();
 sg13g2_decap_8 FILLER_4_751 ();
 sg13g2_decap_4 FILLER_4_758 ();
 sg13g2_fill_1 FILLER_4_762 ();
 sg13g2_fill_2 FILLER_4_789 ();
 sg13g2_fill_1 FILLER_4_799 ();
 sg13g2_fill_1 FILLER_4_826 ();
 sg13g2_fill_1 FILLER_4_921 ();
 sg13g2_fill_2 FILLER_4_936 ();
 sg13g2_fill_1 FILLER_4_967 ();
 sg13g2_fill_1 FILLER_4_973 ();
 sg13g2_decap_4 FILLER_4_978 ();
 sg13g2_fill_2 FILLER_4_982 ();
 sg13g2_decap_8 FILLER_4_994 ();
 sg13g2_decap_8 FILLER_4_1001 ();
 sg13g2_decap_8 FILLER_4_1008 ();
 sg13g2_decap_8 FILLER_4_1015 ();
 sg13g2_fill_1 FILLER_4_1022 ();
 sg13g2_decap_4 FILLER_4_1058 ();
 sg13g2_fill_2 FILLER_4_1062 ();
 sg13g2_decap_8 FILLER_4_1105 ();
 sg13g2_decap_8 FILLER_4_1112 ();
 sg13g2_decap_8 FILLER_4_1119 ();
 sg13g2_decap_8 FILLER_4_1126 ();
 sg13g2_fill_2 FILLER_4_1133 ();
 sg13g2_fill_2 FILLER_4_1143 ();
 sg13g2_fill_2 FILLER_4_1153 ();
 sg13g2_fill_2 FILLER_4_1160 ();
 sg13g2_fill_2 FILLER_4_1178 ();
 sg13g2_fill_1 FILLER_4_1180 ();
 sg13g2_decap_4 FILLER_4_1204 ();
 sg13g2_fill_2 FILLER_4_1208 ();
 sg13g2_decap_8 FILLER_4_1260 ();
 sg13g2_decap_8 FILLER_4_1267 ();
 sg13g2_decap_4 FILLER_4_1274 ();
 sg13g2_fill_2 FILLER_4_1336 ();
 sg13g2_decap_8 FILLER_4_1415 ();
 sg13g2_decap_8 FILLER_4_1422 ();
 sg13g2_decap_4 FILLER_4_1429 ();
 sg13g2_fill_1 FILLER_4_1440 ();
 sg13g2_decap_8 FILLER_4_1456 ();
 sg13g2_decap_4 FILLER_4_1463 ();
 sg13g2_fill_2 FILLER_4_1467 ();
 sg13g2_decap_8 FILLER_4_1519 ();
 sg13g2_decap_8 FILLER_4_1526 ();
 sg13g2_fill_1 FILLER_4_1533 ();
 sg13g2_decap_8 FILLER_4_1564 ();
 sg13g2_decap_4 FILLER_4_1571 ();
 sg13g2_decap_4 FILLER_4_1613 ();
 sg13g2_fill_2 FILLER_4_1630 ();
 sg13g2_fill_1 FILLER_4_1637 ();
 sg13g2_decap_8 FILLER_4_1659 ();
 sg13g2_fill_2 FILLER_4_1666 ();
 sg13g2_fill_1 FILLER_4_1668 ();
 sg13g2_fill_2 FILLER_4_1676 ();
 sg13g2_decap_8 FILLER_4_1686 ();
 sg13g2_decap_8 FILLER_4_1693 ();
 sg13g2_decap_4 FILLER_4_1700 ();
 sg13g2_fill_2 FILLER_4_1704 ();
 sg13g2_fill_2 FILLER_4_1711 ();
 sg13g2_fill_1 FILLER_4_1720 ();
 sg13g2_decap_4 FILLER_4_1747 ();
 sg13g2_fill_2 FILLER_4_1751 ();
 sg13g2_decap_4 FILLER_4_1779 ();
 sg13g2_fill_1 FILLER_4_1783 ();
 sg13g2_decap_8 FILLER_4_1820 ();
 sg13g2_fill_2 FILLER_4_1871 ();
 sg13g2_fill_1 FILLER_4_1873 ();
 sg13g2_fill_1 FILLER_4_1879 ();
 sg13g2_decap_8 FILLER_4_1914 ();
 sg13g2_decap_8 FILLER_4_1921 ();
 sg13g2_decap_4 FILLER_4_1928 ();
 sg13g2_fill_1 FILLER_4_1932 ();
 sg13g2_decap_8 FILLER_4_1949 ();
 sg13g2_decap_8 FILLER_4_1956 ();
 sg13g2_decap_8 FILLER_4_1963 ();
 sg13g2_decap_8 FILLER_4_1970 ();
 sg13g2_fill_1 FILLER_4_1977 ();
 sg13g2_decap_4 FILLER_4_2017 ();
 sg13g2_decap_8 FILLER_4_2033 ();
 sg13g2_fill_1 FILLER_4_2040 ();
 sg13g2_fill_2 FILLER_4_2046 ();
 sg13g2_fill_1 FILLER_4_2048 ();
 sg13g2_fill_1 FILLER_4_2053 ();
 sg13g2_decap_8 FILLER_4_2058 ();
 sg13g2_decap_8 FILLER_4_2065 ();
 sg13g2_decap_8 FILLER_4_2072 ();
 sg13g2_decap_8 FILLER_4_2079 ();
 sg13g2_fill_1 FILLER_4_2086 ();
 sg13g2_fill_2 FILLER_4_2092 ();
 sg13g2_decap_8 FILLER_4_2128 ();
 sg13g2_decap_4 FILLER_4_2135 ();
 sg13g2_fill_1 FILLER_4_2139 ();
 sg13g2_decap_4 FILLER_4_2148 ();
 sg13g2_fill_1 FILLER_4_2152 ();
 sg13g2_decap_4 FILLER_4_2178 ();
 sg13g2_decap_8 FILLER_4_2186 ();
 sg13g2_decap_8 FILLER_4_2193 ();
 sg13g2_decap_8 FILLER_4_2200 ();
 sg13g2_decap_4 FILLER_4_2207 ();
 sg13g2_decap_4 FILLER_4_2220 ();
 sg13g2_decap_8 FILLER_4_2244 ();
 sg13g2_decap_8 FILLER_4_2282 ();
 sg13g2_decap_8 FILLER_4_2289 ();
 sg13g2_decap_8 FILLER_4_2296 ();
 sg13g2_decap_8 FILLER_4_2303 ();
 sg13g2_decap_8 FILLER_4_2310 ();
 sg13g2_fill_1 FILLER_4_2317 ();
 sg13g2_decap_8 FILLER_4_2348 ();
 sg13g2_decap_4 FILLER_4_2355 ();
 sg13g2_fill_2 FILLER_4_2359 ();
 sg13g2_fill_1 FILLER_4_2369 ();
 sg13g2_decap_8 FILLER_4_2385 ();
 sg13g2_decap_8 FILLER_4_2392 ();
 sg13g2_decap_8 FILLER_4_2404 ();
 sg13g2_decap_8 FILLER_4_2411 ();
 sg13g2_fill_1 FILLER_4_2444 ();
 sg13g2_fill_2 FILLER_4_2450 ();
 sg13g2_fill_1 FILLER_4_2452 ();
 sg13g2_fill_2 FILLER_4_2460 ();
 sg13g2_decap_8 FILLER_4_2510 ();
 sg13g2_decap_8 FILLER_4_2517 ();
 sg13g2_decap_8 FILLER_4_2524 ();
 sg13g2_decap_8 FILLER_4_2531 ();
 sg13g2_decap_8 FILLER_4_2538 ();
 sg13g2_decap_8 FILLER_4_2545 ();
 sg13g2_decap_8 FILLER_4_2552 ();
 sg13g2_decap_8 FILLER_4_2559 ();
 sg13g2_decap_8 FILLER_4_2566 ();
 sg13g2_decap_8 FILLER_4_2573 ();
 sg13g2_decap_8 FILLER_4_2580 ();
 sg13g2_decap_8 FILLER_4_2587 ();
 sg13g2_decap_8 FILLER_4_2594 ();
 sg13g2_decap_8 FILLER_4_2601 ();
 sg13g2_decap_8 FILLER_4_2608 ();
 sg13g2_decap_8 FILLER_4_2615 ();
 sg13g2_decap_8 FILLER_4_2622 ();
 sg13g2_decap_8 FILLER_4_2629 ();
 sg13g2_decap_8 FILLER_4_2636 ();
 sg13g2_decap_8 FILLER_4_2643 ();
 sg13g2_decap_8 FILLER_4_2650 ();
 sg13g2_decap_8 FILLER_4_2657 ();
 sg13g2_decap_8 FILLER_4_2664 ();
 sg13g2_decap_8 FILLER_4_2671 ();
 sg13g2_decap_8 FILLER_4_2678 ();
 sg13g2_decap_8 FILLER_4_2685 ();
 sg13g2_decap_8 FILLER_4_2692 ();
 sg13g2_decap_8 FILLER_4_2699 ();
 sg13g2_decap_8 FILLER_4_2706 ();
 sg13g2_decap_8 FILLER_4_2713 ();
 sg13g2_decap_8 FILLER_4_2720 ();
 sg13g2_decap_8 FILLER_4_2727 ();
 sg13g2_decap_8 FILLER_4_2734 ();
 sg13g2_decap_8 FILLER_4_2741 ();
 sg13g2_decap_8 FILLER_4_2748 ();
 sg13g2_decap_8 FILLER_4_2755 ();
 sg13g2_decap_8 FILLER_4_2762 ();
 sg13g2_decap_8 FILLER_4_2769 ();
 sg13g2_decap_8 FILLER_4_2776 ();
 sg13g2_decap_8 FILLER_4_2783 ();
 sg13g2_decap_8 FILLER_4_2790 ();
 sg13g2_decap_8 FILLER_4_2797 ();
 sg13g2_decap_8 FILLER_4_2804 ();
 sg13g2_decap_8 FILLER_4_2811 ();
 sg13g2_decap_8 FILLER_4_2818 ();
 sg13g2_decap_8 FILLER_4_2825 ();
 sg13g2_decap_8 FILLER_4_2832 ();
 sg13g2_decap_8 FILLER_4_2839 ();
 sg13g2_decap_8 FILLER_4_2846 ();
 sg13g2_decap_8 FILLER_4_2853 ();
 sg13g2_decap_8 FILLER_4_2860 ();
 sg13g2_decap_8 FILLER_4_2867 ();
 sg13g2_decap_8 FILLER_4_2874 ();
 sg13g2_decap_8 FILLER_4_2881 ();
 sg13g2_decap_8 FILLER_4_2888 ();
 sg13g2_decap_8 FILLER_4_2895 ();
 sg13g2_decap_8 FILLER_4_2902 ();
 sg13g2_decap_8 FILLER_4_2909 ();
 sg13g2_decap_8 FILLER_4_2916 ();
 sg13g2_decap_8 FILLER_4_2923 ();
 sg13g2_decap_8 FILLER_4_2930 ();
 sg13g2_decap_8 FILLER_4_2937 ();
 sg13g2_decap_8 FILLER_4_2944 ();
 sg13g2_decap_8 FILLER_4_2951 ();
 sg13g2_decap_8 FILLER_4_2958 ();
 sg13g2_decap_8 FILLER_4_2965 ();
 sg13g2_decap_8 FILLER_4_2972 ();
 sg13g2_decap_8 FILLER_4_2979 ();
 sg13g2_decap_8 FILLER_4_2986 ();
 sg13g2_decap_8 FILLER_4_2993 ();
 sg13g2_decap_8 FILLER_4_3000 ();
 sg13g2_decap_8 FILLER_4_3007 ();
 sg13g2_decap_8 FILLER_4_3014 ();
 sg13g2_decap_8 FILLER_4_3021 ();
 sg13g2_decap_8 FILLER_4_3028 ();
 sg13g2_decap_8 FILLER_4_3035 ();
 sg13g2_decap_8 FILLER_4_3042 ();
 sg13g2_decap_8 FILLER_4_3049 ();
 sg13g2_decap_8 FILLER_4_3056 ();
 sg13g2_decap_8 FILLER_4_3063 ();
 sg13g2_decap_8 FILLER_4_3070 ();
 sg13g2_decap_8 FILLER_4_3077 ();
 sg13g2_decap_8 FILLER_4_3084 ();
 sg13g2_decap_8 FILLER_4_3091 ();
 sg13g2_decap_8 FILLER_4_3098 ();
 sg13g2_decap_8 FILLER_4_3105 ();
 sg13g2_decap_8 FILLER_4_3112 ();
 sg13g2_decap_8 FILLER_4_3119 ();
 sg13g2_decap_8 FILLER_4_3126 ();
 sg13g2_decap_8 FILLER_4_3133 ();
 sg13g2_decap_8 FILLER_4_3140 ();
 sg13g2_decap_8 FILLER_4_3147 ();
 sg13g2_decap_8 FILLER_4_3154 ();
 sg13g2_decap_8 FILLER_4_3161 ();
 sg13g2_decap_8 FILLER_4_3168 ();
 sg13g2_decap_8 FILLER_4_3175 ();
 sg13g2_decap_8 FILLER_4_3182 ();
 sg13g2_decap_8 FILLER_4_3189 ();
 sg13g2_decap_8 FILLER_4_3196 ();
 sg13g2_decap_8 FILLER_4_3203 ();
 sg13g2_decap_8 FILLER_4_3210 ();
 sg13g2_decap_8 FILLER_4_3217 ();
 sg13g2_decap_8 FILLER_4_3224 ();
 sg13g2_decap_8 FILLER_4_3231 ();
 sg13g2_decap_8 FILLER_4_3238 ();
 sg13g2_decap_8 FILLER_4_3245 ();
 sg13g2_decap_8 FILLER_4_3252 ();
 sg13g2_decap_8 FILLER_4_3259 ();
 sg13g2_decap_8 FILLER_4_3266 ();
 sg13g2_decap_8 FILLER_4_3273 ();
 sg13g2_decap_8 FILLER_4_3280 ();
 sg13g2_decap_8 FILLER_4_3287 ();
 sg13g2_decap_8 FILLER_4_3294 ();
 sg13g2_decap_8 FILLER_4_3301 ();
 sg13g2_decap_8 FILLER_4_3308 ();
 sg13g2_decap_8 FILLER_4_3315 ();
 sg13g2_decap_8 FILLER_4_3322 ();
 sg13g2_decap_8 FILLER_4_3329 ();
 sg13g2_decap_8 FILLER_4_3336 ();
 sg13g2_decap_8 FILLER_4_3343 ();
 sg13g2_decap_8 FILLER_4_3350 ();
 sg13g2_decap_8 FILLER_4_3357 ();
 sg13g2_decap_8 FILLER_4_3364 ();
 sg13g2_decap_8 FILLER_4_3371 ();
 sg13g2_decap_8 FILLER_4_3378 ();
 sg13g2_decap_8 FILLER_4_3385 ();
 sg13g2_decap_8 FILLER_4_3392 ();
 sg13g2_decap_8 FILLER_4_3399 ();
 sg13g2_decap_8 FILLER_4_3406 ();
 sg13g2_decap_8 FILLER_4_3413 ();
 sg13g2_decap_8 FILLER_4_3420 ();
 sg13g2_decap_8 FILLER_4_3427 ();
 sg13g2_decap_8 FILLER_4_3434 ();
 sg13g2_decap_8 FILLER_4_3441 ();
 sg13g2_decap_8 FILLER_4_3448 ();
 sg13g2_decap_8 FILLER_4_3455 ();
 sg13g2_decap_8 FILLER_4_3462 ();
 sg13g2_decap_8 FILLER_4_3469 ();
 sg13g2_decap_8 FILLER_4_3476 ();
 sg13g2_decap_8 FILLER_4_3483 ();
 sg13g2_decap_8 FILLER_4_3490 ();
 sg13g2_decap_8 FILLER_4_3497 ();
 sg13g2_decap_8 FILLER_4_3504 ();
 sg13g2_decap_8 FILLER_4_3511 ();
 sg13g2_decap_8 FILLER_4_3518 ();
 sg13g2_decap_8 FILLER_4_3525 ();
 sg13g2_decap_8 FILLER_4_3532 ();
 sg13g2_decap_8 FILLER_4_3539 ();
 sg13g2_decap_8 FILLER_4_3546 ();
 sg13g2_decap_8 FILLER_4_3553 ();
 sg13g2_decap_8 FILLER_4_3560 ();
 sg13g2_decap_8 FILLER_4_3567 ();
 sg13g2_decap_4 FILLER_4_3574 ();
 sg13g2_fill_2 FILLER_4_3578 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_fill_1 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_638 ();
 sg13g2_decap_8 FILLER_5_645 ();
 sg13g2_decap_4 FILLER_5_652 ();
 sg13g2_fill_2 FILLER_5_656 ();
 sg13g2_decap_8 FILLER_5_704 ();
 sg13g2_decap_8 FILLER_5_711 ();
 sg13g2_fill_1 FILLER_5_718 ();
 sg13g2_decap_8 FILLER_5_743 ();
 sg13g2_fill_2 FILLER_5_750 ();
 sg13g2_fill_1 FILLER_5_752 ();
 sg13g2_decap_8 FILLER_5_779 ();
 sg13g2_decap_4 FILLER_5_786 ();
 sg13g2_fill_1 FILLER_5_790 ();
 sg13g2_decap_8 FILLER_5_799 ();
 sg13g2_decap_8 FILLER_5_806 ();
 sg13g2_decap_8 FILLER_5_813 ();
 sg13g2_decap_4 FILLER_5_820 ();
 sg13g2_fill_1 FILLER_5_824 ();
 sg13g2_decap_8 FILLER_5_867 ();
 sg13g2_fill_2 FILLER_5_874 ();
 sg13g2_fill_1 FILLER_5_876 ();
 sg13g2_fill_2 FILLER_5_989 ();
 sg13g2_fill_1 FILLER_5_991 ();
 sg13g2_fill_2 FILLER_5_997 ();
 sg13g2_fill_2 FILLER_5_1007 ();
 sg13g2_fill_1 FILLER_5_1009 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_decap_4 FILLER_5_1026 ();
 sg13g2_fill_2 FILLER_5_1030 ();
 sg13g2_decap_4 FILLER_5_1053 ();
 sg13g2_fill_1 FILLER_5_1057 ();
 sg13g2_fill_1 FILLER_5_1062 ();
 sg13g2_decap_8 FILLER_5_1112 ();
 sg13g2_fill_2 FILLER_5_1119 ();
 sg13g2_fill_1 FILLER_5_1147 ();
 sg13g2_decap_4 FILLER_5_1205 ();
 sg13g2_fill_1 FILLER_5_1209 ();
 sg13g2_decap_8 FILLER_5_1263 ();
 sg13g2_decap_8 FILLER_5_1270 ();
 sg13g2_decap_4 FILLER_5_1277 ();
 sg13g2_fill_1 FILLER_5_1289 ();
 sg13g2_decap_8 FILLER_5_1297 ();
 sg13g2_decap_8 FILLER_5_1304 ();
 sg13g2_decap_8 FILLER_5_1311 ();
 sg13g2_fill_1 FILLER_5_1318 ();
 sg13g2_decap_8 FILLER_5_1343 ();
 sg13g2_decap_8 FILLER_5_1350 ();
 sg13g2_decap_8 FILLER_5_1357 ();
 sg13g2_decap_8 FILLER_5_1364 ();
 sg13g2_fill_2 FILLER_5_1371 ();
 sg13g2_fill_2 FILLER_5_1383 ();
 sg13g2_decap_8 FILLER_5_1453 ();
 sg13g2_decap_8 FILLER_5_1460 ();
 sg13g2_decap_8 FILLER_5_1467 ();
 sg13g2_fill_2 FILLER_5_1474 ();
 sg13g2_fill_1 FILLER_5_1476 ();
 sg13g2_decap_8 FILLER_5_1511 ();
 sg13g2_decap_8 FILLER_5_1518 ();
 sg13g2_decap_4 FILLER_5_1525 ();
 sg13g2_fill_1 FILLER_5_1529 ();
 sg13g2_fill_2 FILLER_5_1564 ();
 sg13g2_fill_1 FILLER_5_1566 ();
 sg13g2_fill_1 FILLER_5_1605 ();
 sg13g2_decap_4 FILLER_5_1614 ();
 sg13g2_fill_2 FILLER_5_1618 ();
 sg13g2_decap_8 FILLER_5_1686 ();
 sg13g2_fill_1 FILLER_5_1706 ();
 sg13g2_fill_1 FILLER_5_1735 ();
 sg13g2_decap_8 FILLER_5_1762 ();
 sg13g2_decap_4 FILLER_5_1774 ();
 sg13g2_fill_2 FILLER_5_1778 ();
 sg13g2_decap_4 FILLER_5_1801 ();
 sg13g2_fill_2 FILLER_5_1805 ();
 sg13g2_fill_1 FILLER_5_1815 ();
 sg13g2_decap_8 FILLER_5_1825 ();
 sg13g2_decap_4 FILLER_5_1832 ();
 sg13g2_fill_2 FILLER_5_1836 ();
 sg13g2_decap_8 FILLER_5_1870 ();
 sg13g2_decap_8 FILLER_5_1877 ();
 sg13g2_decap_8 FILLER_5_1884 ();
 sg13g2_decap_4 FILLER_5_1891 ();
 sg13g2_fill_2 FILLER_5_1895 ();
 sg13g2_fill_1 FILLER_5_1923 ();
 sg13g2_decap_8 FILLER_5_1962 ();
 sg13g2_decap_8 FILLER_5_1969 ();
 sg13g2_fill_2 FILLER_5_1976 ();
 sg13g2_fill_1 FILLER_5_1978 ();
 sg13g2_fill_2 FILLER_5_2013 ();
 sg13g2_decap_8 FILLER_5_2067 ();
 sg13g2_decap_8 FILLER_5_2074 ();
 sg13g2_fill_1 FILLER_5_2081 ();
 sg13g2_decap_8 FILLER_5_2121 ();
 sg13g2_decap_8 FILLER_5_2128 ();
 sg13g2_decap_4 FILLER_5_2169 ();
 sg13g2_fill_2 FILLER_5_2173 ();
 sg13g2_decap_8 FILLER_5_2195 ();
 sg13g2_fill_2 FILLER_5_2230 ();
 sg13g2_fill_1 FILLER_5_2232 ();
 sg13g2_fill_2 FILLER_5_2259 ();
 sg13g2_fill_1 FILLER_5_2266 ();
 sg13g2_decap_8 FILLER_5_2275 ();
 sg13g2_decap_8 FILLER_5_2282 ();
 sg13g2_decap_8 FILLER_5_2289 ();
 sg13g2_decap_8 FILLER_5_2296 ();
 sg13g2_fill_2 FILLER_5_2303 ();
 sg13g2_fill_1 FILLER_5_2305 ();
 sg13g2_decap_8 FILLER_5_2341 ();
 sg13g2_decap_4 FILLER_5_2348 ();
 sg13g2_fill_2 FILLER_5_2352 ();
 sg13g2_decap_8 FILLER_5_2358 ();
 sg13g2_decap_8 FILLER_5_2365 ();
 sg13g2_decap_8 FILLER_5_2372 ();
 sg13g2_decap_8 FILLER_5_2379 ();
 sg13g2_decap_8 FILLER_5_2386 ();
 sg13g2_fill_2 FILLER_5_2393 ();
 sg13g2_decap_8 FILLER_5_2418 ();
 sg13g2_decap_4 FILLER_5_2425 ();
 sg13g2_decap_4 FILLER_5_2434 ();
 sg13g2_fill_1 FILLER_5_2438 ();
 sg13g2_fill_1 FILLER_5_2447 ();
 sg13g2_decap_4 FILLER_5_2456 ();
 sg13g2_decap_8 FILLER_5_2499 ();
 sg13g2_decap_8 FILLER_5_2506 ();
 sg13g2_decap_8 FILLER_5_2513 ();
 sg13g2_decap_8 FILLER_5_2520 ();
 sg13g2_decap_8 FILLER_5_2527 ();
 sg13g2_decap_8 FILLER_5_2534 ();
 sg13g2_decap_8 FILLER_5_2541 ();
 sg13g2_decap_8 FILLER_5_2548 ();
 sg13g2_decap_8 FILLER_5_2555 ();
 sg13g2_decap_8 FILLER_5_2562 ();
 sg13g2_decap_8 FILLER_5_2569 ();
 sg13g2_decap_8 FILLER_5_2576 ();
 sg13g2_decap_8 FILLER_5_2583 ();
 sg13g2_decap_8 FILLER_5_2590 ();
 sg13g2_decap_8 FILLER_5_2597 ();
 sg13g2_decap_8 FILLER_5_2604 ();
 sg13g2_decap_8 FILLER_5_2611 ();
 sg13g2_decap_8 FILLER_5_2618 ();
 sg13g2_decap_8 FILLER_5_2625 ();
 sg13g2_decap_8 FILLER_5_2632 ();
 sg13g2_decap_8 FILLER_5_2639 ();
 sg13g2_decap_8 FILLER_5_2646 ();
 sg13g2_decap_8 FILLER_5_2653 ();
 sg13g2_decap_8 FILLER_5_2660 ();
 sg13g2_decap_8 FILLER_5_2667 ();
 sg13g2_decap_8 FILLER_5_2674 ();
 sg13g2_decap_8 FILLER_5_2681 ();
 sg13g2_decap_8 FILLER_5_2688 ();
 sg13g2_decap_8 FILLER_5_2695 ();
 sg13g2_decap_8 FILLER_5_2702 ();
 sg13g2_decap_8 FILLER_5_2709 ();
 sg13g2_decap_8 FILLER_5_2716 ();
 sg13g2_decap_8 FILLER_5_2723 ();
 sg13g2_decap_8 FILLER_5_2730 ();
 sg13g2_decap_8 FILLER_5_2737 ();
 sg13g2_decap_8 FILLER_5_2744 ();
 sg13g2_decap_8 FILLER_5_2751 ();
 sg13g2_decap_8 FILLER_5_2758 ();
 sg13g2_decap_8 FILLER_5_2765 ();
 sg13g2_decap_8 FILLER_5_2772 ();
 sg13g2_decap_8 FILLER_5_2779 ();
 sg13g2_decap_8 FILLER_5_2786 ();
 sg13g2_decap_8 FILLER_5_2793 ();
 sg13g2_decap_8 FILLER_5_2800 ();
 sg13g2_decap_8 FILLER_5_2807 ();
 sg13g2_decap_8 FILLER_5_2814 ();
 sg13g2_decap_8 FILLER_5_2821 ();
 sg13g2_decap_8 FILLER_5_2828 ();
 sg13g2_decap_8 FILLER_5_2835 ();
 sg13g2_decap_8 FILLER_5_2842 ();
 sg13g2_decap_8 FILLER_5_2849 ();
 sg13g2_decap_8 FILLER_5_2856 ();
 sg13g2_decap_8 FILLER_5_2863 ();
 sg13g2_decap_8 FILLER_5_2870 ();
 sg13g2_decap_8 FILLER_5_2877 ();
 sg13g2_decap_8 FILLER_5_2884 ();
 sg13g2_decap_8 FILLER_5_2891 ();
 sg13g2_decap_8 FILLER_5_2898 ();
 sg13g2_decap_8 FILLER_5_2905 ();
 sg13g2_decap_8 FILLER_5_2912 ();
 sg13g2_decap_8 FILLER_5_2919 ();
 sg13g2_decap_8 FILLER_5_2926 ();
 sg13g2_decap_8 FILLER_5_2933 ();
 sg13g2_decap_8 FILLER_5_2940 ();
 sg13g2_decap_8 FILLER_5_2947 ();
 sg13g2_decap_8 FILLER_5_2954 ();
 sg13g2_decap_8 FILLER_5_2961 ();
 sg13g2_decap_8 FILLER_5_2968 ();
 sg13g2_decap_8 FILLER_5_2975 ();
 sg13g2_decap_8 FILLER_5_2982 ();
 sg13g2_decap_8 FILLER_5_2989 ();
 sg13g2_decap_8 FILLER_5_2996 ();
 sg13g2_decap_8 FILLER_5_3003 ();
 sg13g2_decap_8 FILLER_5_3010 ();
 sg13g2_decap_8 FILLER_5_3017 ();
 sg13g2_decap_8 FILLER_5_3024 ();
 sg13g2_decap_8 FILLER_5_3031 ();
 sg13g2_decap_8 FILLER_5_3038 ();
 sg13g2_decap_8 FILLER_5_3045 ();
 sg13g2_decap_8 FILLER_5_3052 ();
 sg13g2_decap_8 FILLER_5_3059 ();
 sg13g2_decap_8 FILLER_5_3066 ();
 sg13g2_decap_8 FILLER_5_3073 ();
 sg13g2_decap_8 FILLER_5_3080 ();
 sg13g2_decap_8 FILLER_5_3087 ();
 sg13g2_decap_8 FILLER_5_3094 ();
 sg13g2_decap_8 FILLER_5_3101 ();
 sg13g2_decap_8 FILLER_5_3108 ();
 sg13g2_decap_8 FILLER_5_3115 ();
 sg13g2_decap_8 FILLER_5_3122 ();
 sg13g2_decap_8 FILLER_5_3129 ();
 sg13g2_decap_8 FILLER_5_3136 ();
 sg13g2_decap_8 FILLER_5_3143 ();
 sg13g2_decap_8 FILLER_5_3150 ();
 sg13g2_decap_8 FILLER_5_3157 ();
 sg13g2_decap_8 FILLER_5_3164 ();
 sg13g2_decap_8 FILLER_5_3171 ();
 sg13g2_decap_8 FILLER_5_3178 ();
 sg13g2_decap_8 FILLER_5_3185 ();
 sg13g2_decap_8 FILLER_5_3192 ();
 sg13g2_decap_8 FILLER_5_3199 ();
 sg13g2_decap_8 FILLER_5_3206 ();
 sg13g2_decap_8 FILLER_5_3213 ();
 sg13g2_decap_8 FILLER_5_3220 ();
 sg13g2_decap_8 FILLER_5_3227 ();
 sg13g2_decap_8 FILLER_5_3234 ();
 sg13g2_decap_8 FILLER_5_3241 ();
 sg13g2_decap_8 FILLER_5_3248 ();
 sg13g2_decap_8 FILLER_5_3255 ();
 sg13g2_decap_8 FILLER_5_3262 ();
 sg13g2_decap_8 FILLER_5_3269 ();
 sg13g2_decap_8 FILLER_5_3276 ();
 sg13g2_decap_8 FILLER_5_3283 ();
 sg13g2_decap_8 FILLER_5_3290 ();
 sg13g2_decap_8 FILLER_5_3297 ();
 sg13g2_decap_8 FILLER_5_3304 ();
 sg13g2_decap_8 FILLER_5_3311 ();
 sg13g2_decap_8 FILLER_5_3318 ();
 sg13g2_decap_8 FILLER_5_3325 ();
 sg13g2_decap_8 FILLER_5_3332 ();
 sg13g2_decap_8 FILLER_5_3339 ();
 sg13g2_decap_8 FILLER_5_3346 ();
 sg13g2_decap_8 FILLER_5_3353 ();
 sg13g2_decap_8 FILLER_5_3360 ();
 sg13g2_decap_8 FILLER_5_3367 ();
 sg13g2_decap_8 FILLER_5_3374 ();
 sg13g2_decap_8 FILLER_5_3381 ();
 sg13g2_decap_8 FILLER_5_3388 ();
 sg13g2_decap_8 FILLER_5_3395 ();
 sg13g2_decap_8 FILLER_5_3402 ();
 sg13g2_decap_8 FILLER_5_3409 ();
 sg13g2_decap_8 FILLER_5_3416 ();
 sg13g2_decap_8 FILLER_5_3423 ();
 sg13g2_decap_8 FILLER_5_3430 ();
 sg13g2_decap_8 FILLER_5_3437 ();
 sg13g2_decap_8 FILLER_5_3444 ();
 sg13g2_decap_8 FILLER_5_3451 ();
 sg13g2_decap_8 FILLER_5_3458 ();
 sg13g2_decap_8 FILLER_5_3465 ();
 sg13g2_decap_8 FILLER_5_3472 ();
 sg13g2_decap_8 FILLER_5_3479 ();
 sg13g2_decap_8 FILLER_5_3486 ();
 sg13g2_decap_8 FILLER_5_3493 ();
 sg13g2_decap_8 FILLER_5_3500 ();
 sg13g2_decap_8 FILLER_5_3507 ();
 sg13g2_decap_8 FILLER_5_3514 ();
 sg13g2_decap_8 FILLER_5_3521 ();
 sg13g2_decap_8 FILLER_5_3528 ();
 sg13g2_decap_8 FILLER_5_3535 ();
 sg13g2_decap_8 FILLER_5_3542 ();
 sg13g2_decap_8 FILLER_5_3549 ();
 sg13g2_decap_8 FILLER_5_3556 ();
 sg13g2_decap_8 FILLER_5_3563 ();
 sg13g2_decap_8 FILLER_5_3570 ();
 sg13g2_fill_2 FILLER_5_3577 ();
 sg13g2_fill_1 FILLER_5_3579 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_4 FILLER_6_553 ();
 sg13g2_fill_1 FILLER_6_557 ();
 sg13g2_fill_1 FILLER_6_574 ();
 sg13g2_fill_2 FILLER_6_580 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_4 FILLER_6_648 ();
 sg13g2_fill_2 FILLER_6_652 ();
 sg13g2_decap_4 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_684 ();
 sg13g2_fill_2 FILLER_6_696 ();
 sg13g2_fill_2 FILLER_6_711 ();
 sg13g2_fill_1 FILLER_6_713 ();
 sg13g2_decap_8 FILLER_6_755 ();
 sg13g2_fill_2 FILLER_6_762 ();
 sg13g2_fill_1 FILLER_6_764 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_861 ();
 sg13g2_fill_1 FILLER_6_868 ();
 sg13g2_decap_8 FILLER_6_899 ();
 sg13g2_decap_4 FILLER_6_910 ();
 sg13g2_fill_1 FILLER_6_914 ();
 sg13g2_decap_4 FILLER_6_920 ();
 sg13g2_fill_2 FILLER_6_924 ();
 sg13g2_decap_8 FILLER_6_934 ();
 sg13g2_fill_2 FILLER_6_941 ();
 sg13g2_fill_1 FILLER_6_943 ();
 sg13g2_fill_2 FILLER_6_983 ();
 sg13g2_fill_2 FILLER_6_990 ();
 sg13g2_decap_8 FILLER_6_1028 ();
 sg13g2_fill_1 FILLER_6_1035 ();
 sg13g2_decap_8 FILLER_6_1105 ();
 sg13g2_decap_8 FILLER_6_1112 ();
 sg13g2_decap_4 FILLER_6_1119 ();
 sg13g2_decap_4 FILLER_6_1157 ();
 sg13g2_decap_8 FILLER_6_1173 ();
 sg13g2_decap_8 FILLER_6_1180 ();
 sg13g2_decap_8 FILLER_6_1187 ();
 sg13g2_decap_8 FILLER_6_1194 ();
 sg13g2_decap_8 FILLER_6_1201 ();
 sg13g2_decap_8 FILLER_6_1208 ();
 sg13g2_decap_4 FILLER_6_1215 ();
 sg13g2_fill_2 FILLER_6_1219 ();
 sg13g2_decap_8 FILLER_6_1303 ();
 sg13g2_decap_8 FILLER_6_1310 ();
 sg13g2_decap_4 FILLER_6_1317 ();
 sg13g2_fill_2 FILLER_6_1321 ();
 sg13g2_decap_8 FILLER_6_1349 ();
 sg13g2_decap_8 FILLER_6_1356 ();
 sg13g2_decap_8 FILLER_6_1363 ();
 sg13g2_fill_1 FILLER_6_1370 ();
 sg13g2_fill_2 FILLER_6_1387 ();
 sg13g2_fill_1 FILLER_6_1389 ();
 sg13g2_decap_4 FILLER_6_1403 ();
 sg13g2_decap_8 FILLER_6_1459 ();
 sg13g2_decap_8 FILLER_6_1466 ();
 sg13g2_decap_8 FILLER_6_1473 ();
 sg13g2_fill_2 FILLER_6_1480 ();
 sg13g2_decap_8 FILLER_6_1507 ();
 sg13g2_decap_4 FILLER_6_1514 ();
 sg13g2_fill_2 FILLER_6_1518 ();
 sg13g2_fill_2 FILLER_6_1574 ();
 sg13g2_decap_8 FILLER_6_1633 ();
 sg13g2_decap_4 FILLER_6_1640 ();
 sg13g2_fill_1 FILLER_6_1644 ();
 sg13g2_fill_1 FILLER_6_1649 ();
 sg13g2_decap_8 FILLER_6_1676 ();
 sg13g2_decap_4 FILLER_6_1683 ();
 sg13g2_decap_4 FILLER_6_1729 ();
 sg13g2_fill_2 FILLER_6_1733 ();
 sg13g2_decap_8 FILLER_6_1740 ();
 sg13g2_decap_4 FILLER_6_1747 ();
 sg13g2_fill_2 FILLER_6_1751 ();
 sg13g2_decap_8 FILLER_6_1756 ();
 sg13g2_decap_8 FILLER_6_1763 ();
 sg13g2_decap_8 FILLER_6_1770 ();
 sg13g2_decap_8 FILLER_6_1777 ();
 sg13g2_decap_8 FILLER_6_1784 ();
 sg13g2_decap_8 FILLER_6_1791 ();
 sg13g2_fill_1 FILLER_6_1798 ();
 sg13g2_decap_8 FILLER_6_1833 ();
 sg13g2_decap_4 FILLER_6_1840 ();
 sg13g2_fill_1 FILLER_6_1844 ();
 sg13g2_decap_8 FILLER_6_1883 ();
 sg13g2_fill_2 FILLER_6_1890 ();
 sg13g2_fill_1 FILLER_6_1892 ();
 sg13g2_decap_8 FILLER_6_1898 ();
 sg13g2_decap_4 FILLER_6_1905 ();
 sg13g2_fill_2 FILLER_6_1909 ();
 sg13g2_fill_1 FILLER_6_1919 ();
 sg13g2_decap_8 FILLER_6_1969 ();
 sg13g2_fill_2 FILLER_6_1976 ();
 sg13g2_decap_8 FILLER_6_2017 ();
 sg13g2_fill_2 FILLER_6_2024 ();
 sg13g2_fill_1 FILLER_6_2026 ();
 sg13g2_fill_2 FILLER_6_2078 ();
 sg13g2_fill_2 FILLER_6_2113 ();
 sg13g2_fill_1 FILLER_6_2115 ();
 sg13g2_decap_8 FILLER_6_2124 ();
 sg13g2_decap_8 FILLER_6_2131 ();
 sg13g2_decap_8 FILLER_6_2138 ();
 sg13g2_decap_8 FILLER_6_2145 ();
 sg13g2_fill_2 FILLER_6_2152 ();
 sg13g2_decap_8 FILLER_6_2161 ();
 sg13g2_fill_2 FILLER_6_2168 ();
 sg13g2_fill_1 FILLER_6_2201 ();
 sg13g2_decap_8 FILLER_6_2306 ();
 sg13g2_decap_8 FILLER_6_2321 ();
 sg13g2_fill_2 FILLER_6_2328 ();
 sg13g2_fill_1 FILLER_6_2330 ();
 sg13g2_decap_4 FILLER_6_2343 ();
 sg13g2_fill_1 FILLER_6_2347 ();
 sg13g2_fill_1 FILLER_6_2365 ();
 sg13g2_fill_2 FILLER_6_2392 ();
 sg13g2_fill_1 FILLER_6_2394 ();
 sg13g2_decap_8 FILLER_6_2421 ();
 sg13g2_decap_4 FILLER_6_2433 ();
 sg13g2_decap_8 FILLER_6_2463 ();
 sg13g2_fill_2 FILLER_6_2470 ();
 sg13g2_fill_1 FILLER_6_2472 ();
 sg13g2_decap_8 FILLER_6_2499 ();
 sg13g2_decap_8 FILLER_6_2506 ();
 sg13g2_fill_2 FILLER_6_2513 ();
 sg13g2_decap_8 FILLER_6_2537 ();
 sg13g2_decap_8 FILLER_6_2544 ();
 sg13g2_decap_8 FILLER_6_2551 ();
 sg13g2_decap_8 FILLER_6_2558 ();
 sg13g2_decap_8 FILLER_6_2565 ();
 sg13g2_decap_8 FILLER_6_2572 ();
 sg13g2_decap_8 FILLER_6_2579 ();
 sg13g2_decap_8 FILLER_6_2586 ();
 sg13g2_decap_8 FILLER_6_2593 ();
 sg13g2_decap_8 FILLER_6_2600 ();
 sg13g2_decap_8 FILLER_6_2607 ();
 sg13g2_decap_8 FILLER_6_2614 ();
 sg13g2_decap_8 FILLER_6_2621 ();
 sg13g2_decap_8 FILLER_6_2628 ();
 sg13g2_decap_8 FILLER_6_2635 ();
 sg13g2_decap_8 FILLER_6_2642 ();
 sg13g2_decap_8 FILLER_6_2649 ();
 sg13g2_decap_8 FILLER_6_2656 ();
 sg13g2_decap_8 FILLER_6_2663 ();
 sg13g2_decap_8 FILLER_6_2670 ();
 sg13g2_decap_8 FILLER_6_2677 ();
 sg13g2_decap_8 FILLER_6_2684 ();
 sg13g2_decap_8 FILLER_6_2691 ();
 sg13g2_decap_8 FILLER_6_2698 ();
 sg13g2_decap_8 FILLER_6_2705 ();
 sg13g2_decap_8 FILLER_6_2712 ();
 sg13g2_decap_8 FILLER_6_2719 ();
 sg13g2_decap_8 FILLER_6_2726 ();
 sg13g2_decap_8 FILLER_6_2733 ();
 sg13g2_decap_8 FILLER_6_2740 ();
 sg13g2_decap_8 FILLER_6_2747 ();
 sg13g2_decap_8 FILLER_6_2754 ();
 sg13g2_decap_8 FILLER_6_2761 ();
 sg13g2_decap_8 FILLER_6_2768 ();
 sg13g2_decap_8 FILLER_6_2775 ();
 sg13g2_decap_8 FILLER_6_2782 ();
 sg13g2_decap_8 FILLER_6_2789 ();
 sg13g2_decap_8 FILLER_6_2796 ();
 sg13g2_decap_8 FILLER_6_2803 ();
 sg13g2_decap_8 FILLER_6_2810 ();
 sg13g2_decap_8 FILLER_6_2817 ();
 sg13g2_decap_8 FILLER_6_2824 ();
 sg13g2_decap_8 FILLER_6_2831 ();
 sg13g2_decap_8 FILLER_6_2838 ();
 sg13g2_decap_8 FILLER_6_2845 ();
 sg13g2_decap_8 FILLER_6_2852 ();
 sg13g2_decap_8 FILLER_6_2859 ();
 sg13g2_decap_8 FILLER_6_2866 ();
 sg13g2_decap_8 FILLER_6_2873 ();
 sg13g2_decap_8 FILLER_6_2880 ();
 sg13g2_decap_8 FILLER_6_2887 ();
 sg13g2_decap_8 FILLER_6_2894 ();
 sg13g2_decap_8 FILLER_6_2901 ();
 sg13g2_decap_8 FILLER_6_2908 ();
 sg13g2_decap_8 FILLER_6_2915 ();
 sg13g2_decap_8 FILLER_6_2922 ();
 sg13g2_decap_8 FILLER_6_2929 ();
 sg13g2_decap_8 FILLER_6_2936 ();
 sg13g2_decap_8 FILLER_6_2943 ();
 sg13g2_decap_8 FILLER_6_2950 ();
 sg13g2_decap_8 FILLER_6_2957 ();
 sg13g2_decap_8 FILLER_6_2964 ();
 sg13g2_decap_8 FILLER_6_2971 ();
 sg13g2_decap_8 FILLER_6_2978 ();
 sg13g2_decap_8 FILLER_6_2985 ();
 sg13g2_decap_8 FILLER_6_2992 ();
 sg13g2_decap_8 FILLER_6_2999 ();
 sg13g2_decap_8 FILLER_6_3006 ();
 sg13g2_decap_8 FILLER_6_3013 ();
 sg13g2_decap_8 FILLER_6_3020 ();
 sg13g2_decap_8 FILLER_6_3027 ();
 sg13g2_decap_8 FILLER_6_3034 ();
 sg13g2_decap_8 FILLER_6_3041 ();
 sg13g2_decap_8 FILLER_6_3048 ();
 sg13g2_decap_8 FILLER_6_3055 ();
 sg13g2_decap_8 FILLER_6_3062 ();
 sg13g2_decap_8 FILLER_6_3069 ();
 sg13g2_decap_8 FILLER_6_3076 ();
 sg13g2_decap_8 FILLER_6_3083 ();
 sg13g2_decap_8 FILLER_6_3090 ();
 sg13g2_decap_8 FILLER_6_3097 ();
 sg13g2_decap_8 FILLER_6_3104 ();
 sg13g2_decap_8 FILLER_6_3111 ();
 sg13g2_decap_8 FILLER_6_3118 ();
 sg13g2_decap_8 FILLER_6_3125 ();
 sg13g2_decap_8 FILLER_6_3132 ();
 sg13g2_decap_8 FILLER_6_3139 ();
 sg13g2_decap_8 FILLER_6_3146 ();
 sg13g2_decap_8 FILLER_6_3153 ();
 sg13g2_decap_8 FILLER_6_3160 ();
 sg13g2_decap_8 FILLER_6_3167 ();
 sg13g2_decap_8 FILLER_6_3174 ();
 sg13g2_decap_8 FILLER_6_3181 ();
 sg13g2_decap_8 FILLER_6_3188 ();
 sg13g2_decap_8 FILLER_6_3195 ();
 sg13g2_decap_8 FILLER_6_3202 ();
 sg13g2_decap_8 FILLER_6_3209 ();
 sg13g2_decap_8 FILLER_6_3216 ();
 sg13g2_decap_8 FILLER_6_3223 ();
 sg13g2_decap_8 FILLER_6_3230 ();
 sg13g2_decap_8 FILLER_6_3237 ();
 sg13g2_decap_8 FILLER_6_3244 ();
 sg13g2_decap_8 FILLER_6_3251 ();
 sg13g2_decap_8 FILLER_6_3258 ();
 sg13g2_decap_8 FILLER_6_3265 ();
 sg13g2_decap_8 FILLER_6_3272 ();
 sg13g2_decap_8 FILLER_6_3279 ();
 sg13g2_decap_8 FILLER_6_3286 ();
 sg13g2_decap_8 FILLER_6_3293 ();
 sg13g2_decap_8 FILLER_6_3300 ();
 sg13g2_decap_8 FILLER_6_3307 ();
 sg13g2_decap_8 FILLER_6_3314 ();
 sg13g2_decap_8 FILLER_6_3321 ();
 sg13g2_decap_8 FILLER_6_3328 ();
 sg13g2_decap_8 FILLER_6_3335 ();
 sg13g2_decap_8 FILLER_6_3342 ();
 sg13g2_decap_8 FILLER_6_3349 ();
 sg13g2_decap_8 FILLER_6_3356 ();
 sg13g2_decap_8 FILLER_6_3363 ();
 sg13g2_decap_8 FILLER_6_3370 ();
 sg13g2_decap_8 FILLER_6_3377 ();
 sg13g2_decap_8 FILLER_6_3384 ();
 sg13g2_decap_8 FILLER_6_3391 ();
 sg13g2_decap_8 FILLER_6_3398 ();
 sg13g2_decap_8 FILLER_6_3405 ();
 sg13g2_decap_8 FILLER_6_3412 ();
 sg13g2_decap_8 FILLER_6_3419 ();
 sg13g2_decap_8 FILLER_6_3426 ();
 sg13g2_decap_8 FILLER_6_3433 ();
 sg13g2_decap_8 FILLER_6_3440 ();
 sg13g2_decap_8 FILLER_6_3447 ();
 sg13g2_decap_8 FILLER_6_3454 ();
 sg13g2_decap_8 FILLER_6_3461 ();
 sg13g2_decap_8 FILLER_6_3468 ();
 sg13g2_decap_8 FILLER_6_3475 ();
 sg13g2_decap_8 FILLER_6_3482 ();
 sg13g2_decap_8 FILLER_6_3489 ();
 sg13g2_decap_8 FILLER_6_3496 ();
 sg13g2_decap_8 FILLER_6_3503 ();
 sg13g2_decap_8 FILLER_6_3510 ();
 sg13g2_decap_8 FILLER_6_3517 ();
 sg13g2_decap_8 FILLER_6_3524 ();
 sg13g2_decap_8 FILLER_6_3531 ();
 sg13g2_decap_8 FILLER_6_3538 ();
 sg13g2_decap_8 FILLER_6_3545 ();
 sg13g2_decap_8 FILLER_6_3552 ();
 sg13g2_decap_8 FILLER_6_3559 ();
 sg13g2_decap_8 FILLER_6_3566 ();
 sg13g2_decap_8 FILLER_6_3573 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_4 FILLER_7_546 ();
 sg13g2_fill_2 FILLER_7_550 ();
 sg13g2_decap_4 FILLER_7_622 ();
 sg13g2_decap_8 FILLER_7_631 ();
 sg13g2_decap_8 FILLER_7_638 ();
 sg13g2_fill_1 FILLER_7_645 ();
 sg13g2_decap_8 FILLER_7_669 ();
 sg13g2_decap_8 FILLER_7_676 ();
 sg13g2_decap_8 FILLER_7_683 ();
 sg13g2_fill_1 FILLER_7_690 ();
 sg13g2_decap_4 FILLER_7_761 ();
 sg13g2_decap_8 FILLER_7_796 ();
 sg13g2_decap_8 FILLER_7_803 ();
 sg13g2_decap_4 FILLER_7_810 ();
 sg13g2_fill_1 FILLER_7_814 ();
 sg13g2_decap_8 FILLER_7_866 ();
 sg13g2_fill_2 FILLER_7_873 ();
 sg13g2_decap_8 FILLER_7_901 ();
 sg13g2_fill_1 FILLER_7_908 ();
 sg13g2_decap_8 FILLER_7_914 ();
 sg13g2_decap_8 FILLER_7_921 ();
 sg13g2_decap_4 FILLER_7_928 ();
 sg13g2_fill_1 FILLER_7_932 ();
 sg13g2_fill_1 FILLER_7_937 ();
 sg13g2_fill_2 FILLER_7_943 ();
 sg13g2_fill_1 FILLER_7_945 ();
 sg13g2_fill_2 FILLER_7_952 ();
 sg13g2_fill_1 FILLER_7_954 ();
 sg13g2_fill_1 FILLER_7_959 ();
 sg13g2_fill_2 FILLER_7_968 ();
 sg13g2_fill_1 FILLER_7_970 ();
 sg13g2_fill_2 FILLER_7_981 ();
 sg13g2_fill_1 FILLER_7_983 ();
 sg13g2_decap_4 FILLER_7_992 ();
 sg13g2_decap_8 FILLER_7_1051 ();
 sg13g2_fill_2 FILLER_7_1058 ();
 sg13g2_decap_8 FILLER_7_1099 ();
 sg13g2_decap_8 FILLER_7_1106 ();
 sg13g2_fill_2 FILLER_7_1113 ();
 sg13g2_fill_1 FILLER_7_1150 ();
 sg13g2_fill_1 FILLER_7_1154 ();
 sg13g2_decap_8 FILLER_7_1158 ();
 sg13g2_decap_8 FILLER_7_1165 ();
 sg13g2_decap_8 FILLER_7_1172 ();
 sg13g2_fill_2 FILLER_7_1179 ();
 sg13g2_fill_1 FILLER_7_1181 ();
 sg13g2_decap_8 FILLER_7_1216 ();
 sg13g2_decap_8 FILLER_7_1223 ();
 sg13g2_fill_1 FILLER_7_1230 ();
 sg13g2_fill_2 FILLER_7_1236 ();
 sg13g2_decap_8 FILLER_7_1264 ();
 sg13g2_decap_8 FILLER_7_1315 ();
 sg13g2_decap_4 FILLER_7_1322 ();
 sg13g2_fill_1 FILLER_7_1326 ();
 sg13g2_decap_8 FILLER_7_1360 ();
 sg13g2_decap_8 FILLER_7_1367 ();
 sg13g2_fill_2 FILLER_7_1374 ();
 sg13g2_fill_1 FILLER_7_1384 ();
 sg13g2_decap_8 FILLER_7_1399 ();
 sg13g2_decap_8 FILLER_7_1406 ();
 sg13g2_decap_8 FILLER_7_1413 ();
 sg13g2_fill_1 FILLER_7_1420 ();
 sg13g2_decap_8 FILLER_7_1452 ();
 sg13g2_fill_1 FILLER_7_1459 ();
 sg13g2_fill_2 FILLER_7_1486 ();
 sg13g2_decap_4 FILLER_7_1514 ();
 sg13g2_fill_2 FILLER_7_1518 ();
 sg13g2_decap_8 FILLER_7_1562 ();
 sg13g2_decap_8 FILLER_7_1569 ();
 sg13g2_fill_1 FILLER_7_1576 ();
 sg13g2_decap_8 FILLER_7_1629 ();
 sg13g2_decap_8 FILLER_7_1636 ();
 sg13g2_fill_2 FILLER_7_1643 ();
 sg13g2_fill_1 FILLER_7_1645 ();
 sg13g2_decap_8 FILLER_7_1677 ();
 sg13g2_decap_8 FILLER_7_1684 ();
 sg13g2_decap_8 FILLER_7_1691 ();
 sg13g2_decap_4 FILLER_7_1698 ();
 sg13g2_fill_2 FILLER_7_1702 ();
 sg13g2_decap_4 FILLER_7_1730 ();
 sg13g2_fill_2 FILLER_7_1738 ();
 sg13g2_fill_1 FILLER_7_1740 ();
 sg13g2_decap_8 FILLER_7_1746 ();
 sg13g2_decap_8 FILLER_7_1782 ();
 sg13g2_fill_1 FILLER_7_1789 ();
 sg13g2_fill_1 FILLER_7_1832 ();
 sg13g2_fill_2 FILLER_7_1859 ();
 sg13g2_fill_1 FILLER_7_1861 ();
 sg13g2_fill_1 FILLER_7_1893 ();
 sg13g2_fill_2 FILLER_7_1928 ();
 sg13g2_fill_1 FILLER_7_1930 ();
 sg13g2_decap_8 FILLER_7_1957 ();
 sg13g2_decap_8 FILLER_7_1964 ();
 sg13g2_decap_8 FILLER_7_1971 ();
 sg13g2_decap_8 FILLER_7_1978 ();
 sg13g2_decap_8 FILLER_7_1985 ();
 sg13g2_decap_4 FILLER_7_1992 ();
 sg13g2_fill_1 FILLER_7_1996 ();
 sg13g2_decap_8 FILLER_7_2007 ();
 sg13g2_decap_8 FILLER_7_2014 ();
 sg13g2_decap_8 FILLER_7_2067 ();
 sg13g2_fill_2 FILLER_7_2074 ();
 sg13g2_decap_8 FILLER_7_2128 ();
 sg13g2_decap_8 FILLER_7_2135 ();
 sg13g2_fill_1 FILLER_7_2142 ();
 sg13g2_decap_4 FILLER_7_2247 ();
 sg13g2_fill_1 FILLER_7_2251 ();
 sg13g2_decap_8 FILLER_7_2260 ();
 sg13g2_decap_8 FILLER_7_2267 ();
 sg13g2_decap_4 FILLER_7_2274 ();
 sg13g2_fill_1 FILLER_7_2278 ();
 sg13g2_fill_2 FILLER_7_2295 ();
 sg13g2_decap_8 FILLER_7_2375 ();
 sg13g2_decap_8 FILLER_7_2387 ();
 sg13g2_decap_4 FILLER_7_2394 ();
 sg13g2_fill_1 FILLER_7_2398 ();
 sg13g2_decap_8 FILLER_7_2448 ();
 sg13g2_decap_8 FILLER_7_2455 ();
 sg13g2_decap_8 FILLER_7_2462 ();
 sg13g2_decap_4 FILLER_7_2469 ();
 sg13g2_decap_8 FILLER_7_2499 ();
 sg13g2_decap_8 FILLER_7_2552 ();
 sg13g2_decap_8 FILLER_7_2559 ();
 sg13g2_decap_8 FILLER_7_2566 ();
 sg13g2_decap_8 FILLER_7_2573 ();
 sg13g2_decap_8 FILLER_7_2580 ();
 sg13g2_decap_8 FILLER_7_2587 ();
 sg13g2_decap_8 FILLER_7_2594 ();
 sg13g2_decap_8 FILLER_7_2601 ();
 sg13g2_decap_8 FILLER_7_2608 ();
 sg13g2_decap_8 FILLER_7_2615 ();
 sg13g2_decap_8 FILLER_7_2622 ();
 sg13g2_decap_8 FILLER_7_2629 ();
 sg13g2_decap_8 FILLER_7_2636 ();
 sg13g2_decap_8 FILLER_7_2643 ();
 sg13g2_decap_8 FILLER_7_2650 ();
 sg13g2_decap_8 FILLER_7_2657 ();
 sg13g2_decap_8 FILLER_7_2664 ();
 sg13g2_decap_8 FILLER_7_2671 ();
 sg13g2_decap_8 FILLER_7_2678 ();
 sg13g2_decap_8 FILLER_7_2685 ();
 sg13g2_decap_8 FILLER_7_2692 ();
 sg13g2_decap_8 FILLER_7_2699 ();
 sg13g2_decap_8 FILLER_7_2706 ();
 sg13g2_decap_8 FILLER_7_2713 ();
 sg13g2_decap_8 FILLER_7_2720 ();
 sg13g2_decap_8 FILLER_7_2727 ();
 sg13g2_decap_8 FILLER_7_2734 ();
 sg13g2_decap_8 FILLER_7_2741 ();
 sg13g2_decap_8 FILLER_7_2748 ();
 sg13g2_decap_8 FILLER_7_2755 ();
 sg13g2_decap_8 FILLER_7_2762 ();
 sg13g2_decap_8 FILLER_7_2769 ();
 sg13g2_decap_8 FILLER_7_2776 ();
 sg13g2_decap_8 FILLER_7_2783 ();
 sg13g2_decap_8 FILLER_7_2790 ();
 sg13g2_decap_8 FILLER_7_2797 ();
 sg13g2_decap_8 FILLER_7_2804 ();
 sg13g2_decap_8 FILLER_7_2811 ();
 sg13g2_decap_8 FILLER_7_2818 ();
 sg13g2_decap_8 FILLER_7_2825 ();
 sg13g2_decap_8 FILLER_7_2832 ();
 sg13g2_decap_8 FILLER_7_2839 ();
 sg13g2_decap_8 FILLER_7_2846 ();
 sg13g2_decap_8 FILLER_7_2853 ();
 sg13g2_decap_8 FILLER_7_2860 ();
 sg13g2_decap_8 FILLER_7_2867 ();
 sg13g2_decap_8 FILLER_7_2874 ();
 sg13g2_decap_8 FILLER_7_2881 ();
 sg13g2_decap_8 FILLER_7_2888 ();
 sg13g2_decap_8 FILLER_7_2895 ();
 sg13g2_decap_8 FILLER_7_2902 ();
 sg13g2_decap_8 FILLER_7_2909 ();
 sg13g2_decap_8 FILLER_7_2916 ();
 sg13g2_decap_8 FILLER_7_2923 ();
 sg13g2_decap_8 FILLER_7_2930 ();
 sg13g2_decap_8 FILLER_7_2937 ();
 sg13g2_decap_8 FILLER_7_2944 ();
 sg13g2_decap_8 FILLER_7_2951 ();
 sg13g2_decap_8 FILLER_7_2958 ();
 sg13g2_decap_8 FILLER_7_2965 ();
 sg13g2_decap_8 FILLER_7_2972 ();
 sg13g2_decap_8 FILLER_7_2979 ();
 sg13g2_decap_8 FILLER_7_2986 ();
 sg13g2_decap_8 FILLER_7_2993 ();
 sg13g2_decap_8 FILLER_7_3000 ();
 sg13g2_decap_8 FILLER_7_3007 ();
 sg13g2_decap_8 FILLER_7_3014 ();
 sg13g2_decap_8 FILLER_7_3021 ();
 sg13g2_decap_8 FILLER_7_3028 ();
 sg13g2_decap_8 FILLER_7_3035 ();
 sg13g2_decap_8 FILLER_7_3042 ();
 sg13g2_decap_8 FILLER_7_3049 ();
 sg13g2_decap_8 FILLER_7_3056 ();
 sg13g2_decap_8 FILLER_7_3063 ();
 sg13g2_decap_8 FILLER_7_3070 ();
 sg13g2_decap_8 FILLER_7_3077 ();
 sg13g2_decap_8 FILLER_7_3084 ();
 sg13g2_decap_8 FILLER_7_3091 ();
 sg13g2_decap_8 FILLER_7_3098 ();
 sg13g2_decap_8 FILLER_7_3105 ();
 sg13g2_decap_8 FILLER_7_3112 ();
 sg13g2_decap_8 FILLER_7_3119 ();
 sg13g2_decap_8 FILLER_7_3126 ();
 sg13g2_decap_8 FILLER_7_3133 ();
 sg13g2_decap_8 FILLER_7_3140 ();
 sg13g2_decap_8 FILLER_7_3147 ();
 sg13g2_decap_8 FILLER_7_3154 ();
 sg13g2_decap_8 FILLER_7_3161 ();
 sg13g2_decap_8 FILLER_7_3168 ();
 sg13g2_decap_8 FILLER_7_3175 ();
 sg13g2_decap_8 FILLER_7_3182 ();
 sg13g2_decap_8 FILLER_7_3189 ();
 sg13g2_decap_8 FILLER_7_3196 ();
 sg13g2_decap_8 FILLER_7_3203 ();
 sg13g2_decap_8 FILLER_7_3210 ();
 sg13g2_decap_8 FILLER_7_3217 ();
 sg13g2_decap_8 FILLER_7_3224 ();
 sg13g2_decap_8 FILLER_7_3231 ();
 sg13g2_decap_8 FILLER_7_3238 ();
 sg13g2_decap_8 FILLER_7_3245 ();
 sg13g2_decap_8 FILLER_7_3252 ();
 sg13g2_decap_8 FILLER_7_3259 ();
 sg13g2_decap_8 FILLER_7_3266 ();
 sg13g2_decap_8 FILLER_7_3273 ();
 sg13g2_decap_8 FILLER_7_3280 ();
 sg13g2_decap_8 FILLER_7_3287 ();
 sg13g2_decap_8 FILLER_7_3294 ();
 sg13g2_decap_8 FILLER_7_3301 ();
 sg13g2_decap_8 FILLER_7_3308 ();
 sg13g2_decap_8 FILLER_7_3315 ();
 sg13g2_decap_8 FILLER_7_3322 ();
 sg13g2_decap_8 FILLER_7_3329 ();
 sg13g2_decap_8 FILLER_7_3336 ();
 sg13g2_decap_8 FILLER_7_3343 ();
 sg13g2_decap_8 FILLER_7_3350 ();
 sg13g2_decap_8 FILLER_7_3357 ();
 sg13g2_decap_8 FILLER_7_3364 ();
 sg13g2_decap_8 FILLER_7_3371 ();
 sg13g2_decap_8 FILLER_7_3378 ();
 sg13g2_decap_8 FILLER_7_3385 ();
 sg13g2_decap_8 FILLER_7_3392 ();
 sg13g2_decap_8 FILLER_7_3399 ();
 sg13g2_decap_8 FILLER_7_3406 ();
 sg13g2_decap_8 FILLER_7_3413 ();
 sg13g2_decap_8 FILLER_7_3420 ();
 sg13g2_decap_8 FILLER_7_3427 ();
 sg13g2_decap_8 FILLER_7_3434 ();
 sg13g2_decap_8 FILLER_7_3441 ();
 sg13g2_decap_8 FILLER_7_3448 ();
 sg13g2_decap_8 FILLER_7_3455 ();
 sg13g2_decap_8 FILLER_7_3462 ();
 sg13g2_decap_8 FILLER_7_3469 ();
 sg13g2_decap_8 FILLER_7_3476 ();
 sg13g2_decap_8 FILLER_7_3483 ();
 sg13g2_decap_8 FILLER_7_3490 ();
 sg13g2_decap_8 FILLER_7_3497 ();
 sg13g2_decap_8 FILLER_7_3504 ();
 sg13g2_decap_8 FILLER_7_3511 ();
 sg13g2_decap_8 FILLER_7_3518 ();
 sg13g2_decap_8 FILLER_7_3525 ();
 sg13g2_decap_8 FILLER_7_3532 ();
 sg13g2_decap_8 FILLER_7_3539 ();
 sg13g2_decap_8 FILLER_7_3546 ();
 sg13g2_decap_8 FILLER_7_3553 ();
 sg13g2_decap_8 FILLER_7_3560 ();
 sg13g2_decap_8 FILLER_7_3567 ();
 sg13g2_decap_4 FILLER_7_3574 ();
 sg13g2_fill_2 FILLER_7_3578 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_fill_2 FILLER_8_539 ();
 sg13g2_fill_1 FILLER_8_541 ();
 sg13g2_fill_1 FILLER_8_589 ();
 sg13g2_decap_8 FILLER_8_606 ();
 sg13g2_decap_4 FILLER_8_613 ();
 sg13g2_fill_2 FILLER_8_617 ();
 sg13g2_decap_4 FILLER_8_678 ();
 sg13g2_fill_2 FILLER_8_708 ();
 sg13g2_fill_1 FILLER_8_736 ();
 sg13g2_decap_4 FILLER_8_757 ();
 sg13g2_fill_2 FILLER_8_761 ();
 sg13g2_decap_8 FILLER_8_804 ();
 sg13g2_decap_8 FILLER_8_811 ();
 sg13g2_fill_2 FILLER_8_818 ();
 sg13g2_fill_1 FILLER_8_820 ();
 sg13g2_decap_8 FILLER_8_865 ();
 sg13g2_decap_8 FILLER_8_872 ();
 sg13g2_decap_8 FILLER_8_879 ();
 sg13g2_fill_2 FILLER_8_886 ();
 sg13g2_fill_1 FILLER_8_888 ();
 sg13g2_decap_8 FILLER_8_974 ();
 sg13g2_decap_8 FILLER_8_981 ();
 sg13g2_decap_8 FILLER_8_988 ();
 sg13g2_decap_8 FILLER_8_995 ();
 sg13g2_fill_1 FILLER_8_1002 ();
 sg13g2_fill_2 FILLER_8_1020 ();
 sg13g2_fill_2 FILLER_8_1048 ();
 sg13g2_fill_1 FILLER_8_1050 ();
 sg13g2_decap_8 FILLER_8_1054 ();
 sg13g2_decap_8 FILLER_8_1061 ();
 sg13g2_fill_2 FILLER_8_1068 ();
 sg13g2_fill_1 FILLER_8_1074 ();
 sg13g2_decap_8 FILLER_8_1101 ();
 sg13g2_decap_4 FILLER_8_1108 ();
 sg13g2_fill_1 FILLER_8_1112 ();
 sg13g2_fill_1 FILLER_8_1234 ();
 sg13g2_decap_8 FILLER_8_1243 ();
 sg13g2_decap_8 FILLER_8_1250 ();
 sg13g2_decap_8 FILLER_8_1257 ();
 sg13g2_decap_8 FILLER_8_1264 ();
 sg13g2_decap_4 FILLER_8_1271 ();
 sg13g2_fill_1 FILLER_8_1275 ();
 sg13g2_decap_4 FILLER_8_1322 ();
 sg13g2_fill_1 FILLER_8_1326 ();
 sg13g2_fill_2 FILLER_8_1366 ();
 sg13g2_fill_1 FILLER_8_1368 ();
 sg13g2_decap_8 FILLER_8_1400 ();
 sg13g2_decap_8 FILLER_8_1407 ();
 sg13g2_decap_8 FILLER_8_1456 ();
 sg13g2_decap_8 FILLER_8_1463 ();
 sg13g2_decap_4 FILLER_8_1470 ();
 sg13g2_decap_8 FILLER_8_1513 ();
 sg13g2_decap_8 FILLER_8_1520 ();
 sg13g2_decap_4 FILLER_8_1527 ();
 sg13g2_decap_8 FILLER_8_1557 ();
 sg13g2_decap_8 FILLER_8_1564 ();
 sg13g2_decap_8 FILLER_8_1571 ();
 sg13g2_decap_8 FILLER_8_1578 ();
 sg13g2_decap_8 FILLER_8_1585 ();
 sg13g2_decap_8 FILLER_8_1618 ();
 sg13g2_decap_8 FILLER_8_1625 ();
 sg13g2_decap_4 FILLER_8_1632 ();
 sg13g2_fill_2 FILLER_8_1678 ();
 sg13g2_fill_1 FILLER_8_1680 ();
 sg13g2_fill_2 FILLER_8_1741 ();
 sg13g2_decap_8 FILLER_8_1763 ();
 sg13g2_fill_1 FILLER_8_1770 ();
 sg13g2_decap_8 FILLER_8_1831 ();
 sg13g2_decap_8 FILLER_8_1838 ();
 sg13g2_decap_8 FILLER_8_1845 ();
 sg13g2_fill_2 FILLER_8_1852 ();
 sg13g2_fill_1 FILLER_8_1854 ();
 sg13g2_fill_2 FILLER_8_1876 ();
 sg13g2_fill_1 FILLER_8_1878 ();
 sg13g2_fill_1 FILLER_8_1913 ();
 sg13g2_fill_2 FILLER_8_1926 ();
 sg13g2_fill_1 FILLER_8_1928 ();
 sg13g2_decap_8 FILLER_8_1955 ();
 sg13g2_decap_8 FILLER_8_1962 ();
 sg13g2_decap_8 FILLER_8_1969 ();
 sg13g2_decap_8 FILLER_8_2014 ();
 sg13g2_decap_8 FILLER_8_2021 ();
 sg13g2_fill_2 FILLER_8_2028 ();
 sg13g2_fill_1 FILLER_8_2030 ();
 sg13g2_fill_2 FILLER_8_2120 ();
 sg13g2_decap_8 FILLER_8_2176 ();
 sg13g2_decap_8 FILLER_8_2183 ();
 sg13g2_decap_8 FILLER_8_2219 ();
 sg13g2_fill_2 FILLER_8_2226 ();
 sg13g2_fill_1 FILLER_8_2228 ();
 sg13g2_fill_1 FILLER_8_2256 ();
 sg13g2_fill_1 FILLER_8_2293 ();
 sg13g2_fill_2 FILLER_8_2306 ();
 sg13g2_fill_1 FILLER_8_2313 ();
 sg13g2_fill_2 FILLER_8_2329 ();
 sg13g2_fill_1 FILLER_8_2331 ();
 sg13g2_decap_4 FILLER_8_2371 ();
 sg13g2_fill_1 FILLER_8_2375 ();
 sg13g2_fill_2 FILLER_8_2384 ();
 sg13g2_fill_1 FILLER_8_2386 ();
 sg13g2_decap_4 FILLER_8_2402 ();
 sg13g2_fill_2 FILLER_8_2440 ();
 sg13g2_fill_1 FILLER_8_2442 ();
 sg13g2_fill_2 FILLER_8_2469 ();
 sg13g2_decap_8 FILLER_8_2499 ();
 sg13g2_decap_8 FILLER_8_2555 ();
 sg13g2_decap_8 FILLER_8_2562 ();
 sg13g2_decap_8 FILLER_8_2569 ();
 sg13g2_decap_8 FILLER_8_2576 ();
 sg13g2_decap_8 FILLER_8_2583 ();
 sg13g2_decap_8 FILLER_8_2590 ();
 sg13g2_decap_8 FILLER_8_2597 ();
 sg13g2_decap_8 FILLER_8_2604 ();
 sg13g2_decap_8 FILLER_8_2611 ();
 sg13g2_decap_8 FILLER_8_2618 ();
 sg13g2_decap_8 FILLER_8_2625 ();
 sg13g2_decap_8 FILLER_8_2632 ();
 sg13g2_decap_8 FILLER_8_2639 ();
 sg13g2_decap_8 FILLER_8_2646 ();
 sg13g2_decap_8 FILLER_8_2653 ();
 sg13g2_decap_8 FILLER_8_2660 ();
 sg13g2_decap_8 FILLER_8_2667 ();
 sg13g2_decap_8 FILLER_8_2674 ();
 sg13g2_decap_8 FILLER_8_2681 ();
 sg13g2_decap_8 FILLER_8_2688 ();
 sg13g2_decap_8 FILLER_8_2695 ();
 sg13g2_decap_8 FILLER_8_2702 ();
 sg13g2_decap_8 FILLER_8_2709 ();
 sg13g2_decap_8 FILLER_8_2716 ();
 sg13g2_decap_8 FILLER_8_2723 ();
 sg13g2_decap_8 FILLER_8_2730 ();
 sg13g2_decap_8 FILLER_8_2737 ();
 sg13g2_decap_8 FILLER_8_2744 ();
 sg13g2_decap_8 FILLER_8_2751 ();
 sg13g2_decap_8 FILLER_8_2758 ();
 sg13g2_decap_8 FILLER_8_2765 ();
 sg13g2_decap_8 FILLER_8_2772 ();
 sg13g2_decap_8 FILLER_8_2779 ();
 sg13g2_decap_8 FILLER_8_2786 ();
 sg13g2_decap_8 FILLER_8_2793 ();
 sg13g2_decap_8 FILLER_8_2800 ();
 sg13g2_decap_8 FILLER_8_2807 ();
 sg13g2_decap_8 FILLER_8_2814 ();
 sg13g2_decap_8 FILLER_8_2821 ();
 sg13g2_decap_8 FILLER_8_2828 ();
 sg13g2_decap_8 FILLER_8_2835 ();
 sg13g2_decap_8 FILLER_8_2842 ();
 sg13g2_decap_8 FILLER_8_2849 ();
 sg13g2_decap_8 FILLER_8_2856 ();
 sg13g2_decap_8 FILLER_8_2863 ();
 sg13g2_decap_8 FILLER_8_2870 ();
 sg13g2_decap_8 FILLER_8_2877 ();
 sg13g2_decap_8 FILLER_8_2884 ();
 sg13g2_decap_8 FILLER_8_2891 ();
 sg13g2_decap_8 FILLER_8_2898 ();
 sg13g2_decap_8 FILLER_8_2905 ();
 sg13g2_decap_8 FILLER_8_2912 ();
 sg13g2_decap_8 FILLER_8_2919 ();
 sg13g2_decap_8 FILLER_8_2926 ();
 sg13g2_decap_8 FILLER_8_2933 ();
 sg13g2_decap_8 FILLER_8_2940 ();
 sg13g2_decap_8 FILLER_8_2947 ();
 sg13g2_decap_8 FILLER_8_2954 ();
 sg13g2_decap_8 FILLER_8_2961 ();
 sg13g2_decap_8 FILLER_8_2968 ();
 sg13g2_decap_8 FILLER_8_2975 ();
 sg13g2_decap_8 FILLER_8_2982 ();
 sg13g2_decap_8 FILLER_8_2989 ();
 sg13g2_decap_8 FILLER_8_2996 ();
 sg13g2_decap_8 FILLER_8_3003 ();
 sg13g2_decap_8 FILLER_8_3010 ();
 sg13g2_decap_8 FILLER_8_3017 ();
 sg13g2_decap_8 FILLER_8_3024 ();
 sg13g2_decap_8 FILLER_8_3031 ();
 sg13g2_decap_8 FILLER_8_3038 ();
 sg13g2_decap_8 FILLER_8_3045 ();
 sg13g2_decap_8 FILLER_8_3052 ();
 sg13g2_decap_8 FILLER_8_3059 ();
 sg13g2_decap_8 FILLER_8_3066 ();
 sg13g2_decap_8 FILLER_8_3073 ();
 sg13g2_decap_8 FILLER_8_3080 ();
 sg13g2_decap_8 FILLER_8_3087 ();
 sg13g2_decap_8 FILLER_8_3094 ();
 sg13g2_decap_8 FILLER_8_3101 ();
 sg13g2_decap_8 FILLER_8_3108 ();
 sg13g2_decap_8 FILLER_8_3115 ();
 sg13g2_decap_8 FILLER_8_3122 ();
 sg13g2_decap_8 FILLER_8_3129 ();
 sg13g2_decap_8 FILLER_8_3136 ();
 sg13g2_decap_8 FILLER_8_3143 ();
 sg13g2_decap_8 FILLER_8_3150 ();
 sg13g2_decap_8 FILLER_8_3157 ();
 sg13g2_decap_8 FILLER_8_3164 ();
 sg13g2_decap_8 FILLER_8_3171 ();
 sg13g2_decap_8 FILLER_8_3178 ();
 sg13g2_decap_8 FILLER_8_3185 ();
 sg13g2_decap_8 FILLER_8_3192 ();
 sg13g2_decap_8 FILLER_8_3199 ();
 sg13g2_decap_8 FILLER_8_3206 ();
 sg13g2_decap_8 FILLER_8_3213 ();
 sg13g2_decap_8 FILLER_8_3220 ();
 sg13g2_decap_8 FILLER_8_3227 ();
 sg13g2_decap_8 FILLER_8_3234 ();
 sg13g2_decap_8 FILLER_8_3241 ();
 sg13g2_decap_8 FILLER_8_3248 ();
 sg13g2_decap_8 FILLER_8_3255 ();
 sg13g2_decap_8 FILLER_8_3262 ();
 sg13g2_decap_8 FILLER_8_3269 ();
 sg13g2_decap_8 FILLER_8_3276 ();
 sg13g2_decap_8 FILLER_8_3283 ();
 sg13g2_decap_8 FILLER_8_3290 ();
 sg13g2_decap_8 FILLER_8_3297 ();
 sg13g2_decap_8 FILLER_8_3304 ();
 sg13g2_decap_8 FILLER_8_3311 ();
 sg13g2_decap_8 FILLER_8_3318 ();
 sg13g2_decap_8 FILLER_8_3325 ();
 sg13g2_decap_8 FILLER_8_3332 ();
 sg13g2_decap_8 FILLER_8_3339 ();
 sg13g2_decap_8 FILLER_8_3346 ();
 sg13g2_decap_8 FILLER_8_3353 ();
 sg13g2_decap_8 FILLER_8_3360 ();
 sg13g2_decap_8 FILLER_8_3367 ();
 sg13g2_decap_8 FILLER_8_3374 ();
 sg13g2_decap_8 FILLER_8_3381 ();
 sg13g2_decap_8 FILLER_8_3388 ();
 sg13g2_decap_8 FILLER_8_3395 ();
 sg13g2_decap_8 FILLER_8_3402 ();
 sg13g2_decap_8 FILLER_8_3409 ();
 sg13g2_decap_8 FILLER_8_3416 ();
 sg13g2_decap_8 FILLER_8_3423 ();
 sg13g2_decap_8 FILLER_8_3430 ();
 sg13g2_decap_8 FILLER_8_3437 ();
 sg13g2_decap_8 FILLER_8_3444 ();
 sg13g2_decap_8 FILLER_8_3451 ();
 sg13g2_decap_8 FILLER_8_3458 ();
 sg13g2_decap_8 FILLER_8_3465 ();
 sg13g2_decap_8 FILLER_8_3472 ();
 sg13g2_decap_8 FILLER_8_3479 ();
 sg13g2_decap_8 FILLER_8_3486 ();
 sg13g2_decap_8 FILLER_8_3493 ();
 sg13g2_decap_8 FILLER_8_3500 ();
 sg13g2_decap_8 FILLER_8_3507 ();
 sg13g2_decap_8 FILLER_8_3514 ();
 sg13g2_decap_8 FILLER_8_3521 ();
 sg13g2_decap_8 FILLER_8_3528 ();
 sg13g2_decap_8 FILLER_8_3535 ();
 sg13g2_decap_8 FILLER_8_3542 ();
 sg13g2_decap_8 FILLER_8_3549 ();
 sg13g2_decap_8 FILLER_8_3556 ();
 sg13g2_decap_8 FILLER_8_3563 ();
 sg13g2_decap_8 FILLER_8_3570 ();
 sg13g2_fill_2 FILLER_8_3577 ();
 sg13g2_fill_1 FILLER_8_3579 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_587 ();
 sg13g2_decap_8 FILLER_9_594 ();
 sg13g2_decap_8 FILLER_9_601 ();
 sg13g2_decap_4 FILLER_9_608 ();
 sg13g2_fill_2 FILLER_9_646 ();
 sg13g2_fill_1 FILLER_9_648 ();
 sg13g2_fill_1 FILLER_9_662 ();
 sg13g2_fill_1 FILLER_9_689 ();
 sg13g2_fill_1 FILLER_9_703 ();
 sg13g2_fill_2 FILLER_9_709 ();
 sg13g2_decap_8 FILLER_9_719 ();
 sg13g2_fill_2 FILLER_9_726 ();
 sg13g2_decap_8 FILLER_9_754 ();
 sg13g2_decap_4 FILLER_9_761 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_4 FILLER_9_855 ();
 sg13g2_fill_1 FILLER_9_859 ();
 sg13g2_fill_1 FILLER_9_890 ();
 sg13g2_fill_1 FILLER_9_956 ();
 sg13g2_fill_2 FILLER_9_975 ();
 sg13g2_decap_8 FILLER_9_984 ();
 sg13g2_decap_8 FILLER_9_991 ();
 sg13g2_fill_1 FILLER_9_998 ();
 sg13g2_fill_2 FILLER_9_1025 ();
 sg13g2_fill_2 FILLER_9_1057 ();
 sg13g2_fill_1 FILLER_9_1064 ();
 sg13g2_fill_2 FILLER_9_1070 ();
 sg13g2_fill_1 FILLER_9_1072 ();
 sg13g2_decap_4 FILLER_9_1113 ();
 sg13g2_fill_1 FILLER_9_1117 ();
 sg13g2_decap_8 FILLER_9_1177 ();
 sg13g2_decap_4 FILLER_9_1184 ();
 sg13g2_fill_1 FILLER_9_1188 ();
 sg13g2_fill_2 FILLER_9_1223 ();
 sg13g2_fill_1 FILLER_9_1225 ();
 sg13g2_decap_8 FILLER_9_1256 ();
 sg13g2_fill_2 FILLER_9_1263 ();
 sg13g2_fill_1 FILLER_9_1265 ();
 sg13g2_fill_1 FILLER_9_1326 ();
 sg13g2_decap_4 FILLER_9_1363 ();
 sg13g2_fill_1 FILLER_9_1367 ();
 sg13g2_decap_4 FILLER_9_1402 ();
 sg13g2_fill_2 FILLER_9_1406 ();
 sg13g2_fill_1 FILLER_9_1425 ();
 sg13g2_decap_4 FILLER_9_1468 ();
 sg13g2_decap_4 FILLER_9_1507 ();
 sg13g2_decap_8 FILLER_9_1563 ();
 sg13g2_decap_8 FILLER_9_1570 ();
 sg13g2_decap_8 FILLER_9_1577 ();
 sg13g2_decap_8 FILLER_9_1584 ();
 sg13g2_fill_2 FILLER_9_1591 ();
 sg13g2_fill_1 FILLER_9_1593 ();
 sg13g2_decap_8 FILLER_9_1626 ();
 sg13g2_decap_8 FILLER_9_1633 ();
 sg13g2_decap_4 FILLER_9_1640 ();
 sg13g2_decap_8 FILLER_9_1706 ();
 sg13g2_decap_8 FILLER_9_1713 ();
 sg13g2_decap_4 FILLER_9_1720 ();
 sg13g2_fill_2 FILLER_9_1724 ();
 sg13g2_fill_1 FILLER_9_1752 ();
 sg13g2_decap_4 FILLER_9_1756 ();
 sg13g2_fill_1 FILLER_9_1760 ();
 sg13g2_decap_8 FILLER_9_1830 ();
 sg13g2_decap_8 FILLER_9_1837 ();
 sg13g2_decap_8 FILLER_9_1844 ();
 sg13g2_decap_4 FILLER_9_1851 ();
 sg13g2_decap_4 FILLER_9_1881 ();
 sg13g2_decap_8 FILLER_9_1916 ();
 sg13g2_fill_2 FILLER_9_1923 ();
 sg13g2_decap_8 FILLER_9_1930 ();
 sg13g2_decap_8 FILLER_9_1937 ();
 sg13g2_decap_8 FILLER_9_1944 ();
 sg13g2_decap_8 FILLER_9_1951 ();
 sg13g2_decap_8 FILLER_9_1958 ();
 sg13g2_decap_8 FILLER_9_1965 ();
 sg13g2_decap_8 FILLER_9_1972 ();
 sg13g2_decap_4 FILLER_9_1979 ();
 sg13g2_fill_1 FILLER_9_2018 ();
 sg13g2_decap_4 FILLER_9_2024 ();
 sg13g2_fill_1 FILLER_9_2028 ();
 sg13g2_decap_8 FILLER_9_2034 ();
 sg13g2_fill_2 FILLER_9_2041 ();
 sg13g2_fill_1 FILLER_9_2043 ();
 sg13g2_decap_8 FILLER_9_2049 ();
 sg13g2_decap_8 FILLER_9_2056 ();
 sg13g2_fill_2 FILLER_9_2063 ();
 sg13g2_decap_8 FILLER_9_2068 ();
 sg13g2_decap_8 FILLER_9_2075 ();
 sg13g2_fill_2 FILLER_9_2082 ();
 sg13g2_decap_4 FILLER_9_2087 ();
 sg13g2_fill_2 FILLER_9_2091 ();
 sg13g2_decap_4 FILLER_9_2098 ();
 sg13g2_fill_1 FILLER_9_2102 ();
 sg13g2_decap_8 FILLER_9_2113 ();
 sg13g2_decap_8 FILLER_9_2120 ();
 sg13g2_decap_8 FILLER_9_2127 ();
 sg13g2_fill_2 FILLER_9_2134 ();
 sg13g2_fill_1 FILLER_9_2136 ();
 sg13g2_decap_8 FILLER_9_2166 ();
 sg13g2_decap_8 FILLER_9_2173 ();
 sg13g2_decap_4 FILLER_9_2180 ();
 sg13g2_fill_2 FILLER_9_2184 ();
 sg13g2_fill_1 FILLER_9_2261 ();
 sg13g2_fill_2 FILLER_9_2288 ();
 sg13g2_fill_1 FILLER_9_2290 ();
 sg13g2_fill_1 FILLER_9_2300 ();
 sg13g2_decap_8 FILLER_9_2309 ();
 sg13g2_decap_8 FILLER_9_2316 ();
 sg13g2_decap_8 FILLER_9_2331 ();
 sg13g2_decap_4 FILLER_9_2369 ();
 sg13g2_fill_2 FILLER_9_2373 ();
 sg13g2_fill_1 FILLER_9_2401 ();
 sg13g2_fill_2 FILLER_9_2436 ();
 sg13g2_decap_8 FILLER_9_2446 ();
 sg13g2_fill_2 FILLER_9_2453 ();
 sg13g2_fill_2 FILLER_9_2507 ();
 sg13g2_fill_1 FILLER_9_2509 ();
 sg13g2_fill_2 FILLER_9_2527 ();
 sg13g2_decap_8 FILLER_9_2581 ();
 sg13g2_decap_8 FILLER_9_2588 ();
 sg13g2_decap_4 FILLER_9_2599 ();
 sg13g2_fill_1 FILLER_9_2603 ();
 sg13g2_decap_8 FILLER_9_2607 ();
 sg13g2_fill_2 FILLER_9_2614 ();
 sg13g2_decap_8 FILLER_9_2620 ();
 sg13g2_decap_8 FILLER_9_2632 ();
 sg13g2_decap_8 FILLER_9_2639 ();
 sg13g2_decap_8 FILLER_9_2646 ();
 sg13g2_decap_8 FILLER_9_2653 ();
 sg13g2_decap_8 FILLER_9_2660 ();
 sg13g2_decap_8 FILLER_9_2667 ();
 sg13g2_decap_8 FILLER_9_2674 ();
 sg13g2_decap_8 FILLER_9_2681 ();
 sg13g2_decap_8 FILLER_9_2688 ();
 sg13g2_decap_8 FILLER_9_2695 ();
 sg13g2_decap_8 FILLER_9_2702 ();
 sg13g2_decap_8 FILLER_9_2709 ();
 sg13g2_decap_8 FILLER_9_2716 ();
 sg13g2_decap_8 FILLER_9_2723 ();
 sg13g2_decap_8 FILLER_9_2730 ();
 sg13g2_decap_8 FILLER_9_2737 ();
 sg13g2_decap_8 FILLER_9_2744 ();
 sg13g2_decap_8 FILLER_9_2751 ();
 sg13g2_decap_8 FILLER_9_2758 ();
 sg13g2_decap_8 FILLER_9_2765 ();
 sg13g2_decap_8 FILLER_9_2772 ();
 sg13g2_decap_8 FILLER_9_2779 ();
 sg13g2_decap_8 FILLER_9_2786 ();
 sg13g2_decap_8 FILLER_9_2793 ();
 sg13g2_decap_8 FILLER_9_2800 ();
 sg13g2_decap_8 FILLER_9_2807 ();
 sg13g2_decap_8 FILLER_9_2814 ();
 sg13g2_decap_8 FILLER_9_2821 ();
 sg13g2_decap_8 FILLER_9_2828 ();
 sg13g2_decap_8 FILLER_9_2835 ();
 sg13g2_decap_8 FILLER_9_2842 ();
 sg13g2_decap_8 FILLER_9_2849 ();
 sg13g2_decap_8 FILLER_9_2856 ();
 sg13g2_decap_8 FILLER_9_2863 ();
 sg13g2_decap_8 FILLER_9_2870 ();
 sg13g2_decap_8 FILLER_9_2877 ();
 sg13g2_decap_8 FILLER_9_2884 ();
 sg13g2_decap_8 FILLER_9_2891 ();
 sg13g2_decap_8 FILLER_9_2898 ();
 sg13g2_decap_8 FILLER_9_2905 ();
 sg13g2_decap_8 FILLER_9_2912 ();
 sg13g2_decap_8 FILLER_9_2919 ();
 sg13g2_decap_8 FILLER_9_2926 ();
 sg13g2_decap_8 FILLER_9_2933 ();
 sg13g2_decap_8 FILLER_9_2940 ();
 sg13g2_decap_8 FILLER_9_2947 ();
 sg13g2_decap_8 FILLER_9_2954 ();
 sg13g2_decap_8 FILLER_9_2961 ();
 sg13g2_decap_8 FILLER_9_2968 ();
 sg13g2_decap_8 FILLER_9_2975 ();
 sg13g2_decap_8 FILLER_9_2982 ();
 sg13g2_decap_8 FILLER_9_2989 ();
 sg13g2_decap_8 FILLER_9_2996 ();
 sg13g2_decap_8 FILLER_9_3003 ();
 sg13g2_decap_8 FILLER_9_3010 ();
 sg13g2_decap_8 FILLER_9_3017 ();
 sg13g2_decap_8 FILLER_9_3024 ();
 sg13g2_decap_8 FILLER_9_3031 ();
 sg13g2_decap_8 FILLER_9_3038 ();
 sg13g2_decap_8 FILLER_9_3045 ();
 sg13g2_decap_8 FILLER_9_3052 ();
 sg13g2_decap_8 FILLER_9_3059 ();
 sg13g2_decap_8 FILLER_9_3066 ();
 sg13g2_decap_8 FILLER_9_3073 ();
 sg13g2_decap_8 FILLER_9_3080 ();
 sg13g2_decap_8 FILLER_9_3087 ();
 sg13g2_decap_8 FILLER_9_3094 ();
 sg13g2_decap_8 FILLER_9_3101 ();
 sg13g2_decap_8 FILLER_9_3108 ();
 sg13g2_decap_8 FILLER_9_3115 ();
 sg13g2_decap_8 FILLER_9_3122 ();
 sg13g2_decap_8 FILLER_9_3129 ();
 sg13g2_decap_8 FILLER_9_3136 ();
 sg13g2_decap_8 FILLER_9_3143 ();
 sg13g2_decap_8 FILLER_9_3150 ();
 sg13g2_decap_8 FILLER_9_3157 ();
 sg13g2_decap_8 FILLER_9_3164 ();
 sg13g2_decap_8 FILLER_9_3171 ();
 sg13g2_decap_8 FILLER_9_3178 ();
 sg13g2_decap_8 FILLER_9_3185 ();
 sg13g2_decap_8 FILLER_9_3192 ();
 sg13g2_decap_8 FILLER_9_3199 ();
 sg13g2_decap_8 FILLER_9_3206 ();
 sg13g2_decap_8 FILLER_9_3213 ();
 sg13g2_decap_8 FILLER_9_3220 ();
 sg13g2_decap_8 FILLER_9_3227 ();
 sg13g2_decap_8 FILLER_9_3234 ();
 sg13g2_decap_8 FILLER_9_3241 ();
 sg13g2_decap_8 FILLER_9_3248 ();
 sg13g2_decap_8 FILLER_9_3255 ();
 sg13g2_decap_8 FILLER_9_3262 ();
 sg13g2_decap_8 FILLER_9_3269 ();
 sg13g2_decap_8 FILLER_9_3276 ();
 sg13g2_decap_8 FILLER_9_3283 ();
 sg13g2_decap_8 FILLER_9_3290 ();
 sg13g2_decap_8 FILLER_9_3297 ();
 sg13g2_decap_8 FILLER_9_3304 ();
 sg13g2_decap_8 FILLER_9_3311 ();
 sg13g2_decap_8 FILLER_9_3318 ();
 sg13g2_decap_8 FILLER_9_3325 ();
 sg13g2_decap_8 FILLER_9_3332 ();
 sg13g2_decap_8 FILLER_9_3339 ();
 sg13g2_decap_8 FILLER_9_3346 ();
 sg13g2_decap_8 FILLER_9_3353 ();
 sg13g2_decap_8 FILLER_9_3360 ();
 sg13g2_decap_8 FILLER_9_3367 ();
 sg13g2_decap_8 FILLER_9_3374 ();
 sg13g2_decap_8 FILLER_9_3381 ();
 sg13g2_decap_8 FILLER_9_3388 ();
 sg13g2_decap_8 FILLER_9_3395 ();
 sg13g2_decap_8 FILLER_9_3402 ();
 sg13g2_decap_8 FILLER_9_3409 ();
 sg13g2_decap_8 FILLER_9_3416 ();
 sg13g2_decap_8 FILLER_9_3423 ();
 sg13g2_decap_8 FILLER_9_3430 ();
 sg13g2_decap_8 FILLER_9_3437 ();
 sg13g2_decap_8 FILLER_9_3444 ();
 sg13g2_decap_8 FILLER_9_3451 ();
 sg13g2_decap_8 FILLER_9_3458 ();
 sg13g2_decap_8 FILLER_9_3465 ();
 sg13g2_decap_8 FILLER_9_3472 ();
 sg13g2_decap_8 FILLER_9_3479 ();
 sg13g2_decap_8 FILLER_9_3486 ();
 sg13g2_decap_8 FILLER_9_3493 ();
 sg13g2_decap_8 FILLER_9_3500 ();
 sg13g2_decap_8 FILLER_9_3507 ();
 sg13g2_decap_8 FILLER_9_3514 ();
 sg13g2_decap_8 FILLER_9_3521 ();
 sg13g2_decap_8 FILLER_9_3528 ();
 sg13g2_decap_8 FILLER_9_3535 ();
 sg13g2_decap_8 FILLER_9_3542 ();
 sg13g2_decap_8 FILLER_9_3549 ();
 sg13g2_decap_8 FILLER_9_3556 ();
 sg13g2_decap_8 FILLER_9_3563 ();
 sg13g2_decap_8 FILLER_9_3570 ();
 sg13g2_fill_2 FILLER_9_3577 ();
 sg13g2_fill_1 FILLER_9_3579 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_104 ();
 sg13g2_decap_8 FILLER_10_111 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_decap_8 FILLER_10_125 ();
 sg13g2_decap_8 FILLER_10_132 ();
 sg13g2_decap_8 FILLER_10_139 ();
 sg13g2_decap_8 FILLER_10_146 ();
 sg13g2_decap_8 FILLER_10_153 ();
 sg13g2_decap_8 FILLER_10_160 ();
 sg13g2_decap_8 FILLER_10_167 ();
 sg13g2_decap_8 FILLER_10_174 ();
 sg13g2_decap_8 FILLER_10_181 ();
 sg13g2_decap_8 FILLER_10_188 ();
 sg13g2_decap_8 FILLER_10_195 ();
 sg13g2_decap_8 FILLER_10_202 ();
 sg13g2_decap_8 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_216 ();
 sg13g2_decap_8 FILLER_10_223 ();
 sg13g2_decap_8 FILLER_10_230 ();
 sg13g2_decap_8 FILLER_10_237 ();
 sg13g2_decap_8 FILLER_10_244 ();
 sg13g2_decap_8 FILLER_10_251 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_decap_8 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_321 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_8 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_10_412 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_decap_8 FILLER_10_426 ();
 sg13g2_decap_8 FILLER_10_433 ();
 sg13g2_decap_8 FILLER_10_440 ();
 sg13g2_decap_8 FILLER_10_447 ();
 sg13g2_decap_8 FILLER_10_454 ();
 sg13g2_decap_8 FILLER_10_461 ();
 sg13g2_decap_8 FILLER_10_468 ();
 sg13g2_decap_8 FILLER_10_475 ();
 sg13g2_decap_8 FILLER_10_482 ();
 sg13g2_decap_8 FILLER_10_489 ();
 sg13g2_decap_8 FILLER_10_496 ();
 sg13g2_fill_1 FILLER_10_503 ();
 sg13g2_decap_4 FILLER_10_512 ();
 sg13g2_fill_1 FILLER_10_516 ();
 sg13g2_decap_8 FILLER_10_535 ();
 sg13g2_decap_8 FILLER_10_542 ();
 sg13g2_decap_4 FILLER_10_549 ();
 sg13g2_decap_8 FILLER_10_576 ();
 sg13g2_decap_8 FILLER_10_583 ();
 sg13g2_decap_8 FILLER_10_590 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_4 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_709 ();
 sg13g2_decap_8 FILLER_10_716 ();
 sg13g2_decap_8 FILLER_10_723 ();
 sg13g2_fill_2 FILLER_10_730 ();
 sg13g2_fill_1 FILLER_10_732 ();
 sg13g2_fill_1 FILLER_10_737 ();
 sg13g2_decap_4 FILLER_10_746 ();
 sg13g2_fill_2 FILLER_10_750 ();
 sg13g2_fill_1 FILLER_10_819 ();
 sg13g2_fill_2 FILLER_10_841 ();
 sg13g2_fill_1 FILLER_10_843 ();
 sg13g2_decap_8 FILLER_10_870 ();
 sg13g2_decap_8 FILLER_10_877 ();
 sg13g2_decap_8 FILLER_10_884 ();
 sg13g2_decap_8 FILLER_10_891 ();
 sg13g2_fill_1 FILLER_10_965 ();
 sg13g2_decap_8 FILLER_10_992 ();
 sg13g2_decap_8 FILLER_10_999 ();
 sg13g2_decap_4 FILLER_10_1006 ();
 sg13g2_decap_8 FILLER_10_1014 ();
 sg13g2_decap_8 FILLER_10_1021 ();
 sg13g2_decap_8 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_10_1035 ();
 sg13g2_fill_2 FILLER_10_1046 ();
 sg13g2_fill_1 FILLER_10_1048 ();
 sg13g2_fill_2 FILLER_10_1088 ();
 sg13g2_decap_8 FILLER_10_1116 ();
 sg13g2_decap_8 FILLER_10_1123 ();
 sg13g2_decap_4 FILLER_10_1130 ();
 sg13g2_fill_2 FILLER_10_1134 ();
 sg13g2_decap_8 FILLER_10_1177 ();
 sg13g2_decap_4 FILLER_10_1184 ();
 sg13g2_fill_2 FILLER_10_1188 ();
 sg13g2_fill_2 FILLER_10_1237 ();
 sg13g2_fill_1 FILLER_10_1239 ();
 sg13g2_decap_8 FILLER_10_1266 ();
 sg13g2_decap_8 FILLER_10_1273 ();
 sg13g2_decap_4 FILLER_10_1280 ();
 sg13g2_fill_1 FILLER_10_1284 ();
 sg13g2_decap_4 FILLER_10_1320 ();
 sg13g2_fill_2 FILLER_10_1324 ();
 sg13g2_decap_8 FILLER_10_1352 ();
 sg13g2_decap_8 FILLER_10_1359 ();
 sg13g2_fill_2 FILLER_10_1366 ();
 sg13g2_fill_1 FILLER_10_1368 ();
 sg13g2_fill_2 FILLER_10_1407 ();
 sg13g2_fill_1 FILLER_10_1409 ();
 sg13g2_fill_2 FILLER_10_1444 ();
 sg13g2_fill_2 FILLER_10_1454 ();
 sg13g2_fill_1 FILLER_10_1456 ();
 sg13g2_decap_8 FILLER_10_1460 ();
 sg13g2_decap_8 FILLER_10_1467 ();
 sg13g2_fill_2 FILLER_10_1474 ();
 sg13g2_fill_1 FILLER_10_1476 ();
 sg13g2_decap_8 FILLER_10_1499 ();
 sg13g2_fill_2 FILLER_10_1506 ();
 sg13g2_decap_8 FILLER_10_1534 ();
 sg13g2_decap_8 FILLER_10_1541 ();
 sg13g2_decap_8 FILLER_10_1548 ();
 sg13g2_decap_8 FILLER_10_1555 ();
 sg13g2_decap_8 FILLER_10_1562 ();
 sg13g2_decap_4 FILLER_10_1569 ();
 sg13g2_fill_1 FILLER_10_1573 ();
 sg13g2_fill_1 FILLER_10_1600 ();
 sg13g2_decap_8 FILLER_10_1632 ();
 sg13g2_decap_8 FILLER_10_1639 ();
 sg13g2_decap_8 FILLER_10_1646 ();
 sg13g2_decap_8 FILLER_10_1653 ();
 sg13g2_decap_8 FILLER_10_1668 ();
 sg13g2_decap_4 FILLER_10_1675 ();
 sg13g2_fill_2 FILLER_10_1679 ();
 sg13g2_decap_8 FILLER_10_1710 ();
 sg13g2_decap_8 FILLER_10_1717 ();
 sg13g2_fill_2 FILLER_10_1724 ();
 sg13g2_fill_1 FILLER_10_1726 ();
 sg13g2_decap_8 FILLER_10_1763 ();
 sg13g2_fill_1 FILLER_10_1770 ();
 sg13g2_decap_4 FILLER_10_1791 ();
 sg13g2_fill_2 FILLER_10_1795 ();
 sg13g2_fill_2 FILLER_10_1805 ();
 sg13g2_decap_8 FILLER_10_1823 ();
 sg13g2_fill_2 FILLER_10_1830 ();
 sg13g2_fill_2 FILLER_10_1861 ();
 sg13g2_decap_8 FILLER_10_1894 ();
 sg13g2_decap_8 FILLER_10_1901 ();
 sg13g2_decap_8 FILLER_10_1908 ();
 sg13g2_decap_8 FILLER_10_1915 ();
 sg13g2_decap_8 FILLER_10_1922 ();
 sg13g2_decap_8 FILLER_10_1929 ();
 sg13g2_decap_8 FILLER_10_1936 ();
 sg13g2_fill_1 FILLER_10_1943 ();
 sg13g2_decap_8 FILLER_10_1975 ();
 sg13g2_decap_8 FILLER_10_1982 ();
 sg13g2_fill_2 FILLER_10_1989 ();
 sg13g2_decap_8 FILLER_10_2025 ();
 sg13g2_decap_8 FILLER_10_2032 ();
 sg13g2_decap_8 FILLER_10_2039 ();
 sg13g2_decap_8 FILLER_10_2046 ();
 sg13g2_decap_4 FILLER_10_2053 ();
 sg13g2_fill_2 FILLER_10_2075 ();
 sg13g2_fill_1 FILLER_10_2077 ();
 sg13g2_decap_4 FILLER_10_2081 ();
 sg13g2_fill_1 FILLER_10_2085 ();
 sg13g2_decap_8 FILLER_10_2098 ();
 sg13g2_decap_8 FILLER_10_2105 ();
 sg13g2_fill_2 FILLER_10_2112 ();
 sg13g2_fill_1 FILLER_10_2114 ();
 sg13g2_fill_2 FILLER_10_2141 ();
 sg13g2_fill_1 FILLER_10_2169 ();
 sg13g2_decap_8 FILLER_10_2175 ();
 sg13g2_decap_4 FILLER_10_2182 ();
 sg13g2_decap_8 FILLER_10_2212 ();
 sg13g2_decap_8 FILLER_10_2219 ();
 sg13g2_fill_2 FILLER_10_2226 ();
 sg13g2_fill_1 FILLER_10_2228 ();
 sg13g2_decap_4 FILLER_10_2238 ();
 sg13g2_fill_1 FILLER_10_2242 ();
 sg13g2_decap_8 FILLER_10_2250 ();
 sg13g2_decap_8 FILLER_10_2257 ();
 sg13g2_decap_8 FILLER_10_2264 ();
 sg13g2_decap_8 FILLER_10_2271 ();
 sg13g2_decap_8 FILLER_10_2278 ();
 sg13g2_decap_8 FILLER_10_2285 ();
 sg13g2_decap_4 FILLER_10_2292 ();
 sg13g2_fill_2 FILLER_10_2296 ();
 sg13g2_decap_8 FILLER_10_2303 ();
 sg13g2_fill_1 FILLER_10_2336 ();
 sg13g2_fill_1 FILLER_10_2341 ();
 sg13g2_decap_8 FILLER_10_2368 ();
 sg13g2_fill_2 FILLER_10_2375 ();
 sg13g2_fill_1 FILLER_10_2377 ();
 sg13g2_decap_8 FILLER_10_2404 ();
 sg13g2_decap_8 FILLER_10_2424 ();
 sg13g2_fill_1 FILLER_10_2431 ();
 sg13g2_decap_8 FILLER_10_2439 ();
 sg13g2_fill_2 FILLER_10_2532 ();
 sg13g2_decap_8 FILLER_10_2565 ();
 sg13g2_decap_8 FILLER_10_2572 ();
 sg13g2_decap_4 FILLER_10_2579 ();
 sg13g2_fill_1 FILLER_10_2583 ();
 sg13g2_decap_8 FILLER_10_2645 ();
 sg13g2_decap_8 FILLER_10_2652 ();
 sg13g2_decap_8 FILLER_10_2659 ();
 sg13g2_decap_8 FILLER_10_2666 ();
 sg13g2_decap_8 FILLER_10_2673 ();
 sg13g2_decap_8 FILLER_10_2680 ();
 sg13g2_decap_8 FILLER_10_2687 ();
 sg13g2_decap_8 FILLER_10_2694 ();
 sg13g2_decap_8 FILLER_10_2701 ();
 sg13g2_decap_8 FILLER_10_2708 ();
 sg13g2_decap_8 FILLER_10_2715 ();
 sg13g2_decap_8 FILLER_10_2722 ();
 sg13g2_decap_8 FILLER_10_2729 ();
 sg13g2_decap_8 FILLER_10_2736 ();
 sg13g2_decap_8 FILLER_10_2743 ();
 sg13g2_decap_8 FILLER_10_2750 ();
 sg13g2_decap_8 FILLER_10_2757 ();
 sg13g2_decap_8 FILLER_10_2764 ();
 sg13g2_decap_8 FILLER_10_2771 ();
 sg13g2_decap_8 FILLER_10_2778 ();
 sg13g2_decap_8 FILLER_10_2785 ();
 sg13g2_decap_8 FILLER_10_2792 ();
 sg13g2_decap_8 FILLER_10_2799 ();
 sg13g2_decap_8 FILLER_10_2806 ();
 sg13g2_decap_8 FILLER_10_2813 ();
 sg13g2_decap_8 FILLER_10_2820 ();
 sg13g2_decap_8 FILLER_10_2827 ();
 sg13g2_decap_8 FILLER_10_2834 ();
 sg13g2_decap_8 FILLER_10_2841 ();
 sg13g2_decap_8 FILLER_10_2848 ();
 sg13g2_decap_8 FILLER_10_2855 ();
 sg13g2_decap_8 FILLER_10_2862 ();
 sg13g2_decap_8 FILLER_10_2869 ();
 sg13g2_decap_8 FILLER_10_2876 ();
 sg13g2_decap_8 FILLER_10_2883 ();
 sg13g2_decap_8 FILLER_10_2890 ();
 sg13g2_decap_8 FILLER_10_2897 ();
 sg13g2_decap_8 FILLER_10_2904 ();
 sg13g2_decap_8 FILLER_10_2911 ();
 sg13g2_decap_8 FILLER_10_2918 ();
 sg13g2_decap_8 FILLER_10_2925 ();
 sg13g2_decap_8 FILLER_10_2932 ();
 sg13g2_decap_8 FILLER_10_2939 ();
 sg13g2_decap_8 FILLER_10_2946 ();
 sg13g2_decap_8 FILLER_10_2953 ();
 sg13g2_decap_8 FILLER_10_2960 ();
 sg13g2_decap_8 FILLER_10_2967 ();
 sg13g2_decap_8 FILLER_10_2974 ();
 sg13g2_decap_8 FILLER_10_2981 ();
 sg13g2_decap_8 FILLER_10_2988 ();
 sg13g2_decap_8 FILLER_10_2995 ();
 sg13g2_decap_8 FILLER_10_3002 ();
 sg13g2_decap_8 FILLER_10_3009 ();
 sg13g2_decap_8 FILLER_10_3016 ();
 sg13g2_decap_8 FILLER_10_3023 ();
 sg13g2_decap_8 FILLER_10_3030 ();
 sg13g2_decap_8 FILLER_10_3037 ();
 sg13g2_decap_8 FILLER_10_3044 ();
 sg13g2_decap_8 FILLER_10_3051 ();
 sg13g2_decap_8 FILLER_10_3058 ();
 sg13g2_decap_8 FILLER_10_3065 ();
 sg13g2_decap_8 FILLER_10_3072 ();
 sg13g2_decap_8 FILLER_10_3079 ();
 sg13g2_decap_8 FILLER_10_3086 ();
 sg13g2_decap_8 FILLER_10_3093 ();
 sg13g2_decap_8 FILLER_10_3100 ();
 sg13g2_decap_8 FILLER_10_3107 ();
 sg13g2_decap_8 FILLER_10_3114 ();
 sg13g2_decap_8 FILLER_10_3121 ();
 sg13g2_decap_8 FILLER_10_3128 ();
 sg13g2_decap_8 FILLER_10_3135 ();
 sg13g2_decap_8 FILLER_10_3142 ();
 sg13g2_decap_8 FILLER_10_3149 ();
 sg13g2_decap_8 FILLER_10_3156 ();
 sg13g2_decap_8 FILLER_10_3163 ();
 sg13g2_decap_8 FILLER_10_3170 ();
 sg13g2_decap_8 FILLER_10_3177 ();
 sg13g2_decap_8 FILLER_10_3184 ();
 sg13g2_decap_8 FILLER_10_3191 ();
 sg13g2_decap_8 FILLER_10_3198 ();
 sg13g2_decap_8 FILLER_10_3205 ();
 sg13g2_decap_8 FILLER_10_3212 ();
 sg13g2_decap_8 FILLER_10_3219 ();
 sg13g2_decap_8 FILLER_10_3226 ();
 sg13g2_decap_8 FILLER_10_3233 ();
 sg13g2_decap_8 FILLER_10_3240 ();
 sg13g2_decap_8 FILLER_10_3247 ();
 sg13g2_decap_8 FILLER_10_3254 ();
 sg13g2_decap_8 FILLER_10_3261 ();
 sg13g2_decap_8 FILLER_10_3268 ();
 sg13g2_decap_8 FILLER_10_3275 ();
 sg13g2_decap_8 FILLER_10_3282 ();
 sg13g2_decap_8 FILLER_10_3289 ();
 sg13g2_decap_8 FILLER_10_3296 ();
 sg13g2_decap_8 FILLER_10_3303 ();
 sg13g2_decap_8 FILLER_10_3310 ();
 sg13g2_decap_8 FILLER_10_3317 ();
 sg13g2_decap_8 FILLER_10_3324 ();
 sg13g2_decap_8 FILLER_10_3331 ();
 sg13g2_decap_8 FILLER_10_3338 ();
 sg13g2_decap_8 FILLER_10_3345 ();
 sg13g2_decap_8 FILLER_10_3352 ();
 sg13g2_decap_8 FILLER_10_3359 ();
 sg13g2_decap_8 FILLER_10_3366 ();
 sg13g2_decap_8 FILLER_10_3373 ();
 sg13g2_decap_8 FILLER_10_3380 ();
 sg13g2_decap_8 FILLER_10_3387 ();
 sg13g2_decap_8 FILLER_10_3394 ();
 sg13g2_decap_8 FILLER_10_3401 ();
 sg13g2_decap_8 FILLER_10_3408 ();
 sg13g2_decap_8 FILLER_10_3415 ();
 sg13g2_decap_8 FILLER_10_3422 ();
 sg13g2_decap_8 FILLER_10_3429 ();
 sg13g2_decap_8 FILLER_10_3436 ();
 sg13g2_decap_8 FILLER_10_3443 ();
 sg13g2_decap_8 FILLER_10_3450 ();
 sg13g2_decap_8 FILLER_10_3457 ();
 sg13g2_decap_8 FILLER_10_3464 ();
 sg13g2_decap_8 FILLER_10_3471 ();
 sg13g2_decap_8 FILLER_10_3478 ();
 sg13g2_decap_8 FILLER_10_3485 ();
 sg13g2_decap_8 FILLER_10_3492 ();
 sg13g2_decap_8 FILLER_10_3499 ();
 sg13g2_decap_8 FILLER_10_3506 ();
 sg13g2_decap_8 FILLER_10_3513 ();
 sg13g2_decap_8 FILLER_10_3520 ();
 sg13g2_decap_8 FILLER_10_3527 ();
 sg13g2_decap_8 FILLER_10_3534 ();
 sg13g2_decap_8 FILLER_10_3541 ();
 sg13g2_decap_8 FILLER_10_3548 ();
 sg13g2_decap_8 FILLER_10_3555 ();
 sg13g2_decap_8 FILLER_10_3562 ();
 sg13g2_decap_8 FILLER_10_3569 ();
 sg13g2_decap_4 FILLER_10_3576 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_4 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_108 ();
 sg13g2_decap_8 FILLER_11_115 ();
 sg13g2_fill_2 FILLER_11_122 ();
 sg13g2_fill_1 FILLER_11_124 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_fill_2 FILLER_11_179 ();
 sg13g2_fill_1 FILLER_11_181 ();
 sg13g2_decap_8 FILLER_11_199 ();
 sg13g2_decap_8 FILLER_11_206 ();
 sg13g2_decap_8 FILLER_11_213 ();
 sg13g2_decap_8 FILLER_11_220 ();
 sg13g2_decap_8 FILLER_11_227 ();
 sg13g2_decap_8 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_241 ();
 sg13g2_decap_8 FILLER_11_248 ();
 sg13g2_decap_8 FILLER_11_255 ();
 sg13g2_decap_8 FILLER_11_262 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_283 ();
 sg13g2_decap_4 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_431 ();
 sg13g2_decap_8 FILLER_11_438 ();
 sg13g2_decap_8 FILLER_11_445 ();
 sg13g2_decap_8 FILLER_11_452 ();
 sg13g2_decap_8 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_466 ();
 sg13g2_decap_8 FILLER_11_473 ();
 sg13g2_decap_8 FILLER_11_480 ();
 sg13g2_decap_8 FILLER_11_487 ();
 sg13g2_decap_8 FILLER_11_494 ();
 sg13g2_fill_2 FILLER_11_527 ();
 sg13g2_fill_2 FILLER_11_542 ();
 sg13g2_fill_1 FILLER_11_544 ();
 sg13g2_decap_4 FILLER_11_592 ();
 sg13g2_decap_8 FILLER_11_640 ();
 sg13g2_decap_8 FILLER_11_647 ();
 sg13g2_fill_2 FILLER_11_654 ();
 sg13g2_decap_8 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_fill_1 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_753 ();
 sg13g2_fill_2 FILLER_11_760 ();
 sg13g2_fill_2 FILLER_11_775 ();
 sg13g2_fill_1 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_786 ();
 sg13g2_decap_8 FILLER_11_793 ();
 sg13g2_fill_2 FILLER_11_800 ();
 sg13g2_fill_2 FILLER_11_807 ();
 sg13g2_fill_1 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_822 ();
 sg13g2_fill_2 FILLER_11_829 ();
 sg13g2_decap_8 FILLER_11_836 ();
 sg13g2_decap_4 FILLER_11_843 ();
 sg13g2_fill_1 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_916 ();
 sg13g2_fill_2 FILLER_11_923 ();
 sg13g2_decap_8 FILLER_11_933 ();
 sg13g2_fill_2 FILLER_11_945 ();
 sg13g2_fill_1 FILLER_11_947 ();
 sg13g2_fill_1 FILLER_11_1000 ();
 sg13g2_decap_8 FILLER_11_1006 ();
 sg13g2_decap_8 FILLER_11_1013 ();
 sg13g2_decap_4 FILLER_11_1020 ();
 sg13g2_fill_1 FILLER_11_1024 ();
 sg13g2_decap_4 FILLER_11_1031 ();
 sg13g2_fill_1 FILLER_11_1035 ();
 sg13g2_decap_8 FILLER_11_1041 ();
 sg13g2_decap_8 FILLER_11_1051 ();
 sg13g2_fill_2 FILLER_11_1058 ();
 sg13g2_decap_4 FILLER_11_1064 ();
 sg13g2_fill_2 FILLER_11_1078 ();
 sg13g2_decap_8 FILLER_11_1092 ();
 sg13g2_fill_2 FILLER_11_1099 ();
 sg13g2_decap_8 FILLER_11_1109 ();
 sg13g2_decap_8 FILLER_11_1116 ();
 sg13g2_decap_4 FILLER_11_1123 ();
 sg13g2_fill_2 FILLER_11_1127 ();
 sg13g2_fill_1 FILLER_11_1160 ();
 sg13g2_decap_8 FILLER_11_1175 ();
 sg13g2_decap_8 FILLER_11_1182 ();
 sg13g2_decap_4 FILLER_11_1189 ();
 sg13g2_fill_2 FILLER_11_1193 ();
 sg13g2_fill_1 FILLER_11_1234 ();
 sg13g2_fill_2 FILLER_11_1243 ();
 sg13g2_fill_2 FILLER_11_1261 ();
 sg13g2_decap_8 FILLER_11_1276 ();
 sg13g2_fill_2 FILLER_11_1283 ();
 sg13g2_fill_1 FILLER_11_1285 ();
 sg13g2_decap_8 FILLER_11_1312 ();
 sg13g2_fill_2 FILLER_11_1319 ();
 sg13g2_decap_8 FILLER_11_1347 ();
 sg13g2_decap_8 FILLER_11_1354 ();
 sg13g2_decap_8 FILLER_11_1361 ();
 sg13g2_decap_4 FILLER_11_1368 ();
 sg13g2_fill_1 FILLER_11_1372 ();
 sg13g2_decap_4 FILLER_11_1376 ();
 sg13g2_fill_2 FILLER_11_1380 ();
 sg13g2_decap_8 FILLER_11_1416 ();
 sg13g2_fill_2 FILLER_11_1423 ();
 sg13g2_fill_1 FILLER_11_1425 ();
 sg13g2_fill_2 FILLER_11_1431 ();
 sg13g2_decap_4 FILLER_11_1438 ();
 sg13g2_decap_8 FILLER_11_1446 ();
 sg13g2_fill_1 FILLER_11_1453 ();
 sg13g2_decap_4 FILLER_11_1467 ();
 sg13g2_decap_8 FILLER_11_1505 ();
 sg13g2_decap_8 FILLER_11_1512 ();
 sg13g2_decap_4 FILLER_11_1545 ();
 sg13g2_fill_2 FILLER_11_1549 ();
 sg13g2_decap_4 FILLER_11_1554 ();
 sg13g2_fill_2 FILLER_11_1558 ();
 sg13g2_decap_4 FILLER_11_1564 ();
 sg13g2_fill_1 FILLER_11_1568 ();
 sg13g2_decap_4 FILLER_11_1643 ();
 sg13g2_decap_8 FILLER_11_1651 ();
 sg13g2_decap_8 FILLER_11_1658 ();
 sg13g2_fill_1 FILLER_11_1665 ();
 sg13g2_decap_8 FILLER_11_1670 ();
 sg13g2_fill_2 FILLER_11_1677 ();
 sg13g2_fill_1 FILLER_11_1684 ();
 sg13g2_decap_8 FILLER_11_1696 ();
 sg13g2_decap_8 FILLER_11_1703 ();
 sg13g2_decap_8 FILLER_11_1710 ();
 sg13g2_decap_8 FILLER_11_1717 ();
 sg13g2_decap_4 FILLER_11_1724 ();
 sg13g2_fill_1 FILLER_11_1770 ();
 sg13g2_decap_8 FILLER_11_1823 ();
 sg13g2_decap_8 FILLER_11_1830 ();
 sg13g2_decap_8 FILLER_11_1837 ();
 sg13g2_decap_8 FILLER_11_1844 ();
 sg13g2_fill_1 FILLER_11_1851 ();
 sg13g2_decap_8 FILLER_11_1855 ();
 sg13g2_decap_8 FILLER_11_1862 ();
 sg13g2_decap_8 FILLER_11_1869 ();
 sg13g2_decap_8 FILLER_11_1876 ();
 sg13g2_decap_8 FILLER_11_1883 ();
 sg13g2_decap_8 FILLER_11_1890 ();
 sg13g2_decap_8 FILLER_11_1897 ();
 sg13g2_fill_1 FILLER_11_1904 ();
 sg13g2_fill_1 FILLER_11_1934 ();
 sg13g2_decap_8 FILLER_11_1972 ();
 sg13g2_decap_8 FILLER_11_1979 ();
 sg13g2_decap_8 FILLER_11_2031 ();
 sg13g2_fill_1 FILLER_11_2038 ();
 sg13g2_decap_4 FILLER_11_2068 ();
 sg13g2_fill_1 FILLER_11_2072 ();
 sg13g2_decap_8 FILLER_11_2144 ();
 sg13g2_fill_1 FILLER_11_2151 ();
 sg13g2_fill_2 FILLER_11_2181 ();
 sg13g2_fill_1 FILLER_11_2183 ();
 sg13g2_decap_8 FILLER_11_2210 ();
 sg13g2_decap_8 FILLER_11_2217 ();
 sg13g2_decap_8 FILLER_11_2224 ();
 sg13g2_fill_1 FILLER_11_2231 ();
 sg13g2_decap_4 FILLER_11_2284 ();
 sg13g2_fill_1 FILLER_11_2288 ();
 sg13g2_fill_1 FILLER_11_2294 ();
 sg13g2_decap_4 FILLER_11_2321 ();
 sg13g2_fill_2 FILLER_11_2325 ();
 sg13g2_fill_2 FILLER_11_2335 ();
 sg13g2_fill_2 FILLER_11_2350 ();
 sg13g2_decap_8 FILLER_11_2378 ();
 sg13g2_decap_8 FILLER_11_2385 ();
 sg13g2_decap_4 FILLER_11_2392 ();
 sg13g2_decap_8 FILLER_11_2430 ();
 sg13g2_decap_8 FILLER_11_2437 ();
 sg13g2_decap_8 FILLER_11_2444 ();
 sg13g2_decap_4 FILLER_11_2451 ();
 sg13g2_decap_8 FILLER_11_2481 ();
 sg13g2_decap_8 FILLER_11_2488 ();
 sg13g2_decap_8 FILLER_11_2495 ();
 sg13g2_decap_8 FILLER_11_2502 ();
 sg13g2_decap_8 FILLER_11_2509 ();
 sg13g2_decap_4 FILLER_11_2516 ();
 sg13g2_fill_2 FILLER_11_2520 ();
 sg13g2_fill_2 FILLER_11_2553 ();
 sg13g2_decap_8 FILLER_11_2654 ();
 sg13g2_decap_8 FILLER_11_2661 ();
 sg13g2_decap_8 FILLER_11_2668 ();
 sg13g2_decap_8 FILLER_11_2675 ();
 sg13g2_decap_8 FILLER_11_2682 ();
 sg13g2_decap_8 FILLER_11_2689 ();
 sg13g2_decap_8 FILLER_11_2696 ();
 sg13g2_decap_8 FILLER_11_2703 ();
 sg13g2_decap_8 FILLER_11_2710 ();
 sg13g2_decap_8 FILLER_11_2717 ();
 sg13g2_decap_8 FILLER_11_2724 ();
 sg13g2_decap_8 FILLER_11_2731 ();
 sg13g2_decap_8 FILLER_11_2738 ();
 sg13g2_decap_8 FILLER_11_2745 ();
 sg13g2_decap_8 FILLER_11_2752 ();
 sg13g2_decap_8 FILLER_11_2759 ();
 sg13g2_decap_8 FILLER_11_2766 ();
 sg13g2_decap_8 FILLER_11_2773 ();
 sg13g2_decap_8 FILLER_11_2780 ();
 sg13g2_decap_8 FILLER_11_2787 ();
 sg13g2_decap_8 FILLER_11_2794 ();
 sg13g2_decap_8 FILLER_11_2801 ();
 sg13g2_decap_8 FILLER_11_2808 ();
 sg13g2_decap_8 FILLER_11_2815 ();
 sg13g2_decap_8 FILLER_11_2822 ();
 sg13g2_decap_8 FILLER_11_2829 ();
 sg13g2_decap_8 FILLER_11_2836 ();
 sg13g2_decap_8 FILLER_11_2843 ();
 sg13g2_decap_8 FILLER_11_2850 ();
 sg13g2_decap_8 FILLER_11_2857 ();
 sg13g2_decap_8 FILLER_11_2864 ();
 sg13g2_decap_8 FILLER_11_2871 ();
 sg13g2_decap_8 FILLER_11_2878 ();
 sg13g2_decap_8 FILLER_11_2885 ();
 sg13g2_decap_8 FILLER_11_2892 ();
 sg13g2_decap_8 FILLER_11_2899 ();
 sg13g2_decap_8 FILLER_11_2906 ();
 sg13g2_decap_8 FILLER_11_2913 ();
 sg13g2_decap_8 FILLER_11_2920 ();
 sg13g2_decap_8 FILLER_11_2927 ();
 sg13g2_decap_8 FILLER_11_2934 ();
 sg13g2_decap_8 FILLER_11_2941 ();
 sg13g2_decap_8 FILLER_11_2948 ();
 sg13g2_decap_8 FILLER_11_2955 ();
 sg13g2_decap_8 FILLER_11_2962 ();
 sg13g2_decap_8 FILLER_11_2969 ();
 sg13g2_decap_8 FILLER_11_2976 ();
 sg13g2_decap_8 FILLER_11_2983 ();
 sg13g2_decap_8 FILLER_11_2990 ();
 sg13g2_decap_8 FILLER_11_2997 ();
 sg13g2_decap_8 FILLER_11_3004 ();
 sg13g2_decap_8 FILLER_11_3011 ();
 sg13g2_decap_8 FILLER_11_3018 ();
 sg13g2_decap_8 FILLER_11_3025 ();
 sg13g2_decap_8 FILLER_11_3032 ();
 sg13g2_decap_8 FILLER_11_3039 ();
 sg13g2_decap_8 FILLER_11_3046 ();
 sg13g2_decap_8 FILLER_11_3053 ();
 sg13g2_decap_8 FILLER_11_3060 ();
 sg13g2_decap_8 FILLER_11_3067 ();
 sg13g2_decap_8 FILLER_11_3074 ();
 sg13g2_decap_8 FILLER_11_3081 ();
 sg13g2_decap_8 FILLER_11_3088 ();
 sg13g2_decap_8 FILLER_11_3095 ();
 sg13g2_decap_8 FILLER_11_3102 ();
 sg13g2_decap_8 FILLER_11_3109 ();
 sg13g2_decap_8 FILLER_11_3116 ();
 sg13g2_decap_8 FILLER_11_3123 ();
 sg13g2_decap_8 FILLER_11_3130 ();
 sg13g2_decap_8 FILLER_11_3137 ();
 sg13g2_decap_8 FILLER_11_3144 ();
 sg13g2_decap_8 FILLER_11_3151 ();
 sg13g2_decap_8 FILLER_11_3158 ();
 sg13g2_decap_8 FILLER_11_3165 ();
 sg13g2_decap_8 FILLER_11_3172 ();
 sg13g2_decap_8 FILLER_11_3179 ();
 sg13g2_decap_8 FILLER_11_3186 ();
 sg13g2_decap_8 FILLER_11_3193 ();
 sg13g2_decap_8 FILLER_11_3200 ();
 sg13g2_decap_8 FILLER_11_3207 ();
 sg13g2_decap_8 FILLER_11_3214 ();
 sg13g2_decap_8 FILLER_11_3221 ();
 sg13g2_decap_8 FILLER_11_3228 ();
 sg13g2_decap_8 FILLER_11_3235 ();
 sg13g2_decap_8 FILLER_11_3242 ();
 sg13g2_decap_8 FILLER_11_3249 ();
 sg13g2_decap_8 FILLER_11_3256 ();
 sg13g2_decap_8 FILLER_11_3263 ();
 sg13g2_decap_8 FILLER_11_3270 ();
 sg13g2_decap_8 FILLER_11_3277 ();
 sg13g2_decap_8 FILLER_11_3284 ();
 sg13g2_decap_8 FILLER_11_3291 ();
 sg13g2_decap_8 FILLER_11_3298 ();
 sg13g2_decap_8 FILLER_11_3305 ();
 sg13g2_decap_8 FILLER_11_3312 ();
 sg13g2_decap_8 FILLER_11_3319 ();
 sg13g2_decap_8 FILLER_11_3326 ();
 sg13g2_decap_8 FILLER_11_3333 ();
 sg13g2_decap_8 FILLER_11_3340 ();
 sg13g2_decap_8 FILLER_11_3347 ();
 sg13g2_decap_8 FILLER_11_3354 ();
 sg13g2_decap_8 FILLER_11_3361 ();
 sg13g2_decap_8 FILLER_11_3368 ();
 sg13g2_decap_8 FILLER_11_3375 ();
 sg13g2_decap_8 FILLER_11_3382 ();
 sg13g2_decap_8 FILLER_11_3389 ();
 sg13g2_decap_8 FILLER_11_3396 ();
 sg13g2_decap_8 FILLER_11_3403 ();
 sg13g2_decap_8 FILLER_11_3410 ();
 sg13g2_decap_8 FILLER_11_3417 ();
 sg13g2_decap_8 FILLER_11_3424 ();
 sg13g2_decap_8 FILLER_11_3431 ();
 sg13g2_decap_8 FILLER_11_3438 ();
 sg13g2_decap_8 FILLER_11_3445 ();
 sg13g2_decap_8 FILLER_11_3452 ();
 sg13g2_decap_8 FILLER_11_3459 ();
 sg13g2_decap_8 FILLER_11_3466 ();
 sg13g2_decap_8 FILLER_11_3473 ();
 sg13g2_decap_8 FILLER_11_3480 ();
 sg13g2_decap_8 FILLER_11_3487 ();
 sg13g2_decap_8 FILLER_11_3494 ();
 sg13g2_decap_8 FILLER_11_3501 ();
 sg13g2_decap_8 FILLER_11_3508 ();
 sg13g2_decap_8 FILLER_11_3515 ();
 sg13g2_decap_8 FILLER_11_3522 ();
 sg13g2_decap_8 FILLER_11_3529 ();
 sg13g2_decap_8 FILLER_11_3536 ();
 sg13g2_decap_8 FILLER_11_3543 ();
 sg13g2_decap_8 FILLER_11_3550 ();
 sg13g2_decap_8 FILLER_11_3557 ();
 sg13g2_decap_8 FILLER_11_3564 ();
 sg13g2_decap_8 FILLER_11_3571 ();
 sg13g2_fill_2 FILLER_11_3578 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_fill_2 FILLER_12_49 ();
 sg13g2_fill_1 FILLER_12_51 ();
 sg13g2_fill_2 FILLER_12_55 ();
 sg13g2_decap_8 FILLER_12_62 ();
 sg13g2_decap_8 FILLER_12_69 ();
 sg13g2_decap_4 FILLER_12_76 ();
 sg13g2_decap_4 FILLER_12_122 ();
 sg13g2_decap_8 FILLER_12_152 ();
 sg13g2_decap_8 FILLER_12_159 ();
 sg13g2_decap_4 FILLER_12_166 ();
 sg13g2_fill_2 FILLER_12_170 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_4 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_218 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_4 FILLER_12_266 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_fill_1 FILLER_12_279 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_fill_2 FILLER_12_323 ();
 sg13g2_fill_1 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_4 FILLER_12_394 ();
 sg13g2_fill_2 FILLER_12_398 ();
 sg13g2_decap_8 FILLER_12_426 ();
 sg13g2_decap_8 FILLER_12_433 ();
 sg13g2_decap_8 FILLER_12_440 ();
 sg13g2_decap_8 FILLER_12_447 ();
 sg13g2_decap_8 FILLER_12_454 ();
 sg13g2_decap_8 FILLER_12_461 ();
 sg13g2_decap_8 FILLER_12_468 ();
 sg13g2_decap_8 FILLER_12_475 ();
 sg13g2_decap_4 FILLER_12_482 ();
 sg13g2_fill_1 FILLER_12_486 ();
 sg13g2_fill_1 FILLER_12_539 ();
 sg13g2_decap_4 FILLER_12_592 ();
 sg13g2_fill_2 FILLER_12_596 ();
 sg13g2_decap_8 FILLER_12_636 ();
 sg13g2_decap_8 FILLER_12_643 ();
 sg13g2_decap_8 FILLER_12_650 ();
 sg13g2_decap_8 FILLER_12_657 ();
 sg13g2_fill_1 FILLER_12_668 ();
 sg13g2_decap_8 FILLER_12_674 ();
 sg13g2_decap_4 FILLER_12_681 ();
 sg13g2_fill_1 FILLER_12_685 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_4 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_fill_1 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_796 ();
 sg13g2_decap_4 FILLER_12_803 ();
 sg13g2_decap_4 FILLER_12_810 ();
 sg13g2_decap_8 FILLER_12_845 ();
 sg13g2_fill_1 FILLER_12_852 ();
 sg13g2_decap_4 FILLER_12_856 ();
 sg13g2_fill_2 FILLER_12_860 ();
 sg13g2_fill_2 FILLER_12_896 ();
 sg13g2_decap_8 FILLER_12_924 ();
 sg13g2_decap_8 FILLER_12_931 ();
 sg13g2_decap_4 FILLER_12_938 ();
 sg13g2_decap_8 FILLER_12_946 ();
 sg13g2_decap_8 FILLER_12_953 ();
 sg13g2_decap_4 FILLER_12_960 ();
 sg13g2_fill_2 FILLER_12_964 ();
 sg13g2_fill_1 FILLER_12_970 ();
 sg13g2_decap_4 FILLER_12_1062 ();
 sg13g2_fill_2 FILLER_12_1066 ();
 sg13g2_fill_1 FILLER_12_1073 ();
 sg13g2_decap_8 FILLER_12_1082 ();
 sg13g2_decap_8 FILLER_12_1089 ();
 sg13g2_decap_8 FILLER_12_1096 ();
 sg13g2_fill_1 FILLER_12_1103 ();
 sg13g2_fill_1 FILLER_12_1156 ();
 sg13g2_decap_8 FILLER_12_1183 ();
 sg13g2_decap_8 FILLER_12_1190 ();
 sg13g2_decap_8 FILLER_12_1197 ();
 sg13g2_decap_4 FILLER_12_1208 ();
 sg13g2_fill_1 FILLER_12_1212 ();
 sg13g2_fill_2 FILLER_12_1218 ();
 sg13g2_fill_2 FILLER_12_1230 ();
 sg13g2_fill_2 FILLER_12_1236 ();
 sg13g2_fill_1 FILLER_12_1238 ();
 sg13g2_decap_8 FILLER_12_1285 ();
 sg13g2_fill_2 FILLER_12_1292 ();
 sg13g2_fill_1 FILLER_12_1294 ();
 sg13g2_decap_8 FILLER_12_1302 ();
 sg13g2_decap_4 FILLER_12_1309 ();
 sg13g2_fill_2 FILLER_12_1313 ();
 sg13g2_decap_8 FILLER_12_1323 ();
 sg13g2_decap_4 FILLER_12_1330 ();
 sg13g2_decap_8 FILLER_12_1360 ();
 sg13g2_fill_1 FILLER_12_1367 ();
 sg13g2_fill_2 FILLER_12_1394 ();
 sg13g2_fill_1 FILLER_12_1396 ();
 sg13g2_fill_2 FILLER_12_1454 ();
 sg13g2_fill_1 FILLER_12_1456 ();
 sg13g2_decap_4 FILLER_12_1464 ();
 sg13g2_fill_1 FILLER_12_1468 ();
 sg13g2_fill_1 FILLER_12_1482 ();
 sg13g2_decap_8 FILLER_12_1509 ();
 sg13g2_decap_4 FILLER_12_1516 ();
 sg13g2_fill_2 FILLER_12_1520 ();
 sg13g2_fill_1 FILLER_12_1574 ();
 sg13g2_fill_2 FILLER_12_1583 ();
 sg13g2_decap_8 FILLER_12_1593 ();
 sg13g2_decap_8 FILLER_12_1600 ();
 sg13g2_fill_1 FILLER_12_1607 ();
 sg13g2_fill_1 FILLER_12_1623 ();
 sg13g2_decap_4 FILLER_12_1632 ();
 sg13g2_decap_8 FILLER_12_1662 ();
 sg13g2_decap_4 FILLER_12_1669 ();
 sg13g2_fill_1 FILLER_12_1673 ();
 sg13g2_fill_2 FILLER_12_1682 ();
 sg13g2_fill_2 FILLER_12_1714 ();
 sg13g2_fill_1 FILLER_12_1721 ();
 sg13g2_decap_4 FILLER_12_1748 ();
 sg13g2_fill_1 FILLER_12_1752 ();
 sg13g2_decap_8 FILLER_12_1761 ();
 sg13g2_fill_2 FILLER_12_1768 ();
 sg13g2_fill_1 FILLER_12_1770 ();
 sg13g2_decap_8 FILLER_12_1823 ();
 sg13g2_fill_2 FILLER_12_1830 ();
 sg13g2_fill_1 FILLER_12_1832 ();
 sg13g2_decap_8 FILLER_12_1867 ();
 sg13g2_fill_2 FILLER_12_1874 ();
 sg13g2_fill_2 FILLER_12_1936 ();
 sg13g2_fill_2 FILLER_12_1976 ();
 sg13g2_fill_1 FILLER_12_2038 ();
 sg13g2_decap_8 FILLER_12_2056 ();
 sg13g2_fill_2 FILLER_12_2063 ();
 sg13g2_decap_8 FILLER_12_2094 ();
 sg13g2_decap_8 FILLER_12_2101 ();
 sg13g2_fill_2 FILLER_12_2108 ();
 sg13g2_decap_8 FILLER_12_2135 ();
 sg13g2_fill_2 FILLER_12_2142 ();
 sg13g2_fill_1 FILLER_12_2144 ();
 sg13g2_fill_1 FILLER_12_2171 ();
 sg13g2_decap_8 FILLER_12_2212 ();
 sg13g2_decap_8 FILLER_12_2219 ();
 sg13g2_decap_4 FILLER_12_2226 ();
 sg13g2_fill_1 FILLER_12_2230 ();
 sg13g2_decap_4 FILLER_12_2283 ();
 sg13g2_fill_1 FILLER_12_2325 ();
 sg13g2_decap_8 FILLER_12_2357 ();
 sg13g2_decap_8 FILLER_12_2364 ();
 sg13g2_decap_4 FILLER_12_2371 ();
 sg13g2_decap_8 FILLER_12_2379 ();
 sg13g2_fill_1 FILLER_12_2386 ();
 sg13g2_fill_2 FILLER_12_2421 ();
 sg13g2_fill_1 FILLER_12_2423 ();
 sg13g2_decap_8 FILLER_12_2428 ();
 sg13g2_decap_8 FILLER_12_2435 ();
 sg13g2_decap_8 FILLER_12_2481 ();
 sg13g2_decap_8 FILLER_12_2488 ();
 sg13g2_decap_8 FILLER_12_2495 ();
 sg13g2_decap_8 FILLER_12_2502 ();
 sg13g2_fill_2 FILLER_12_2509 ();
 sg13g2_fill_1 FILLER_12_2511 ();
 sg13g2_decap_4 FILLER_12_2515 ();
 sg13g2_fill_2 FILLER_12_2519 ();
 sg13g2_decap_4 FILLER_12_2537 ();
 sg13g2_fill_2 FILLER_12_2549 ();
 sg13g2_fill_2 FILLER_12_2562 ();
 sg13g2_fill_1 FILLER_12_2564 ();
 sg13g2_decap_8 FILLER_12_2569 ();
 sg13g2_decap_8 FILLER_12_2576 ();
 sg13g2_decap_4 FILLER_12_2583 ();
 sg13g2_decap_8 FILLER_12_2594 ();
 sg13g2_decap_8 FILLER_12_2601 ();
 sg13g2_fill_2 FILLER_12_2608 ();
 sg13g2_decap_4 FILLER_12_2614 ();
 sg13g2_decap_8 FILLER_12_2662 ();
 sg13g2_decap_8 FILLER_12_2669 ();
 sg13g2_decap_8 FILLER_12_2676 ();
 sg13g2_decap_8 FILLER_12_2683 ();
 sg13g2_decap_8 FILLER_12_2690 ();
 sg13g2_decap_8 FILLER_12_2697 ();
 sg13g2_decap_8 FILLER_12_2704 ();
 sg13g2_decap_8 FILLER_12_2711 ();
 sg13g2_decap_8 FILLER_12_2718 ();
 sg13g2_decap_8 FILLER_12_2725 ();
 sg13g2_decap_8 FILLER_12_2732 ();
 sg13g2_decap_8 FILLER_12_2739 ();
 sg13g2_decap_8 FILLER_12_2746 ();
 sg13g2_decap_8 FILLER_12_2753 ();
 sg13g2_decap_8 FILLER_12_2760 ();
 sg13g2_decap_8 FILLER_12_2767 ();
 sg13g2_decap_8 FILLER_12_2774 ();
 sg13g2_decap_8 FILLER_12_2781 ();
 sg13g2_decap_8 FILLER_12_2788 ();
 sg13g2_decap_8 FILLER_12_2795 ();
 sg13g2_decap_8 FILLER_12_2802 ();
 sg13g2_decap_8 FILLER_12_2809 ();
 sg13g2_decap_8 FILLER_12_2816 ();
 sg13g2_decap_8 FILLER_12_2823 ();
 sg13g2_decap_8 FILLER_12_2830 ();
 sg13g2_decap_8 FILLER_12_2837 ();
 sg13g2_decap_8 FILLER_12_2844 ();
 sg13g2_decap_8 FILLER_12_2851 ();
 sg13g2_decap_8 FILLER_12_2858 ();
 sg13g2_decap_8 FILLER_12_2865 ();
 sg13g2_decap_8 FILLER_12_2872 ();
 sg13g2_decap_8 FILLER_12_2879 ();
 sg13g2_decap_8 FILLER_12_2886 ();
 sg13g2_decap_8 FILLER_12_2893 ();
 sg13g2_decap_8 FILLER_12_2900 ();
 sg13g2_decap_8 FILLER_12_2907 ();
 sg13g2_decap_8 FILLER_12_2914 ();
 sg13g2_decap_8 FILLER_12_2921 ();
 sg13g2_decap_8 FILLER_12_2928 ();
 sg13g2_decap_8 FILLER_12_2935 ();
 sg13g2_decap_8 FILLER_12_2942 ();
 sg13g2_decap_8 FILLER_12_2949 ();
 sg13g2_decap_8 FILLER_12_2956 ();
 sg13g2_decap_8 FILLER_12_2963 ();
 sg13g2_decap_8 FILLER_12_2970 ();
 sg13g2_decap_8 FILLER_12_2977 ();
 sg13g2_decap_8 FILLER_12_2984 ();
 sg13g2_decap_8 FILLER_12_2991 ();
 sg13g2_decap_8 FILLER_12_2998 ();
 sg13g2_decap_8 FILLER_12_3005 ();
 sg13g2_decap_8 FILLER_12_3012 ();
 sg13g2_decap_8 FILLER_12_3019 ();
 sg13g2_decap_8 FILLER_12_3026 ();
 sg13g2_decap_8 FILLER_12_3033 ();
 sg13g2_decap_8 FILLER_12_3040 ();
 sg13g2_decap_8 FILLER_12_3047 ();
 sg13g2_decap_8 FILLER_12_3054 ();
 sg13g2_decap_8 FILLER_12_3061 ();
 sg13g2_decap_8 FILLER_12_3068 ();
 sg13g2_decap_8 FILLER_12_3075 ();
 sg13g2_decap_8 FILLER_12_3082 ();
 sg13g2_decap_8 FILLER_12_3089 ();
 sg13g2_decap_8 FILLER_12_3096 ();
 sg13g2_decap_8 FILLER_12_3103 ();
 sg13g2_decap_8 FILLER_12_3110 ();
 sg13g2_decap_8 FILLER_12_3117 ();
 sg13g2_decap_8 FILLER_12_3124 ();
 sg13g2_decap_8 FILLER_12_3131 ();
 sg13g2_decap_8 FILLER_12_3138 ();
 sg13g2_decap_8 FILLER_12_3145 ();
 sg13g2_decap_8 FILLER_12_3152 ();
 sg13g2_decap_8 FILLER_12_3159 ();
 sg13g2_decap_8 FILLER_12_3166 ();
 sg13g2_decap_8 FILLER_12_3173 ();
 sg13g2_decap_8 FILLER_12_3180 ();
 sg13g2_decap_8 FILLER_12_3187 ();
 sg13g2_decap_8 FILLER_12_3194 ();
 sg13g2_decap_8 FILLER_12_3201 ();
 sg13g2_decap_8 FILLER_12_3208 ();
 sg13g2_decap_8 FILLER_12_3215 ();
 sg13g2_decap_8 FILLER_12_3222 ();
 sg13g2_decap_8 FILLER_12_3229 ();
 sg13g2_decap_8 FILLER_12_3236 ();
 sg13g2_decap_8 FILLER_12_3243 ();
 sg13g2_decap_8 FILLER_12_3250 ();
 sg13g2_decap_8 FILLER_12_3257 ();
 sg13g2_decap_8 FILLER_12_3264 ();
 sg13g2_decap_8 FILLER_12_3271 ();
 sg13g2_decap_8 FILLER_12_3278 ();
 sg13g2_decap_8 FILLER_12_3285 ();
 sg13g2_decap_8 FILLER_12_3292 ();
 sg13g2_decap_8 FILLER_12_3299 ();
 sg13g2_decap_8 FILLER_12_3306 ();
 sg13g2_decap_8 FILLER_12_3313 ();
 sg13g2_decap_8 FILLER_12_3320 ();
 sg13g2_decap_8 FILLER_12_3327 ();
 sg13g2_decap_8 FILLER_12_3334 ();
 sg13g2_decap_8 FILLER_12_3341 ();
 sg13g2_decap_8 FILLER_12_3348 ();
 sg13g2_decap_8 FILLER_12_3355 ();
 sg13g2_decap_8 FILLER_12_3362 ();
 sg13g2_decap_8 FILLER_12_3369 ();
 sg13g2_decap_8 FILLER_12_3376 ();
 sg13g2_decap_8 FILLER_12_3383 ();
 sg13g2_decap_8 FILLER_12_3390 ();
 sg13g2_decap_8 FILLER_12_3397 ();
 sg13g2_decap_8 FILLER_12_3404 ();
 sg13g2_decap_8 FILLER_12_3411 ();
 sg13g2_decap_8 FILLER_12_3418 ();
 sg13g2_decap_8 FILLER_12_3425 ();
 sg13g2_decap_8 FILLER_12_3432 ();
 sg13g2_decap_8 FILLER_12_3439 ();
 sg13g2_decap_8 FILLER_12_3446 ();
 sg13g2_decap_8 FILLER_12_3453 ();
 sg13g2_decap_8 FILLER_12_3460 ();
 sg13g2_decap_8 FILLER_12_3467 ();
 sg13g2_decap_8 FILLER_12_3474 ();
 sg13g2_decap_8 FILLER_12_3481 ();
 sg13g2_decap_8 FILLER_12_3488 ();
 sg13g2_decap_8 FILLER_12_3495 ();
 sg13g2_decap_8 FILLER_12_3502 ();
 sg13g2_decap_8 FILLER_12_3509 ();
 sg13g2_decap_8 FILLER_12_3516 ();
 sg13g2_decap_8 FILLER_12_3523 ();
 sg13g2_decap_8 FILLER_12_3530 ();
 sg13g2_decap_8 FILLER_12_3537 ();
 sg13g2_decap_8 FILLER_12_3544 ();
 sg13g2_decap_8 FILLER_12_3551 ();
 sg13g2_decap_8 FILLER_12_3558 ();
 sg13g2_decap_8 FILLER_12_3565 ();
 sg13g2_decap_8 FILLER_12_3572 ();
 sg13g2_fill_1 FILLER_12_3579 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_fill_2 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_4 FILLER_13_217 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_248 ();
 sg13g2_fill_1 FILLER_13_255 ();
 sg13g2_decap_8 FILLER_13_316 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_fill_1 FILLER_13_374 ();
 sg13g2_fill_2 FILLER_13_401 ();
 sg13g2_decap_8 FILLER_13_432 ();
 sg13g2_decap_8 FILLER_13_439 ();
 sg13g2_decap_8 FILLER_13_446 ();
 sg13g2_decap_8 FILLER_13_453 ();
 sg13g2_decap_8 FILLER_13_460 ();
 sg13g2_decap_8 FILLER_13_467 ();
 sg13g2_decap_8 FILLER_13_474 ();
 sg13g2_decap_8 FILLER_13_481 ();
 sg13g2_decap_8 FILLER_13_488 ();
 sg13g2_decap_8 FILLER_13_495 ();
 sg13g2_decap_8 FILLER_13_502 ();
 sg13g2_fill_1 FILLER_13_509 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_fill_2 FILLER_13_546 ();
 sg13g2_decap_4 FILLER_13_583 ();
 sg13g2_fill_1 FILLER_13_587 ();
 sg13g2_fill_2 FILLER_13_608 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_fill_2 FILLER_13_651 ();
 sg13g2_fill_2 FILLER_13_717 ();
 sg13g2_fill_1 FILLER_13_719 ();
 sg13g2_decap_4 FILLER_13_725 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_decap_4 FILLER_13_774 ();
 sg13g2_fill_1 FILLER_13_778 ();
 sg13g2_decap_8 FILLER_13_843 ();
 sg13g2_decap_8 FILLER_13_850 ();
 sg13g2_fill_2 FILLER_13_857 ();
 sg13g2_fill_1 FILLER_13_863 ();
 sg13g2_fill_1 FILLER_13_892 ();
 sg13g2_decap_4 FILLER_13_897 ();
 sg13g2_fill_1 FILLER_13_901 ();
 sg13g2_decap_8 FILLER_13_941 ();
 sg13g2_decap_4 FILLER_13_948 ();
 sg13g2_fill_2 FILLER_13_952 ();
 sg13g2_fill_1 FILLER_13_957 ();
 sg13g2_decap_8 FILLER_13_963 ();
 sg13g2_decap_4 FILLER_13_970 ();
 sg13g2_decap_4 FILLER_13_977 ();
 sg13g2_fill_1 FILLER_13_981 ();
 sg13g2_fill_1 FILLER_13_990 ();
 sg13g2_fill_1 FILLER_13_999 ();
 sg13g2_fill_2 FILLER_13_1057 ();
 sg13g2_decap_8 FILLER_13_1067 ();
 sg13g2_fill_1 FILLER_13_1074 ();
 sg13g2_decap_4 FILLER_13_1080 ();
 sg13g2_decap_8 FILLER_13_1188 ();
 sg13g2_fill_1 FILLER_13_1195 ();
 sg13g2_decap_8 FILLER_13_1222 ();
 sg13g2_decap_8 FILLER_13_1229 ();
 sg13g2_decap_8 FILLER_13_1236 ();
 sg13g2_decap_8 FILLER_13_1243 ();
 sg13g2_fill_2 FILLER_13_1250 ();
 sg13g2_fill_1 FILLER_13_1252 ();
 sg13g2_fill_2 FILLER_13_1287 ();
 sg13g2_fill_1 FILLER_13_1310 ();
 sg13g2_decap_8 FILLER_13_1337 ();
 sg13g2_decap_4 FILLER_13_1344 ();
 sg13g2_fill_2 FILLER_13_1348 ();
 sg13g2_decap_8 FILLER_13_1354 ();
 sg13g2_decap_4 FILLER_13_1361 ();
 sg13g2_fill_2 FILLER_13_1365 ();
 sg13g2_fill_2 FILLER_13_1393 ();
 sg13g2_fill_1 FILLER_13_1395 ();
 sg13g2_fill_2 FILLER_13_1435 ();
 sg13g2_decap_8 FILLER_13_1473 ();
 sg13g2_fill_2 FILLER_13_1480 ();
 sg13g2_fill_1 FILLER_13_1482 ();
 sg13g2_decap_8 FILLER_13_1517 ();
 sg13g2_decap_8 FILLER_13_1524 ();
 sg13g2_decap_4 FILLER_13_1531 ();
 sg13g2_fill_2 FILLER_13_1547 ();
 sg13g2_fill_1 FILLER_13_1575 ();
 sg13g2_fill_2 FILLER_13_1602 ();
 sg13g2_decap_8 FILLER_13_1625 ();
 sg13g2_fill_2 FILLER_13_1632 ();
 sg13g2_fill_1 FILLER_13_1634 ();
 sg13g2_decap_8 FILLER_13_1730 ();
 sg13g2_fill_1 FILLER_13_1750 ();
 sg13g2_decap_8 FILLER_13_1758 ();
 sg13g2_decap_8 FILLER_13_1765 ();
 sg13g2_decap_8 FILLER_13_1772 ();
 sg13g2_decap_8 FILLER_13_1805 ();
 sg13g2_decap_8 FILLER_13_1812 ();
 sg13g2_decap_8 FILLER_13_1819 ();
 sg13g2_fill_1 FILLER_13_1826 ();
 sg13g2_fill_1 FILLER_13_1913 ();
 sg13g2_fill_1 FILLER_13_1939 ();
 sg13g2_decap_4 FILLER_13_1977 ();
 sg13g2_fill_2 FILLER_13_1981 ();
 sg13g2_decap_8 FILLER_13_2098 ();
 sg13g2_decap_4 FILLER_13_2105 ();
 sg13g2_fill_2 FILLER_13_2109 ();
 sg13g2_decap_4 FILLER_13_2115 ();
 sg13g2_decap_8 FILLER_13_2145 ();
 sg13g2_fill_2 FILLER_13_2152 ();
 sg13g2_fill_1 FILLER_13_2154 ();
 sg13g2_decap_4 FILLER_13_2187 ();
 sg13g2_fill_1 FILLER_13_2191 ();
 sg13g2_fill_2 FILLER_13_2213 ();
 sg13g2_fill_1 FILLER_13_2267 ();
 sg13g2_decap_8 FILLER_13_2281 ();
 sg13g2_decap_8 FILLER_13_2288 ();
 sg13g2_fill_2 FILLER_13_2295 ();
 sg13g2_fill_1 FILLER_13_2297 ();
 sg13g2_decap_8 FILLER_13_2310 ();
 sg13g2_fill_2 FILLER_13_2317 ();
 sg13g2_fill_1 FILLER_13_2319 ();
 sg13g2_fill_1 FILLER_13_2324 ();
 sg13g2_fill_2 FILLER_13_2346 ();
 sg13g2_fill_2 FILLER_13_2356 ();
 sg13g2_fill_1 FILLER_13_2366 ();
 sg13g2_fill_1 FILLER_13_2447 ();
 sg13g2_decap_8 FILLER_13_2479 ();
 sg13g2_decap_8 FILLER_13_2486 ();
 sg13g2_fill_1 FILLER_13_2493 ();
 sg13g2_fill_2 FILLER_13_2498 ();
 sg13g2_fill_2 FILLER_13_2526 ();
 sg13g2_fill_2 FILLER_13_2549 ();
 sg13g2_decap_8 FILLER_13_2559 ();
 sg13g2_decap_8 FILLER_13_2566 ();
 sg13g2_fill_2 FILLER_13_2599 ();
 sg13g2_fill_1 FILLER_13_2601 ();
 sg13g2_decap_8 FILLER_13_2606 ();
 sg13g2_fill_1 FILLER_13_2634 ();
 sg13g2_decap_8 FILLER_13_2669 ();
 sg13g2_decap_8 FILLER_13_2676 ();
 sg13g2_decap_8 FILLER_13_2683 ();
 sg13g2_decap_8 FILLER_13_2690 ();
 sg13g2_decap_8 FILLER_13_2697 ();
 sg13g2_decap_8 FILLER_13_2704 ();
 sg13g2_decap_8 FILLER_13_2711 ();
 sg13g2_decap_8 FILLER_13_2718 ();
 sg13g2_decap_8 FILLER_13_2725 ();
 sg13g2_decap_8 FILLER_13_2732 ();
 sg13g2_decap_8 FILLER_13_2739 ();
 sg13g2_decap_8 FILLER_13_2746 ();
 sg13g2_decap_8 FILLER_13_2753 ();
 sg13g2_decap_8 FILLER_13_2760 ();
 sg13g2_decap_8 FILLER_13_2767 ();
 sg13g2_decap_8 FILLER_13_2774 ();
 sg13g2_decap_8 FILLER_13_2781 ();
 sg13g2_decap_8 FILLER_13_2788 ();
 sg13g2_decap_8 FILLER_13_2795 ();
 sg13g2_decap_8 FILLER_13_2802 ();
 sg13g2_decap_8 FILLER_13_2809 ();
 sg13g2_decap_8 FILLER_13_2816 ();
 sg13g2_decap_8 FILLER_13_2823 ();
 sg13g2_decap_8 FILLER_13_2830 ();
 sg13g2_decap_8 FILLER_13_2837 ();
 sg13g2_decap_8 FILLER_13_2844 ();
 sg13g2_decap_8 FILLER_13_2851 ();
 sg13g2_decap_8 FILLER_13_2858 ();
 sg13g2_decap_8 FILLER_13_2865 ();
 sg13g2_decap_8 FILLER_13_2872 ();
 sg13g2_decap_8 FILLER_13_2879 ();
 sg13g2_decap_8 FILLER_13_2886 ();
 sg13g2_decap_8 FILLER_13_2893 ();
 sg13g2_decap_8 FILLER_13_2900 ();
 sg13g2_decap_8 FILLER_13_2907 ();
 sg13g2_decap_8 FILLER_13_2914 ();
 sg13g2_decap_8 FILLER_13_2921 ();
 sg13g2_decap_8 FILLER_13_2928 ();
 sg13g2_decap_8 FILLER_13_2935 ();
 sg13g2_decap_8 FILLER_13_2942 ();
 sg13g2_decap_8 FILLER_13_2949 ();
 sg13g2_decap_8 FILLER_13_2956 ();
 sg13g2_decap_8 FILLER_13_2963 ();
 sg13g2_decap_8 FILLER_13_2970 ();
 sg13g2_decap_8 FILLER_13_2977 ();
 sg13g2_decap_8 FILLER_13_2984 ();
 sg13g2_decap_8 FILLER_13_2991 ();
 sg13g2_decap_8 FILLER_13_2998 ();
 sg13g2_decap_8 FILLER_13_3005 ();
 sg13g2_decap_8 FILLER_13_3012 ();
 sg13g2_decap_8 FILLER_13_3019 ();
 sg13g2_decap_8 FILLER_13_3026 ();
 sg13g2_decap_8 FILLER_13_3033 ();
 sg13g2_decap_8 FILLER_13_3040 ();
 sg13g2_decap_8 FILLER_13_3047 ();
 sg13g2_decap_8 FILLER_13_3054 ();
 sg13g2_decap_8 FILLER_13_3061 ();
 sg13g2_decap_8 FILLER_13_3068 ();
 sg13g2_decap_8 FILLER_13_3075 ();
 sg13g2_decap_8 FILLER_13_3082 ();
 sg13g2_decap_8 FILLER_13_3089 ();
 sg13g2_decap_8 FILLER_13_3096 ();
 sg13g2_decap_8 FILLER_13_3103 ();
 sg13g2_decap_8 FILLER_13_3110 ();
 sg13g2_decap_8 FILLER_13_3117 ();
 sg13g2_decap_8 FILLER_13_3124 ();
 sg13g2_decap_8 FILLER_13_3131 ();
 sg13g2_decap_8 FILLER_13_3138 ();
 sg13g2_decap_8 FILLER_13_3145 ();
 sg13g2_decap_8 FILLER_13_3152 ();
 sg13g2_decap_8 FILLER_13_3159 ();
 sg13g2_decap_8 FILLER_13_3166 ();
 sg13g2_decap_8 FILLER_13_3173 ();
 sg13g2_decap_8 FILLER_13_3180 ();
 sg13g2_decap_8 FILLER_13_3187 ();
 sg13g2_decap_8 FILLER_13_3194 ();
 sg13g2_decap_8 FILLER_13_3201 ();
 sg13g2_decap_8 FILLER_13_3208 ();
 sg13g2_decap_8 FILLER_13_3215 ();
 sg13g2_decap_8 FILLER_13_3222 ();
 sg13g2_decap_8 FILLER_13_3229 ();
 sg13g2_decap_8 FILLER_13_3236 ();
 sg13g2_decap_8 FILLER_13_3243 ();
 sg13g2_decap_8 FILLER_13_3250 ();
 sg13g2_decap_8 FILLER_13_3257 ();
 sg13g2_decap_8 FILLER_13_3264 ();
 sg13g2_decap_8 FILLER_13_3271 ();
 sg13g2_decap_8 FILLER_13_3278 ();
 sg13g2_decap_8 FILLER_13_3285 ();
 sg13g2_decap_8 FILLER_13_3292 ();
 sg13g2_decap_8 FILLER_13_3299 ();
 sg13g2_decap_8 FILLER_13_3306 ();
 sg13g2_decap_8 FILLER_13_3313 ();
 sg13g2_decap_8 FILLER_13_3320 ();
 sg13g2_decap_8 FILLER_13_3327 ();
 sg13g2_decap_8 FILLER_13_3334 ();
 sg13g2_decap_8 FILLER_13_3341 ();
 sg13g2_decap_8 FILLER_13_3348 ();
 sg13g2_decap_8 FILLER_13_3355 ();
 sg13g2_decap_8 FILLER_13_3362 ();
 sg13g2_decap_8 FILLER_13_3369 ();
 sg13g2_decap_8 FILLER_13_3376 ();
 sg13g2_decap_8 FILLER_13_3383 ();
 sg13g2_decap_8 FILLER_13_3390 ();
 sg13g2_decap_8 FILLER_13_3397 ();
 sg13g2_decap_8 FILLER_13_3404 ();
 sg13g2_decap_8 FILLER_13_3411 ();
 sg13g2_decap_8 FILLER_13_3418 ();
 sg13g2_decap_8 FILLER_13_3425 ();
 sg13g2_decap_8 FILLER_13_3432 ();
 sg13g2_decap_8 FILLER_13_3439 ();
 sg13g2_decap_8 FILLER_13_3446 ();
 sg13g2_decap_8 FILLER_13_3453 ();
 sg13g2_decap_8 FILLER_13_3460 ();
 sg13g2_decap_8 FILLER_13_3467 ();
 sg13g2_decap_8 FILLER_13_3474 ();
 sg13g2_decap_8 FILLER_13_3481 ();
 sg13g2_decap_8 FILLER_13_3488 ();
 sg13g2_decap_8 FILLER_13_3495 ();
 sg13g2_decap_8 FILLER_13_3502 ();
 sg13g2_decap_8 FILLER_13_3509 ();
 sg13g2_decap_8 FILLER_13_3516 ();
 sg13g2_decap_8 FILLER_13_3523 ();
 sg13g2_decap_8 FILLER_13_3530 ();
 sg13g2_decap_8 FILLER_13_3537 ();
 sg13g2_decap_8 FILLER_13_3544 ();
 sg13g2_decap_8 FILLER_13_3551 ();
 sg13g2_decap_8 FILLER_13_3558 ();
 sg13g2_decap_8 FILLER_13_3565 ();
 sg13g2_decap_8 FILLER_13_3572 ();
 sg13g2_fill_1 FILLER_13_3579 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_32 ();
 sg13g2_fill_1 FILLER_14_72 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_130 ();
 sg13g2_fill_2 FILLER_14_162 ();
 sg13g2_fill_1 FILLER_14_168 ();
 sg13g2_decap_4 FILLER_14_205 ();
 sg13g2_fill_1 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_236 ();
 sg13g2_decap_4 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_247 ();
 sg13g2_decap_4 FILLER_14_252 ();
 sg13g2_fill_2 FILLER_14_256 ();
 sg13g2_fill_1 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_4 FILLER_14_322 ();
 sg13g2_fill_1 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_551 ();
 sg13g2_fill_1 FILLER_14_558 ();
 sg13g2_fill_2 FILLER_14_573 ();
 sg13g2_fill_1 FILLER_14_575 ();
 sg13g2_decap_8 FILLER_14_583 ();
 sg13g2_decap_8 FILLER_14_590 ();
 sg13g2_fill_2 FILLER_14_597 ();
 sg13g2_fill_2 FILLER_14_612 ();
 sg13g2_decap_8 FILLER_14_737 ();
 sg13g2_decap_4 FILLER_14_744 ();
 sg13g2_fill_1 FILLER_14_815 ();
 sg13g2_decap_4 FILLER_14_820 ();
 sg13g2_fill_1 FILLER_14_824 ();
 sg13g2_fill_2 FILLER_14_841 ();
 sg13g2_fill_1 FILLER_14_843 ();
 sg13g2_decap_4 FILLER_14_870 ();
 sg13g2_fill_2 FILLER_14_874 ();
 sg13g2_fill_2 FILLER_14_902 ();
 sg13g2_fill_1 FILLER_14_904 ();
 sg13g2_fill_2 FILLER_14_935 ();
 sg13g2_fill_1 FILLER_14_948 ();
 sg13g2_decap_4 FILLER_14_980 ();
 sg13g2_fill_1 FILLER_14_984 ();
 sg13g2_fill_1 FILLER_14_989 ();
 sg13g2_decap_4 FILLER_14_995 ();
 sg13g2_fill_2 FILLER_14_999 ();
 sg13g2_decap_4 FILLER_14_1009 ();
 sg13g2_fill_2 FILLER_14_1021 ();
 sg13g2_fill_1 FILLER_14_1023 ();
 sg13g2_fill_2 FILLER_14_1045 ();
 sg13g2_fill_1 FILLER_14_1047 ();
 sg13g2_decap_8 FILLER_14_1082 ();
 sg13g2_decap_4 FILLER_14_1115 ();
 sg13g2_fill_2 FILLER_14_1148 ();
 sg13g2_fill_2 FILLER_14_1183 ();
 sg13g2_fill_2 FILLER_14_1192 ();
 sg13g2_decap_4 FILLER_14_1227 ();
 sg13g2_fill_2 FILLER_14_1231 ();
 sg13g2_decap_8 FILLER_14_1238 ();
 sg13g2_decap_8 FILLER_14_1245 ();
 sg13g2_decap_4 FILLER_14_1252 ();
 sg13g2_fill_1 FILLER_14_1256 ();
 sg13g2_fill_1 FILLER_14_1288 ();
 sg13g2_fill_2 FILLER_14_1343 ();
 sg13g2_fill_1 FILLER_14_1345 ();
 sg13g2_fill_1 FILLER_14_1367 ();
 sg13g2_fill_1 FILLER_14_1397 ();
 sg13g2_decap_4 FILLER_14_1405 ();
 sg13g2_fill_2 FILLER_14_1417 ();
 sg13g2_fill_2 FILLER_14_1424 ();
 sg13g2_decap_8 FILLER_14_1478 ();
 sg13g2_fill_2 FILLER_14_1485 ();
 sg13g2_fill_1 FILLER_14_1487 ();
 sg13g2_fill_2 FILLER_14_1493 ();
 sg13g2_decap_4 FILLER_14_1521 ();
 sg13g2_fill_2 FILLER_14_1538 ();
 sg13g2_decap_8 FILLER_14_1548 ();
 sg13g2_fill_2 FILLER_14_1585 ();
 sg13g2_fill_1 FILLER_14_1621 ();
 sg13g2_decap_4 FILLER_14_1630 ();
 sg13g2_decap_4 FILLER_14_1660 ();
 sg13g2_fill_1 FILLER_14_1690 ();
 sg13g2_fill_1 FILLER_14_1694 ();
 sg13g2_fill_2 FILLER_14_1699 ();
 sg13g2_fill_1 FILLER_14_1701 ();
 sg13g2_fill_1 FILLER_14_1715 ();
 sg13g2_decap_4 FILLER_14_1732 ();
 sg13g2_decap_4 FILLER_14_1757 ();
 sg13g2_decap_8 FILLER_14_1787 ();
 sg13g2_decap_8 FILLER_14_1794 ();
 sg13g2_decap_8 FILLER_14_1801 ();
 sg13g2_decap_4 FILLER_14_1808 ();
 sg13g2_fill_1 FILLER_14_1812 ();
 sg13g2_fill_1 FILLER_14_1852 ();
 sg13g2_fill_2 FILLER_14_1878 ();
 sg13g2_fill_1 FILLER_14_1880 ();
 sg13g2_decap_8 FILLER_14_1904 ();
 sg13g2_decap_8 FILLER_14_1911 ();
 sg13g2_fill_2 FILLER_14_1918 ();
 sg13g2_fill_1 FILLER_14_1923 ();
 sg13g2_fill_2 FILLER_14_1937 ();
 sg13g2_decap_8 FILLER_14_1967 ();
 sg13g2_decap_8 FILLER_14_1974 ();
 sg13g2_decap_8 FILLER_14_1981 ();
 sg13g2_decap_4 FILLER_14_1988 ();
 sg13g2_fill_2 FILLER_14_1992 ();
 sg13g2_decap_8 FILLER_14_2041 ();
 sg13g2_decap_8 FILLER_14_2048 ();
 sg13g2_fill_2 FILLER_14_2055 ();
 sg13g2_fill_1 FILLER_14_2057 ();
 sg13g2_decap_8 FILLER_14_2075 ();
 sg13g2_decap_8 FILLER_14_2090 ();
 sg13g2_decap_8 FILLER_14_2097 ();
 sg13g2_decap_4 FILLER_14_2104 ();
 sg13g2_decap_8 FILLER_14_2113 ();
 sg13g2_fill_2 FILLER_14_2120 ();
 sg13g2_fill_1 FILLER_14_2122 ();
 sg13g2_decap_8 FILLER_14_2138 ();
 sg13g2_decap_8 FILLER_14_2145 ();
 sg13g2_decap_8 FILLER_14_2152 ();
 sg13g2_decap_8 FILLER_14_2159 ();
 sg13g2_fill_1 FILLER_14_2166 ();
 sg13g2_fill_2 FILLER_14_2176 ();
 sg13g2_decap_8 FILLER_14_2212 ();
 sg13g2_decap_8 FILLER_14_2219 ();
 sg13g2_decap_4 FILLER_14_2230 ();
 sg13g2_fill_1 FILLER_14_2253 ();
 sg13g2_decap_8 FILLER_14_2279 ();
 sg13g2_fill_2 FILLER_14_2286 ();
 sg13g2_fill_1 FILLER_14_2288 ();
 sg13g2_decap_4 FILLER_14_2402 ();
 sg13g2_fill_2 FILLER_14_2406 ();
 sg13g2_decap_4 FILLER_14_2411 ();
 sg13g2_fill_2 FILLER_14_2422 ();
 sg13g2_fill_2 FILLER_14_2464 ();
 sg13g2_fill_1 FILLER_14_2466 ();
 sg13g2_decap_8 FILLER_14_2475 ();
 sg13g2_fill_2 FILLER_14_2482 ();
 sg13g2_fill_2 FILLER_14_2562 ();
 sg13g2_fill_1 FILLER_14_2564 ();
 sg13g2_fill_1 FILLER_14_2569 ();
 sg13g2_decap_4 FILLER_14_2664 ();
 sg13g2_fill_1 FILLER_14_2668 ();
 sg13g2_decap_8 FILLER_14_2695 ();
 sg13g2_decap_8 FILLER_14_2702 ();
 sg13g2_decap_8 FILLER_14_2709 ();
 sg13g2_decap_8 FILLER_14_2716 ();
 sg13g2_decap_8 FILLER_14_2723 ();
 sg13g2_decap_8 FILLER_14_2730 ();
 sg13g2_decap_8 FILLER_14_2737 ();
 sg13g2_decap_8 FILLER_14_2744 ();
 sg13g2_decap_8 FILLER_14_2751 ();
 sg13g2_decap_8 FILLER_14_2758 ();
 sg13g2_decap_8 FILLER_14_2765 ();
 sg13g2_decap_8 FILLER_14_2772 ();
 sg13g2_decap_8 FILLER_14_2779 ();
 sg13g2_decap_8 FILLER_14_2786 ();
 sg13g2_decap_8 FILLER_14_2793 ();
 sg13g2_decap_8 FILLER_14_2800 ();
 sg13g2_decap_8 FILLER_14_2807 ();
 sg13g2_decap_8 FILLER_14_2814 ();
 sg13g2_decap_8 FILLER_14_2821 ();
 sg13g2_decap_8 FILLER_14_2828 ();
 sg13g2_decap_8 FILLER_14_2835 ();
 sg13g2_decap_8 FILLER_14_2842 ();
 sg13g2_decap_8 FILLER_14_2849 ();
 sg13g2_decap_8 FILLER_14_2856 ();
 sg13g2_decap_8 FILLER_14_2863 ();
 sg13g2_decap_8 FILLER_14_2870 ();
 sg13g2_decap_8 FILLER_14_2877 ();
 sg13g2_decap_8 FILLER_14_2884 ();
 sg13g2_decap_8 FILLER_14_2891 ();
 sg13g2_decap_8 FILLER_14_2898 ();
 sg13g2_decap_8 FILLER_14_2905 ();
 sg13g2_decap_8 FILLER_14_2912 ();
 sg13g2_decap_8 FILLER_14_2919 ();
 sg13g2_decap_8 FILLER_14_2926 ();
 sg13g2_decap_8 FILLER_14_2933 ();
 sg13g2_decap_8 FILLER_14_2940 ();
 sg13g2_decap_8 FILLER_14_2947 ();
 sg13g2_decap_8 FILLER_14_2954 ();
 sg13g2_decap_8 FILLER_14_2961 ();
 sg13g2_decap_8 FILLER_14_2968 ();
 sg13g2_decap_8 FILLER_14_2975 ();
 sg13g2_decap_8 FILLER_14_2982 ();
 sg13g2_decap_8 FILLER_14_2989 ();
 sg13g2_decap_8 FILLER_14_2996 ();
 sg13g2_decap_8 FILLER_14_3003 ();
 sg13g2_decap_8 FILLER_14_3010 ();
 sg13g2_decap_8 FILLER_14_3017 ();
 sg13g2_decap_8 FILLER_14_3024 ();
 sg13g2_decap_8 FILLER_14_3031 ();
 sg13g2_decap_8 FILLER_14_3038 ();
 sg13g2_decap_8 FILLER_14_3045 ();
 sg13g2_decap_8 FILLER_14_3052 ();
 sg13g2_decap_8 FILLER_14_3059 ();
 sg13g2_decap_8 FILLER_14_3066 ();
 sg13g2_decap_8 FILLER_14_3073 ();
 sg13g2_decap_8 FILLER_14_3080 ();
 sg13g2_decap_8 FILLER_14_3087 ();
 sg13g2_decap_8 FILLER_14_3094 ();
 sg13g2_decap_8 FILLER_14_3101 ();
 sg13g2_decap_8 FILLER_14_3108 ();
 sg13g2_decap_8 FILLER_14_3115 ();
 sg13g2_decap_8 FILLER_14_3122 ();
 sg13g2_decap_8 FILLER_14_3129 ();
 sg13g2_decap_8 FILLER_14_3136 ();
 sg13g2_decap_8 FILLER_14_3143 ();
 sg13g2_decap_8 FILLER_14_3150 ();
 sg13g2_decap_8 FILLER_14_3157 ();
 sg13g2_decap_8 FILLER_14_3164 ();
 sg13g2_decap_8 FILLER_14_3171 ();
 sg13g2_decap_8 FILLER_14_3178 ();
 sg13g2_decap_8 FILLER_14_3185 ();
 sg13g2_decap_8 FILLER_14_3192 ();
 sg13g2_decap_8 FILLER_14_3199 ();
 sg13g2_decap_8 FILLER_14_3206 ();
 sg13g2_decap_8 FILLER_14_3213 ();
 sg13g2_decap_8 FILLER_14_3220 ();
 sg13g2_decap_8 FILLER_14_3227 ();
 sg13g2_decap_8 FILLER_14_3234 ();
 sg13g2_decap_8 FILLER_14_3241 ();
 sg13g2_decap_8 FILLER_14_3248 ();
 sg13g2_decap_8 FILLER_14_3255 ();
 sg13g2_decap_8 FILLER_14_3262 ();
 sg13g2_decap_8 FILLER_14_3269 ();
 sg13g2_decap_8 FILLER_14_3276 ();
 sg13g2_decap_8 FILLER_14_3283 ();
 sg13g2_decap_8 FILLER_14_3290 ();
 sg13g2_decap_8 FILLER_14_3297 ();
 sg13g2_decap_8 FILLER_14_3304 ();
 sg13g2_decap_8 FILLER_14_3311 ();
 sg13g2_decap_8 FILLER_14_3318 ();
 sg13g2_decap_8 FILLER_14_3325 ();
 sg13g2_decap_8 FILLER_14_3332 ();
 sg13g2_decap_8 FILLER_14_3339 ();
 sg13g2_decap_8 FILLER_14_3346 ();
 sg13g2_decap_8 FILLER_14_3353 ();
 sg13g2_decap_8 FILLER_14_3360 ();
 sg13g2_decap_8 FILLER_14_3367 ();
 sg13g2_decap_8 FILLER_14_3374 ();
 sg13g2_decap_8 FILLER_14_3381 ();
 sg13g2_decap_8 FILLER_14_3388 ();
 sg13g2_decap_8 FILLER_14_3395 ();
 sg13g2_decap_8 FILLER_14_3402 ();
 sg13g2_decap_8 FILLER_14_3409 ();
 sg13g2_decap_8 FILLER_14_3416 ();
 sg13g2_decap_8 FILLER_14_3423 ();
 sg13g2_decap_8 FILLER_14_3430 ();
 sg13g2_decap_8 FILLER_14_3437 ();
 sg13g2_decap_8 FILLER_14_3444 ();
 sg13g2_decap_8 FILLER_14_3451 ();
 sg13g2_decap_8 FILLER_14_3458 ();
 sg13g2_decap_8 FILLER_14_3465 ();
 sg13g2_decap_8 FILLER_14_3472 ();
 sg13g2_decap_8 FILLER_14_3479 ();
 sg13g2_decap_8 FILLER_14_3486 ();
 sg13g2_decap_8 FILLER_14_3493 ();
 sg13g2_decap_8 FILLER_14_3500 ();
 sg13g2_decap_8 FILLER_14_3507 ();
 sg13g2_decap_8 FILLER_14_3514 ();
 sg13g2_decap_8 FILLER_14_3521 ();
 sg13g2_decap_8 FILLER_14_3528 ();
 sg13g2_decap_8 FILLER_14_3535 ();
 sg13g2_decap_8 FILLER_14_3542 ();
 sg13g2_decap_8 FILLER_14_3549 ();
 sg13g2_decap_8 FILLER_14_3556 ();
 sg13g2_decap_8 FILLER_14_3563 ();
 sg13g2_decap_8 FILLER_14_3570 ();
 sg13g2_fill_2 FILLER_14_3577 ();
 sg13g2_fill_1 FILLER_14_3579 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_73 ();
 sg13g2_decap_8 FILLER_15_80 ();
 sg13g2_decap_8 FILLER_15_129 ();
 sg13g2_fill_1 FILLER_15_136 ();
 sg13g2_fill_2 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_200 ();
 sg13g2_fill_1 FILLER_15_202 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_decap_4 FILLER_15_298 ();
 sg13g2_fill_2 FILLER_15_302 ();
 sg13g2_decap_4 FILLER_15_320 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_432 ();
 sg13g2_decap_8 FILLER_15_439 ();
 sg13g2_decap_8 FILLER_15_446 ();
 sg13g2_decap_8 FILLER_15_453 ();
 sg13g2_decap_8 FILLER_15_460 ();
 sg13g2_decap_8 FILLER_15_467 ();
 sg13g2_decap_8 FILLER_15_474 ();
 sg13g2_decap_8 FILLER_15_481 ();
 sg13g2_decap_4 FILLER_15_488 ();
 sg13g2_decap_4 FILLER_15_557 ();
 sg13g2_fill_1 FILLER_15_561 ();
 sg13g2_fill_1 FILLER_15_570 ();
 sg13g2_decap_8 FILLER_15_579 ();
 sg13g2_decap_8 FILLER_15_586 ();
 sg13g2_decap_8 FILLER_15_593 ();
 sg13g2_decap_8 FILLER_15_600 ();
 sg13g2_decap_8 FILLER_15_607 ();
 sg13g2_decap_4 FILLER_15_614 ();
 sg13g2_fill_1 FILLER_15_618 ();
 sg13g2_fill_1 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_643 ();
 sg13g2_decap_8 FILLER_15_650 ();
 sg13g2_fill_1 FILLER_15_670 ();
 sg13g2_decap_8 FILLER_15_684 ();
 sg13g2_decap_4 FILLER_15_691 ();
 sg13g2_fill_2 FILLER_15_695 ();
 sg13g2_fill_2 FILLER_15_702 ();
 sg13g2_fill_1 FILLER_15_704 ();
 sg13g2_decap_8 FILLER_15_713 ();
 sg13g2_decap_8 FILLER_15_720 ();
 sg13g2_decap_8 FILLER_15_727 ();
 sg13g2_decap_4 FILLER_15_734 ();
 sg13g2_fill_1 FILLER_15_738 ();
 sg13g2_fill_1 FILLER_15_804 ();
 sg13g2_decap_8 FILLER_15_821 ();
 sg13g2_decap_8 FILLER_15_828 ();
 sg13g2_decap_8 FILLER_15_835 ();
 sg13g2_decap_8 FILLER_15_880 ();
 sg13g2_decap_8 FILLER_15_891 ();
 sg13g2_decap_8 FILLER_15_898 ();
 sg13g2_decap_8 FILLER_15_905 ();
 sg13g2_decap_8 FILLER_15_912 ();
 sg13g2_decap_4 FILLER_15_919 ();
 sg13g2_fill_2 FILLER_15_978 ();
 sg13g2_decap_8 FILLER_15_1006 ();
 sg13g2_decap_8 FILLER_15_1013 ();
 sg13g2_fill_2 FILLER_15_1020 ();
 sg13g2_decap_8 FILLER_15_1053 ();
 sg13g2_decap_8 FILLER_15_1060 ();
 sg13g2_fill_2 FILLER_15_1097 ();
 sg13g2_fill_1 FILLER_15_1099 ();
 sg13g2_decap_8 FILLER_15_1108 ();
 sg13g2_decap_8 FILLER_15_1115 ();
 sg13g2_decap_8 FILLER_15_1122 ();
 sg13g2_decap_8 FILLER_15_1171 ();
 sg13g2_decap_8 FILLER_15_1178 ();
 sg13g2_decap_8 FILLER_15_1185 ();
 sg13g2_decap_8 FILLER_15_1192 ();
 sg13g2_fill_2 FILLER_15_1199 ();
 sg13g2_fill_1 FILLER_15_1201 ();
 sg13g2_fill_2 FILLER_15_1234 ();
 sg13g2_fill_1 FILLER_15_1236 ();
 sg13g2_decap_8 FILLER_15_1241 ();
 sg13g2_decap_8 FILLER_15_1248 ();
 sg13g2_fill_1 FILLER_15_1255 ();
 sg13g2_fill_2 FILLER_15_1290 ();
 sg13g2_fill_1 FILLER_15_1292 ();
 sg13g2_decap_4 FILLER_15_1301 ();
 sg13g2_fill_2 FILLER_15_1305 ();
 sg13g2_fill_1 FILLER_15_1341 ();
 sg13g2_fill_2 FILLER_15_1368 ();
 sg13g2_fill_1 FILLER_15_1370 ();
 sg13g2_decap_8 FILLER_15_1394 ();
 sg13g2_decap_8 FILLER_15_1401 ();
 sg13g2_decap_8 FILLER_15_1408 ();
 sg13g2_decap_8 FILLER_15_1415 ();
 sg13g2_decap_4 FILLER_15_1422 ();
 sg13g2_fill_1 FILLER_15_1426 ();
 sg13g2_decap_8 FILLER_15_1465 ();
 sg13g2_decap_8 FILLER_15_1472 ();
 sg13g2_decap_8 FILLER_15_1479 ();
 sg13g2_fill_1 FILLER_15_1486 ();
 sg13g2_decap_8 FILLER_15_1497 ();
 sg13g2_decap_8 FILLER_15_1504 ();
 sg13g2_decap_8 FILLER_15_1511 ();
 sg13g2_fill_1 FILLER_15_1518 ();
 sg13g2_fill_2 FILLER_15_1548 ();
 sg13g2_fill_1 FILLER_15_1554 ();
 sg13g2_decap_8 FILLER_15_1559 ();
 sg13g2_decap_4 FILLER_15_1566 ();
 sg13g2_fill_2 FILLER_15_1574 ();
 sg13g2_fill_2 FILLER_15_1584 ();
 sg13g2_fill_1 FILLER_15_1586 ();
 sg13g2_fill_2 FILLER_15_1591 ();
 sg13g2_fill_1 FILLER_15_1593 ();
 sg13g2_decap_4 FILLER_15_1603 ();
 sg13g2_decap_4 FILLER_15_1622 ();
 sg13g2_fill_1 FILLER_15_1626 ();
 sg13g2_decap_8 FILLER_15_1632 ();
 sg13g2_decap_4 FILLER_15_1639 ();
 sg13g2_fill_2 FILLER_15_1643 ();
 sg13g2_decap_8 FILLER_15_1649 ();
 sg13g2_decap_4 FILLER_15_1656 ();
 sg13g2_decap_8 FILLER_15_1665 ();
 sg13g2_fill_2 FILLER_15_1672 ();
 sg13g2_fill_1 FILLER_15_1682 ();
 sg13g2_decap_8 FILLER_15_1765 ();
 sg13g2_fill_2 FILLER_15_1772 ();
 sg13g2_fill_1 FILLER_15_1774 ();
 sg13g2_decap_4 FILLER_15_1809 ();
 sg13g2_fill_1 FILLER_15_1813 ();
 sg13g2_fill_2 FILLER_15_1839 ();
 sg13g2_fill_2 FILLER_15_1844 ();
 sg13g2_fill_2 FILLER_15_1859 ();
 sg13g2_fill_1 FILLER_15_1861 ();
 sg13g2_decap_8 FILLER_15_1870 ();
 sg13g2_fill_2 FILLER_15_1877 ();
 sg13g2_fill_1 FILLER_15_1879 ();
 sg13g2_decap_8 FILLER_15_1885 ();
 sg13g2_decap_8 FILLER_15_1892 ();
 sg13g2_decap_8 FILLER_15_1899 ();
 sg13g2_decap_8 FILLER_15_1906 ();
 sg13g2_decap_8 FILLER_15_1913 ();
 sg13g2_decap_8 FILLER_15_1920 ();
 sg13g2_decap_8 FILLER_15_1927 ();
 sg13g2_fill_1 FILLER_15_1960 ();
 sg13g2_decap_8 FILLER_15_1969 ();
 sg13g2_decap_8 FILLER_15_1976 ();
 sg13g2_decap_8 FILLER_15_1983 ();
 sg13g2_decap_8 FILLER_15_1990 ();
 sg13g2_decap_8 FILLER_15_1997 ();
 sg13g2_fill_1 FILLER_15_2004 ();
 sg13g2_fill_2 FILLER_15_2018 ();
 sg13g2_decap_8 FILLER_15_2036 ();
 sg13g2_decap_8 FILLER_15_2043 ();
 sg13g2_decap_4 FILLER_15_2050 ();
 sg13g2_fill_1 FILLER_15_2054 ();
 sg13g2_decap_8 FILLER_15_2081 ();
 sg13g2_fill_1 FILLER_15_2122 ();
 sg13g2_fill_2 FILLER_15_2149 ();
 sg13g2_decap_8 FILLER_15_2156 ();
 sg13g2_decap_8 FILLER_15_2163 ();
 sg13g2_fill_2 FILLER_15_2170 ();
 sg13g2_fill_1 FILLER_15_2172 ();
 sg13g2_decap_4 FILLER_15_2230 ();
 sg13g2_fill_2 FILLER_15_2234 ();
 sg13g2_fill_2 FILLER_15_2239 ();
 sg13g2_fill_1 FILLER_15_2241 ();
 sg13g2_fill_2 FILLER_15_2247 ();
 sg13g2_fill_2 FILLER_15_2253 ();
 sg13g2_fill_1 FILLER_15_2255 ();
 sg13g2_decap_8 FILLER_15_2259 ();
 sg13g2_fill_1 FILLER_15_2266 ();
 sg13g2_decap_4 FILLER_15_2275 ();
 sg13g2_fill_2 FILLER_15_2279 ();
 sg13g2_decap_8 FILLER_15_2285 ();
 sg13g2_fill_1 FILLER_15_2292 ();
 sg13g2_fill_2 FILLER_15_2307 ();
 sg13g2_decap_4 FILLER_15_2366 ();
 sg13g2_decap_8 FILLER_15_2396 ();
 sg13g2_decap_8 FILLER_15_2403 ();
 sg13g2_fill_2 FILLER_15_2410 ();
 sg13g2_decap_8 FILLER_15_2441 ();
 sg13g2_fill_2 FILLER_15_2448 ();
 sg13g2_decap_8 FILLER_15_2455 ();
 sg13g2_decap_8 FILLER_15_2462 ();
 sg13g2_decap_8 FILLER_15_2469 ();
 sg13g2_decap_8 FILLER_15_2476 ();
 sg13g2_decap_8 FILLER_15_2483 ();
 sg13g2_fill_1 FILLER_15_2490 ();
 sg13g2_fill_2 FILLER_15_2517 ();
 sg13g2_fill_1 FILLER_15_2519 ();
 sg13g2_decap_4 FILLER_15_2524 ();
 sg13g2_fill_2 FILLER_15_2528 ();
 sg13g2_decap_4 FILLER_15_2655 ();
 sg13g2_fill_1 FILLER_15_2659 ();
 sg13g2_decap_4 FILLER_15_2664 ();
 sg13g2_decap_8 FILLER_15_2694 ();
 sg13g2_decap_8 FILLER_15_2701 ();
 sg13g2_decap_8 FILLER_15_2708 ();
 sg13g2_decap_8 FILLER_15_2715 ();
 sg13g2_decap_8 FILLER_15_2722 ();
 sg13g2_decap_8 FILLER_15_2729 ();
 sg13g2_decap_8 FILLER_15_2736 ();
 sg13g2_decap_8 FILLER_15_2743 ();
 sg13g2_decap_8 FILLER_15_2750 ();
 sg13g2_decap_8 FILLER_15_2757 ();
 sg13g2_decap_8 FILLER_15_2764 ();
 sg13g2_decap_8 FILLER_15_2771 ();
 sg13g2_decap_8 FILLER_15_2778 ();
 sg13g2_decap_8 FILLER_15_2785 ();
 sg13g2_decap_8 FILLER_15_2792 ();
 sg13g2_decap_8 FILLER_15_2799 ();
 sg13g2_decap_8 FILLER_15_2806 ();
 sg13g2_decap_8 FILLER_15_2813 ();
 sg13g2_decap_8 FILLER_15_2820 ();
 sg13g2_decap_8 FILLER_15_2827 ();
 sg13g2_decap_8 FILLER_15_2834 ();
 sg13g2_decap_8 FILLER_15_2841 ();
 sg13g2_decap_8 FILLER_15_2848 ();
 sg13g2_decap_8 FILLER_15_2855 ();
 sg13g2_decap_8 FILLER_15_2862 ();
 sg13g2_decap_8 FILLER_15_2869 ();
 sg13g2_decap_8 FILLER_15_2876 ();
 sg13g2_decap_8 FILLER_15_2883 ();
 sg13g2_decap_8 FILLER_15_2890 ();
 sg13g2_decap_8 FILLER_15_2897 ();
 sg13g2_decap_8 FILLER_15_2904 ();
 sg13g2_decap_8 FILLER_15_2911 ();
 sg13g2_decap_8 FILLER_15_2918 ();
 sg13g2_decap_8 FILLER_15_2925 ();
 sg13g2_decap_8 FILLER_15_2932 ();
 sg13g2_decap_8 FILLER_15_2939 ();
 sg13g2_decap_8 FILLER_15_2946 ();
 sg13g2_decap_8 FILLER_15_2953 ();
 sg13g2_decap_8 FILLER_15_2960 ();
 sg13g2_decap_8 FILLER_15_2967 ();
 sg13g2_decap_8 FILLER_15_2974 ();
 sg13g2_decap_8 FILLER_15_2981 ();
 sg13g2_decap_8 FILLER_15_2988 ();
 sg13g2_decap_8 FILLER_15_2995 ();
 sg13g2_decap_8 FILLER_15_3002 ();
 sg13g2_decap_8 FILLER_15_3009 ();
 sg13g2_decap_8 FILLER_15_3016 ();
 sg13g2_decap_8 FILLER_15_3023 ();
 sg13g2_decap_8 FILLER_15_3030 ();
 sg13g2_decap_8 FILLER_15_3037 ();
 sg13g2_decap_8 FILLER_15_3044 ();
 sg13g2_decap_8 FILLER_15_3051 ();
 sg13g2_decap_8 FILLER_15_3058 ();
 sg13g2_decap_8 FILLER_15_3065 ();
 sg13g2_decap_8 FILLER_15_3072 ();
 sg13g2_decap_8 FILLER_15_3079 ();
 sg13g2_decap_8 FILLER_15_3086 ();
 sg13g2_decap_8 FILLER_15_3093 ();
 sg13g2_decap_8 FILLER_15_3100 ();
 sg13g2_decap_8 FILLER_15_3107 ();
 sg13g2_decap_8 FILLER_15_3114 ();
 sg13g2_decap_8 FILLER_15_3121 ();
 sg13g2_decap_8 FILLER_15_3128 ();
 sg13g2_decap_8 FILLER_15_3135 ();
 sg13g2_decap_8 FILLER_15_3142 ();
 sg13g2_decap_8 FILLER_15_3149 ();
 sg13g2_decap_8 FILLER_15_3156 ();
 sg13g2_decap_8 FILLER_15_3163 ();
 sg13g2_decap_8 FILLER_15_3170 ();
 sg13g2_decap_8 FILLER_15_3177 ();
 sg13g2_decap_8 FILLER_15_3184 ();
 sg13g2_decap_8 FILLER_15_3191 ();
 sg13g2_decap_8 FILLER_15_3198 ();
 sg13g2_decap_8 FILLER_15_3205 ();
 sg13g2_decap_8 FILLER_15_3212 ();
 sg13g2_decap_8 FILLER_15_3219 ();
 sg13g2_decap_8 FILLER_15_3226 ();
 sg13g2_decap_8 FILLER_15_3233 ();
 sg13g2_decap_8 FILLER_15_3240 ();
 sg13g2_decap_8 FILLER_15_3247 ();
 sg13g2_decap_8 FILLER_15_3254 ();
 sg13g2_decap_8 FILLER_15_3261 ();
 sg13g2_decap_8 FILLER_15_3268 ();
 sg13g2_decap_8 FILLER_15_3275 ();
 sg13g2_decap_8 FILLER_15_3282 ();
 sg13g2_decap_8 FILLER_15_3289 ();
 sg13g2_decap_8 FILLER_15_3296 ();
 sg13g2_decap_8 FILLER_15_3303 ();
 sg13g2_decap_8 FILLER_15_3310 ();
 sg13g2_decap_8 FILLER_15_3317 ();
 sg13g2_decap_8 FILLER_15_3324 ();
 sg13g2_decap_8 FILLER_15_3331 ();
 sg13g2_decap_8 FILLER_15_3338 ();
 sg13g2_decap_8 FILLER_15_3345 ();
 sg13g2_decap_8 FILLER_15_3352 ();
 sg13g2_decap_8 FILLER_15_3359 ();
 sg13g2_decap_8 FILLER_15_3366 ();
 sg13g2_decap_8 FILLER_15_3373 ();
 sg13g2_decap_8 FILLER_15_3380 ();
 sg13g2_decap_8 FILLER_15_3387 ();
 sg13g2_decap_8 FILLER_15_3394 ();
 sg13g2_decap_8 FILLER_15_3401 ();
 sg13g2_decap_8 FILLER_15_3408 ();
 sg13g2_decap_8 FILLER_15_3415 ();
 sg13g2_decap_8 FILLER_15_3422 ();
 sg13g2_decap_8 FILLER_15_3429 ();
 sg13g2_decap_8 FILLER_15_3436 ();
 sg13g2_decap_8 FILLER_15_3443 ();
 sg13g2_decap_8 FILLER_15_3450 ();
 sg13g2_decap_8 FILLER_15_3457 ();
 sg13g2_decap_8 FILLER_15_3464 ();
 sg13g2_decap_8 FILLER_15_3471 ();
 sg13g2_decap_8 FILLER_15_3478 ();
 sg13g2_decap_8 FILLER_15_3485 ();
 sg13g2_decap_8 FILLER_15_3492 ();
 sg13g2_decap_8 FILLER_15_3499 ();
 sg13g2_decap_8 FILLER_15_3506 ();
 sg13g2_decap_8 FILLER_15_3513 ();
 sg13g2_decap_8 FILLER_15_3520 ();
 sg13g2_decap_8 FILLER_15_3527 ();
 sg13g2_decap_8 FILLER_15_3534 ();
 sg13g2_decap_8 FILLER_15_3541 ();
 sg13g2_decap_8 FILLER_15_3548 ();
 sg13g2_decap_8 FILLER_15_3555 ();
 sg13g2_decap_8 FILLER_15_3562 ();
 sg13g2_decap_8 FILLER_15_3569 ();
 sg13g2_decap_4 FILLER_15_3576 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_52 ();
 sg13g2_fill_1 FILLER_16_54 ();
 sg13g2_decap_8 FILLER_16_65 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_decap_8 FILLER_16_79 ();
 sg13g2_decap_8 FILLER_16_129 ();
 sg13g2_decap_8 FILLER_16_136 ();
 sg13g2_decap_8 FILLER_16_143 ();
 sg13g2_decap_8 FILLER_16_150 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_fill_2 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_fill_2 FILLER_16_231 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_decap_4 FILLER_16_278 ();
 sg13g2_fill_2 FILLER_16_292 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_fill_2 FILLER_16_312 ();
 sg13g2_fill_1 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_fill_1 FILLER_16_348 ();
 sg13g2_decap_4 FILLER_16_390 ();
 sg13g2_fill_1 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_16_435 ();
 sg13g2_decap_8 FILLER_16_442 ();
 sg13g2_decap_8 FILLER_16_449 ();
 sg13g2_decap_8 FILLER_16_456 ();
 sg13g2_decap_8 FILLER_16_463 ();
 sg13g2_decap_8 FILLER_16_470 ();
 sg13g2_decap_8 FILLER_16_477 ();
 sg13g2_fill_1 FILLER_16_484 ();
 sg13g2_fill_2 FILLER_16_531 ();
 sg13g2_decap_8 FILLER_16_585 ();
 sg13g2_decap_8 FILLER_16_592 ();
 sg13g2_decap_8 FILLER_16_599 ();
 sg13g2_decap_8 FILLER_16_606 ();
 sg13g2_decap_4 FILLER_16_613 ();
 sg13g2_decap_4 FILLER_16_633 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_fill_2 FILLER_16_658 ();
 sg13g2_fill_2 FILLER_16_668 ();
 sg13g2_fill_1 FILLER_16_670 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_4 FILLER_16_730 ();
 sg13g2_decap_4 FILLER_16_738 ();
 sg13g2_fill_1 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_fill_1 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_799 ();
 sg13g2_decap_8 FILLER_16_806 ();
 sg13g2_decap_8 FILLER_16_813 ();
 sg13g2_decap_8 FILLER_16_820 ();
 sg13g2_decap_4 FILLER_16_827 ();
 sg13g2_fill_2 FILLER_16_831 ();
 sg13g2_decap_8 FILLER_16_896 ();
 sg13g2_decap_8 FILLER_16_903 ();
 sg13g2_decap_8 FILLER_16_910 ();
 sg13g2_fill_2 FILLER_16_917 ();
 sg13g2_fill_2 FILLER_16_953 ();
 sg13g2_fill_1 FILLER_16_1000 ();
 sg13g2_decap_4 FILLER_16_1027 ();
 sg13g2_fill_2 FILLER_16_1031 ();
 sg13g2_decap_8 FILLER_16_1059 ();
 sg13g2_decap_8 FILLER_16_1066 ();
 sg13g2_decap_8 FILLER_16_1073 ();
 sg13g2_fill_1 FILLER_16_1080 ();
 sg13g2_decap_8 FILLER_16_1090 ();
 sg13g2_decap_8 FILLER_16_1097 ();
 sg13g2_decap_8 FILLER_16_1104 ();
 sg13g2_decap_8 FILLER_16_1111 ();
 sg13g2_decap_8 FILLER_16_1118 ();
 sg13g2_decap_8 FILLER_16_1125 ();
 sg13g2_decap_8 FILLER_16_1164 ();
 sg13g2_decap_8 FILLER_16_1171 ();
 sg13g2_decap_8 FILLER_16_1178 ();
 sg13g2_decap_8 FILLER_16_1185 ();
 sg13g2_decap_8 FILLER_16_1192 ();
 sg13g2_decap_8 FILLER_16_1199 ();
 sg13g2_decap_8 FILLER_16_1245 ();
 sg13g2_decap_8 FILLER_16_1252 ();
 sg13g2_decap_8 FILLER_16_1259 ();
 sg13g2_decap_8 FILLER_16_1266 ();
 sg13g2_decap_8 FILLER_16_1273 ();
 sg13g2_fill_2 FILLER_16_1280 ();
 sg13g2_fill_2 FILLER_16_1316 ();
 sg13g2_fill_1 FILLER_16_1344 ();
 sg13g2_decap_8 FILLER_16_1401 ();
 sg13g2_decap_8 FILLER_16_1408 ();
 sg13g2_decap_8 FILLER_16_1415 ();
 sg13g2_decap_8 FILLER_16_1422 ();
 sg13g2_decap_4 FILLER_16_1429 ();
 sg13g2_fill_2 FILLER_16_1433 ();
 sg13g2_decap_8 FILLER_16_1461 ();
 sg13g2_decap_4 FILLER_16_1468 ();
 sg13g2_fill_2 FILLER_16_1472 ();
 sg13g2_decap_8 FILLER_16_1500 ();
 sg13g2_decap_4 FILLER_16_1507 ();
 sg13g2_fill_1 FILLER_16_1511 ();
 sg13g2_fill_1 FILLER_16_1553 ();
 sg13g2_decap_4 FILLER_16_1585 ();
 sg13g2_fill_1 FILLER_16_1589 ();
 sg13g2_decap_4 FILLER_16_1593 ();
 sg13g2_decap_8 FILLER_16_1605 ();
 sg13g2_decap_8 FILLER_16_1620 ();
 sg13g2_decap_8 FILLER_16_1627 ();
 sg13g2_fill_1 FILLER_16_1634 ();
 sg13g2_decap_8 FILLER_16_1640 ();
 sg13g2_decap_4 FILLER_16_1647 ();
 sg13g2_fill_1 FILLER_16_1651 ();
 sg13g2_decap_4 FILLER_16_1690 ();
 sg13g2_fill_2 FILLER_16_1698 ();
 sg13g2_fill_1 FILLER_16_1700 ();
 sg13g2_fill_2 FILLER_16_1727 ();
 sg13g2_decap_8 FILLER_16_1763 ();
 sg13g2_fill_2 FILLER_16_1770 ();
 sg13g2_decap_8 FILLER_16_1776 ();
 sg13g2_decap_4 FILLER_16_1783 ();
 sg13g2_fill_2 FILLER_16_1787 ();
 sg13g2_fill_2 FILLER_16_1801 ();
 sg13g2_decap_8 FILLER_16_1819 ();
 sg13g2_decap_8 FILLER_16_1826 ();
 sg13g2_decap_4 FILLER_16_1833 ();
 sg13g2_fill_1 FILLER_16_1845 ();
 sg13g2_decap_8 FILLER_16_1880 ();
 sg13g2_decap_4 FILLER_16_1887 ();
 sg13g2_fill_1 FILLER_16_1891 ();
 sg13g2_decap_8 FILLER_16_1918 ();
 sg13g2_decap_8 FILLER_16_1981 ();
 sg13g2_decap_8 FILLER_16_1988 ();
 sg13g2_decap_8 FILLER_16_1995 ();
 sg13g2_decap_4 FILLER_16_2002 ();
 sg13g2_decap_4 FILLER_16_2050 ();
 sg13g2_fill_1 FILLER_16_2054 ();
 sg13g2_decap_8 FILLER_16_2088 ();
 sg13g2_fill_1 FILLER_16_2095 ();
 sg13g2_fill_1 FILLER_16_2134 ();
 sg13g2_fill_2 FILLER_16_2171 ();
 sg13g2_fill_2 FILLER_16_2199 ();
 sg13g2_fill_1 FILLER_16_2201 ();
 sg13g2_decap_8 FILLER_16_2219 ();
 sg13g2_decap_4 FILLER_16_2226 ();
 sg13g2_decap_8 FILLER_16_2261 ();
 sg13g2_fill_2 FILLER_16_2268 ();
 sg13g2_fill_1 FILLER_16_2270 ();
 sg13g2_decap_8 FILLER_16_2297 ();
 sg13g2_decap_8 FILLER_16_2304 ();
 sg13g2_decap_4 FILLER_16_2311 ();
 sg13g2_fill_2 FILLER_16_2318 ();
 sg13g2_fill_1 FILLER_16_2320 ();
 sg13g2_decap_8 FILLER_16_2360 ();
 sg13g2_decap_8 FILLER_16_2367 ();
 sg13g2_decap_8 FILLER_16_2374 ();
 sg13g2_decap_8 FILLER_16_2385 ();
 sg13g2_decap_4 FILLER_16_2392 ();
 sg13g2_decap_8 FILLER_16_2442 ();
 sg13g2_fill_2 FILLER_16_2449 ();
 sg13g2_fill_1 FILLER_16_2451 ();
 sg13g2_fill_1 FILLER_16_2481 ();
 sg13g2_decap_8 FILLER_16_2516 ();
 sg13g2_fill_1 FILLER_16_2523 ();
 sg13g2_decap_8 FILLER_16_2529 ();
 sg13g2_fill_2 FILLER_16_2536 ();
 sg13g2_fill_1 FILLER_16_2542 ();
 sg13g2_decap_4 FILLER_16_2561 ();
 sg13g2_fill_2 FILLER_16_2565 ();
 sg13g2_decap_8 FILLER_16_2601 ();
 sg13g2_fill_1 FILLER_16_2608 ();
 sg13g2_decap_8 FILLER_16_2613 ();
 sg13g2_fill_2 FILLER_16_2620 ();
 sg13g2_decap_4 FILLER_16_2627 ();
 sg13g2_fill_1 FILLER_16_2634 ();
 sg13g2_fill_1 FILLER_16_2639 ();
 sg13g2_fill_2 FILLER_16_2648 ();
 sg13g2_fill_2 FILLER_16_2676 ();
 sg13g2_fill_1 FILLER_16_2678 ();
 sg13g2_decap_4 FILLER_16_2687 ();
 sg13g2_fill_2 FILLER_16_2691 ();
 sg13g2_decap_8 FILLER_16_2729 ();
 sg13g2_decap_8 FILLER_16_2736 ();
 sg13g2_decap_8 FILLER_16_2743 ();
 sg13g2_decap_8 FILLER_16_2750 ();
 sg13g2_decap_8 FILLER_16_2757 ();
 sg13g2_decap_8 FILLER_16_2764 ();
 sg13g2_decap_8 FILLER_16_2771 ();
 sg13g2_decap_8 FILLER_16_2778 ();
 sg13g2_decap_8 FILLER_16_2785 ();
 sg13g2_decap_8 FILLER_16_2792 ();
 sg13g2_decap_8 FILLER_16_2799 ();
 sg13g2_decap_8 FILLER_16_2806 ();
 sg13g2_decap_8 FILLER_16_2813 ();
 sg13g2_decap_8 FILLER_16_2820 ();
 sg13g2_decap_8 FILLER_16_2827 ();
 sg13g2_decap_8 FILLER_16_2834 ();
 sg13g2_decap_8 FILLER_16_2841 ();
 sg13g2_decap_8 FILLER_16_2848 ();
 sg13g2_decap_8 FILLER_16_2855 ();
 sg13g2_decap_8 FILLER_16_2862 ();
 sg13g2_decap_8 FILLER_16_2869 ();
 sg13g2_decap_8 FILLER_16_2876 ();
 sg13g2_decap_8 FILLER_16_2883 ();
 sg13g2_decap_8 FILLER_16_2890 ();
 sg13g2_decap_8 FILLER_16_2897 ();
 sg13g2_decap_8 FILLER_16_2904 ();
 sg13g2_decap_8 FILLER_16_2911 ();
 sg13g2_decap_8 FILLER_16_2918 ();
 sg13g2_decap_8 FILLER_16_2925 ();
 sg13g2_decap_8 FILLER_16_2932 ();
 sg13g2_decap_8 FILLER_16_2939 ();
 sg13g2_decap_8 FILLER_16_2946 ();
 sg13g2_decap_8 FILLER_16_2953 ();
 sg13g2_decap_8 FILLER_16_2960 ();
 sg13g2_decap_8 FILLER_16_2967 ();
 sg13g2_decap_8 FILLER_16_2974 ();
 sg13g2_decap_8 FILLER_16_2981 ();
 sg13g2_decap_8 FILLER_16_2988 ();
 sg13g2_decap_8 FILLER_16_2995 ();
 sg13g2_decap_8 FILLER_16_3002 ();
 sg13g2_decap_8 FILLER_16_3009 ();
 sg13g2_decap_8 FILLER_16_3016 ();
 sg13g2_decap_8 FILLER_16_3023 ();
 sg13g2_decap_8 FILLER_16_3030 ();
 sg13g2_decap_8 FILLER_16_3037 ();
 sg13g2_decap_8 FILLER_16_3044 ();
 sg13g2_decap_8 FILLER_16_3051 ();
 sg13g2_decap_8 FILLER_16_3058 ();
 sg13g2_decap_8 FILLER_16_3065 ();
 sg13g2_decap_8 FILLER_16_3072 ();
 sg13g2_decap_8 FILLER_16_3079 ();
 sg13g2_decap_8 FILLER_16_3086 ();
 sg13g2_decap_8 FILLER_16_3093 ();
 sg13g2_decap_8 FILLER_16_3100 ();
 sg13g2_decap_8 FILLER_16_3107 ();
 sg13g2_decap_8 FILLER_16_3114 ();
 sg13g2_decap_8 FILLER_16_3121 ();
 sg13g2_decap_8 FILLER_16_3128 ();
 sg13g2_decap_8 FILLER_16_3135 ();
 sg13g2_decap_8 FILLER_16_3142 ();
 sg13g2_decap_8 FILLER_16_3149 ();
 sg13g2_decap_8 FILLER_16_3156 ();
 sg13g2_decap_8 FILLER_16_3163 ();
 sg13g2_decap_8 FILLER_16_3170 ();
 sg13g2_decap_8 FILLER_16_3177 ();
 sg13g2_decap_8 FILLER_16_3184 ();
 sg13g2_decap_8 FILLER_16_3191 ();
 sg13g2_decap_8 FILLER_16_3198 ();
 sg13g2_decap_8 FILLER_16_3205 ();
 sg13g2_decap_8 FILLER_16_3212 ();
 sg13g2_decap_8 FILLER_16_3219 ();
 sg13g2_decap_8 FILLER_16_3226 ();
 sg13g2_decap_8 FILLER_16_3233 ();
 sg13g2_decap_8 FILLER_16_3240 ();
 sg13g2_decap_8 FILLER_16_3247 ();
 sg13g2_decap_8 FILLER_16_3254 ();
 sg13g2_decap_8 FILLER_16_3261 ();
 sg13g2_decap_8 FILLER_16_3268 ();
 sg13g2_decap_8 FILLER_16_3275 ();
 sg13g2_decap_8 FILLER_16_3282 ();
 sg13g2_decap_8 FILLER_16_3289 ();
 sg13g2_decap_8 FILLER_16_3296 ();
 sg13g2_decap_8 FILLER_16_3303 ();
 sg13g2_decap_8 FILLER_16_3310 ();
 sg13g2_decap_8 FILLER_16_3317 ();
 sg13g2_decap_8 FILLER_16_3324 ();
 sg13g2_decap_8 FILLER_16_3331 ();
 sg13g2_decap_8 FILLER_16_3338 ();
 sg13g2_decap_8 FILLER_16_3345 ();
 sg13g2_decap_8 FILLER_16_3352 ();
 sg13g2_decap_8 FILLER_16_3359 ();
 sg13g2_decap_8 FILLER_16_3366 ();
 sg13g2_decap_8 FILLER_16_3373 ();
 sg13g2_decap_8 FILLER_16_3380 ();
 sg13g2_decap_8 FILLER_16_3387 ();
 sg13g2_decap_8 FILLER_16_3394 ();
 sg13g2_decap_8 FILLER_16_3401 ();
 sg13g2_decap_8 FILLER_16_3408 ();
 sg13g2_decap_8 FILLER_16_3415 ();
 sg13g2_decap_8 FILLER_16_3422 ();
 sg13g2_decap_8 FILLER_16_3429 ();
 sg13g2_decap_8 FILLER_16_3436 ();
 sg13g2_decap_8 FILLER_16_3443 ();
 sg13g2_decap_8 FILLER_16_3450 ();
 sg13g2_decap_8 FILLER_16_3457 ();
 sg13g2_decap_8 FILLER_16_3464 ();
 sg13g2_decap_8 FILLER_16_3471 ();
 sg13g2_decap_8 FILLER_16_3478 ();
 sg13g2_decap_8 FILLER_16_3485 ();
 sg13g2_decap_8 FILLER_16_3492 ();
 sg13g2_decap_8 FILLER_16_3499 ();
 sg13g2_decap_8 FILLER_16_3506 ();
 sg13g2_decap_8 FILLER_16_3513 ();
 sg13g2_decap_8 FILLER_16_3520 ();
 sg13g2_decap_8 FILLER_16_3527 ();
 sg13g2_decap_8 FILLER_16_3534 ();
 sg13g2_decap_8 FILLER_16_3541 ();
 sg13g2_decap_8 FILLER_16_3548 ();
 sg13g2_decap_8 FILLER_16_3555 ();
 sg13g2_decap_8 FILLER_16_3562 ();
 sg13g2_decap_8 FILLER_16_3569 ();
 sg13g2_decap_4 FILLER_16_3576 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_4 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_113 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_4 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_decap_4 FILLER_17_187 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_fill_1 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_decap_4 FILLER_17_316 ();
 sg13g2_fill_2 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_fill_2 FILLER_17_362 ();
 sg13g2_fill_1 FILLER_17_364 ();
 sg13g2_fill_2 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_432 ();
 sg13g2_fill_2 FILLER_17_439 ();
 sg13g2_fill_1 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_446 ();
 sg13g2_decap_4 FILLER_17_453 ();
 sg13g2_fill_2 FILLER_17_457 ();
 sg13g2_decap_4 FILLER_17_465 ();
 sg13g2_fill_2 FILLER_17_477 ();
 sg13g2_fill_1 FILLER_17_479 ();
 sg13g2_fill_1 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_517 ();
 sg13g2_decap_4 FILLER_17_524 ();
 sg13g2_fill_2 FILLER_17_528 ();
 sg13g2_decap_8 FILLER_17_590 ();
 sg13g2_decap_4 FILLER_17_597 ();
 sg13g2_fill_1 FILLER_17_601 ();
 sg13g2_decap_4 FILLER_17_605 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_4 FILLER_17_686 ();
 sg13g2_fill_1 FILLER_17_729 ();
 sg13g2_decap_4 FILLER_17_782 ();
 sg13g2_fill_2 FILLER_17_799 ();
 sg13g2_decap_4 FILLER_17_827 ();
 sg13g2_fill_1 FILLER_17_831 ();
 sg13g2_decap_8 FILLER_17_865 ();
 sg13g2_decap_8 FILLER_17_872 ();
 sg13g2_decap_8 FILLER_17_879 ();
 sg13g2_decap_8 FILLER_17_886 ();
 sg13g2_decap_8 FILLER_17_893 ();
 sg13g2_fill_2 FILLER_17_900 ();
 sg13g2_decap_8 FILLER_17_906 ();
 sg13g2_decap_8 FILLER_17_913 ();
 sg13g2_decap_8 FILLER_17_920 ();
 sg13g2_decap_8 FILLER_17_927 ();
 sg13g2_fill_1 FILLER_17_947 ();
 sg13g2_decap_8 FILLER_17_953 ();
 sg13g2_fill_2 FILLER_17_960 ();
 sg13g2_fill_1 FILLER_17_962 ();
 sg13g2_decap_8 FILLER_17_1004 ();
 sg13g2_fill_1 FILLER_17_1011 ();
 sg13g2_fill_2 FILLER_17_1016 ();
 sg13g2_decap_4 FILLER_17_1044 ();
 sg13g2_fill_1 FILLER_17_1048 ();
 sg13g2_fill_1 FILLER_17_1075 ();
 sg13g2_decap_4 FILLER_17_1079 ();
 sg13g2_decap_8 FILLER_17_1116 ();
 sg13g2_fill_2 FILLER_17_1123 ();
 sg13g2_fill_1 FILLER_17_1125 ();
 sg13g2_fill_1 FILLER_17_1185 ();
 sg13g2_fill_2 FILLER_17_1212 ();
 sg13g2_fill_1 FILLER_17_1214 ();
 sg13g2_decap_8 FILLER_17_1258 ();
 sg13g2_decap_8 FILLER_17_1265 ();
 sg13g2_decap_8 FILLER_17_1272 ();
 sg13g2_decap_8 FILLER_17_1290 ();
 sg13g2_decap_8 FILLER_17_1297 ();
 sg13g2_decap_8 FILLER_17_1304 ();
 sg13g2_fill_1 FILLER_17_1311 ();
 sg13g2_fill_1 FILLER_17_1364 ();
 sg13g2_decap_8 FILLER_17_1370 ();
 sg13g2_decap_8 FILLER_17_1403 ();
 sg13g2_decap_8 FILLER_17_1410 ();
 sg13g2_fill_2 FILLER_17_1417 ();
 sg13g2_decap_8 FILLER_17_1445 ();
 sg13g2_decap_8 FILLER_17_1452 ();
 sg13g2_decap_8 FILLER_17_1459 ();
 sg13g2_decap_4 FILLER_17_1466 ();
 sg13g2_fill_1 FILLER_17_1470 ();
 sg13g2_fill_2 FILLER_17_1574 ();
 sg13g2_fill_1 FILLER_17_1630 ();
 sg13g2_fill_2 FILLER_17_1654 ();
 sg13g2_fill_1 FILLER_17_1656 ();
 sg13g2_fill_2 FILLER_17_1665 ();
 sg13g2_fill_1 FILLER_17_1667 ();
 sg13g2_decap_8 FILLER_17_1698 ();
 sg13g2_decap_8 FILLER_17_1705 ();
 sg13g2_fill_1 FILLER_17_1716 ();
 sg13g2_decap_8 FILLER_17_1759 ();
 sg13g2_decap_8 FILLER_17_1766 ();
 sg13g2_decap_8 FILLER_17_1773 ();
 sg13g2_fill_1 FILLER_17_1780 ();
 sg13g2_decap_8 FILLER_17_1818 ();
 sg13g2_decap_4 FILLER_17_1825 ();
 sg13g2_fill_1 FILLER_17_1829 ();
 sg13g2_fill_2 FILLER_17_1843 ();
 sg13g2_fill_1 FILLER_17_1845 ();
 sg13g2_decap_4 FILLER_17_1883 ();
 sg13g2_decap_4 FILLER_17_1913 ();
 sg13g2_fill_1 FILLER_17_1917 ();
 sg13g2_fill_2 FILLER_17_1952 ();
 sg13g2_decap_8 FILLER_17_1990 ();
 sg13g2_fill_1 FILLER_17_1997 ();
 sg13g2_decap_8 FILLER_17_2040 ();
 sg13g2_decap_4 FILLER_17_2089 ();
 sg13g2_decap_4 FILLER_17_2140 ();
 sg13g2_fill_2 FILLER_17_2144 ();
 sg13g2_decap_4 FILLER_17_2150 ();
 sg13g2_fill_2 FILLER_17_2154 ();
 sg13g2_fill_1 FILLER_17_2164 ();
 sg13g2_decap_8 FILLER_17_2173 ();
 sg13g2_fill_2 FILLER_17_2214 ();
 sg13g2_fill_1 FILLER_17_2216 ();
 sg13g2_decap_8 FILLER_17_2309 ();
 sg13g2_decap_4 FILLER_17_2316 ();
 sg13g2_fill_2 FILLER_17_2320 ();
 sg13g2_decap_8 FILLER_17_2355 ();
 sg13g2_fill_2 FILLER_17_2414 ();
 sg13g2_decap_8 FILLER_17_2435 ();
 sg13g2_fill_1 FILLER_17_2442 ();
 sg13g2_decap_8 FILLER_17_2486 ();
 sg13g2_decap_4 FILLER_17_2497 ();
 sg13g2_fill_2 FILLER_17_2505 ();
 sg13g2_fill_2 FILLER_17_2543 ();
 sg13g2_decap_8 FILLER_17_2550 ();
 sg13g2_decap_8 FILLER_17_2557 ();
 sg13g2_decap_8 FILLER_17_2564 ();
 sg13g2_decap_8 FILLER_17_2571 ();
 sg13g2_decap_8 FILLER_17_2578 ();
 sg13g2_decap_8 FILLER_17_2585 ();
 sg13g2_decap_8 FILLER_17_2592 ();
 sg13g2_decap_4 FILLER_17_2599 ();
 sg13g2_fill_1 FILLER_17_2603 ();
 sg13g2_fill_1 FILLER_17_2608 ();
 sg13g2_fill_2 FILLER_17_2622 ();
 sg13g2_fill_1 FILLER_17_2624 ();
 sg13g2_fill_2 FILLER_17_2682 ();
 sg13g2_fill_1 FILLER_17_2684 ();
 sg13g2_decap_8 FILLER_17_2720 ();
 sg13g2_decap_8 FILLER_17_2727 ();
 sg13g2_decap_8 FILLER_17_2734 ();
 sg13g2_decap_8 FILLER_17_2741 ();
 sg13g2_decap_8 FILLER_17_2748 ();
 sg13g2_decap_8 FILLER_17_2755 ();
 sg13g2_decap_8 FILLER_17_2762 ();
 sg13g2_decap_8 FILLER_17_2769 ();
 sg13g2_decap_8 FILLER_17_2776 ();
 sg13g2_decap_8 FILLER_17_2783 ();
 sg13g2_decap_8 FILLER_17_2790 ();
 sg13g2_decap_8 FILLER_17_2797 ();
 sg13g2_decap_8 FILLER_17_2804 ();
 sg13g2_decap_8 FILLER_17_2811 ();
 sg13g2_decap_8 FILLER_17_2818 ();
 sg13g2_decap_8 FILLER_17_2825 ();
 sg13g2_decap_8 FILLER_17_2832 ();
 sg13g2_decap_8 FILLER_17_2839 ();
 sg13g2_decap_8 FILLER_17_2846 ();
 sg13g2_decap_8 FILLER_17_2853 ();
 sg13g2_decap_8 FILLER_17_2860 ();
 sg13g2_decap_8 FILLER_17_2867 ();
 sg13g2_decap_8 FILLER_17_2874 ();
 sg13g2_decap_8 FILLER_17_2881 ();
 sg13g2_decap_8 FILLER_17_2888 ();
 sg13g2_decap_8 FILLER_17_2895 ();
 sg13g2_decap_8 FILLER_17_2902 ();
 sg13g2_decap_8 FILLER_17_2909 ();
 sg13g2_decap_8 FILLER_17_2916 ();
 sg13g2_decap_8 FILLER_17_2923 ();
 sg13g2_decap_8 FILLER_17_2930 ();
 sg13g2_decap_8 FILLER_17_2937 ();
 sg13g2_decap_8 FILLER_17_2944 ();
 sg13g2_decap_8 FILLER_17_2951 ();
 sg13g2_decap_8 FILLER_17_2958 ();
 sg13g2_decap_8 FILLER_17_2965 ();
 sg13g2_decap_8 FILLER_17_2972 ();
 sg13g2_decap_8 FILLER_17_2979 ();
 sg13g2_decap_8 FILLER_17_2986 ();
 sg13g2_decap_8 FILLER_17_2993 ();
 sg13g2_decap_8 FILLER_17_3000 ();
 sg13g2_decap_8 FILLER_17_3007 ();
 sg13g2_decap_8 FILLER_17_3014 ();
 sg13g2_decap_8 FILLER_17_3021 ();
 sg13g2_decap_8 FILLER_17_3028 ();
 sg13g2_decap_8 FILLER_17_3035 ();
 sg13g2_decap_8 FILLER_17_3042 ();
 sg13g2_decap_8 FILLER_17_3049 ();
 sg13g2_decap_8 FILLER_17_3056 ();
 sg13g2_decap_8 FILLER_17_3063 ();
 sg13g2_decap_8 FILLER_17_3070 ();
 sg13g2_decap_8 FILLER_17_3077 ();
 sg13g2_decap_8 FILLER_17_3084 ();
 sg13g2_decap_8 FILLER_17_3091 ();
 sg13g2_decap_8 FILLER_17_3098 ();
 sg13g2_decap_8 FILLER_17_3105 ();
 sg13g2_decap_8 FILLER_17_3112 ();
 sg13g2_decap_8 FILLER_17_3119 ();
 sg13g2_decap_8 FILLER_17_3126 ();
 sg13g2_decap_8 FILLER_17_3133 ();
 sg13g2_decap_8 FILLER_17_3140 ();
 sg13g2_decap_8 FILLER_17_3147 ();
 sg13g2_decap_8 FILLER_17_3154 ();
 sg13g2_decap_8 FILLER_17_3161 ();
 sg13g2_decap_8 FILLER_17_3168 ();
 sg13g2_decap_8 FILLER_17_3175 ();
 sg13g2_decap_8 FILLER_17_3182 ();
 sg13g2_decap_8 FILLER_17_3189 ();
 sg13g2_decap_8 FILLER_17_3196 ();
 sg13g2_decap_8 FILLER_17_3203 ();
 sg13g2_decap_8 FILLER_17_3210 ();
 sg13g2_decap_8 FILLER_17_3217 ();
 sg13g2_decap_8 FILLER_17_3224 ();
 sg13g2_decap_8 FILLER_17_3231 ();
 sg13g2_decap_8 FILLER_17_3238 ();
 sg13g2_decap_8 FILLER_17_3245 ();
 sg13g2_decap_8 FILLER_17_3252 ();
 sg13g2_decap_8 FILLER_17_3259 ();
 sg13g2_decap_8 FILLER_17_3266 ();
 sg13g2_decap_8 FILLER_17_3273 ();
 sg13g2_decap_8 FILLER_17_3280 ();
 sg13g2_decap_8 FILLER_17_3287 ();
 sg13g2_decap_8 FILLER_17_3294 ();
 sg13g2_decap_8 FILLER_17_3301 ();
 sg13g2_decap_8 FILLER_17_3308 ();
 sg13g2_decap_8 FILLER_17_3315 ();
 sg13g2_decap_8 FILLER_17_3322 ();
 sg13g2_decap_8 FILLER_17_3329 ();
 sg13g2_decap_8 FILLER_17_3336 ();
 sg13g2_decap_8 FILLER_17_3343 ();
 sg13g2_decap_8 FILLER_17_3350 ();
 sg13g2_decap_8 FILLER_17_3357 ();
 sg13g2_decap_8 FILLER_17_3364 ();
 sg13g2_decap_8 FILLER_17_3371 ();
 sg13g2_decap_8 FILLER_17_3378 ();
 sg13g2_decap_8 FILLER_17_3385 ();
 sg13g2_decap_8 FILLER_17_3392 ();
 sg13g2_decap_8 FILLER_17_3399 ();
 sg13g2_decap_8 FILLER_17_3406 ();
 sg13g2_decap_8 FILLER_17_3413 ();
 sg13g2_decap_8 FILLER_17_3420 ();
 sg13g2_decap_8 FILLER_17_3427 ();
 sg13g2_decap_8 FILLER_17_3434 ();
 sg13g2_decap_8 FILLER_17_3441 ();
 sg13g2_decap_8 FILLER_17_3448 ();
 sg13g2_decap_8 FILLER_17_3455 ();
 sg13g2_decap_8 FILLER_17_3462 ();
 sg13g2_decap_8 FILLER_17_3469 ();
 sg13g2_decap_8 FILLER_17_3476 ();
 sg13g2_decap_8 FILLER_17_3483 ();
 sg13g2_decap_8 FILLER_17_3490 ();
 sg13g2_decap_8 FILLER_17_3497 ();
 sg13g2_decap_8 FILLER_17_3504 ();
 sg13g2_decap_8 FILLER_17_3511 ();
 sg13g2_decap_8 FILLER_17_3518 ();
 sg13g2_decap_8 FILLER_17_3525 ();
 sg13g2_decap_8 FILLER_17_3532 ();
 sg13g2_decap_8 FILLER_17_3539 ();
 sg13g2_decap_8 FILLER_17_3546 ();
 sg13g2_decap_8 FILLER_17_3553 ();
 sg13g2_decap_8 FILLER_17_3560 ();
 sg13g2_decap_8 FILLER_17_3567 ();
 sg13g2_decap_4 FILLER_17_3574 ();
 sg13g2_fill_2 FILLER_17_3578 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_73 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_fill_2 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_fill_2 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_283 ();
 sg13g2_fill_2 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_fill_2 FILLER_18_317 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_357 ();
 sg13g2_decap_4 FILLER_18_364 ();
 sg13g2_fill_1 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_fill_2 FILLER_18_457 ();
 sg13g2_fill_1 FILLER_18_488 ();
 sg13g2_decap_8 FILLER_18_499 ();
 sg13g2_decap_8 FILLER_18_506 ();
 sg13g2_decap_8 FILLER_18_513 ();
 sg13g2_fill_2 FILLER_18_520 ();
 sg13g2_fill_1 FILLER_18_522 ();
 sg13g2_decap_4 FILLER_18_590 ();
 sg13g2_fill_2 FILLER_18_628 ();
 sg13g2_fill_1 FILLER_18_630 ();
 sg13g2_fill_2 FILLER_18_665 ();
 sg13g2_fill_1 FILLER_18_667 ();
 sg13g2_decap_4 FILLER_18_720 ();
 sg13g2_fill_1 FILLER_18_758 ();
 sg13g2_fill_1 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_792 ();
 sg13g2_decap_4 FILLER_18_799 ();
 sg13g2_fill_2 FILLER_18_803 ();
 sg13g2_decap_4 FILLER_18_831 ();
 sg13g2_fill_1 FILLER_18_835 ();
 sg13g2_fill_1 FILLER_18_841 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_decap_4 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_18_927 ();
 sg13g2_decap_4 FILLER_18_934 ();
 sg13g2_decap_8 FILLER_18_946 ();
 sg13g2_decap_8 FILLER_18_953 ();
 sg13g2_decap_8 FILLER_18_960 ();
 sg13g2_decap_8 FILLER_18_967 ();
 sg13g2_decap_8 FILLER_18_974 ();
 sg13g2_decap_8 FILLER_18_981 ();
 sg13g2_decap_8 FILLER_18_1014 ();
 sg13g2_decap_8 FILLER_18_1021 ();
 sg13g2_fill_2 FILLER_18_1028 ();
 sg13g2_fill_1 FILLER_18_1062 ();
 sg13g2_fill_1 FILLER_18_1089 ();
 sg13g2_decap_4 FILLER_18_1182 ();
 sg13g2_fill_2 FILLER_18_1219 ();
 sg13g2_decap_4 FILLER_18_1278 ();
 sg13g2_fill_2 FILLER_18_1285 ();
 sg13g2_fill_1 FILLER_18_1313 ();
 sg13g2_decap_8 FILLER_18_1322 ();
 sg13g2_decap_8 FILLER_18_1338 ();
 sg13g2_decap_8 FILLER_18_1345 ();
 sg13g2_fill_1 FILLER_18_1352 ();
 sg13g2_decap_8 FILLER_18_1379 ();
 sg13g2_decap_8 FILLER_18_1386 ();
 sg13g2_decap_8 FILLER_18_1393 ();
 sg13g2_decap_4 FILLER_18_1400 ();
 sg13g2_decap_8 FILLER_18_1433 ();
 sg13g2_decap_8 FILLER_18_1440 ();
 sg13g2_decap_4 FILLER_18_1447 ();
 sg13g2_fill_1 FILLER_18_1451 ();
 sg13g2_decap_4 FILLER_18_1457 ();
 sg13g2_fill_1 FILLER_18_1461 ();
 sg13g2_fill_1 FILLER_18_1493 ();
 sg13g2_decap_8 FILLER_18_1504 ();
 sg13g2_decap_8 FILLER_18_1511 ();
 sg13g2_fill_2 FILLER_18_1518 ();
 sg13g2_fill_1 FILLER_18_1520 ();
 sg13g2_decap_4 FILLER_18_1567 ();
 sg13g2_decap_8 FILLER_18_1574 ();
 sg13g2_fill_1 FILLER_18_1581 ();
 sg13g2_decap_8 FILLER_18_1620 ();
 sg13g2_decap_4 FILLER_18_1627 ();
 sg13g2_fill_1 FILLER_18_1631 ();
 sg13g2_fill_1 FILLER_18_1658 ();
 sg13g2_decap_4 FILLER_18_1667 ();
 sg13g2_decap_8 FILLER_18_1708 ();
 sg13g2_decap_4 FILLER_18_1715 ();
 sg13g2_fill_1 FILLER_18_1719 ();
 sg13g2_fill_2 FILLER_18_1725 ();
 sg13g2_fill_1 FILLER_18_1727 ();
 sg13g2_fill_2 FILLER_18_1733 ();
 sg13g2_fill_1 FILLER_18_1735 ();
 sg13g2_fill_2 FILLER_18_1741 ();
 sg13g2_fill_1 FILLER_18_1743 ();
 sg13g2_decap_8 FILLER_18_1770 ();
 sg13g2_decap_4 FILLER_18_1777 ();
 sg13g2_decap_4 FILLER_18_1889 ();
 sg13g2_fill_1 FILLER_18_1893 ();
 sg13g2_fill_1 FILLER_18_1924 ();
 sg13g2_fill_2 FILLER_18_1930 ();
 sg13g2_decap_8 FILLER_18_1944 ();
 sg13g2_decap_8 FILLER_18_1977 ();
 sg13g2_decap_8 FILLER_18_1984 ();
 sg13g2_decap_8 FILLER_18_1991 ();
 sg13g2_fill_2 FILLER_18_1998 ();
 sg13g2_fill_1 FILLER_18_2000 ();
 sg13g2_fill_2 FILLER_18_2053 ();
 sg13g2_decap_8 FILLER_18_2078 ();
 sg13g2_decap_8 FILLER_18_2085 ();
 sg13g2_decap_4 FILLER_18_2092 ();
 sg13g2_fill_2 FILLER_18_2096 ();
 sg13g2_fill_2 FILLER_18_2106 ();
 sg13g2_decap_8 FILLER_18_2139 ();
 sg13g2_decap_8 FILLER_18_2146 ();
 sg13g2_decap_8 FILLER_18_2153 ();
 sg13g2_decap_8 FILLER_18_2160 ();
 sg13g2_decap_4 FILLER_18_2167 ();
 sg13g2_fill_1 FILLER_18_2171 ();
 sg13g2_decap_8 FILLER_18_2180 ();
 sg13g2_decap_8 FILLER_18_2187 ();
 sg13g2_fill_1 FILLER_18_2194 ();
 sg13g2_fill_2 FILLER_18_2204 ();
 sg13g2_fill_2 FILLER_18_2236 ();
 sg13g2_fill_1 FILLER_18_2238 ();
 sg13g2_fill_2 FILLER_18_2252 ();
 sg13g2_fill_1 FILLER_18_2254 ();
 sg13g2_decap_8 FILLER_18_2263 ();
 sg13g2_decap_8 FILLER_18_2270 ();
 sg13g2_fill_2 FILLER_18_2277 ();
 sg13g2_fill_1 FILLER_18_2279 ();
 sg13g2_fill_2 FILLER_18_2284 ();
 sg13g2_decap_8 FILLER_18_2338 ();
 sg13g2_fill_1 FILLER_18_2345 ();
 sg13g2_decap_4 FILLER_18_2356 ();
 sg13g2_fill_2 FILLER_18_2360 ();
 sg13g2_decap_8 FILLER_18_2388 ();
 sg13g2_decap_4 FILLER_18_2395 ();
 sg13g2_fill_2 FILLER_18_2403 ();
 sg13g2_fill_2 FILLER_18_2408 ();
 sg13g2_fill_1 FILLER_18_2410 ();
 sg13g2_decap_8 FILLER_18_2426 ();
 sg13g2_decap_8 FILLER_18_2433 ();
 sg13g2_decap_8 FILLER_18_2440 ();
 sg13g2_decap_8 FILLER_18_2447 ();
 sg13g2_decap_4 FILLER_18_2458 ();
 sg13g2_fill_2 FILLER_18_2462 ();
 sg13g2_decap_8 FILLER_18_2482 ();
 sg13g2_fill_1 FILLER_18_2489 ();
 sg13g2_decap_4 FILLER_18_2525 ();
 sg13g2_fill_1 FILLER_18_2529 ();
 sg13g2_decap_8 FILLER_18_2567 ();
 sg13g2_fill_2 FILLER_18_2574 ();
 sg13g2_fill_2 FILLER_18_2592 ();
 sg13g2_fill_2 FILLER_18_2675 ();
 sg13g2_decap_8 FILLER_18_2715 ();
 sg13g2_decap_8 FILLER_18_2722 ();
 sg13g2_decap_8 FILLER_18_2729 ();
 sg13g2_decap_8 FILLER_18_2736 ();
 sg13g2_decap_8 FILLER_18_2743 ();
 sg13g2_decap_8 FILLER_18_2750 ();
 sg13g2_decap_8 FILLER_18_2757 ();
 sg13g2_decap_8 FILLER_18_2764 ();
 sg13g2_decap_8 FILLER_18_2771 ();
 sg13g2_decap_8 FILLER_18_2778 ();
 sg13g2_decap_8 FILLER_18_2785 ();
 sg13g2_decap_8 FILLER_18_2792 ();
 sg13g2_decap_8 FILLER_18_2799 ();
 sg13g2_decap_8 FILLER_18_2806 ();
 sg13g2_decap_8 FILLER_18_2813 ();
 sg13g2_decap_8 FILLER_18_2820 ();
 sg13g2_decap_8 FILLER_18_2827 ();
 sg13g2_decap_8 FILLER_18_2834 ();
 sg13g2_decap_8 FILLER_18_2841 ();
 sg13g2_decap_8 FILLER_18_2848 ();
 sg13g2_decap_8 FILLER_18_2855 ();
 sg13g2_decap_8 FILLER_18_2862 ();
 sg13g2_decap_8 FILLER_18_2869 ();
 sg13g2_decap_8 FILLER_18_2876 ();
 sg13g2_decap_8 FILLER_18_2883 ();
 sg13g2_decap_8 FILLER_18_2890 ();
 sg13g2_decap_8 FILLER_18_2897 ();
 sg13g2_decap_8 FILLER_18_2904 ();
 sg13g2_decap_8 FILLER_18_2911 ();
 sg13g2_decap_8 FILLER_18_2918 ();
 sg13g2_decap_8 FILLER_18_2925 ();
 sg13g2_decap_8 FILLER_18_2932 ();
 sg13g2_decap_8 FILLER_18_2939 ();
 sg13g2_decap_8 FILLER_18_2946 ();
 sg13g2_decap_8 FILLER_18_2953 ();
 sg13g2_decap_8 FILLER_18_2960 ();
 sg13g2_decap_8 FILLER_18_2967 ();
 sg13g2_decap_8 FILLER_18_2974 ();
 sg13g2_decap_8 FILLER_18_2981 ();
 sg13g2_decap_8 FILLER_18_2988 ();
 sg13g2_decap_8 FILLER_18_2995 ();
 sg13g2_decap_8 FILLER_18_3002 ();
 sg13g2_decap_8 FILLER_18_3009 ();
 sg13g2_decap_8 FILLER_18_3016 ();
 sg13g2_decap_8 FILLER_18_3023 ();
 sg13g2_decap_8 FILLER_18_3030 ();
 sg13g2_decap_8 FILLER_18_3037 ();
 sg13g2_decap_8 FILLER_18_3044 ();
 sg13g2_decap_8 FILLER_18_3051 ();
 sg13g2_decap_8 FILLER_18_3058 ();
 sg13g2_decap_8 FILLER_18_3065 ();
 sg13g2_decap_8 FILLER_18_3072 ();
 sg13g2_decap_8 FILLER_18_3079 ();
 sg13g2_decap_8 FILLER_18_3086 ();
 sg13g2_decap_8 FILLER_18_3093 ();
 sg13g2_decap_8 FILLER_18_3100 ();
 sg13g2_decap_8 FILLER_18_3107 ();
 sg13g2_decap_8 FILLER_18_3114 ();
 sg13g2_decap_8 FILLER_18_3121 ();
 sg13g2_decap_8 FILLER_18_3128 ();
 sg13g2_decap_8 FILLER_18_3135 ();
 sg13g2_decap_8 FILLER_18_3142 ();
 sg13g2_decap_8 FILLER_18_3149 ();
 sg13g2_decap_8 FILLER_18_3156 ();
 sg13g2_decap_8 FILLER_18_3163 ();
 sg13g2_decap_8 FILLER_18_3170 ();
 sg13g2_decap_8 FILLER_18_3177 ();
 sg13g2_decap_8 FILLER_18_3184 ();
 sg13g2_decap_8 FILLER_18_3191 ();
 sg13g2_decap_8 FILLER_18_3198 ();
 sg13g2_decap_8 FILLER_18_3205 ();
 sg13g2_decap_8 FILLER_18_3212 ();
 sg13g2_decap_8 FILLER_18_3219 ();
 sg13g2_decap_8 FILLER_18_3226 ();
 sg13g2_decap_8 FILLER_18_3233 ();
 sg13g2_decap_8 FILLER_18_3240 ();
 sg13g2_decap_8 FILLER_18_3247 ();
 sg13g2_decap_8 FILLER_18_3254 ();
 sg13g2_decap_8 FILLER_18_3261 ();
 sg13g2_decap_8 FILLER_18_3268 ();
 sg13g2_decap_8 FILLER_18_3275 ();
 sg13g2_decap_8 FILLER_18_3282 ();
 sg13g2_decap_8 FILLER_18_3289 ();
 sg13g2_decap_8 FILLER_18_3296 ();
 sg13g2_decap_8 FILLER_18_3303 ();
 sg13g2_decap_8 FILLER_18_3310 ();
 sg13g2_decap_8 FILLER_18_3317 ();
 sg13g2_decap_8 FILLER_18_3324 ();
 sg13g2_decap_8 FILLER_18_3331 ();
 sg13g2_decap_8 FILLER_18_3338 ();
 sg13g2_decap_8 FILLER_18_3345 ();
 sg13g2_decap_8 FILLER_18_3352 ();
 sg13g2_decap_8 FILLER_18_3359 ();
 sg13g2_decap_8 FILLER_18_3366 ();
 sg13g2_decap_8 FILLER_18_3373 ();
 sg13g2_decap_8 FILLER_18_3380 ();
 sg13g2_decap_8 FILLER_18_3387 ();
 sg13g2_decap_8 FILLER_18_3394 ();
 sg13g2_decap_8 FILLER_18_3401 ();
 sg13g2_decap_8 FILLER_18_3408 ();
 sg13g2_decap_8 FILLER_18_3415 ();
 sg13g2_decap_8 FILLER_18_3422 ();
 sg13g2_decap_8 FILLER_18_3429 ();
 sg13g2_decap_8 FILLER_18_3436 ();
 sg13g2_decap_8 FILLER_18_3443 ();
 sg13g2_decap_8 FILLER_18_3450 ();
 sg13g2_decap_8 FILLER_18_3457 ();
 sg13g2_decap_8 FILLER_18_3464 ();
 sg13g2_decap_8 FILLER_18_3471 ();
 sg13g2_decap_8 FILLER_18_3478 ();
 sg13g2_decap_8 FILLER_18_3485 ();
 sg13g2_decap_8 FILLER_18_3492 ();
 sg13g2_decap_8 FILLER_18_3499 ();
 sg13g2_decap_8 FILLER_18_3506 ();
 sg13g2_decap_8 FILLER_18_3513 ();
 sg13g2_decap_8 FILLER_18_3520 ();
 sg13g2_decap_8 FILLER_18_3527 ();
 sg13g2_decap_8 FILLER_18_3534 ();
 sg13g2_decap_8 FILLER_18_3541 ();
 sg13g2_decap_8 FILLER_18_3548 ();
 sg13g2_decap_8 FILLER_18_3555 ();
 sg13g2_decap_8 FILLER_18_3562 ();
 sg13g2_decap_8 FILLER_18_3569 ();
 sg13g2_decap_4 FILLER_18_3576 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_29 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_204 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_fill_2 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_220 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_decap_4 FILLER_19_261 ();
 sg13g2_fill_2 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_271 ();
 sg13g2_fill_1 FILLER_19_298 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_fill_2 FILLER_19_349 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_362 ();
 sg13g2_fill_2 FILLER_19_373 ();
 sg13g2_fill_1 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_405 ();
 sg13g2_fill_2 FILLER_19_412 ();
 sg13g2_fill_1 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_503 ();
 sg13g2_decap_8 FILLER_19_510 ();
 sg13g2_decap_8 FILLER_19_543 ();
 sg13g2_decap_8 FILLER_19_550 ();
 sg13g2_decap_4 FILLER_19_557 ();
 sg13g2_fill_2 FILLER_19_587 ();
 sg13g2_fill_2 FILLER_19_596 ();
 sg13g2_fill_2 FILLER_19_624 ();
 sg13g2_decap_8 FILLER_19_657 ();
 sg13g2_decap_4 FILLER_19_664 ();
 sg13g2_fill_1 FILLER_19_668 ();
 sg13g2_fill_2 FILLER_19_702 ();
 sg13g2_fill_2 FILLER_19_735 ();
 sg13g2_fill_1 FILLER_19_737 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_fill_2 FILLER_19_756 ();
 sg13g2_decap_4 FILLER_19_766 ();
 sg13g2_fill_1 FILLER_19_770 ();
 sg13g2_fill_1 FILLER_19_786 ();
 sg13g2_decap_8 FILLER_19_795 ();
 sg13g2_decap_8 FILLER_19_802 ();
 sg13g2_fill_2 FILLER_19_809 ();
 sg13g2_fill_1 FILLER_19_811 ();
 sg13g2_fill_1 FILLER_19_816 ();
 sg13g2_fill_2 FILLER_19_821 ();
 sg13g2_fill_2 FILLER_19_849 ();
 sg13g2_fill_1 FILLER_19_858 ();
 sg13g2_decap_8 FILLER_19_869 ();
 sg13g2_fill_2 FILLER_19_880 ();
 sg13g2_fill_1 FILLER_19_882 ();
 sg13g2_fill_2 FILLER_19_912 ();
 sg13g2_decap_4 FILLER_19_932 ();
 sg13g2_fill_1 FILLER_19_936 ();
 sg13g2_fill_2 FILLER_19_941 ();
 sg13g2_fill_1 FILLER_19_943 ();
 sg13g2_decap_8 FILLER_19_970 ();
 sg13g2_decap_8 FILLER_19_977 ();
 sg13g2_fill_2 FILLER_19_984 ();
 sg13g2_fill_1 FILLER_19_986 ();
 sg13g2_fill_2 FILLER_19_996 ();
 sg13g2_fill_1 FILLER_19_998 ();
 sg13g2_decap_8 FILLER_19_1008 ();
 sg13g2_fill_2 FILLER_19_1015 ();
 sg13g2_fill_1 FILLER_19_1017 ();
 sg13g2_fill_2 FILLER_19_1047 ();
 sg13g2_decap_8 FILLER_19_1056 ();
 sg13g2_fill_1 FILLER_19_1096 ();
 sg13g2_decap_8 FILLER_19_1123 ();
 sg13g2_fill_2 FILLER_19_1130 ();
 sg13g2_fill_1 FILLER_19_1132 ();
 sg13g2_fill_1 FILLER_19_1141 ();
 sg13g2_decap_8 FILLER_19_1164 ();
 sg13g2_decap_4 FILLER_19_1171 ();
 sg13g2_decap_4 FILLER_19_1211 ();
 sg13g2_fill_2 FILLER_19_1215 ();
 sg13g2_decap_8 FILLER_19_1256 ();
 sg13g2_decap_8 FILLER_19_1263 ();
 sg13g2_decap_8 FILLER_19_1270 ();
 sg13g2_decap_4 FILLER_19_1277 ();
 sg13g2_fill_1 FILLER_19_1281 ();
 sg13g2_fill_1 FILLER_19_1285 ();
 sg13g2_fill_1 FILLER_19_1290 ();
 sg13g2_decap_8 FILLER_19_1320 ();
 sg13g2_decap_8 FILLER_19_1327 ();
 sg13g2_decap_8 FILLER_19_1334 ();
 sg13g2_decap_8 FILLER_19_1341 ();
 sg13g2_decap_4 FILLER_19_1348 ();
 sg13g2_fill_2 FILLER_19_1352 ();
 sg13g2_fill_2 FILLER_19_1380 ();
 sg13g2_decap_8 FILLER_19_1385 ();
 sg13g2_decap_8 FILLER_19_1392 ();
 sg13g2_fill_2 FILLER_19_1399 ();
 sg13g2_fill_1 FILLER_19_1401 ();
 sg13g2_decap_4 FILLER_19_1467 ();
 sg13g2_fill_2 FILLER_19_1471 ();
 sg13g2_decap_8 FILLER_19_1477 ();
 sg13g2_fill_1 FILLER_19_1484 ();
 sg13g2_fill_1 FILLER_19_1489 ();
 sg13g2_decap_8 FILLER_19_1495 ();
 sg13g2_fill_2 FILLER_19_1502 ();
 sg13g2_fill_1 FILLER_19_1504 ();
 sg13g2_decap_8 FILLER_19_1513 ();
 sg13g2_decap_4 FILLER_19_1520 ();
 sg13g2_fill_1 FILLER_19_1524 ();
 sg13g2_fill_2 FILLER_19_1529 ();
 sg13g2_decap_8 FILLER_19_1562 ();
 sg13g2_decap_8 FILLER_19_1569 ();
 sg13g2_decap_8 FILLER_19_1576 ();
 sg13g2_decap_8 FILLER_19_1583 ();
 sg13g2_decap_4 FILLER_19_1590 ();
 sg13g2_decap_8 FILLER_19_1599 ();
 sg13g2_decap_8 FILLER_19_1611 ();
 sg13g2_decap_8 FILLER_19_1618 ();
 sg13g2_decap_8 FILLER_19_1625 ();
 sg13g2_decap_4 FILLER_19_1632 ();
 sg13g2_decap_8 FILLER_19_1662 ();
 sg13g2_decap_4 FILLER_19_1669 ();
 sg13g2_fill_2 FILLER_19_1673 ();
 sg13g2_decap_4 FILLER_19_1679 ();
 sg13g2_fill_1 FILLER_19_1709 ();
 sg13g2_fill_2 FILLER_19_1722 ();
 sg13g2_decap_8 FILLER_19_1732 ();
 sg13g2_decap_8 FILLER_19_1739 ();
 sg13g2_decap_8 FILLER_19_1746 ();
 sg13g2_decap_8 FILLER_19_1753 ();
 sg13g2_decap_8 FILLER_19_1760 ();
 sg13g2_decap_4 FILLER_19_1767 ();
 sg13g2_decap_4 FILLER_19_1781 ();
 sg13g2_fill_2 FILLER_19_1785 ();
 sg13g2_fill_2 FILLER_19_1790 ();
 sg13g2_fill_1 FILLER_19_1809 ();
 sg13g2_decap_8 FILLER_19_1836 ();
 sg13g2_fill_1 FILLER_19_1843 ();
 sg13g2_fill_1 FILLER_19_1848 ();
 sg13g2_decap_8 FILLER_19_1854 ();
 sg13g2_fill_2 FILLER_19_1861 ();
 sg13g2_decap_8 FILLER_19_1889 ();
 sg13g2_decap_8 FILLER_19_1896 ();
 sg13g2_fill_2 FILLER_19_1907 ();
 sg13g2_decap_8 FILLER_19_1935 ();
 sg13g2_decap_4 FILLER_19_1942 ();
 sg13g2_decap_8 FILLER_19_1987 ();
 sg13g2_decap_8 FILLER_19_1994 ();
 sg13g2_fill_1 FILLER_19_2001 ();
 sg13g2_decap_8 FILLER_19_2051 ();
 sg13g2_decap_8 FILLER_19_2058 ();
 sg13g2_decap_8 FILLER_19_2065 ();
 sg13g2_decap_8 FILLER_19_2072 ();
 sg13g2_decap_8 FILLER_19_2079 ();
 sg13g2_fill_1 FILLER_19_2086 ();
 sg13g2_decap_8 FILLER_19_2129 ();
 sg13g2_fill_1 FILLER_19_2136 ();
 sg13g2_decap_8 FILLER_19_2168 ();
 sg13g2_decap_4 FILLER_19_2175 ();
 sg13g2_fill_1 FILLER_19_2179 ();
 sg13g2_fill_2 FILLER_19_2196 ();
 sg13g2_decap_8 FILLER_19_2203 ();
 sg13g2_decap_4 FILLER_19_2210 ();
 sg13g2_fill_2 FILLER_19_2214 ();
 sg13g2_decap_8 FILLER_19_2220 ();
 sg13g2_decap_8 FILLER_19_2227 ();
 sg13g2_decap_8 FILLER_19_2234 ();
 sg13g2_fill_2 FILLER_19_2245 ();
 sg13g2_decap_4 FILLER_19_2302 ();
 sg13g2_fill_1 FILLER_19_2306 ();
 sg13g2_fill_1 FILLER_19_2336 ();
 sg13g2_fill_2 FILLER_19_2341 ();
 sg13g2_fill_1 FILLER_19_2343 ();
 sg13g2_decap_8 FILLER_19_2380 ();
 sg13g2_decap_8 FILLER_19_2387 ();
 sg13g2_fill_2 FILLER_19_2394 ();
 sg13g2_decap_8 FILLER_19_2422 ();
 sg13g2_decap_8 FILLER_19_2429 ();
 sg13g2_decap_4 FILLER_19_2436 ();
 sg13g2_fill_2 FILLER_19_2440 ();
 sg13g2_decap_8 FILLER_19_2468 ();
 sg13g2_decap_8 FILLER_19_2475 ();
 sg13g2_decap_4 FILLER_19_2482 ();
 sg13g2_decap_8 FILLER_19_2538 ();
 sg13g2_decap_8 FILLER_19_2545 ();
 sg13g2_fill_1 FILLER_19_2552 ();
 sg13g2_decap_8 FILLER_19_2647 ();
 sg13g2_fill_2 FILLER_19_2659 ();
 sg13g2_decap_8 FILLER_19_2737 ();
 sg13g2_decap_8 FILLER_19_2744 ();
 sg13g2_decap_8 FILLER_19_2751 ();
 sg13g2_decap_8 FILLER_19_2758 ();
 sg13g2_decap_8 FILLER_19_2765 ();
 sg13g2_decap_8 FILLER_19_2772 ();
 sg13g2_decap_8 FILLER_19_2779 ();
 sg13g2_decap_8 FILLER_19_2786 ();
 sg13g2_decap_8 FILLER_19_2793 ();
 sg13g2_decap_8 FILLER_19_2800 ();
 sg13g2_decap_8 FILLER_19_2807 ();
 sg13g2_decap_8 FILLER_19_2814 ();
 sg13g2_decap_8 FILLER_19_2821 ();
 sg13g2_decap_8 FILLER_19_2828 ();
 sg13g2_decap_8 FILLER_19_2835 ();
 sg13g2_decap_8 FILLER_19_2842 ();
 sg13g2_decap_8 FILLER_19_2849 ();
 sg13g2_decap_8 FILLER_19_2856 ();
 sg13g2_decap_8 FILLER_19_2863 ();
 sg13g2_decap_8 FILLER_19_2870 ();
 sg13g2_decap_8 FILLER_19_2877 ();
 sg13g2_decap_8 FILLER_19_2884 ();
 sg13g2_decap_8 FILLER_19_2891 ();
 sg13g2_decap_8 FILLER_19_2898 ();
 sg13g2_decap_8 FILLER_19_2905 ();
 sg13g2_decap_8 FILLER_19_2912 ();
 sg13g2_decap_8 FILLER_19_2919 ();
 sg13g2_decap_8 FILLER_19_2926 ();
 sg13g2_decap_8 FILLER_19_2933 ();
 sg13g2_decap_8 FILLER_19_2940 ();
 sg13g2_decap_8 FILLER_19_2947 ();
 sg13g2_decap_8 FILLER_19_2954 ();
 sg13g2_decap_8 FILLER_19_2961 ();
 sg13g2_decap_8 FILLER_19_2968 ();
 sg13g2_decap_8 FILLER_19_2975 ();
 sg13g2_decap_8 FILLER_19_2982 ();
 sg13g2_decap_8 FILLER_19_2989 ();
 sg13g2_decap_8 FILLER_19_2996 ();
 sg13g2_decap_8 FILLER_19_3003 ();
 sg13g2_decap_8 FILLER_19_3010 ();
 sg13g2_decap_8 FILLER_19_3017 ();
 sg13g2_decap_8 FILLER_19_3024 ();
 sg13g2_decap_8 FILLER_19_3031 ();
 sg13g2_decap_8 FILLER_19_3038 ();
 sg13g2_decap_8 FILLER_19_3045 ();
 sg13g2_decap_8 FILLER_19_3052 ();
 sg13g2_decap_8 FILLER_19_3059 ();
 sg13g2_decap_8 FILLER_19_3066 ();
 sg13g2_decap_8 FILLER_19_3073 ();
 sg13g2_decap_8 FILLER_19_3080 ();
 sg13g2_decap_8 FILLER_19_3087 ();
 sg13g2_decap_8 FILLER_19_3094 ();
 sg13g2_decap_8 FILLER_19_3101 ();
 sg13g2_decap_8 FILLER_19_3108 ();
 sg13g2_decap_8 FILLER_19_3115 ();
 sg13g2_decap_8 FILLER_19_3122 ();
 sg13g2_decap_8 FILLER_19_3129 ();
 sg13g2_decap_8 FILLER_19_3136 ();
 sg13g2_decap_8 FILLER_19_3143 ();
 sg13g2_decap_8 FILLER_19_3150 ();
 sg13g2_decap_8 FILLER_19_3157 ();
 sg13g2_decap_8 FILLER_19_3164 ();
 sg13g2_decap_8 FILLER_19_3171 ();
 sg13g2_decap_8 FILLER_19_3178 ();
 sg13g2_decap_8 FILLER_19_3185 ();
 sg13g2_decap_8 FILLER_19_3192 ();
 sg13g2_decap_8 FILLER_19_3199 ();
 sg13g2_decap_8 FILLER_19_3206 ();
 sg13g2_decap_8 FILLER_19_3213 ();
 sg13g2_decap_8 FILLER_19_3220 ();
 sg13g2_decap_8 FILLER_19_3227 ();
 sg13g2_decap_8 FILLER_19_3234 ();
 sg13g2_decap_8 FILLER_19_3241 ();
 sg13g2_decap_8 FILLER_19_3248 ();
 sg13g2_decap_8 FILLER_19_3255 ();
 sg13g2_decap_8 FILLER_19_3262 ();
 sg13g2_decap_8 FILLER_19_3269 ();
 sg13g2_decap_8 FILLER_19_3276 ();
 sg13g2_decap_8 FILLER_19_3283 ();
 sg13g2_decap_8 FILLER_19_3290 ();
 sg13g2_decap_8 FILLER_19_3297 ();
 sg13g2_decap_8 FILLER_19_3304 ();
 sg13g2_decap_8 FILLER_19_3311 ();
 sg13g2_decap_8 FILLER_19_3318 ();
 sg13g2_decap_8 FILLER_19_3325 ();
 sg13g2_decap_8 FILLER_19_3332 ();
 sg13g2_decap_8 FILLER_19_3339 ();
 sg13g2_decap_8 FILLER_19_3346 ();
 sg13g2_decap_8 FILLER_19_3353 ();
 sg13g2_decap_8 FILLER_19_3360 ();
 sg13g2_decap_8 FILLER_19_3367 ();
 sg13g2_decap_8 FILLER_19_3374 ();
 sg13g2_decap_8 FILLER_19_3381 ();
 sg13g2_decap_8 FILLER_19_3388 ();
 sg13g2_decap_8 FILLER_19_3395 ();
 sg13g2_decap_8 FILLER_19_3402 ();
 sg13g2_decap_8 FILLER_19_3409 ();
 sg13g2_decap_8 FILLER_19_3416 ();
 sg13g2_decap_8 FILLER_19_3423 ();
 sg13g2_decap_8 FILLER_19_3430 ();
 sg13g2_decap_8 FILLER_19_3437 ();
 sg13g2_decap_8 FILLER_19_3444 ();
 sg13g2_decap_8 FILLER_19_3451 ();
 sg13g2_decap_8 FILLER_19_3458 ();
 sg13g2_decap_8 FILLER_19_3465 ();
 sg13g2_decap_8 FILLER_19_3472 ();
 sg13g2_decap_8 FILLER_19_3479 ();
 sg13g2_decap_8 FILLER_19_3486 ();
 sg13g2_decap_8 FILLER_19_3493 ();
 sg13g2_decap_8 FILLER_19_3500 ();
 sg13g2_decap_8 FILLER_19_3507 ();
 sg13g2_decap_8 FILLER_19_3514 ();
 sg13g2_decap_8 FILLER_19_3521 ();
 sg13g2_decap_8 FILLER_19_3528 ();
 sg13g2_decap_8 FILLER_19_3535 ();
 sg13g2_decap_8 FILLER_19_3542 ();
 sg13g2_decap_8 FILLER_19_3549 ();
 sg13g2_decap_8 FILLER_19_3556 ();
 sg13g2_decap_8 FILLER_19_3563 ();
 sg13g2_decap_8 FILLER_19_3570 ();
 sg13g2_fill_2 FILLER_19_3577 ();
 sg13g2_fill_1 FILLER_19_3579 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_211 ();
 sg13g2_fill_1 FILLER_20_223 ();
 sg13g2_decap_4 FILLER_20_253 ();
 sg13g2_fill_1 FILLER_20_319 ();
 sg13g2_decap_4 FILLER_20_325 ();
 sg13g2_fill_1 FILLER_20_329 ();
 sg13g2_fill_1 FILLER_20_334 ();
 sg13g2_decap_4 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_fill_2 FILLER_20_409 ();
 sg13g2_fill_2 FILLER_20_472 ();
 sg13g2_decap_4 FILLER_20_513 ();
 sg13g2_fill_2 FILLER_20_517 ();
 sg13g2_decap_8 FILLER_20_545 ();
 sg13g2_decap_8 FILLER_20_552 ();
 sg13g2_fill_1 FILLER_20_559 ();
 sg13g2_decap_8 FILLER_20_576 ();
 sg13g2_decap_8 FILLER_20_583 ();
 sg13g2_decap_8 FILLER_20_646 ();
 sg13g2_decap_8 FILLER_20_653 ();
 sg13g2_decap_8 FILLER_20_660 ();
 sg13g2_fill_2 FILLER_20_667 ();
 sg13g2_decap_8 FILLER_20_702 ();
 sg13g2_decap_8 FILLER_20_709 ();
 sg13g2_decap_8 FILLER_20_716 ();
 sg13g2_decap_4 FILLER_20_723 ();
 sg13g2_fill_1 FILLER_20_727 ();
 sg13g2_fill_1 FILLER_20_783 ();
 sg13g2_decap_8 FILLER_20_792 ();
 sg13g2_decap_8 FILLER_20_799 ();
 sg13g2_fill_1 FILLER_20_832 ();
 sg13g2_decap_8 FILLER_20_837 ();
 sg13g2_fill_2 FILLER_20_875 ();
 sg13g2_fill_1 FILLER_20_877 ();
 sg13g2_decap_8 FILLER_20_999 ();
 sg13g2_decap_8 FILLER_20_1006 ();
 sg13g2_decap_8 FILLER_20_1013 ();
 sg13g2_fill_2 FILLER_20_1020 ();
 sg13g2_fill_1 FILLER_20_1022 ();
 sg13g2_decap_8 FILLER_20_1056 ();
 sg13g2_decap_8 FILLER_20_1063 ();
 sg13g2_decap_4 FILLER_20_1083 ();
 sg13g2_fill_2 FILLER_20_1087 ();
 sg13g2_decap_4 FILLER_20_1125 ();
 sg13g2_decap_8 FILLER_20_1160 ();
 sg13g2_decap_8 FILLER_20_1167 ();
 sg13g2_decap_8 FILLER_20_1174 ();
 sg13g2_decap_4 FILLER_20_1181 ();
 sg13g2_fill_2 FILLER_20_1185 ();
 sg13g2_decap_8 FILLER_20_1216 ();
 sg13g2_decap_4 FILLER_20_1223 ();
 sg13g2_fill_1 FILLER_20_1227 ();
 sg13g2_decap_4 FILLER_20_1260 ();
 sg13g2_fill_1 FILLER_20_1264 ();
 sg13g2_fill_2 FILLER_20_1272 ();
 sg13g2_fill_1 FILLER_20_1274 ();
 sg13g2_fill_2 FILLER_20_1301 ();
 sg13g2_decap_8 FILLER_20_1334 ();
 sg13g2_decap_8 FILLER_20_1341 ();
 sg13g2_fill_2 FILLER_20_1348 ();
 sg13g2_decap_4 FILLER_20_1405 ();
 sg13g2_fill_2 FILLER_20_1409 ();
 sg13g2_fill_1 FILLER_20_1450 ();
 sg13g2_fill_2 FILLER_20_1456 ();
 sg13g2_decap_8 FILLER_20_1466 ();
 sg13g2_fill_1 FILLER_20_1473 ();
 sg13g2_decap_8 FILLER_20_1478 ();
 sg13g2_fill_1 FILLER_20_1485 ();
 sg13g2_decap_4 FILLER_20_1489 ();
 sg13g2_fill_2 FILLER_20_1493 ();
 sg13g2_decap_4 FILLER_20_1502 ();
 sg13g2_fill_2 FILLER_20_1506 ();
 sg13g2_decap_8 FILLER_20_1513 ();
 sg13g2_decap_8 FILLER_20_1520 ();
 sg13g2_decap_8 FILLER_20_1527 ();
 sg13g2_fill_2 FILLER_20_1534 ();
 sg13g2_decap_8 FILLER_20_1562 ();
 sg13g2_decap_8 FILLER_20_1569 ();
 sg13g2_decap_4 FILLER_20_1576 ();
 sg13g2_fill_2 FILLER_20_1580 ();
 sg13g2_fill_2 FILLER_20_1594 ();
 sg13g2_fill_1 FILLER_20_1604 ();
 sg13g2_decap_8 FILLER_20_1634 ();
 sg13g2_fill_1 FILLER_20_1641 ();
 sg13g2_decap_8 FILLER_20_1672 ();
 sg13g2_decap_8 FILLER_20_1679 ();
 sg13g2_decap_8 FILLER_20_1686 ();
 sg13g2_fill_1 FILLER_20_1693 ();
 sg13g2_fill_2 FILLER_20_1698 ();
 sg13g2_decap_8 FILLER_20_1739 ();
 sg13g2_decap_4 FILLER_20_1746 ();
 sg13g2_fill_1 FILLER_20_1750 ();
 sg13g2_decap_8 FILLER_20_1790 ();
 sg13g2_fill_1 FILLER_20_1797 ();
 sg13g2_decap_8 FILLER_20_1811 ();
 sg13g2_decap_8 FILLER_20_1818 ();
 sg13g2_decap_8 FILLER_20_1825 ();
 sg13g2_decap_8 FILLER_20_1832 ();
 sg13g2_decap_8 FILLER_20_1839 ();
 sg13g2_decap_8 FILLER_20_1846 ();
 sg13g2_decap_8 FILLER_20_1853 ();
 sg13g2_decap_8 FILLER_20_1860 ();
 sg13g2_fill_2 FILLER_20_1867 ();
 sg13g2_fill_1 FILLER_20_1873 ();
 sg13g2_fill_2 FILLER_20_1878 ();
 sg13g2_fill_1 FILLER_20_1888 ();
 sg13g2_decap_8 FILLER_20_1892 ();
 sg13g2_decap_8 FILLER_20_1899 ();
 sg13g2_decap_8 FILLER_20_1906 ();
 sg13g2_decap_8 FILLER_20_1913 ();
 sg13g2_decap_8 FILLER_20_1920 ();
 sg13g2_decap_8 FILLER_20_1927 ();
 sg13g2_decap_4 FILLER_20_1934 ();
 sg13g2_fill_2 FILLER_20_1938 ();
 sg13g2_decap_8 FILLER_20_1996 ();
 sg13g2_fill_2 FILLER_20_2003 ();
 sg13g2_fill_1 FILLER_20_2005 ();
 sg13g2_decap_8 FILLER_20_2039 ();
 sg13g2_decap_8 FILLER_20_2046 ();
 sg13g2_decap_8 FILLER_20_2053 ();
 sg13g2_decap_8 FILLER_20_2060 ();
 sg13g2_decap_4 FILLER_20_2067 ();
 sg13g2_fill_1 FILLER_20_2128 ();
 sg13g2_fill_2 FILLER_20_2155 ();
 sg13g2_decap_4 FILLER_20_2183 ();
 sg13g2_decap_8 FILLER_20_2213 ();
 sg13g2_decap_8 FILLER_20_2220 ();
 sg13g2_decap_8 FILLER_20_2227 ();
 sg13g2_decap_4 FILLER_20_2234 ();
 sg13g2_fill_1 FILLER_20_2238 ();
 sg13g2_decap_4 FILLER_20_2275 ();
 sg13g2_decap_8 FILLER_20_2318 ();
 sg13g2_fill_2 FILLER_20_2325 ();
 sg13g2_fill_1 FILLER_20_2327 ();
 sg13g2_fill_2 FILLER_20_2354 ();
 sg13g2_decap_8 FILLER_20_2382 ();
 sg13g2_decap_8 FILLER_20_2389 ();
 sg13g2_decap_8 FILLER_20_2396 ();
 sg13g2_decap_8 FILLER_20_2403 ();
 sg13g2_fill_2 FILLER_20_2410 ();
 sg13g2_fill_1 FILLER_20_2412 ();
 sg13g2_decap_8 FILLER_20_2418 ();
 sg13g2_decap_4 FILLER_20_2425 ();
 sg13g2_decap_4 FILLER_20_2434 ();
 sg13g2_decap_8 FILLER_20_2542 ();
 sg13g2_decap_4 FILLER_20_2559 ();
 sg13g2_decap_8 FILLER_20_2567 ();
 sg13g2_fill_2 FILLER_20_2574 ();
 sg13g2_fill_1 FILLER_20_2576 ();
 sg13g2_fill_2 FILLER_20_2605 ();
 sg13g2_decap_8 FILLER_20_2641 ();
 sg13g2_decap_8 FILLER_20_2648 ();
 sg13g2_decap_4 FILLER_20_2655 ();
 sg13g2_fill_2 FILLER_20_2659 ();
 sg13g2_fill_2 FILLER_20_2665 ();
 sg13g2_fill_1 FILLER_20_2696 ();
 sg13g2_decap_8 FILLER_20_2726 ();
 sg13g2_decap_8 FILLER_20_2733 ();
 sg13g2_decap_8 FILLER_20_2740 ();
 sg13g2_decap_8 FILLER_20_2747 ();
 sg13g2_decap_8 FILLER_20_2754 ();
 sg13g2_decap_8 FILLER_20_2761 ();
 sg13g2_decap_8 FILLER_20_2768 ();
 sg13g2_decap_8 FILLER_20_2775 ();
 sg13g2_decap_8 FILLER_20_2782 ();
 sg13g2_decap_8 FILLER_20_2789 ();
 sg13g2_decap_8 FILLER_20_2796 ();
 sg13g2_decap_8 FILLER_20_2803 ();
 sg13g2_decap_8 FILLER_20_2810 ();
 sg13g2_decap_8 FILLER_20_2817 ();
 sg13g2_decap_8 FILLER_20_2824 ();
 sg13g2_decap_8 FILLER_20_2831 ();
 sg13g2_decap_8 FILLER_20_2838 ();
 sg13g2_decap_8 FILLER_20_2845 ();
 sg13g2_decap_8 FILLER_20_2852 ();
 sg13g2_decap_8 FILLER_20_2859 ();
 sg13g2_decap_8 FILLER_20_2866 ();
 sg13g2_decap_8 FILLER_20_2873 ();
 sg13g2_decap_8 FILLER_20_2880 ();
 sg13g2_decap_8 FILLER_20_2887 ();
 sg13g2_decap_8 FILLER_20_2894 ();
 sg13g2_decap_8 FILLER_20_2901 ();
 sg13g2_decap_8 FILLER_20_2908 ();
 sg13g2_decap_8 FILLER_20_2915 ();
 sg13g2_decap_8 FILLER_20_2922 ();
 sg13g2_decap_8 FILLER_20_2929 ();
 sg13g2_decap_8 FILLER_20_2936 ();
 sg13g2_decap_8 FILLER_20_2943 ();
 sg13g2_decap_8 FILLER_20_2950 ();
 sg13g2_decap_8 FILLER_20_2957 ();
 sg13g2_decap_8 FILLER_20_2964 ();
 sg13g2_decap_8 FILLER_20_2971 ();
 sg13g2_decap_8 FILLER_20_2978 ();
 sg13g2_decap_8 FILLER_20_2985 ();
 sg13g2_decap_8 FILLER_20_2992 ();
 sg13g2_decap_8 FILLER_20_2999 ();
 sg13g2_decap_8 FILLER_20_3006 ();
 sg13g2_decap_8 FILLER_20_3013 ();
 sg13g2_decap_8 FILLER_20_3020 ();
 sg13g2_decap_8 FILLER_20_3027 ();
 sg13g2_decap_8 FILLER_20_3034 ();
 sg13g2_decap_8 FILLER_20_3041 ();
 sg13g2_decap_8 FILLER_20_3048 ();
 sg13g2_decap_8 FILLER_20_3055 ();
 sg13g2_decap_8 FILLER_20_3062 ();
 sg13g2_decap_8 FILLER_20_3069 ();
 sg13g2_decap_8 FILLER_20_3076 ();
 sg13g2_decap_8 FILLER_20_3083 ();
 sg13g2_decap_8 FILLER_20_3090 ();
 sg13g2_decap_8 FILLER_20_3097 ();
 sg13g2_decap_8 FILLER_20_3104 ();
 sg13g2_decap_8 FILLER_20_3111 ();
 sg13g2_decap_8 FILLER_20_3118 ();
 sg13g2_decap_8 FILLER_20_3125 ();
 sg13g2_decap_8 FILLER_20_3132 ();
 sg13g2_decap_8 FILLER_20_3139 ();
 sg13g2_decap_8 FILLER_20_3146 ();
 sg13g2_decap_8 FILLER_20_3153 ();
 sg13g2_decap_8 FILLER_20_3160 ();
 sg13g2_decap_8 FILLER_20_3167 ();
 sg13g2_decap_8 FILLER_20_3174 ();
 sg13g2_decap_8 FILLER_20_3181 ();
 sg13g2_decap_8 FILLER_20_3188 ();
 sg13g2_decap_8 FILLER_20_3195 ();
 sg13g2_decap_8 FILLER_20_3202 ();
 sg13g2_decap_8 FILLER_20_3209 ();
 sg13g2_decap_8 FILLER_20_3216 ();
 sg13g2_decap_8 FILLER_20_3223 ();
 sg13g2_decap_8 FILLER_20_3230 ();
 sg13g2_decap_8 FILLER_20_3237 ();
 sg13g2_decap_8 FILLER_20_3244 ();
 sg13g2_decap_8 FILLER_20_3251 ();
 sg13g2_decap_8 FILLER_20_3258 ();
 sg13g2_decap_8 FILLER_20_3265 ();
 sg13g2_decap_8 FILLER_20_3272 ();
 sg13g2_decap_8 FILLER_20_3279 ();
 sg13g2_decap_8 FILLER_20_3286 ();
 sg13g2_decap_8 FILLER_20_3293 ();
 sg13g2_decap_8 FILLER_20_3300 ();
 sg13g2_decap_8 FILLER_20_3307 ();
 sg13g2_decap_8 FILLER_20_3314 ();
 sg13g2_decap_8 FILLER_20_3321 ();
 sg13g2_decap_8 FILLER_20_3328 ();
 sg13g2_decap_8 FILLER_20_3335 ();
 sg13g2_decap_8 FILLER_20_3342 ();
 sg13g2_decap_8 FILLER_20_3349 ();
 sg13g2_decap_8 FILLER_20_3356 ();
 sg13g2_decap_8 FILLER_20_3363 ();
 sg13g2_decap_8 FILLER_20_3370 ();
 sg13g2_decap_8 FILLER_20_3377 ();
 sg13g2_decap_8 FILLER_20_3384 ();
 sg13g2_decap_8 FILLER_20_3391 ();
 sg13g2_decap_8 FILLER_20_3398 ();
 sg13g2_decap_8 FILLER_20_3405 ();
 sg13g2_decap_8 FILLER_20_3412 ();
 sg13g2_decap_8 FILLER_20_3419 ();
 sg13g2_decap_8 FILLER_20_3426 ();
 sg13g2_decap_8 FILLER_20_3433 ();
 sg13g2_decap_8 FILLER_20_3440 ();
 sg13g2_decap_8 FILLER_20_3447 ();
 sg13g2_decap_8 FILLER_20_3454 ();
 sg13g2_decap_8 FILLER_20_3461 ();
 sg13g2_decap_8 FILLER_20_3468 ();
 sg13g2_decap_8 FILLER_20_3475 ();
 sg13g2_decap_8 FILLER_20_3482 ();
 sg13g2_decap_8 FILLER_20_3489 ();
 sg13g2_decap_8 FILLER_20_3496 ();
 sg13g2_decap_8 FILLER_20_3503 ();
 sg13g2_decap_8 FILLER_20_3510 ();
 sg13g2_decap_8 FILLER_20_3517 ();
 sg13g2_decap_8 FILLER_20_3524 ();
 sg13g2_decap_8 FILLER_20_3531 ();
 sg13g2_decap_8 FILLER_20_3538 ();
 sg13g2_decap_8 FILLER_20_3545 ();
 sg13g2_decap_8 FILLER_20_3552 ();
 sg13g2_decap_8 FILLER_20_3559 ();
 sg13g2_decap_8 FILLER_20_3566 ();
 sg13g2_decap_8 FILLER_20_3573 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_fill_1 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_decap_8 FILLER_21_68 ();
 sg13g2_decap_8 FILLER_21_75 ();
 sg13g2_fill_2 FILLER_21_82 ();
 sg13g2_fill_2 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_204 ();
 sg13g2_decap_4 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_4 FILLER_21_256 ();
 sg13g2_fill_2 FILLER_21_324 ();
 sg13g2_fill_1 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_fill_2 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_356 ();
 sg13g2_fill_2 FILLER_21_387 ();
 sg13g2_fill_1 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_406 ();
 sg13g2_fill_2 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_fill_2 FILLER_21_448 ();
 sg13g2_fill_1 FILLER_21_450 ();
 sg13g2_fill_1 FILLER_21_455 ();
 sg13g2_fill_2 FILLER_21_477 ();
 sg13g2_fill_1 FILLER_21_479 ();
 sg13g2_decap_8 FILLER_21_485 ();
 sg13g2_decap_4 FILLER_21_492 ();
 sg13g2_decap_4 FILLER_21_501 ();
 sg13g2_decap_8 FILLER_21_513 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_4 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_594 ();
 sg13g2_decap_8 FILLER_21_601 ();
 sg13g2_decap_8 FILLER_21_608 ();
 sg13g2_fill_2 FILLER_21_615 ();
 sg13g2_decap_8 FILLER_21_625 ();
 sg13g2_decap_8 FILLER_21_632 ();
 sg13g2_decap_8 FILLER_21_639 ();
 sg13g2_decap_8 FILLER_21_646 ();
 sg13g2_fill_1 FILLER_21_653 ();
 sg13g2_decap_8 FILLER_21_657 ();
 sg13g2_decap_4 FILLER_21_664 ();
 sg13g2_decap_8 FILLER_21_694 ();
 sg13g2_decap_8 FILLER_21_701 ();
 sg13g2_decap_8 FILLER_21_708 ();
 sg13g2_fill_1 FILLER_21_715 ();
 sg13g2_fill_1 FILLER_21_720 ();
 sg13g2_fill_2 FILLER_21_755 ();
 sg13g2_fill_2 FILLER_21_791 ();
 sg13g2_fill_1 FILLER_21_793 ();
 sg13g2_decap_8 FILLER_21_824 ();
 sg13g2_decap_8 FILLER_21_831 ();
 sg13g2_decap_8 FILLER_21_838 ();
 sg13g2_decap_4 FILLER_21_845 ();
 sg13g2_fill_2 FILLER_21_930 ();
 sg13g2_fill_1 FILLER_21_932 ();
 sg13g2_decap_8 FILLER_21_963 ();
 sg13g2_fill_2 FILLER_21_970 ();
 sg13g2_decap_8 FILLER_21_1005 ();
 sg13g2_decap_8 FILLER_21_1012 ();
 sg13g2_decap_4 FILLER_21_1019 ();
 sg13g2_fill_1 FILLER_21_1023 ();
 sg13g2_decap_4 FILLER_21_1053 ();
 sg13g2_fill_2 FILLER_21_1057 ();
 sg13g2_decap_8 FILLER_21_1093 ();
 sg13g2_fill_1 FILLER_21_1103 ();
 sg13g2_fill_2 FILLER_21_1137 ();
 sg13g2_decap_8 FILLER_21_1165 ();
 sg13g2_decap_8 FILLER_21_1172 ();
 sg13g2_decap_8 FILLER_21_1179 ();
 sg13g2_decap_4 FILLER_21_1186 ();
 sg13g2_fill_2 FILLER_21_1190 ();
 sg13g2_decap_4 FILLER_21_1218 ();
 sg13g2_fill_2 FILLER_21_1222 ();
 sg13g2_decap_8 FILLER_21_1283 ();
 sg13g2_fill_1 FILLER_21_1293 ();
 sg13g2_fill_2 FILLER_21_1310 ();
 sg13g2_fill_1 FILLER_21_1312 ();
 sg13g2_decap_8 FILLER_21_1335 ();
 sg13g2_fill_2 FILLER_21_1368 ();
 sg13g2_fill_2 FILLER_21_1388 ();
 sg13g2_decap_4 FILLER_21_1394 ();
 sg13g2_fill_2 FILLER_21_1416 ();
 sg13g2_fill_1 FILLER_21_1418 ();
 sg13g2_decap_8 FILLER_21_1445 ();
 sg13g2_decap_4 FILLER_21_1452 ();
 sg13g2_fill_2 FILLER_21_1456 ();
 sg13g2_fill_1 FILLER_21_1518 ();
 sg13g2_decap_4 FILLER_21_1527 ();
 sg13g2_fill_1 FILLER_21_1531 ();
 sg13g2_decap_8 FILLER_21_1558 ();
 sg13g2_decap_8 FILLER_21_1565 ();
 sg13g2_decap_4 FILLER_21_1572 ();
 sg13g2_fill_1 FILLER_21_1576 ();
 sg13g2_fill_1 FILLER_21_1633 ();
 sg13g2_decap_8 FILLER_21_1660 ();
 sg13g2_decap_8 FILLER_21_1667 ();
 sg13g2_decap_8 FILLER_21_1674 ();
 sg13g2_decap_4 FILLER_21_1681 ();
 sg13g2_fill_2 FILLER_21_1685 ();
 sg13g2_decap_8 FILLER_21_1734 ();
 sg13g2_decap_4 FILLER_21_1741 ();
 sg13g2_fill_2 FILLER_21_1745 ();
 sg13g2_decap_8 FILLER_21_1792 ();
 sg13g2_fill_1 FILLER_21_1803 ();
 sg13g2_decap_8 FILLER_21_1830 ();
 sg13g2_decap_4 FILLER_21_1837 ();
 sg13g2_fill_2 FILLER_21_1841 ();
 sg13g2_decap_8 FILLER_21_1852 ();
 sg13g2_decap_4 FILLER_21_1859 ();
 sg13g2_fill_2 FILLER_21_1863 ();
 sg13g2_decap_8 FILLER_21_1900 ();
 sg13g2_decap_4 FILLER_21_1907 ();
 sg13g2_fill_2 FILLER_21_1911 ();
 sg13g2_fill_2 FILLER_21_1932 ();
 sg13g2_fill_2 FILLER_21_1947 ();
 sg13g2_fill_1 FILLER_21_1963 ();
 sg13g2_decap_8 FILLER_21_1993 ();
 sg13g2_decap_8 FILLER_21_2000 ();
 sg13g2_decap_4 FILLER_21_2007 ();
 sg13g2_decap_8 FILLER_21_2047 ();
 sg13g2_fill_2 FILLER_21_2054 ();
 sg13g2_fill_1 FILLER_21_2092 ();
 sg13g2_fill_2 FILLER_21_2124 ();
 sg13g2_fill_1 FILLER_21_2126 ();
 sg13g2_fill_1 FILLER_21_2179 ();
 sg13g2_decap_8 FILLER_21_2214 ();
 sg13g2_decap_8 FILLER_21_2221 ();
 sg13g2_fill_1 FILLER_21_2228 ();
 sg13g2_fill_2 FILLER_21_2288 ();
 sg13g2_decap_8 FILLER_21_2294 ();
 sg13g2_fill_2 FILLER_21_2301 ();
 sg13g2_decap_8 FILLER_21_2306 ();
 sg13g2_decap_8 FILLER_21_2313 ();
 sg13g2_decap_8 FILLER_21_2320 ();
 sg13g2_decap_8 FILLER_21_2327 ();
 sg13g2_fill_2 FILLER_21_2334 ();
 sg13g2_fill_1 FILLER_21_2336 ();
 sg13g2_decap_8 FILLER_21_2371 ();
 sg13g2_decap_8 FILLER_21_2378 ();
 sg13g2_decap_8 FILLER_21_2385 ();
 sg13g2_decap_8 FILLER_21_2392 ();
 sg13g2_fill_2 FILLER_21_2399 ();
 sg13g2_fill_1 FILLER_21_2401 ();
 sg13g2_fill_2 FILLER_21_2433 ();
 sg13g2_fill_1 FILLER_21_2435 ();
 sg13g2_fill_2 FILLER_21_2444 ();
 sg13g2_decap_8 FILLER_21_2472 ();
 sg13g2_decap_8 FILLER_21_2479 ();
 sg13g2_decap_8 FILLER_21_2486 ();
 sg13g2_decap_8 FILLER_21_2493 ();
 sg13g2_fill_1 FILLER_21_2500 ();
 sg13g2_fill_2 FILLER_21_2558 ();
 sg13g2_fill_1 FILLER_21_2560 ();
 sg13g2_fill_2 FILLER_21_2587 ();
 sg13g2_decap_8 FILLER_21_2628 ();
 sg13g2_decap_8 FILLER_21_2635 ();
 sg13g2_decap_8 FILLER_21_2642 ();
 sg13g2_decap_8 FILLER_21_2649 ();
 sg13g2_decap_8 FILLER_21_2656 ();
 sg13g2_fill_1 FILLER_21_2663 ();
 sg13g2_decap_4 FILLER_21_2716 ();
 sg13g2_fill_2 FILLER_21_2720 ();
 sg13g2_decap_8 FILLER_21_2726 ();
 sg13g2_decap_8 FILLER_21_2733 ();
 sg13g2_decap_8 FILLER_21_2740 ();
 sg13g2_decap_8 FILLER_21_2747 ();
 sg13g2_decap_8 FILLER_21_2754 ();
 sg13g2_decap_8 FILLER_21_2761 ();
 sg13g2_decap_8 FILLER_21_2768 ();
 sg13g2_decap_8 FILLER_21_2775 ();
 sg13g2_decap_8 FILLER_21_2782 ();
 sg13g2_decap_8 FILLER_21_2789 ();
 sg13g2_decap_8 FILLER_21_2796 ();
 sg13g2_decap_8 FILLER_21_2803 ();
 sg13g2_decap_8 FILLER_21_2810 ();
 sg13g2_decap_8 FILLER_21_2817 ();
 sg13g2_decap_8 FILLER_21_2824 ();
 sg13g2_decap_8 FILLER_21_2831 ();
 sg13g2_decap_8 FILLER_21_2838 ();
 sg13g2_decap_8 FILLER_21_2845 ();
 sg13g2_decap_8 FILLER_21_2852 ();
 sg13g2_decap_8 FILLER_21_2859 ();
 sg13g2_decap_8 FILLER_21_2866 ();
 sg13g2_decap_8 FILLER_21_2873 ();
 sg13g2_decap_8 FILLER_21_2880 ();
 sg13g2_decap_8 FILLER_21_2887 ();
 sg13g2_decap_8 FILLER_21_2894 ();
 sg13g2_decap_8 FILLER_21_2901 ();
 sg13g2_decap_8 FILLER_21_2908 ();
 sg13g2_decap_8 FILLER_21_2915 ();
 sg13g2_decap_8 FILLER_21_2922 ();
 sg13g2_decap_8 FILLER_21_2929 ();
 sg13g2_decap_8 FILLER_21_2936 ();
 sg13g2_decap_8 FILLER_21_2943 ();
 sg13g2_decap_8 FILLER_21_2950 ();
 sg13g2_decap_8 FILLER_21_2957 ();
 sg13g2_decap_8 FILLER_21_2964 ();
 sg13g2_decap_8 FILLER_21_2971 ();
 sg13g2_decap_8 FILLER_21_2978 ();
 sg13g2_decap_8 FILLER_21_2985 ();
 sg13g2_decap_8 FILLER_21_2992 ();
 sg13g2_decap_8 FILLER_21_2999 ();
 sg13g2_decap_8 FILLER_21_3006 ();
 sg13g2_decap_8 FILLER_21_3013 ();
 sg13g2_decap_8 FILLER_21_3020 ();
 sg13g2_decap_8 FILLER_21_3027 ();
 sg13g2_decap_8 FILLER_21_3034 ();
 sg13g2_decap_8 FILLER_21_3041 ();
 sg13g2_decap_8 FILLER_21_3048 ();
 sg13g2_decap_8 FILLER_21_3055 ();
 sg13g2_decap_8 FILLER_21_3062 ();
 sg13g2_decap_8 FILLER_21_3069 ();
 sg13g2_decap_8 FILLER_21_3076 ();
 sg13g2_decap_8 FILLER_21_3083 ();
 sg13g2_decap_8 FILLER_21_3090 ();
 sg13g2_decap_8 FILLER_21_3097 ();
 sg13g2_decap_8 FILLER_21_3104 ();
 sg13g2_decap_8 FILLER_21_3111 ();
 sg13g2_decap_8 FILLER_21_3118 ();
 sg13g2_decap_8 FILLER_21_3125 ();
 sg13g2_decap_8 FILLER_21_3132 ();
 sg13g2_decap_8 FILLER_21_3139 ();
 sg13g2_decap_8 FILLER_21_3146 ();
 sg13g2_decap_8 FILLER_21_3153 ();
 sg13g2_decap_8 FILLER_21_3160 ();
 sg13g2_decap_8 FILLER_21_3167 ();
 sg13g2_decap_8 FILLER_21_3174 ();
 sg13g2_decap_8 FILLER_21_3181 ();
 sg13g2_decap_8 FILLER_21_3188 ();
 sg13g2_decap_8 FILLER_21_3195 ();
 sg13g2_decap_8 FILLER_21_3202 ();
 sg13g2_decap_8 FILLER_21_3209 ();
 sg13g2_decap_8 FILLER_21_3216 ();
 sg13g2_decap_8 FILLER_21_3223 ();
 sg13g2_decap_8 FILLER_21_3230 ();
 sg13g2_decap_8 FILLER_21_3237 ();
 sg13g2_decap_8 FILLER_21_3244 ();
 sg13g2_decap_8 FILLER_21_3251 ();
 sg13g2_decap_8 FILLER_21_3258 ();
 sg13g2_decap_8 FILLER_21_3265 ();
 sg13g2_decap_8 FILLER_21_3272 ();
 sg13g2_decap_8 FILLER_21_3279 ();
 sg13g2_decap_8 FILLER_21_3286 ();
 sg13g2_decap_8 FILLER_21_3293 ();
 sg13g2_decap_8 FILLER_21_3300 ();
 sg13g2_decap_8 FILLER_21_3307 ();
 sg13g2_decap_8 FILLER_21_3314 ();
 sg13g2_decap_8 FILLER_21_3321 ();
 sg13g2_decap_8 FILLER_21_3328 ();
 sg13g2_decap_8 FILLER_21_3335 ();
 sg13g2_decap_8 FILLER_21_3342 ();
 sg13g2_decap_8 FILLER_21_3349 ();
 sg13g2_decap_8 FILLER_21_3356 ();
 sg13g2_decap_8 FILLER_21_3363 ();
 sg13g2_decap_8 FILLER_21_3370 ();
 sg13g2_decap_8 FILLER_21_3377 ();
 sg13g2_decap_8 FILLER_21_3384 ();
 sg13g2_decap_8 FILLER_21_3391 ();
 sg13g2_decap_8 FILLER_21_3398 ();
 sg13g2_decap_8 FILLER_21_3405 ();
 sg13g2_decap_8 FILLER_21_3412 ();
 sg13g2_decap_8 FILLER_21_3419 ();
 sg13g2_decap_8 FILLER_21_3426 ();
 sg13g2_decap_8 FILLER_21_3433 ();
 sg13g2_decap_8 FILLER_21_3440 ();
 sg13g2_decap_8 FILLER_21_3447 ();
 sg13g2_decap_8 FILLER_21_3454 ();
 sg13g2_decap_8 FILLER_21_3461 ();
 sg13g2_decap_8 FILLER_21_3468 ();
 sg13g2_decap_8 FILLER_21_3475 ();
 sg13g2_decap_8 FILLER_21_3482 ();
 sg13g2_decap_8 FILLER_21_3489 ();
 sg13g2_decap_8 FILLER_21_3496 ();
 sg13g2_decap_8 FILLER_21_3503 ();
 sg13g2_decap_8 FILLER_21_3510 ();
 sg13g2_decap_8 FILLER_21_3517 ();
 sg13g2_decap_8 FILLER_21_3524 ();
 sg13g2_decap_8 FILLER_21_3531 ();
 sg13g2_decap_8 FILLER_21_3538 ();
 sg13g2_decap_8 FILLER_21_3545 ();
 sg13g2_decap_8 FILLER_21_3552 ();
 sg13g2_decap_8 FILLER_21_3559 ();
 sg13g2_decap_8 FILLER_21_3566 ();
 sg13g2_decap_8 FILLER_21_3573 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_73 ();
 sg13g2_decap_8 FILLER_22_80 ();
 sg13g2_decap_8 FILLER_22_87 ();
 sg13g2_fill_2 FILLER_22_94 ();
 sg13g2_fill_1 FILLER_22_111 ();
 sg13g2_decap_8 FILLER_22_146 ();
 sg13g2_decap_8 FILLER_22_153 ();
 sg13g2_decap_8 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_decap_4 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_decap_8 FILLER_22_251 ();
 sg13g2_decap_8 FILLER_22_258 ();
 sg13g2_decap_4 FILLER_22_265 ();
 sg13g2_fill_2 FILLER_22_295 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_fill_2 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_353 ();
 sg13g2_fill_2 FILLER_22_360 ();
 sg13g2_fill_1 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_452 ();
 sg13g2_fill_2 FILLER_22_485 ();
 sg13g2_fill_1 FILLER_22_487 ();
 sg13g2_decap_8 FILLER_22_506 ();
 sg13g2_decap_8 FILLER_22_513 ();
 sg13g2_fill_1 FILLER_22_520 ();
 sg13g2_decap_4 FILLER_22_551 ();
 sg13g2_fill_1 FILLER_22_555 ();
 sg13g2_fill_1 FILLER_22_569 ();
 sg13g2_decap_8 FILLER_22_596 ();
 sg13g2_decap_4 FILLER_22_603 ();
 sg13g2_decap_8 FILLER_22_633 ();
 sg13g2_fill_2 FILLER_22_640 ();
 sg13g2_fill_2 FILLER_22_652 ();
 sg13g2_decap_8 FILLER_22_680 ();
 sg13g2_decap_4 FILLER_22_687 ();
 sg13g2_decap_8 FILLER_22_696 ();
 sg13g2_fill_2 FILLER_22_703 ();
 sg13g2_fill_2 FILLER_22_770 ();
 sg13g2_decap_4 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_811 ();
 sg13g2_decap_8 FILLER_22_818 ();
 sg13g2_decap_8 FILLER_22_825 ();
 sg13g2_decap_8 FILLER_22_832 ();
 sg13g2_fill_2 FILLER_22_839 ();
 sg13g2_fill_1 FILLER_22_841 ();
 sg13g2_fill_2 FILLER_22_856 ();
 sg13g2_fill_1 FILLER_22_869 ();
 sg13g2_fill_1 FILLER_22_879 ();
 sg13g2_decap_8 FILLER_22_893 ();
 sg13g2_decap_8 FILLER_22_903 ();
 sg13g2_decap_4 FILLER_22_910 ();
 sg13g2_fill_1 FILLER_22_914 ();
 sg13g2_decap_8 FILLER_22_919 ();
 sg13g2_decap_4 FILLER_22_956 ();
 sg13g2_fill_1 FILLER_22_960 ();
 sg13g2_decap_8 FILLER_22_1059 ();
 sg13g2_decap_4 FILLER_22_1066 ();
 sg13g2_fill_1 FILLER_22_1070 ();
 sg13g2_decap_8 FILLER_22_1103 ();
 sg13g2_decap_8 FILLER_22_1110 ();
 sg13g2_decap_8 FILLER_22_1117 ();
 sg13g2_fill_2 FILLER_22_1124 ();
 sg13g2_fill_1 FILLER_22_1126 ();
 sg13g2_decap_8 FILLER_22_1165 ();
 sg13g2_decap_4 FILLER_22_1172 ();
 sg13g2_decap_8 FILLER_22_1220 ();
 sg13g2_decap_8 FILLER_22_1227 ();
 sg13g2_decap_8 FILLER_22_1234 ();
 sg13g2_fill_2 FILLER_22_1241 ();
 sg13g2_fill_1 FILLER_22_1243 ();
 sg13g2_fill_2 FILLER_22_1258 ();
 sg13g2_fill_1 FILLER_22_1260 ();
 sg13g2_decap_8 FILLER_22_1287 ();
 sg13g2_decap_4 FILLER_22_1294 ();
 sg13g2_decap_8 FILLER_22_1306 ();
 sg13g2_decap_4 FILLER_22_1313 ();
 sg13g2_fill_2 FILLER_22_1338 ();
 sg13g2_fill_2 FILLER_22_1350 ();
 sg13g2_fill_1 FILLER_22_1352 ();
 sg13g2_fill_1 FILLER_22_1362 ();
 sg13g2_decap_8 FILLER_22_1368 ();
 sg13g2_fill_2 FILLER_22_1375 ();
 sg13g2_fill_1 FILLER_22_1377 ();
 sg13g2_fill_1 FILLER_22_1388 ();
 sg13g2_decap_4 FILLER_22_1397 ();
 sg13g2_fill_1 FILLER_22_1401 ();
 sg13g2_decap_4 FILLER_22_1407 ();
 sg13g2_fill_2 FILLER_22_1411 ();
 sg13g2_fill_2 FILLER_22_1421 ();
 sg13g2_fill_1 FILLER_22_1423 ();
 sg13g2_fill_1 FILLER_22_1434 ();
 sg13g2_decap_8 FILLER_22_1450 ();
 sg13g2_decap_8 FILLER_22_1457 ();
 sg13g2_fill_2 FILLER_22_1464 ();
 sg13g2_fill_1 FILLER_22_1466 ();
 sg13g2_decap_4 FILLER_22_1519 ();
 sg13g2_decap_8 FILLER_22_1536 ();
 sg13g2_decap_4 FILLER_22_1543 ();
 sg13g2_decap_8 FILLER_22_1551 ();
 sg13g2_decap_8 FILLER_22_1558 ();
 sg13g2_fill_1 FILLER_22_1565 ();
 sg13g2_decap_8 FILLER_22_1602 ();
 sg13g2_decap_8 FILLER_22_1609 ();
 sg13g2_fill_2 FILLER_22_1616 ();
 sg13g2_decap_4 FILLER_22_1622 ();
 sg13g2_decap_8 FILLER_22_1655 ();
 sg13g2_fill_2 FILLER_22_1662 ();
 sg13g2_fill_1 FILLER_22_1664 ();
 sg13g2_fill_2 FILLER_22_1691 ();
 sg13g2_fill_2 FILLER_22_1724 ();
 sg13g2_decap_4 FILLER_22_1739 ();
 sg13g2_fill_2 FILLER_22_1743 ();
 sg13g2_decap_8 FILLER_22_1819 ();
 sg13g2_decap_8 FILLER_22_1826 ();
 sg13g2_fill_2 FILLER_22_1859 ();
 sg13g2_decap_4 FILLER_22_1938 ();
 sg13g2_fill_2 FILLER_22_1942 ();
 sg13g2_fill_2 FILLER_22_1947 ();
 sg13g2_fill_1 FILLER_22_1967 ();
 sg13g2_decap_8 FILLER_22_1994 ();
 sg13g2_decap_8 FILLER_22_2001 ();
 sg13g2_fill_2 FILLER_22_2008 ();
 sg13g2_fill_1 FILLER_22_2010 ();
 sg13g2_decap_8 FILLER_22_2037 ();
 sg13g2_decap_8 FILLER_22_2044 ();
 sg13g2_decap_8 FILLER_22_2051 ();
 sg13g2_decap_4 FILLER_22_2058 ();
 sg13g2_fill_1 FILLER_22_2062 ();
 sg13g2_decap_8 FILLER_22_2115 ();
 sg13g2_decap_8 FILLER_22_2122 ();
 sg13g2_decap_4 FILLER_22_2129 ();
 sg13g2_decap_4 FILLER_22_2164 ();
 sg13g2_fill_1 FILLER_22_2168 ();
 sg13g2_fill_1 FILLER_22_2173 ();
 sg13g2_fill_1 FILLER_22_2231 ();
 sg13g2_decap_8 FILLER_22_2271 ();
 sg13g2_decap_8 FILLER_22_2278 ();
 sg13g2_decap_8 FILLER_22_2285 ();
 sg13g2_decap_4 FILLER_22_2292 ();
 sg13g2_fill_1 FILLER_22_2296 ();
 sg13g2_fill_1 FILLER_22_2302 ();
 sg13g2_decap_8 FILLER_22_2310 ();
 sg13g2_decap_8 FILLER_22_2317 ();
 sg13g2_decap_8 FILLER_22_2324 ();
 sg13g2_decap_8 FILLER_22_2331 ();
 sg13g2_decap_8 FILLER_22_2390 ();
 sg13g2_decap_8 FILLER_22_2483 ();
 sg13g2_decap_4 FILLER_22_2490 ();
 sg13g2_decap_8 FILLER_22_2528 ();
 sg13g2_fill_1 FILLER_22_2535 ();
 sg13g2_decap_8 FILLER_22_2562 ();
 sg13g2_decap_8 FILLER_22_2569 ();
 sg13g2_decap_8 FILLER_22_2576 ();
 sg13g2_fill_2 FILLER_22_2583 ();
 sg13g2_fill_1 FILLER_22_2585 ();
 sg13g2_fill_2 FILLER_22_2624 ();
 sg13g2_decap_8 FILLER_22_2630 ();
 sg13g2_decap_8 FILLER_22_2663 ();
 sg13g2_fill_2 FILLER_22_2670 ();
 sg13g2_fill_1 FILLER_22_2672 ();
 sg13g2_fill_1 FILLER_22_2678 ();
 sg13g2_decap_8 FILLER_22_2705 ();
 sg13g2_decap_8 FILLER_22_2712 ();
 sg13g2_decap_8 FILLER_22_2719 ();
 sg13g2_decap_8 FILLER_22_2726 ();
 sg13g2_decap_8 FILLER_22_2733 ();
 sg13g2_decap_8 FILLER_22_2740 ();
 sg13g2_decap_8 FILLER_22_2747 ();
 sg13g2_decap_8 FILLER_22_2754 ();
 sg13g2_decap_8 FILLER_22_2761 ();
 sg13g2_decap_8 FILLER_22_2768 ();
 sg13g2_decap_8 FILLER_22_2775 ();
 sg13g2_decap_8 FILLER_22_2782 ();
 sg13g2_decap_8 FILLER_22_2789 ();
 sg13g2_decap_8 FILLER_22_2796 ();
 sg13g2_decap_8 FILLER_22_2803 ();
 sg13g2_decap_8 FILLER_22_2810 ();
 sg13g2_decap_8 FILLER_22_2817 ();
 sg13g2_decap_8 FILLER_22_2824 ();
 sg13g2_decap_8 FILLER_22_2831 ();
 sg13g2_fill_2 FILLER_22_2838 ();
 sg13g2_decap_8 FILLER_22_2866 ();
 sg13g2_decap_8 FILLER_22_2873 ();
 sg13g2_decap_8 FILLER_22_2880 ();
 sg13g2_decap_8 FILLER_22_2887 ();
 sg13g2_decap_8 FILLER_22_2894 ();
 sg13g2_decap_4 FILLER_22_2901 ();
 sg13g2_fill_1 FILLER_22_2910 ();
 sg13g2_decap_8 FILLER_22_2921 ();
 sg13g2_decap_8 FILLER_22_2928 ();
 sg13g2_decap_8 FILLER_22_2935 ();
 sg13g2_decap_8 FILLER_22_2942 ();
 sg13g2_decap_8 FILLER_22_2949 ();
 sg13g2_decap_8 FILLER_22_2956 ();
 sg13g2_decap_8 FILLER_22_2963 ();
 sg13g2_decap_8 FILLER_22_2970 ();
 sg13g2_decap_8 FILLER_22_2977 ();
 sg13g2_decap_8 FILLER_22_2984 ();
 sg13g2_decap_8 FILLER_22_2991 ();
 sg13g2_decap_8 FILLER_22_2998 ();
 sg13g2_decap_8 FILLER_22_3005 ();
 sg13g2_decap_8 FILLER_22_3012 ();
 sg13g2_decap_8 FILLER_22_3019 ();
 sg13g2_decap_8 FILLER_22_3026 ();
 sg13g2_decap_8 FILLER_22_3033 ();
 sg13g2_decap_8 FILLER_22_3040 ();
 sg13g2_decap_8 FILLER_22_3047 ();
 sg13g2_decap_8 FILLER_22_3054 ();
 sg13g2_decap_8 FILLER_22_3061 ();
 sg13g2_decap_8 FILLER_22_3068 ();
 sg13g2_decap_8 FILLER_22_3075 ();
 sg13g2_decap_8 FILLER_22_3082 ();
 sg13g2_decap_8 FILLER_22_3089 ();
 sg13g2_decap_8 FILLER_22_3096 ();
 sg13g2_decap_8 FILLER_22_3103 ();
 sg13g2_decap_8 FILLER_22_3110 ();
 sg13g2_decap_8 FILLER_22_3117 ();
 sg13g2_decap_8 FILLER_22_3124 ();
 sg13g2_decap_8 FILLER_22_3131 ();
 sg13g2_decap_8 FILLER_22_3138 ();
 sg13g2_decap_8 FILLER_22_3145 ();
 sg13g2_decap_8 FILLER_22_3152 ();
 sg13g2_decap_8 FILLER_22_3159 ();
 sg13g2_decap_8 FILLER_22_3166 ();
 sg13g2_decap_8 FILLER_22_3173 ();
 sg13g2_decap_8 FILLER_22_3180 ();
 sg13g2_decap_8 FILLER_22_3187 ();
 sg13g2_decap_8 FILLER_22_3194 ();
 sg13g2_decap_8 FILLER_22_3201 ();
 sg13g2_decap_8 FILLER_22_3208 ();
 sg13g2_decap_8 FILLER_22_3215 ();
 sg13g2_decap_8 FILLER_22_3222 ();
 sg13g2_decap_8 FILLER_22_3229 ();
 sg13g2_decap_8 FILLER_22_3236 ();
 sg13g2_decap_8 FILLER_22_3243 ();
 sg13g2_decap_8 FILLER_22_3250 ();
 sg13g2_decap_8 FILLER_22_3257 ();
 sg13g2_decap_8 FILLER_22_3264 ();
 sg13g2_decap_8 FILLER_22_3271 ();
 sg13g2_decap_8 FILLER_22_3278 ();
 sg13g2_decap_8 FILLER_22_3285 ();
 sg13g2_decap_8 FILLER_22_3292 ();
 sg13g2_decap_8 FILLER_22_3299 ();
 sg13g2_decap_8 FILLER_22_3306 ();
 sg13g2_decap_8 FILLER_22_3313 ();
 sg13g2_decap_8 FILLER_22_3320 ();
 sg13g2_decap_8 FILLER_22_3327 ();
 sg13g2_decap_8 FILLER_22_3334 ();
 sg13g2_decap_8 FILLER_22_3341 ();
 sg13g2_decap_8 FILLER_22_3348 ();
 sg13g2_decap_8 FILLER_22_3355 ();
 sg13g2_decap_8 FILLER_22_3362 ();
 sg13g2_decap_8 FILLER_22_3369 ();
 sg13g2_decap_8 FILLER_22_3376 ();
 sg13g2_decap_8 FILLER_22_3383 ();
 sg13g2_decap_8 FILLER_22_3390 ();
 sg13g2_decap_8 FILLER_22_3397 ();
 sg13g2_decap_8 FILLER_22_3404 ();
 sg13g2_decap_8 FILLER_22_3411 ();
 sg13g2_decap_8 FILLER_22_3418 ();
 sg13g2_decap_8 FILLER_22_3425 ();
 sg13g2_decap_8 FILLER_22_3432 ();
 sg13g2_decap_8 FILLER_22_3439 ();
 sg13g2_decap_8 FILLER_22_3446 ();
 sg13g2_decap_8 FILLER_22_3453 ();
 sg13g2_decap_8 FILLER_22_3460 ();
 sg13g2_decap_8 FILLER_22_3467 ();
 sg13g2_decap_8 FILLER_22_3474 ();
 sg13g2_decap_8 FILLER_22_3481 ();
 sg13g2_decap_8 FILLER_22_3488 ();
 sg13g2_decap_8 FILLER_22_3495 ();
 sg13g2_decap_8 FILLER_22_3502 ();
 sg13g2_decap_8 FILLER_22_3509 ();
 sg13g2_decap_8 FILLER_22_3516 ();
 sg13g2_decap_8 FILLER_22_3523 ();
 sg13g2_decap_8 FILLER_22_3530 ();
 sg13g2_decap_8 FILLER_22_3537 ();
 sg13g2_decap_8 FILLER_22_3544 ();
 sg13g2_decap_8 FILLER_22_3551 ();
 sg13g2_decap_8 FILLER_22_3558 ();
 sg13g2_decap_8 FILLER_22_3565 ();
 sg13g2_decap_8 FILLER_22_3572 ();
 sg13g2_fill_1 FILLER_22_3579 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_37 ();
 sg13g2_decap_8 FILLER_23_64 ();
 sg13g2_decap_8 FILLER_23_71 ();
 sg13g2_decap_8 FILLER_23_78 ();
 sg13g2_decap_8 FILLER_23_85 ();
 sg13g2_decap_8 FILLER_23_92 ();
 sg13g2_decap_8 FILLER_23_99 ();
 sg13g2_fill_2 FILLER_23_106 ();
 sg13g2_fill_2 FILLER_23_136 ();
 sg13g2_decap_8 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_202 ();
 sg13g2_decap_8 FILLER_23_209 ();
 sg13g2_fill_2 FILLER_23_216 ();
 sg13g2_fill_1 FILLER_23_218 ();
 sg13g2_fill_2 FILLER_23_222 ();
 sg13g2_decap_8 FILLER_23_250 ();
 sg13g2_decap_8 FILLER_23_257 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_fill_2 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_fill_2 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_decap_4 FILLER_23_358 ();
 sg13g2_fill_2 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_fill_2 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_482 ();
 sg13g2_decap_8 FILLER_23_509 ();
 sg13g2_decap_8 FILLER_23_516 ();
 sg13g2_fill_2 FILLER_23_523 ();
 sg13g2_fill_1 FILLER_23_525 ();
 sg13g2_fill_1 FILLER_23_534 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_fill_2 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_4 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_decap_8 FILLER_23_690 ();
 sg13g2_decap_4 FILLER_23_697 ();
 sg13g2_fill_2 FILLER_23_730 ();
 sg13g2_decap_4 FILLER_23_736 ();
 sg13g2_fill_2 FILLER_23_740 ();
 sg13g2_decap_8 FILLER_23_746 ();
 sg13g2_fill_1 FILLER_23_753 ();
 sg13g2_fill_1 FILLER_23_762 ();
 sg13g2_decap_8 FILLER_23_766 ();
 sg13g2_fill_2 FILLER_23_773 ();
 sg13g2_fill_1 FILLER_23_775 ();
 sg13g2_decap_8 FILLER_23_780 ();
 sg13g2_decap_4 FILLER_23_787 ();
 sg13g2_fill_1 FILLER_23_791 ();
 sg13g2_decap_4 FILLER_23_796 ();
 sg13g2_fill_2 FILLER_23_800 ();
 sg13g2_fill_2 FILLER_23_828 ();
 sg13g2_fill_1 FILLER_23_860 ();
 sg13g2_decap_4 FILLER_23_887 ();
 sg13g2_decap_8 FILLER_23_904 ();
 sg13g2_fill_2 FILLER_23_911 ();
 sg13g2_decap_4 FILLER_23_920 ();
 sg13g2_decap_8 FILLER_23_932 ();
 sg13g2_decap_8 FILLER_23_939 ();
 sg13g2_decap_8 FILLER_23_946 ();
 sg13g2_decap_8 FILLER_23_953 ();
 sg13g2_decap_4 FILLER_23_960 ();
 sg13g2_fill_2 FILLER_23_964 ();
 sg13g2_decap_8 FILLER_23_1000 ();
 sg13g2_decap_8 FILLER_23_1007 ();
 sg13g2_decap_8 FILLER_23_1014 ();
 sg13g2_decap_4 FILLER_23_1021 ();
 sg13g2_decap_8 FILLER_23_1051 ();
 sg13g2_decap_8 FILLER_23_1058 ();
 sg13g2_decap_8 FILLER_23_1065 ();
 sg13g2_decap_8 FILLER_23_1072 ();
 sg13g2_decap_4 FILLER_23_1079 ();
 sg13g2_fill_1 FILLER_23_1083 ();
 sg13g2_fill_2 FILLER_23_1092 ();
 sg13g2_fill_2 FILLER_23_1130 ();
 sg13g2_fill_1 FILLER_23_1164 ();
 sg13g2_decap_8 FILLER_23_1177 ();
 sg13g2_decap_8 FILLER_23_1218 ();
 sg13g2_decap_8 FILLER_23_1225 ();
 sg13g2_fill_1 FILLER_23_1232 ();
 sg13g2_fill_2 FILLER_23_1236 ();
 sg13g2_fill_1 FILLER_23_1238 ();
 sg13g2_decap_4 FILLER_23_1242 ();
 sg13g2_fill_2 FILLER_23_1246 ();
 sg13g2_fill_2 FILLER_23_1253 ();
 sg13g2_decap_4 FILLER_23_1258 ();
 sg13g2_fill_1 FILLER_23_1262 ();
 sg13g2_decap_4 FILLER_23_1292 ();
 sg13g2_fill_2 FILLER_23_1296 ();
 sg13g2_decap_8 FILLER_23_1302 ();
 sg13g2_fill_2 FILLER_23_1369 ();
 sg13g2_decap_4 FILLER_23_1397 ();
 sg13g2_fill_2 FILLER_23_1401 ();
 sg13g2_decap_4 FILLER_23_1429 ();
 sg13g2_decap_4 FILLER_23_1459 ();
 sg13g2_fill_2 FILLER_23_1463 ();
 sg13g2_fill_2 FILLER_23_1491 ();
 sg13g2_decap_4 FILLER_23_1532 ();
 sg13g2_fill_1 FILLER_23_1562 ();
 sg13g2_fill_1 FILLER_23_1607 ();
 sg13g2_decap_4 FILLER_23_1613 ();
 sg13g2_fill_1 FILLER_23_1617 ();
 sg13g2_fill_1 FILLER_23_1651 ();
 sg13g2_decap_8 FILLER_23_1682 ();
 sg13g2_fill_2 FILLER_23_1692 ();
 sg13g2_fill_1 FILLER_23_1701 ();
 sg13g2_decap_8 FILLER_23_1737 ();
 sg13g2_fill_2 FILLER_23_1744 ();
 sg13g2_fill_1 FILLER_23_1746 ();
 sg13g2_decap_8 FILLER_23_1778 ();
 sg13g2_fill_2 FILLER_23_1785 ();
 sg13g2_fill_1 FILLER_23_1813 ();
 sg13g2_fill_2 FILLER_23_1822 ();
 sg13g2_fill_2 FILLER_23_1827 ();
 sg13g2_fill_1 FILLER_23_1829 ();
 sg13g2_fill_1 FILLER_23_1870 ();
 sg13g2_fill_2 FILLER_23_1945 ();
 sg13g2_fill_1 FILLER_23_1947 ();
 sg13g2_decap_8 FILLER_23_1993 ();
 sg13g2_decap_4 FILLER_23_2000 ();
 sg13g2_fill_2 FILLER_23_2069 ();
 sg13g2_fill_1 FILLER_23_2071 ();
 sg13g2_decap_8 FILLER_23_2118 ();
 sg13g2_decap_8 FILLER_23_2125 ();
 sg13g2_fill_1 FILLER_23_2132 ();
 sg13g2_decap_8 FILLER_23_2168 ();
 sg13g2_decap_4 FILLER_23_2175 ();
 sg13g2_fill_2 FILLER_23_2179 ();
 sg13g2_decap_4 FILLER_23_2238 ();
 sg13g2_decap_8 FILLER_23_2268 ();
 sg13g2_fill_2 FILLER_23_2275 ();
 sg13g2_decap_8 FILLER_23_2306 ();
 sg13g2_decap_8 FILLER_23_2313 ();
 sg13g2_decap_8 FILLER_23_2320 ();
 sg13g2_fill_1 FILLER_23_2327 ();
 sg13g2_decap_8 FILLER_23_2479 ();
 sg13g2_decap_8 FILLER_23_2486 ();
 sg13g2_decap_8 FILLER_23_2493 ();
 sg13g2_decap_4 FILLER_23_2500 ();
 sg13g2_fill_1 FILLER_23_2504 ();
 sg13g2_decap_8 FILLER_23_2583 ();
 sg13g2_decap_8 FILLER_23_2590 ();
 sg13g2_fill_2 FILLER_23_2597 ();
 sg13g2_fill_1 FILLER_23_2599 ();
 sg13g2_decap_8 FILLER_23_2605 ();
 sg13g2_decap_8 FILLER_23_2661 ();
 sg13g2_decap_4 FILLER_23_2668 ();
 sg13g2_fill_2 FILLER_23_2672 ();
 sg13g2_decap_8 FILLER_23_2708 ();
 sg13g2_decap_8 FILLER_23_2715 ();
 sg13g2_decap_8 FILLER_23_2722 ();
 sg13g2_decap_8 FILLER_23_2729 ();
 sg13g2_decap_8 FILLER_23_2736 ();
 sg13g2_decap_8 FILLER_23_2743 ();
 sg13g2_decap_8 FILLER_23_2750 ();
 sg13g2_decap_8 FILLER_23_2757 ();
 sg13g2_decap_8 FILLER_23_2764 ();
 sg13g2_decap_8 FILLER_23_2771 ();
 sg13g2_decap_8 FILLER_23_2778 ();
 sg13g2_decap_8 FILLER_23_2785 ();
 sg13g2_decap_8 FILLER_23_2792 ();
 sg13g2_decap_8 FILLER_23_2799 ();
 sg13g2_decap_8 FILLER_23_2806 ();
 sg13g2_decap_8 FILLER_23_2813 ();
 sg13g2_decap_4 FILLER_23_2820 ();
 sg13g2_fill_2 FILLER_23_2824 ();
 sg13g2_decap_4 FILLER_23_2834 ();
 sg13g2_fill_1 FILLER_23_2838 ();
 sg13g2_decap_8 FILLER_23_2878 ();
 sg13g2_decap_8 FILLER_23_2885 ();
 sg13g2_decap_4 FILLER_23_2892 ();
 sg13g2_fill_1 FILLER_23_2896 ();
 sg13g2_decap_8 FILLER_23_2930 ();
 sg13g2_decap_8 FILLER_23_2937 ();
 sg13g2_decap_8 FILLER_23_2944 ();
 sg13g2_fill_2 FILLER_23_2951 ();
 sg13g2_fill_1 FILLER_23_2953 ();
 sg13g2_decap_8 FILLER_23_2962 ();
 sg13g2_decap_8 FILLER_23_2969 ();
 sg13g2_decap_8 FILLER_23_2976 ();
 sg13g2_decap_8 FILLER_23_2983 ();
 sg13g2_decap_8 FILLER_23_2990 ();
 sg13g2_decap_8 FILLER_23_2997 ();
 sg13g2_decap_4 FILLER_23_3004 ();
 sg13g2_decap_8 FILLER_23_3013 ();
 sg13g2_decap_8 FILLER_23_3020 ();
 sg13g2_decap_8 FILLER_23_3027 ();
 sg13g2_decap_8 FILLER_23_3034 ();
 sg13g2_decap_8 FILLER_23_3041 ();
 sg13g2_decap_8 FILLER_23_3048 ();
 sg13g2_decap_8 FILLER_23_3083 ();
 sg13g2_decap_8 FILLER_23_3090 ();
 sg13g2_decap_8 FILLER_23_3097 ();
 sg13g2_decap_8 FILLER_23_3104 ();
 sg13g2_decap_8 FILLER_23_3111 ();
 sg13g2_decap_8 FILLER_23_3118 ();
 sg13g2_decap_8 FILLER_23_3125 ();
 sg13g2_decap_8 FILLER_23_3132 ();
 sg13g2_decap_8 FILLER_23_3139 ();
 sg13g2_decap_8 FILLER_23_3146 ();
 sg13g2_decap_8 FILLER_23_3153 ();
 sg13g2_decap_8 FILLER_23_3160 ();
 sg13g2_decap_8 FILLER_23_3167 ();
 sg13g2_decap_8 FILLER_23_3174 ();
 sg13g2_decap_8 FILLER_23_3181 ();
 sg13g2_decap_8 FILLER_23_3188 ();
 sg13g2_decap_8 FILLER_23_3195 ();
 sg13g2_decap_8 FILLER_23_3202 ();
 sg13g2_decap_8 FILLER_23_3209 ();
 sg13g2_decap_8 FILLER_23_3216 ();
 sg13g2_decap_8 FILLER_23_3223 ();
 sg13g2_decap_8 FILLER_23_3230 ();
 sg13g2_decap_8 FILLER_23_3237 ();
 sg13g2_decap_8 FILLER_23_3244 ();
 sg13g2_decap_8 FILLER_23_3251 ();
 sg13g2_decap_8 FILLER_23_3258 ();
 sg13g2_decap_8 FILLER_23_3265 ();
 sg13g2_decap_8 FILLER_23_3272 ();
 sg13g2_decap_8 FILLER_23_3279 ();
 sg13g2_decap_8 FILLER_23_3286 ();
 sg13g2_decap_8 FILLER_23_3293 ();
 sg13g2_decap_8 FILLER_23_3300 ();
 sg13g2_decap_8 FILLER_23_3307 ();
 sg13g2_decap_8 FILLER_23_3314 ();
 sg13g2_decap_8 FILLER_23_3321 ();
 sg13g2_decap_8 FILLER_23_3328 ();
 sg13g2_decap_8 FILLER_23_3335 ();
 sg13g2_decap_8 FILLER_23_3342 ();
 sg13g2_decap_8 FILLER_23_3349 ();
 sg13g2_decap_8 FILLER_23_3356 ();
 sg13g2_decap_8 FILLER_23_3363 ();
 sg13g2_decap_8 FILLER_23_3370 ();
 sg13g2_decap_8 FILLER_23_3377 ();
 sg13g2_decap_8 FILLER_23_3384 ();
 sg13g2_decap_8 FILLER_23_3391 ();
 sg13g2_decap_8 FILLER_23_3398 ();
 sg13g2_decap_8 FILLER_23_3405 ();
 sg13g2_decap_8 FILLER_23_3412 ();
 sg13g2_decap_8 FILLER_23_3419 ();
 sg13g2_decap_8 FILLER_23_3426 ();
 sg13g2_decap_8 FILLER_23_3433 ();
 sg13g2_decap_8 FILLER_23_3440 ();
 sg13g2_decap_8 FILLER_23_3447 ();
 sg13g2_decap_8 FILLER_23_3454 ();
 sg13g2_decap_8 FILLER_23_3461 ();
 sg13g2_decap_8 FILLER_23_3468 ();
 sg13g2_decap_8 FILLER_23_3475 ();
 sg13g2_decap_8 FILLER_23_3482 ();
 sg13g2_decap_8 FILLER_23_3489 ();
 sg13g2_decap_8 FILLER_23_3496 ();
 sg13g2_decap_8 FILLER_23_3503 ();
 sg13g2_decap_8 FILLER_23_3510 ();
 sg13g2_decap_8 FILLER_23_3517 ();
 sg13g2_decap_8 FILLER_23_3524 ();
 sg13g2_decap_8 FILLER_23_3531 ();
 sg13g2_decap_8 FILLER_23_3538 ();
 sg13g2_decap_8 FILLER_23_3545 ();
 sg13g2_decap_8 FILLER_23_3552 ();
 sg13g2_decap_8 FILLER_23_3559 ();
 sg13g2_decap_8 FILLER_23_3566 ();
 sg13g2_decap_8 FILLER_23_3573 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_decap_8 FILLER_24_90 ();
 sg13g2_decap_4 FILLER_24_97 ();
 sg13g2_fill_2 FILLER_24_101 ();
 sg13g2_decap_8 FILLER_24_142 ();
 sg13g2_fill_2 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_decap_8 FILLER_24_260 ();
 sg13g2_fill_2 FILLER_24_267 ();
 sg13g2_fill_1 FILLER_24_269 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_decap_4 FILLER_24_333 ();
 sg13g2_fill_2 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_4 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_475 ();
 sg13g2_fill_1 FILLER_24_477 ();
 sg13g2_fill_2 FILLER_24_506 ();
 sg13g2_decap_8 FILLER_24_534 ();
 sg13g2_decap_8 FILLER_24_541 ();
 sg13g2_fill_2 FILLER_24_548 ();
 sg13g2_decap_8 FILLER_24_671 ();
 sg13g2_decap_8 FILLER_24_678 ();
 sg13g2_decap_8 FILLER_24_685 ();
 sg13g2_decap_8 FILLER_24_692 ();
 sg13g2_decap_4 FILLER_24_699 ();
 sg13g2_fill_1 FILLER_24_703 ();
 sg13g2_fill_2 FILLER_24_709 ();
 sg13g2_fill_1 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_716 ();
 sg13g2_decap_8 FILLER_24_723 ();
 sg13g2_decap_8 FILLER_24_730 ();
 sg13g2_decap_8 FILLER_24_737 ();
 sg13g2_fill_2 FILLER_24_744 ();
 sg13g2_fill_1 FILLER_24_746 ();
 sg13g2_decap_8 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_758 ();
 sg13g2_decap_4 FILLER_24_791 ();
 sg13g2_fill_2 FILLER_24_847 ();
 sg13g2_fill_2 FILLER_24_870 ();
 sg13g2_fill_1 FILLER_24_876 ();
 sg13g2_fill_2 FILLER_24_885 ();
 sg13g2_decap_4 FILLER_24_944 ();
 sg13g2_fill_1 FILLER_24_948 ();
 sg13g2_fill_2 FILLER_24_959 ();
 sg13g2_decap_8 FILLER_24_1002 ();
 sg13g2_decap_8 FILLER_24_1009 ();
 sg13g2_decap_8 FILLER_24_1016 ();
 sg13g2_decap_8 FILLER_24_1023 ();
 sg13g2_decap_4 FILLER_24_1033 ();
 sg13g2_decap_8 FILLER_24_1063 ();
 sg13g2_decap_8 FILLER_24_1070 ();
 sg13g2_decap_8 FILLER_24_1103 ();
 sg13g2_fill_2 FILLER_24_1110 ();
 sg13g2_fill_1 FILLER_24_1164 ();
 sg13g2_fill_2 FILLER_24_1217 ();
 sg13g2_fill_1 FILLER_24_1219 ();
 sg13g2_fill_1 FILLER_24_1223 ();
 sg13g2_decap_4 FILLER_24_1257 ();
 sg13g2_fill_1 FILLER_24_1372 ();
 sg13g2_fill_2 FILLER_24_1393 ();
 sg13g2_fill_1 FILLER_24_1395 ();
 sg13g2_fill_2 FILLER_24_1448 ();
 sg13g2_fill_1 FILLER_24_1450 ();
 sg13g2_decap_8 FILLER_24_1459 ();
 sg13g2_decap_8 FILLER_24_1466 ();
 sg13g2_fill_2 FILLER_24_1473 ();
 sg13g2_fill_1 FILLER_24_1475 ();
 sg13g2_decap_4 FILLER_24_1480 ();
 sg13g2_fill_1 FILLER_24_1484 ();
 sg13g2_decap_4 FILLER_24_1489 ();
 sg13g2_fill_2 FILLER_24_1493 ();
 sg13g2_fill_2 FILLER_24_1499 ();
 sg13g2_decap_4 FILLER_24_1535 ();
 sg13g2_decap_8 FILLER_24_1653 ();
 sg13g2_fill_2 FILLER_24_1660 ();
 sg13g2_fill_1 FILLER_24_1662 ();
 sg13g2_decap_8 FILLER_24_1667 ();
 sg13g2_decap_8 FILLER_24_1674 ();
 sg13g2_decap_8 FILLER_24_1681 ();
 sg13g2_fill_2 FILLER_24_1688 ();
 sg13g2_decap_8 FILLER_24_1693 ();
 sg13g2_decap_4 FILLER_24_1700 ();
 sg13g2_decap_8 FILLER_24_1707 ();
 sg13g2_decap_8 FILLER_24_1714 ();
 sg13g2_fill_1 FILLER_24_1721 ();
 sg13g2_decap_4 FILLER_24_1726 ();
 sg13g2_fill_2 FILLER_24_1730 ();
 sg13g2_fill_2 FILLER_24_1750 ();
 sg13g2_decap_8 FILLER_24_1773 ();
 sg13g2_decap_8 FILLER_24_1780 ();
 sg13g2_decap_8 FILLER_24_1787 ();
 sg13g2_decap_8 FILLER_24_1794 ();
 sg13g2_fill_2 FILLER_24_1801 ();
 sg13g2_fill_2 FILLER_24_1876 ();
 sg13g2_fill_1 FILLER_24_1878 ();
 sg13g2_decap_4 FILLER_24_1954 ();
 sg13g2_decap_8 FILLER_24_1992 ();
 sg13g2_decap_8 FILLER_24_1999 ();
 sg13g2_fill_1 FILLER_24_2006 ();
 sg13g2_fill_1 FILLER_24_2011 ();
 sg13g2_decap_8 FILLER_24_2049 ();
 sg13g2_decap_8 FILLER_24_2056 ();
 sg13g2_decap_8 FILLER_24_2063 ();
 sg13g2_fill_2 FILLER_24_2070 ();
 sg13g2_decap_8 FILLER_24_2129 ();
 sg13g2_decap_4 FILLER_24_2136 ();
 sg13g2_fill_2 FILLER_24_2140 ();
 sg13g2_decap_8 FILLER_24_2168 ();
 sg13g2_decap_8 FILLER_24_2175 ();
 sg13g2_decap_4 FILLER_24_2182 ();
 sg13g2_fill_2 FILLER_24_2186 ();
 sg13g2_decap_8 FILLER_24_2226 ();
 sg13g2_decap_8 FILLER_24_2233 ();
 sg13g2_decap_8 FILLER_24_2240 ();
 sg13g2_decap_8 FILLER_24_2299 ();
 sg13g2_decap_4 FILLER_24_2306 ();
 sg13g2_fill_1 FILLER_24_2310 ();
 sg13g2_decap_8 FILLER_24_2319 ();
 sg13g2_decap_8 FILLER_24_2326 ();
 sg13g2_decap_4 FILLER_24_2333 ();
 sg13g2_decap_8 FILLER_24_2394 ();
 sg13g2_decap_8 FILLER_24_2401 ();
 sg13g2_fill_2 FILLER_24_2408 ();
 sg13g2_decap_8 FILLER_24_2414 ();
 sg13g2_fill_1 FILLER_24_2421 ();
 sg13g2_decap_8 FILLER_24_2473 ();
 sg13g2_decap_8 FILLER_24_2480 ();
 sg13g2_decap_8 FILLER_24_2487 ();
 sg13g2_decap_4 FILLER_24_2494 ();
 sg13g2_fill_1 FILLER_24_2498 ();
 sg13g2_decap_8 FILLER_24_2564 ();
 sg13g2_decap_8 FILLER_24_2571 ();
 sg13g2_decap_8 FILLER_24_2578 ();
 sg13g2_decap_8 FILLER_24_2585 ();
 sg13g2_decap_8 FILLER_24_2592 ();
 sg13g2_fill_1 FILLER_24_2599 ();
 sg13g2_decap_8 FILLER_24_2626 ();
 sg13g2_fill_2 FILLER_24_2633 ();
 sg13g2_fill_1 FILLER_24_2635 ();
 sg13g2_decap_8 FILLER_24_2672 ();
 sg13g2_decap_8 FILLER_24_2722 ();
 sg13g2_decap_8 FILLER_24_2729 ();
 sg13g2_decap_8 FILLER_24_2736 ();
 sg13g2_decap_8 FILLER_24_2743 ();
 sg13g2_decap_8 FILLER_24_2750 ();
 sg13g2_decap_8 FILLER_24_2757 ();
 sg13g2_decap_8 FILLER_24_2764 ();
 sg13g2_decap_8 FILLER_24_2771 ();
 sg13g2_decap_8 FILLER_24_2778 ();
 sg13g2_decap_8 FILLER_24_2785 ();
 sg13g2_decap_8 FILLER_24_2792 ();
 sg13g2_decap_8 FILLER_24_2799 ();
 sg13g2_decap_8 FILLER_24_2806 ();
 sg13g2_fill_2 FILLER_24_2813 ();
 sg13g2_fill_1 FILLER_24_2815 ();
 sg13g2_fill_2 FILLER_24_2829 ();
 sg13g2_decap_4 FILLER_24_2883 ();
 sg13g2_fill_1 FILLER_24_2887 ();
 sg13g2_decap_8 FILLER_24_2939 ();
 sg13g2_fill_2 FILLER_24_2946 ();
 sg13g2_fill_1 FILLER_24_2948 ();
 sg13g2_decap_8 FILLER_24_2974 ();
 sg13g2_decap_8 FILLER_24_2981 ();
 sg13g2_decap_8 FILLER_24_2988 ();
 sg13g2_fill_2 FILLER_24_2995 ();
 sg13g2_fill_1 FILLER_24_2997 ();
 sg13g2_decap_8 FILLER_24_3026 ();
 sg13g2_decap_8 FILLER_24_3033 ();
 sg13g2_decap_8 FILLER_24_3040 ();
 sg13g2_decap_4 FILLER_24_3047 ();
 sg13g2_fill_1 FILLER_24_3051 ();
 sg13g2_fill_2 FILLER_24_3072 ();
 sg13g2_fill_1 FILLER_24_3074 ();
 sg13g2_decap_8 FILLER_24_3101 ();
 sg13g2_decap_8 FILLER_24_3108 ();
 sg13g2_decap_8 FILLER_24_3115 ();
 sg13g2_decap_8 FILLER_24_3122 ();
 sg13g2_fill_2 FILLER_24_3129 ();
 sg13g2_fill_2 FILLER_24_3135 ();
 sg13g2_fill_1 FILLER_24_3137 ();
 sg13g2_decap_8 FILLER_24_3143 ();
 sg13g2_decap_8 FILLER_24_3150 ();
 sg13g2_decap_8 FILLER_24_3157 ();
 sg13g2_decap_8 FILLER_24_3164 ();
 sg13g2_decap_8 FILLER_24_3171 ();
 sg13g2_decap_8 FILLER_24_3178 ();
 sg13g2_decap_8 FILLER_24_3185 ();
 sg13g2_decap_8 FILLER_24_3192 ();
 sg13g2_decap_8 FILLER_24_3199 ();
 sg13g2_decap_8 FILLER_24_3206 ();
 sg13g2_decap_8 FILLER_24_3213 ();
 sg13g2_decap_8 FILLER_24_3220 ();
 sg13g2_decap_8 FILLER_24_3227 ();
 sg13g2_decap_8 FILLER_24_3234 ();
 sg13g2_decap_8 FILLER_24_3241 ();
 sg13g2_decap_8 FILLER_24_3248 ();
 sg13g2_decap_8 FILLER_24_3255 ();
 sg13g2_decap_8 FILLER_24_3262 ();
 sg13g2_decap_8 FILLER_24_3269 ();
 sg13g2_decap_8 FILLER_24_3276 ();
 sg13g2_decap_8 FILLER_24_3283 ();
 sg13g2_decap_8 FILLER_24_3290 ();
 sg13g2_decap_8 FILLER_24_3297 ();
 sg13g2_decap_8 FILLER_24_3304 ();
 sg13g2_decap_8 FILLER_24_3311 ();
 sg13g2_decap_8 FILLER_24_3318 ();
 sg13g2_decap_8 FILLER_24_3325 ();
 sg13g2_decap_8 FILLER_24_3332 ();
 sg13g2_decap_8 FILLER_24_3339 ();
 sg13g2_decap_8 FILLER_24_3346 ();
 sg13g2_decap_8 FILLER_24_3353 ();
 sg13g2_decap_8 FILLER_24_3360 ();
 sg13g2_decap_8 FILLER_24_3367 ();
 sg13g2_decap_8 FILLER_24_3374 ();
 sg13g2_decap_8 FILLER_24_3381 ();
 sg13g2_decap_8 FILLER_24_3388 ();
 sg13g2_decap_8 FILLER_24_3395 ();
 sg13g2_decap_8 FILLER_24_3402 ();
 sg13g2_decap_8 FILLER_24_3409 ();
 sg13g2_decap_8 FILLER_24_3416 ();
 sg13g2_decap_8 FILLER_24_3423 ();
 sg13g2_decap_8 FILLER_24_3430 ();
 sg13g2_decap_8 FILLER_24_3437 ();
 sg13g2_decap_8 FILLER_24_3444 ();
 sg13g2_decap_8 FILLER_24_3451 ();
 sg13g2_decap_8 FILLER_24_3458 ();
 sg13g2_decap_8 FILLER_24_3465 ();
 sg13g2_decap_8 FILLER_24_3472 ();
 sg13g2_decap_8 FILLER_24_3479 ();
 sg13g2_decap_8 FILLER_24_3486 ();
 sg13g2_decap_8 FILLER_24_3493 ();
 sg13g2_decap_8 FILLER_24_3500 ();
 sg13g2_decap_8 FILLER_24_3507 ();
 sg13g2_decap_8 FILLER_24_3514 ();
 sg13g2_decap_8 FILLER_24_3521 ();
 sg13g2_decap_8 FILLER_24_3528 ();
 sg13g2_decap_8 FILLER_24_3535 ();
 sg13g2_decap_8 FILLER_24_3542 ();
 sg13g2_decap_8 FILLER_24_3549 ();
 sg13g2_decap_8 FILLER_24_3556 ();
 sg13g2_decap_8 FILLER_24_3563 ();
 sg13g2_decap_8 FILLER_24_3570 ();
 sg13g2_fill_2 FILLER_24_3577 ();
 sg13g2_fill_1 FILLER_24_3579 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_4 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_decap_4 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_decap_8 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_256 ();
 sg13g2_decap_8 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_4 FILLER_25_392 ();
 sg13g2_fill_2 FILLER_25_396 ();
 sg13g2_fill_2 FILLER_25_450 ();
 sg13g2_decap_4 FILLER_25_457 ();
 sg13g2_fill_2 FILLER_25_466 ();
 sg13g2_fill_1 FILLER_25_468 ();
 sg13g2_decap_8 FILLER_25_477 ();
 sg13g2_decap_8 FILLER_25_484 ();
 sg13g2_decap_8 FILLER_25_491 ();
 sg13g2_decap_8 FILLER_25_498 ();
 sg13g2_decap_8 FILLER_25_505 ();
 sg13g2_decap_4 FILLER_25_597 ();
 sg13g2_fill_2 FILLER_25_601 ();
 sg13g2_fill_1 FILLER_25_655 ();
 sg13g2_decap_8 FILLER_25_659 ();
 sg13g2_decap_8 FILLER_25_666 ();
 sg13g2_fill_1 FILLER_25_673 ();
 sg13g2_decap_4 FILLER_25_734 ();
 sg13g2_fill_1 FILLER_25_738 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_4 FILLER_25_777 ();
 sg13g2_fill_2 FILLER_25_781 ();
 sg13g2_decap_4 FILLER_25_809 ();
 sg13g2_fill_1 FILLER_25_853 ();
 sg13g2_decap_8 FILLER_25_870 ();
 sg13g2_decap_4 FILLER_25_903 ();
 sg13g2_fill_1 FILLER_25_907 ();
 sg13g2_decap_8 FILLER_25_912 ();
 sg13g2_fill_1 FILLER_25_919 ();
 sg13g2_decap_8 FILLER_25_1011 ();
 sg13g2_decap_8 FILLER_25_1018 ();
 sg13g2_decap_8 FILLER_25_1025 ();
 sg13g2_decap_4 FILLER_25_1032 ();
 sg13g2_decap_8 FILLER_25_1060 ();
 sg13g2_fill_2 FILLER_25_1067 ();
 sg13g2_fill_1 FILLER_25_1083 ();
 sg13g2_decap_8 FILLER_25_1113 ();
 sg13g2_fill_2 FILLER_25_1120 ();
 sg13g2_decap_4 FILLER_25_1151 ();
 sg13g2_decap_8 FILLER_25_1165 ();
 sg13g2_decap_8 FILLER_25_1172 ();
 sg13g2_decap_4 FILLER_25_1179 ();
 sg13g2_fill_2 FILLER_25_1183 ();
 sg13g2_fill_2 FILLER_25_1193 ();
 sg13g2_fill_1 FILLER_25_1195 ();
 sg13g2_fill_1 FILLER_25_1203 ();
 sg13g2_fill_2 FILLER_25_1270 ();
 sg13g2_decap_8 FILLER_25_1282 ();
 sg13g2_decap_8 FILLER_25_1289 ();
 sg13g2_decap_8 FILLER_25_1296 ();
 sg13g2_decap_8 FILLER_25_1303 ();
 sg13g2_decap_8 FILLER_25_1310 ();
 sg13g2_decap_8 FILLER_25_1317 ();
 sg13g2_decap_8 FILLER_25_1384 ();
 sg13g2_decap_8 FILLER_25_1391 ();
 sg13g2_decap_8 FILLER_25_1398 ();
 sg13g2_decap_4 FILLER_25_1405 ();
 sg13g2_fill_2 FILLER_25_1412 ();
 sg13g2_decap_8 FILLER_25_1422 ();
 sg13g2_decap_4 FILLER_25_1429 ();
 sg13g2_decap_4 FILLER_25_1437 ();
 sg13g2_fill_2 FILLER_25_1441 ();
 sg13g2_decap_4 FILLER_25_1448 ();
 sg13g2_fill_2 FILLER_25_1452 ();
 sg13g2_decap_4 FILLER_25_1480 ();
 sg13g2_fill_1 FILLER_25_1484 ();
 sg13g2_fill_1 FILLER_25_1586 ();
 sg13g2_fill_2 FILLER_25_1617 ();
 sg13g2_fill_2 FILLER_25_1664 ();
 sg13g2_fill_2 FILLER_25_1671 ();
 sg13g2_decap_4 FILLER_25_1713 ();
 sg13g2_fill_2 FILLER_25_1717 ();
 sg13g2_decap_8 FILLER_25_1740 ();
 sg13g2_fill_1 FILLER_25_1747 ();
 sg13g2_decap_8 FILLER_25_1756 ();
 sg13g2_decap_8 FILLER_25_1763 ();
 sg13g2_fill_2 FILLER_25_1770 ();
 sg13g2_fill_1 FILLER_25_1772 ();
 sg13g2_decap_8 FILLER_25_1777 ();
 sg13g2_decap_8 FILLER_25_1787 ();
 sg13g2_decap_4 FILLER_25_1802 ();
 sg13g2_fill_1 FILLER_25_1806 ();
 sg13g2_fill_2 FILLER_25_1838 ();
 sg13g2_decap_8 FILLER_25_1883 ();
 sg13g2_decap_8 FILLER_25_1890 ();
 sg13g2_fill_2 FILLER_25_1897 ();
 sg13g2_fill_1 FILLER_25_1899 ();
 sg13g2_decap_8 FILLER_25_1904 ();
 sg13g2_decap_4 FILLER_25_1911 ();
 sg13g2_decap_8 FILLER_25_1941 ();
 sg13g2_decap_4 FILLER_25_1948 ();
 sg13g2_fill_1 FILLER_25_1952 ();
 sg13g2_decap_8 FILLER_25_1979 ();
 sg13g2_decap_8 FILLER_25_1986 ();
 sg13g2_decap_8 FILLER_25_1993 ();
 sg13g2_decap_8 FILLER_25_2052 ();
 sg13g2_decap_8 FILLER_25_2059 ();
 sg13g2_decap_8 FILLER_25_2066 ();
 sg13g2_fill_1 FILLER_25_2073 ();
 sg13g2_decap_8 FILLER_25_2126 ();
 sg13g2_decap_4 FILLER_25_2133 ();
 sg13g2_decap_8 FILLER_25_2171 ();
 sg13g2_decap_8 FILLER_25_2178 ();
 sg13g2_decap_4 FILLER_25_2185 ();
 sg13g2_decap_8 FILLER_25_2226 ();
 sg13g2_fill_1 FILLER_25_2233 ();
 sg13g2_decap_8 FILLER_25_2321 ();
 sg13g2_decap_8 FILLER_25_2328 ();
 sg13g2_decap_4 FILLER_25_2343 ();
 sg13g2_fill_1 FILLER_25_2353 ();
 sg13g2_decap_8 FILLER_25_2380 ();
 sg13g2_decap_8 FILLER_25_2387 ();
 sg13g2_decap_8 FILLER_25_2394 ();
 sg13g2_decap_8 FILLER_25_2409 ();
 sg13g2_decap_8 FILLER_25_2416 ();
 sg13g2_decap_8 FILLER_25_2423 ();
 sg13g2_decap_8 FILLER_25_2476 ();
 sg13g2_decap_8 FILLER_25_2483 ();
 sg13g2_decap_8 FILLER_25_2490 ();
 sg13g2_decap_4 FILLER_25_2497 ();
 sg13g2_decap_8 FILLER_25_2537 ();
 sg13g2_decap_4 FILLER_25_2544 ();
 sg13g2_fill_2 FILLER_25_2548 ();
 sg13g2_decap_8 FILLER_25_2555 ();
 sg13g2_fill_2 FILLER_25_2562 ();
 sg13g2_decap_4 FILLER_25_2572 ();
 sg13g2_fill_2 FILLER_25_2576 ();
 sg13g2_decap_4 FILLER_25_2630 ();
 sg13g2_fill_2 FILLER_25_2634 ();
 sg13g2_decap_8 FILLER_25_2662 ();
 sg13g2_decap_8 FILLER_25_2669 ();
 sg13g2_fill_2 FILLER_25_2676 ();
 sg13g2_fill_2 FILLER_25_2707 ();
 sg13g2_fill_1 FILLER_25_2709 ();
 sg13g2_decap_8 FILLER_25_2771 ();
 sg13g2_decap_8 FILLER_25_2778 ();
 sg13g2_decap_8 FILLER_25_2785 ();
 sg13g2_fill_2 FILLER_25_2833 ();
 sg13g2_fill_1 FILLER_25_2835 ();
 sg13g2_fill_2 FILLER_25_2883 ();
 sg13g2_fill_2 FILLER_25_2961 ();
 sg13g2_fill_2 FILLER_25_2989 ();
 sg13g2_fill_1 FILLER_25_2991 ();
 sg13g2_decap_4 FILLER_25_3036 ();
 sg13g2_decap_8 FILLER_25_3112 ();
 sg13g2_decap_4 FILLER_25_3119 ();
 sg13g2_fill_2 FILLER_25_3123 ();
 sg13g2_fill_1 FILLER_25_3134 ();
 sg13g2_decap_8 FILLER_25_3151 ();
 sg13g2_decap_8 FILLER_25_3158 ();
 sg13g2_decap_8 FILLER_25_3165 ();
 sg13g2_decap_8 FILLER_25_3172 ();
 sg13g2_decap_8 FILLER_25_3179 ();
 sg13g2_decap_8 FILLER_25_3186 ();
 sg13g2_decap_8 FILLER_25_3193 ();
 sg13g2_decap_8 FILLER_25_3200 ();
 sg13g2_decap_8 FILLER_25_3207 ();
 sg13g2_decap_8 FILLER_25_3214 ();
 sg13g2_decap_8 FILLER_25_3221 ();
 sg13g2_decap_8 FILLER_25_3228 ();
 sg13g2_decap_8 FILLER_25_3235 ();
 sg13g2_decap_8 FILLER_25_3242 ();
 sg13g2_decap_8 FILLER_25_3249 ();
 sg13g2_decap_8 FILLER_25_3256 ();
 sg13g2_decap_8 FILLER_25_3263 ();
 sg13g2_decap_8 FILLER_25_3270 ();
 sg13g2_decap_8 FILLER_25_3277 ();
 sg13g2_decap_8 FILLER_25_3284 ();
 sg13g2_decap_8 FILLER_25_3291 ();
 sg13g2_decap_8 FILLER_25_3298 ();
 sg13g2_decap_8 FILLER_25_3305 ();
 sg13g2_decap_8 FILLER_25_3312 ();
 sg13g2_decap_8 FILLER_25_3319 ();
 sg13g2_decap_8 FILLER_25_3326 ();
 sg13g2_decap_8 FILLER_25_3333 ();
 sg13g2_decap_8 FILLER_25_3340 ();
 sg13g2_decap_8 FILLER_25_3347 ();
 sg13g2_decap_8 FILLER_25_3354 ();
 sg13g2_decap_8 FILLER_25_3361 ();
 sg13g2_decap_8 FILLER_25_3368 ();
 sg13g2_decap_8 FILLER_25_3375 ();
 sg13g2_decap_8 FILLER_25_3382 ();
 sg13g2_decap_8 FILLER_25_3389 ();
 sg13g2_decap_8 FILLER_25_3396 ();
 sg13g2_decap_8 FILLER_25_3403 ();
 sg13g2_decap_8 FILLER_25_3410 ();
 sg13g2_decap_8 FILLER_25_3417 ();
 sg13g2_decap_8 FILLER_25_3424 ();
 sg13g2_decap_8 FILLER_25_3431 ();
 sg13g2_decap_8 FILLER_25_3438 ();
 sg13g2_decap_8 FILLER_25_3445 ();
 sg13g2_decap_8 FILLER_25_3452 ();
 sg13g2_decap_8 FILLER_25_3459 ();
 sg13g2_decap_8 FILLER_25_3466 ();
 sg13g2_decap_8 FILLER_25_3473 ();
 sg13g2_decap_8 FILLER_25_3480 ();
 sg13g2_decap_8 FILLER_25_3487 ();
 sg13g2_decap_8 FILLER_25_3494 ();
 sg13g2_decap_8 FILLER_25_3501 ();
 sg13g2_decap_8 FILLER_25_3508 ();
 sg13g2_decap_8 FILLER_25_3515 ();
 sg13g2_decap_8 FILLER_25_3522 ();
 sg13g2_decap_8 FILLER_25_3529 ();
 sg13g2_decap_8 FILLER_25_3536 ();
 sg13g2_decap_8 FILLER_25_3543 ();
 sg13g2_decap_8 FILLER_25_3550 ();
 sg13g2_decap_8 FILLER_25_3557 ();
 sg13g2_decap_8 FILLER_25_3564 ();
 sg13g2_decap_8 FILLER_25_3571 ();
 sg13g2_fill_2 FILLER_25_3578 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_4 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_57 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_4 FILLER_26_105 ();
 sg13g2_fill_1 FILLER_26_109 ();
 sg13g2_decap_4 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_152 ();
 sg13g2_decap_4 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_183 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_decap_4 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_decap_4 FILLER_26_302 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_decap_4 FILLER_26_341 ();
 sg13g2_decap_8 FILLER_26_353 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_decap_4 FILLER_26_388 ();
 sg13g2_fill_1 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_26_405 ();
 sg13g2_decap_4 FILLER_26_419 ();
 sg13g2_decap_4 FILLER_26_439 ();
 sg13g2_fill_1 FILLER_26_443 ();
 sg13g2_decap_4 FILLER_26_464 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_4 FILLER_26_490 ();
 sg13g2_fill_1 FILLER_26_494 ();
 sg13g2_decap_4 FILLER_26_526 ();
 sg13g2_fill_2 FILLER_26_534 ();
 sg13g2_decap_4 FILLER_26_568 ();
 sg13g2_decap_4 FILLER_26_582 ();
 sg13g2_fill_2 FILLER_26_622 ();
 sg13g2_fill_2 FILLER_26_637 ();
 sg13g2_fill_1 FILLER_26_639 ();
 sg13g2_decap_4 FILLER_26_676 ();
 sg13g2_fill_1 FILLER_26_680 ();
 sg13g2_decap_8 FILLER_26_738 ();
 sg13g2_decap_8 FILLER_26_745 ();
 sg13g2_decap_8 FILLER_26_752 ();
 sg13g2_fill_1 FILLER_26_759 ();
 sg13g2_fill_2 FILLER_26_786 ();
 sg13g2_fill_1 FILLER_26_788 ();
 sg13g2_decap_8 FILLER_26_815 ();
 sg13g2_decap_8 FILLER_26_822 ();
 sg13g2_decap_8 FILLER_26_829 ();
 sg13g2_fill_1 FILLER_26_836 ();
 sg13g2_decap_4 FILLER_26_841 ();
 sg13g2_fill_1 FILLER_26_845 ();
 sg13g2_fill_2 FILLER_26_857 ();
 sg13g2_decap_8 FILLER_26_896 ();
 sg13g2_decap_8 FILLER_26_903 ();
 sg13g2_decap_4 FILLER_26_910 ();
 sg13g2_decap_8 FILLER_26_946 ();
 sg13g2_fill_2 FILLER_26_953 ();
 sg13g2_fill_1 FILLER_26_955 ();
 sg13g2_fill_2 FILLER_26_1008 ();
 sg13g2_fill_1 FILLER_26_1010 ();
 sg13g2_decap_8 FILLER_26_1016 ();
 sg13g2_decap_4 FILLER_26_1023 ();
 sg13g2_decap_4 FILLER_26_1035 ();
 sg13g2_decap_4 FILLER_26_1104 ();
 sg13g2_fill_1 FILLER_26_1108 ();
 sg13g2_decap_8 FILLER_26_1145 ();
 sg13g2_decap_8 FILLER_26_1152 ();
 sg13g2_decap_8 FILLER_26_1159 ();
 sg13g2_decap_8 FILLER_26_1166 ();
 sg13g2_decap_8 FILLER_26_1173 ();
 sg13g2_decap_8 FILLER_26_1180 ();
 sg13g2_decap_8 FILLER_26_1187 ();
 sg13g2_decap_4 FILLER_26_1194 ();
 sg13g2_fill_2 FILLER_26_1208 ();
 sg13g2_fill_2 FILLER_26_1262 ();
 sg13g2_fill_2 FILLER_26_1269 ();
 sg13g2_decap_8 FILLER_26_1279 ();
 sg13g2_decap_8 FILLER_26_1286 ();
 sg13g2_decap_4 FILLER_26_1293 ();
 sg13g2_decap_8 FILLER_26_1323 ();
 sg13g2_fill_1 FILLER_26_1330 ();
 sg13g2_decap_8 FILLER_26_1336 ();
 sg13g2_fill_1 FILLER_26_1347 ();
 sg13g2_decap_8 FILLER_26_1378 ();
 sg13g2_decap_8 FILLER_26_1385 ();
 sg13g2_decap_8 FILLER_26_1392 ();
 sg13g2_decap_8 FILLER_26_1399 ();
 sg13g2_fill_2 FILLER_26_1406 ();
 sg13g2_fill_1 FILLER_26_1413 ();
 sg13g2_decap_4 FILLER_26_1419 ();
 sg13g2_decap_8 FILLER_26_1426 ();
 sg13g2_fill_2 FILLER_26_1433 ();
 sg13g2_fill_1 FILLER_26_1435 ();
 sg13g2_decap_8 FILLER_26_1440 ();
 sg13g2_fill_2 FILLER_26_1452 ();
 sg13g2_fill_1 FILLER_26_1454 ();
 sg13g2_decap_8 FILLER_26_1485 ();
 sg13g2_decap_8 FILLER_26_1492 ();
 sg13g2_decap_4 FILLER_26_1499 ();
 sg13g2_fill_1 FILLER_26_1503 ();
 sg13g2_decap_8 FILLER_26_1507 ();
 sg13g2_fill_2 FILLER_26_1514 ();
 sg13g2_decap_8 FILLER_26_1520 ();
 sg13g2_decap_4 FILLER_26_1527 ();
 sg13g2_decap_8 FILLER_26_1541 ();
 sg13g2_decap_4 FILLER_26_1548 ();
 sg13g2_fill_1 FILLER_26_1552 ();
 sg13g2_fill_1 FILLER_26_1566 ();
 sg13g2_decap_8 FILLER_26_1583 ();
 sg13g2_decap_8 FILLER_26_1590 ();
 sg13g2_fill_1 FILLER_26_1597 ();
 sg13g2_decap_8 FILLER_26_1602 ();
 sg13g2_decap_8 FILLER_26_1609 ();
 sg13g2_decap_8 FILLER_26_1616 ();
 sg13g2_fill_2 FILLER_26_1623 ();
 sg13g2_fill_1 FILLER_26_1625 ();
 sg13g2_decap_8 FILLER_26_1652 ();
 sg13g2_fill_2 FILLER_26_1659 ();
 sg13g2_decap_4 FILLER_26_1674 ();
 sg13g2_fill_2 FILLER_26_1678 ();
 sg13g2_decap_8 FILLER_26_1739 ();
 sg13g2_decap_8 FILLER_26_1746 ();
 sg13g2_decap_4 FILLER_26_1753 ();
 sg13g2_decap_8 FILLER_26_1827 ();
 sg13g2_fill_2 FILLER_26_1834 ();
 sg13g2_fill_1 FILLER_26_1851 ();
 sg13g2_fill_2 FILLER_26_1868 ();
 sg13g2_decap_8 FILLER_26_1878 ();
 sg13g2_decap_8 FILLER_26_1937 ();
 sg13g2_decap_4 FILLER_26_1944 ();
 sg13g2_fill_2 FILLER_26_1948 ();
 sg13g2_fill_1 FILLER_26_1976 ();
 sg13g2_decap_8 FILLER_26_1981 ();
 sg13g2_decap_8 FILLER_26_1988 ();
 sg13g2_decap_4 FILLER_26_1995 ();
 sg13g2_fill_2 FILLER_26_1999 ();
 sg13g2_decap_8 FILLER_26_2050 ();
 sg13g2_decap_8 FILLER_26_2057 ();
 sg13g2_decap_8 FILLER_26_2064 ();
 sg13g2_fill_2 FILLER_26_2071 ();
 sg13g2_decap_4 FILLER_26_2188 ();
 sg13g2_decap_4 FILLER_26_2232 ();
 sg13g2_fill_2 FILLER_26_2236 ();
 sg13g2_fill_2 FILLER_26_2302 ();
 sg13g2_fill_1 FILLER_26_2304 ();
 sg13g2_decap_4 FILLER_26_2318 ();
 sg13g2_fill_1 FILLER_26_2322 ();
 sg13g2_fill_2 FILLER_26_2366 ();
 sg13g2_fill_1 FILLER_26_2368 ();
 sg13g2_decap_8 FILLER_26_2403 ();
 sg13g2_fill_2 FILLER_26_2410 ();
 sg13g2_fill_1 FILLER_26_2412 ();
 sg13g2_fill_1 FILLER_26_2444 ();
 sg13g2_decap_8 FILLER_26_2451 ();
 sg13g2_fill_2 FILLER_26_2458 ();
 sg13g2_fill_1 FILLER_26_2460 ();
 sg13g2_fill_2 FILLER_26_2467 ();
 sg13g2_decap_8 FILLER_26_2477 ();
 sg13g2_fill_2 FILLER_26_2484 ();
 sg13g2_fill_1 FILLER_26_2486 ();
 sg13g2_decap_8 FILLER_26_2517 ();
 sg13g2_decap_8 FILLER_26_2524 ();
 sg13g2_decap_4 FILLER_26_2531 ();
 sg13g2_fill_2 FILLER_26_2535 ();
 sg13g2_decap_8 FILLER_26_2563 ();
 sg13g2_decap_8 FILLER_26_2570 ();
 sg13g2_decap_4 FILLER_26_2577 ();
 sg13g2_fill_1 FILLER_26_2581 ();
 sg13g2_decap_4 FILLER_26_2634 ();
 sg13g2_fill_2 FILLER_26_2638 ();
 sg13g2_decap_8 FILLER_26_2666 ();
 sg13g2_decap_8 FILLER_26_2673 ();
 sg13g2_fill_2 FILLER_26_2680 ();
 sg13g2_fill_1 FILLER_26_2682 ();
 sg13g2_decap_4 FILLER_26_2745 ();
 sg13g2_fill_1 FILLER_26_2788 ();
 sg13g2_decap_8 FILLER_26_2841 ();
 sg13g2_fill_2 FILLER_26_2848 ();
 sg13g2_fill_2 FILLER_26_2877 ();
 sg13g2_decap_4 FILLER_26_2884 ();
 sg13g2_fill_1 FILLER_26_2888 ();
 sg13g2_decap_8 FILLER_26_2939 ();
 sg13g2_fill_2 FILLER_26_2946 ();
 sg13g2_decap_8 FILLER_26_2987 ();
 sg13g2_fill_2 FILLER_26_2994 ();
 sg13g2_fill_1 FILLER_26_2996 ();
 sg13g2_fill_2 FILLER_26_3036 ();
 sg13g2_fill_1 FILLER_26_3038 ();
 sg13g2_fill_2 FILLER_26_3081 ();
 sg13g2_fill_2 FILLER_26_3117 ();
 sg13g2_fill_1 FILLER_26_3119 ();
 sg13g2_decap_8 FILLER_26_3162 ();
 sg13g2_decap_8 FILLER_26_3169 ();
 sg13g2_decap_8 FILLER_26_3176 ();
 sg13g2_decap_8 FILLER_26_3183 ();
 sg13g2_decap_8 FILLER_26_3190 ();
 sg13g2_decap_8 FILLER_26_3197 ();
 sg13g2_decap_8 FILLER_26_3204 ();
 sg13g2_decap_8 FILLER_26_3211 ();
 sg13g2_decap_8 FILLER_26_3218 ();
 sg13g2_decap_8 FILLER_26_3225 ();
 sg13g2_decap_8 FILLER_26_3232 ();
 sg13g2_decap_8 FILLER_26_3239 ();
 sg13g2_decap_8 FILLER_26_3246 ();
 sg13g2_decap_8 FILLER_26_3253 ();
 sg13g2_decap_8 FILLER_26_3260 ();
 sg13g2_decap_8 FILLER_26_3267 ();
 sg13g2_decap_8 FILLER_26_3274 ();
 sg13g2_decap_8 FILLER_26_3281 ();
 sg13g2_decap_8 FILLER_26_3288 ();
 sg13g2_decap_8 FILLER_26_3295 ();
 sg13g2_decap_8 FILLER_26_3302 ();
 sg13g2_decap_8 FILLER_26_3309 ();
 sg13g2_decap_8 FILLER_26_3316 ();
 sg13g2_decap_8 FILLER_26_3323 ();
 sg13g2_decap_8 FILLER_26_3330 ();
 sg13g2_decap_8 FILLER_26_3337 ();
 sg13g2_decap_8 FILLER_26_3344 ();
 sg13g2_decap_8 FILLER_26_3351 ();
 sg13g2_decap_8 FILLER_26_3358 ();
 sg13g2_decap_8 FILLER_26_3365 ();
 sg13g2_decap_8 FILLER_26_3372 ();
 sg13g2_decap_8 FILLER_26_3379 ();
 sg13g2_decap_8 FILLER_26_3386 ();
 sg13g2_decap_8 FILLER_26_3393 ();
 sg13g2_decap_8 FILLER_26_3400 ();
 sg13g2_decap_8 FILLER_26_3407 ();
 sg13g2_decap_8 FILLER_26_3414 ();
 sg13g2_decap_8 FILLER_26_3421 ();
 sg13g2_decap_8 FILLER_26_3428 ();
 sg13g2_decap_8 FILLER_26_3435 ();
 sg13g2_decap_8 FILLER_26_3442 ();
 sg13g2_decap_8 FILLER_26_3449 ();
 sg13g2_decap_8 FILLER_26_3456 ();
 sg13g2_decap_8 FILLER_26_3463 ();
 sg13g2_decap_8 FILLER_26_3470 ();
 sg13g2_decap_8 FILLER_26_3477 ();
 sg13g2_decap_8 FILLER_26_3484 ();
 sg13g2_decap_8 FILLER_26_3491 ();
 sg13g2_decap_8 FILLER_26_3498 ();
 sg13g2_decap_8 FILLER_26_3505 ();
 sg13g2_decap_8 FILLER_26_3512 ();
 sg13g2_decap_8 FILLER_26_3519 ();
 sg13g2_decap_8 FILLER_26_3526 ();
 sg13g2_decap_8 FILLER_26_3533 ();
 sg13g2_decap_8 FILLER_26_3540 ();
 sg13g2_decap_8 FILLER_26_3547 ();
 sg13g2_decap_8 FILLER_26_3554 ();
 sg13g2_decap_8 FILLER_26_3561 ();
 sg13g2_decap_8 FILLER_26_3568 ();
 sg13g2_decap_4 FILLER_26_3575 ();
 sg13g2_fill_1 FILLER_26_3579 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_4 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_178 ();
 sg13g2_decap_4 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_decap_4 FILLER_27_220 ();
 sg13g2_decap_8 FILLER_27_250 ();
 sg13g2_decap_8 FILLER_27_257 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_decap_8 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_353 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_fill_2 FILLER_27_413 ();
 sg13g2_fill_2 FILLER_27_441 ();
 sg13g2_fill_1 FILLER_27_443 ();
 sg13g2_fill_2 FILLER_27_457 ();
 sg13g2_decap_8 FILLER_27_472 ();
 sg13g2_fill_2 FILLER_27_479 ();
 sg13g2_fill_1 FILLER_27_481 ();
 sg13g2_fill_1 FILLER_27_487 ();
 sg13g2_decap_4 FILLER_27_522 ();
 sg13g2_fill_1 FILLER_27_526 ();
 sg13g2_decap_4 FILLER_27_582 ();
 sg13g2_fill_1 FILLER_27_586 ();
 sg13g2_decap_4 FILLER_27_628 ();
 sg13g2_fill_1 FILLER_27_632 ();
 sg13g2_decap_4 FILLER_27_641 ();
 sg13g2_fill_2 FILLER_27_645 ();
 sg13g2_decap_8 FILLER_27_699 ();
 sg13g2_fill_1 FILLER_27_738 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_4 FILLER_27_840 ();
 sg13g2_fill_2 FILLER_27_900 ();
 sg13g2_decap_8 FILLER_27_942 ();
 sg13g2_decap_8 FILLER_27_949 ();
 sg13g2_fill_1 FILLER_27_956 ();
 sg13g2_decap_4 FILLER_27_996 ();
 sg13g2_decap_4 FILLER_27_1010 ();
 sg13g2_decap_4 FILLER_27_1089 ();
 sg13g2_fill_1 FILLER_27_1093 ();
 sg13g2_fill_1 FILLER_27_1120 ();
 sg13g2_decap_8 FILLER_27_1150 ();
 sg13g2_decap_8 FILLER_27_1157 ();
 sg13g2_decap_8 FILLER_27_1164 ();
 sg13g2_decap_8 FILLER_27_1171 ();
 sg13g2_fill_1 FILLER_27_1178 ();
 sg13g2_decap_8 FILLER_27_1184 ();
 sg13g2_fill_2 FILLER_27_1191 ();
 sg13g2_fill_1 FILLER_27_1193 ();
 sg13g2_decap_8 FILLER_27_1222 ();
 sg13g2_fill_2 FILLER_27_1229 ();
 sg13g2_decap_8 FILLER_27_1236 ();
 sg13g2_decap_8 FILLER_27_1243 ();
 sg13g2_fill_2 FILLER_27_1250 ();
 sg13g2_fill_1 FILLER_27_1252 ();
 sg13g2_decap_4 FILLER_27_1282 ();
 sg13g2_fill_2 FILLER_27_1286 ();
 sg13g2_decap_8 FILLER_27_1293 ();
 sg13g2_fill_2 FILLER_27_1300 ();
 sg13g2_fill_1 FILLER_27_1302 ();
 sg13g2_fill_1 FILLER_27_1311 ();
 sg13g2_decap_8 FILLER_27_1338 ();
 sg13g2_decap_8 FILLER_27_1345 ();
 sg13g2_decap_4 FILLER_27_1352 ();
 sg13g2_decap_4 FILLER_27_1389 ();
 sg13g2_fill_2 FILLER_27_1393 ();
 sg13g2_decap_8 FILLER_27_1477 ();
 sg13g2_decap_4 FILLER_27_1484 ();
 sg13g2_fill_1 FILLER_27_1488 ();
 sg13g2_decap_8 FILLER_27_1493 ();
 sg13g2_fill_2 FILLER_27_1500 ();
 sg13g2_fill_1 FILLER_27_1509 ();
 sg13g2_decap_8 FILLER_27_1513 ();
 sg13g2_fill_2 FILLER_27_1520 ();
 sg13g2_decap_8 FILLER_27_1527 ();
 sg13g2_decap_4 FILLER_27_1534 ();
 sg13g2_fill_1 FILLER_27_1538 ();
 sg13g2_decap_4 FILLER_27_1549 ();
 sg13g2_fill_2 FILLER_27_1562 ();
 sg13g2_fill_2 FILLER_27_1569 ();
 sg13g2_fill_1 FILLER_27_1571 ();
 sg13g2_decap_4 FILLER_27_1580 ();
 sg13g2_decap_4 FILLER_27_1589 ();
 sg13g2_decap_8 FILLER_27_1597 ();
 sg13g2_fill_2 FILLER_27_1604 ();
 sg13g2_decap_8 FILLER_27_1609 ();
 sg13g2_decap_8 FILLER_27_1616 ();
 sg13g2_fill_2 FILLER_27_1623 ();
 sg13g2_fill_2 FILLER_27_1633 ();
 sg13g2_fill_1 FILLER_27_1635 ();
 sg13g2_decap_4 FILLER_27_1662 ();
 sg13g2_decap_8 FILLER_27_1679 ();
 sg13g2_fill_2 FILLER_27_1694 ();
 sg13g2_fill_1 FILLER_27_1696 ();
 sg13g2_decap_4 FILLER_27_1747 ();
 sg13g2_fill_1 FILLER_27_1751 ();
 sg13g2_fill_2 FILLER_27_1802 ();
 sg13g2_fill_2 FILLER_27_1809 ();
 sg13g2_decap_8 FILLER_27_1824 ();
 sg13g2_decap_8 FILLER_27_1831 ();
 sg13g2_decap_8 FILLER_27_1838 ();
 sg13g2_decap_8 FILLER_27_1845 ();
 sg13g2_fill_2 FILLER_27_1852 ();
 sg13g2_fill_1 FILLER_27_1854 ();
 sg13g2_decap_8 FILLER_27_1881 ();
 sg13g2_decap_4 FILLER_27_1888 ();
 sg13g2_fill_1 FILLER_27_1892 ();
 sg13g2_decap_8 FILLER_27_1949 ();
 sg13g2_decap_4 FILLER_27_1956 ();
 sg13g2_fill_1 FILLER_27_1960 ();
 sg13g2_decap_8 FILLER_27_1969 ();
 sg13g2_decap_8 FILLER_27_1976 ();
 sg13g2_decap_8 FILLER_27_1983 ();
 sg13g2_fill_1 FILLER_27_1990 ();
 sg13g2_fill_2 FILLER_27_1999 ();
 sg13g2_decap_8 FILLER_27_2053 ();
 sg13g2_decap_8 FILLER_27_2060 ();
 sg13g2_decap_8 FILLER_27_2067 ();
 sg13g2_fill_1 FILLER_27_2074 ();
 sg13g2_decap_8 FILLER_27_2120 ();
 sg13g2_decap_8 FILLER_27_2127 ();
 sg13g2_decap_8 FILLER_27_2134 ();
 sg13g2_decap_8 FILLER_27_2173 ();
 sg13g2_decap_8 FILLER_27_2180 ();
 sg13g2_decap_4 FILLER_27_2187 ();
 sg13g2_fill_1 FILLER_27_2191 ();
 sg13g2_decap_8 FILLER_27_2224 ();
 sg13g2_decap_8 FILLER_27_2231 ();
 sg13g2_fill_2 FILLER_27_2238 ();
 sg13g2_decap_8 FILLER_27_2246 ();
 sg13g2_decap_4 FILLER_27_2253 ();
 sg13g2_fill_1 FILLER_27_2257 ();
 sg13g2_decap_8 FILLER_27_2290 ();
 sg13g2_decap_4 FILLER_27_2297 ();
 sg13g2_fill_1 FILLER_27_2301 ();
 sg13g2_fill_2 FILLER_27_2341 ();
 sg13g2_decap_8 FILLER_27_2401 ();
 sg13g2_decap_8 FILLER_27_2408 ();
 sg13g2_fill_2 FILLER_27_2415 ();
 sg13g2_fill_1 FILLER_27_2417 ();
 sg13g2_decap_8 FILLER_27_2449 ();
 sg13g2_decap_8 FILLER_27_2456 ();
 sg13g2_decap_8 FILLER_27_2463 ();
 sg13g2_decap_8 FILLER_27_2470 ();
 sg13g2_fill_1 FILLER_27_2477 ();
 sg13g2_decap_8 FILLER_27_2522 ();
 sg13g2_decap_8 FILLER_27_2529 ();
 sg13g2_fill_2 FILLER_27_2536 ();
 sg13g2_fill_1 FILLER_27_2538 ();
 sg13g2_decap_8 FILLER_27_2565 ();
 sg13g2_fill_2 FILLER_27_2572 ();
 sg13g2_fill_2 FILLER_27_2579 ();
 sg13g2_decap_8 FILLER_27_2615 ();
 sg13g2_decap_8 FILLER_27_2622 ();
 sg13g2_decap_8 FILLER_27_2632 ();
 sg13g2_fill_2 FILLER_27_2639 ();
 sg13g2_decap_8 FILLER_27_2667 ();
 sg13g2_decap_4 FILLER_27_2674 ();
 sg13g2_fill_1 FILLER_27_2715 ();
 sg13g2_decap_8 FILLER_27_2725 ();
 sg13g2_decap_8 FILLER_27_2732 ();
 sg13g2_decap_4 FILLER_27_2739 ();
 sg13g2_fill_1 FILLER_27_2743 ();
 sg13g2_fill_1 FILLER_27_2791 ();
 sg13g2_decap_8 FILLER_27_2826 ();
 sg13g2_fill_2 FILLER_27_2833 ();
 sg13g2_fill_1 FILLER_27_2835 ();
 sg13g2_fill_1 FILLER_27_2869 ();
 sg13g2_decap_8 FILLER_27_2875 ();
 sg13g2_decap_8 FILLER_27_2882 ();
 sg13g2_decap_8 FILLER_27_2889 ();
 sg13g2_decap_4 FILLER_27_2896 ();
 sg13g2_decap_8 FILLER_27_2932 ();
 sg13g2_decap_8 FILLER_27_2939 ();
 sg13g2_decap_8 FILLER_27_2946 ();
 sg13g2_fill_2 FILLER_27_2953 ();
 sg13g2_decap_8 FILLER_27_2994 ();
 sg13g2_fill_1 FILLER_27_3001 ();
 sg13g2_fill_2 FILLER_27_3044 ();
 sg13g2_fill_2 FILLER_27_3059 ();
 sg13g2_fill_1 FILLER_27_3061 ();
 sg13g2_decap_8 FILLER_27_3107 ();
 sg13g2_decap_8 FILLER_27_3188 ();
 sg13g2_decap_8 FILLER_27_3195 ();
 sg13g2_decap_8 FILLER_27_3202 ();
 sg13g2_decap_8 FILLER_27_3209 ();
 sg13g2_decap_8 FILLER_27_3216 ();
 sg13g2_decap_8 FILLER_27_3223 ();
 sg13g2_decap_8 FILLER_27_3230 ();
 sg13g2_decap_8 FILLER_27_3237 ();
 sg13g2_decap_8 FILLER_27_3244 ();
 sg13g2_decap_8 FILLER_27_3251 ();
 sg13g2_decap_8 FILLER_27_3258 ();
 sg13g2_decap_8 FILLER_27_3265 ();
 sg13g2_decap_8 FILLER_27_3272 ();
 sg13g2_decap_8 FILLER_27_3279 ();
 sg13g2_decap_8 FILLER_27_3286 ();
 sg13g2_decap_8 FILLER_27_3293 ();
 sg13g2_decap_8 FILLER_27_3300 ();
 sg13g2_decap_8 FILLER_27_3307 ();
 sg13g2_decap_8 FILLER_27_3314 ();
 sg13g2_decap_8 FILLER_27_3321 ();
 sg13g2_decap_8 FILLER_27_3328 ();
 sg13g2_decap_8 FILLER_27_3335 ();
 sg13g2_decap_8 FILLER_27_3342 ();
 sg13g2_decap_8 FILLER_27_3349 ();
 sg13g2_decap_8 FILLER_27_3356 ();
 sg13g2_decap_8 FILLER_27_3363 ();
 sg13g2_decap_8 FILLER_27_3370 ();
 sg13g2_decap_8 FILLER_27_3377 ();
 sg13g2_decap_8 FILLER_27_3384 ();
 sg13g2_decap_8 FILLER_27_3391 ();
 sg13g2_decap_8 FILLER_27_3398 ();
 sg13g2_decap_8 FILLER_27_3405 ();
 sg13g2_decap_8 FILLER_27_3412 ();
 sg13g2_decap_8 FILLER_27_3419 ();
 sg13g2_decap_8 FILLER_27_3426 ();
 sg13g2_decap_8 FILLER_27_3433 ();
 sg13g2_decap_8 FILLER_27_3440 ();
 sg13g2_decap_8 FILLER_27_3447 ();
 sg13g2_decap_8 FILLER_27_3454 ();
 sg13g2_decap_8 FILLER_27_3461 ();
 sg13g2_decap_8 FILLER_27_3468 ();
 sg13g2_decap_8 FILLER_27_3475 ();
 sg13g2_decap_8 FILLER_27_3482 ();
 sg13g2_decap_8 FILLER_27_3489 ();
 sg13g2_decap_8 FILLER_27_3496 ();
 sg13g2_decap_8 FILLER_27_3503 ();
 sg13g2_decap_8 FILLER_27_3510 ();
 sg13g2_decap_8 FILLER_27_3517 ();
 sg13g2_decap_8 FILLER_27_3524 ();
 sg13g2_decap_8 FILLER_27_3531 ();
 sg13g2_decap_8 FILLER_27_3538 ();
 sg13g2_decap_8 FILLER_27_3545 ();
 sg13g2_decap_8 FILLER_27_3552 ();
 sg13g2_decap_8 FILLER_27_3559 ();
 sg13g2_decap_8 FILLER_27_3566 ();
 sg13g2_decap_8 FILLER_27_3573 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_37 ();
 sg13g2_decap_8 FILLER_28_76 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_decap_8 FILLER_28_97 ();
 sg13g2_decap_4 FILLER_28_104 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_147 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_255 ();
 sg13g2_decap_8 FILLER_28_262 ();
 sg13g2_decap_8 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_333 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_4 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_390 ();
 sg13g2_fill_2 FILLER_28_417 ();
 sg13g2_fill_1 FILLER_28_419 ();
 sg13g2_decap_8 FILLER_28_521 ();
 sg13g2_decap_4 FILLER_28_528 ();
 sg13g2_fill_1 FILLER_28_573 ();
 sg13g2_decap_4 FILLER_28_584 ();
 sg13g2_fill_1 FILLER_28_588 ();
 sg13g2_fill_1 FILLER_28_593 ();
 sg13g2_decap_8 FILLER_28_643 ();
 sg13g2_decap_8 FILLER_28_650 ();
 sg13g2_decap_8 FILLER_28_657 ();
 sg13g2_decap_8 FILLER_28_664 ();
 sg13g2_fill_1 FILLER_28_671 ();
 sg13g2_fill_1 FILLER_28_704 ();
 sg13g2_fill_1 FILLER_28_747 ();
 sg13g2_fill_2 FILLER_28_779 ();
 sg13g2_fill_1 FILLER_28_781 ();
 sg13g2_decap_8 FILLER_28_830 ();
 sg13g2_decap_8 FILLER_28_837 ();
 sg13g2_decap_8 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_fill_2 FILLER_28_858 ();
 sg13g2_fill_1 FILLER_28_860 ();
 sg13g2_fill_2 FILLER_28_913 ();
 sg13g2_decap_8 FILLER_28_946 ();
 sg13g2_decap_4 FILLER_28_953 ();
 sg13g2_fill_2 FILLER_28_957 ();
 sg13g2_fill_2 FILLER_28_964 ();
 sg13g2_decap_8 FILLER_28_997 ();
 sg13g2_decap_4 FILLER_28_1033 ();
 sg13g2_fill_1 FILLER_28_1071 ();
 sg13g2_fill_2 FILLER_28_1087 ();
 sg13g2_fill_1 FILLER_28_1089 ();
 sg13g2_fill_2 FILLER_28_1098 ();
 sg13g2_decap_8 FILLER_28_1125 ();
 sg13g2_decap_8 FILLER_28_1132 ();
 sg13g2_decap_8 FILLER_28_1139 ();
 sg13g2_fill_1 FILLER_28_1146 ();
 sg13g2_decap_8 FILLER_28_1173 ();
 sg13g2_decap_4 FILLER_28_1180 ();
 sg13g2_fill_2 FILLER_28_1184 ();
 sg13g2_decap_8 FILLER_28_1241 ();
 sg13g2_decap_8 FILLER_28_1248 ();
 sg13g2_fill_1 FILLER_28_1255 ();
 sg13g2_decap_8 FILLER_28_1289 ();
 sg13g2_decap_8 FILLER_28_1341 ();
 sg13g2_decap_8 FILLER_28_1348 ();
 sg13g2_decap_4 FILLER_28_1355 ();
 sg13g2_fill_2 FILLER_28_1381 ();
 sg13g2_fill_1 FILLER_28_1383 ();
 sg13g2_decap_8 FILLER_28_1414 ();
 sg13g2_fill_1 FILLER_28_1421 ();
 sg13g2_fill_2 FILLER_28_1448 ();
 sg13g2_fill_1 FILLER_28_1450 ();
 sg13g2_fill_2 FILLER_28_1455 ();
 sg13g2_fill_1 FILLER_28_1457 ();
 sg13g2_decap_8 FILLER_28_1462 ();
 sg13g2_decap_8 FILLER_28_1469 ();
 sg13g2_fill_2 FILLER_28_1528 ();
 sg13g2_decap_8 FILLER_28_1535 ();
 sg13g2_fill_2 FILLER_28_1576 ();
 sg13g2_fill_2 FILLER_28_1630 ();
 sg13g2_fill_1 FILLER_28_1648 ();
 sg13g2_decap_8 FILLER_28_1683 ();
 sg13g2_decap_8 FILLER_28_1690 ();
 sg13g2_decap_4 FILLER_28_1697 ();
 sg13g2_fill_1 FILLER_28_1701 ();
 sg13g2_decap_8 FILLER_28_1741 ();
 sg13g2_decap_4 FILLER_28_1748 ();
 sg13g2_fill_2 FILLER_28_1778 ();
 sg13g2_decap_8 FILLER_28_1832 ();
 sg13g2_decap_8 FILLER_28_1839 ();
 sg13g2_decap_8 FILLER_28_1846 ();
 sg13g2_decap_8 FILLER_28_1879 ();
 sg13g2_fill_1 FILLER_28_1886 ();
 sg13g2_decap_8 FILLER_28_1895 ();
 sg13g2_decap_8 FILLER_28_1902 ();
 sg13g2_fill_2 FILLER_28_1909 ();
 sg13g2_decap_8 FILLER_28_1937 ();
 sg13g2_fill_2 FILLER_28_1944 ();
 sg13g2_fill_1 FILLER_28_1946 ();
 sg13g2_decap_8 FILLER_28_1953 ();
 sg13g2_fill_2 FILLER_28_1960 ();
 sg13g2_decap_8 FILLER_28_1988 ();
 sg13g2_decap_4 FILLER_28_1995 ();
 sg13g2_fill_2 FILLER_28_2051 ();
 sg13g2_decap_8 FILLER_28_2061 ();
 sg13g2_decap_8 FILLER_28_2068 ();
 sg13g2_decap_8 FILLER_28_2075 ();
 sg13g2_decap_8 FILLER_28_2082 ();
 sg13g2_decap_4 FILLER_28_2089 ();
 sg13g2_fill_2 FILLER_28_2093 ();
 sg13g2_decap_8 FILLER_28_2107 ();
 sg13g2_decap_8 FILLER_28_2114 ();
 sg13g2_decap_8 FILLER_28_2121 ();
 sg13g2_decap_4 FILLER_28_2128 ();
 sg13g2_fill_1 FILLER_28_2132 ();
 sg13g2_decap_8 FILLER_28_2182 ();
 sg13g2_decap_4 FILLER_28_2189 ();
 sg13g2_decap_4 FILLER_28_2219 ();
 sg13g2_decap_8 FILLER_28_2231 ();
 sg13g2_decap_8 FILLER_28_2238 ();
 sg13g2_decap_8 FILLER_28_2245 ();
 sg13g2_decap_8 FILLER_28_2252 ();
 sg13g2_decap_8 FILLER_28_2259 ();
 sg13g2_decap_8 FILLER_28_2277 ();
 sg13g2_decap_8 FILLER_28_2284 ();
 sg13g2_decap_8 FILLER_28_2291 ();
 sg13g2_decap_8 FILLER_28_2298 ();
 sg13g2_fill_1 FILLER_28_2409 ();
 sg13g2_decap_8 FILLER_28_2452 ();
 sg13g2_decap_8 FILLER_28_2459 ();
 sg13g2_decap_4 FILLER_28_2466 ();
 sg13g2_fill_1 FILLER_28_2470 ();
 sg13g2_decap_4 FILLER_28_2533 ();
 sg13g2_fill_1 FILLER_28_2537 ();
 sg13g2_decap_8 FILLER_28_2616 ();
 sg13g2_decap_8 FILLER_28_2662 ();
 sg13g2_decap_8 FILLER_28_2669 ();
 sg13g2_decap_8 FILLER_28_2676 ();
 sg13g2_decap_4 FILLER_28_2683 ();
 sg13g2_decap_4 FILLER_28_2717 ();
 sg13g2_decap_4 FILLER_28_2747 ();
 sg13g2_decap_8 FILLER_28_2792 ();
 sg13g2_fill_2 FILLER_28_2799 ();
 sg13g2_fill_1 FILLER_28_2801 ();
 sg13g2_decap_8 FILLER_28_2854 ();
 sg13g2_fill_2 FILLER_28_2861 ();
 sg13g2_fill_1 FILLER_28_2880 ();
 sg13g2_decap_8 FILLER_28_2888 ();
 sg13g2_decap_8 FILLER_28_2895 ();
 sg13g2_fill_2 FILLER_28_2902 ();
 sg13g2_fill_1 FILLER_28_2908 ();
 sg13g2_decap_8 FILLER_28_2927 ();
 sg13g2_decap_8 FILLER_28_2934 ();
 sg13g2_decap_4 FILLER_28_2941 ();
 sg13g2_decap_8 FILLER_28_2952 ();
 sg13g2_decap_4 FILLER_28_2959 ();
 sg13g2_fill_1 FILLER_28_2963 ();
 sg13g2_fill_2 FILLER_28_2976 ();
 sg13g2_fill_1 FILLER_28_2978 ();
 sg13g2_decap_8 FILLER_28_2987 ();
 sg13g2_decap_8 FILLER_28_2994 ();
 sg13g2_fill_2 FILLER_28_3001 ();
 sg13g2_fill_2 FILLER_28_3012 ();
 sg13g2_decap_8 FILLER_28_3026 ();
 sg13g2_decap_8 FILLER_28_3033 ();
 sg13g2_decap_8 FILLER_28_3040 ();
 sg13g2_decap_4 FILLER_28_3047 ();
 sg13g2_fill_1 FILLER_28_3051 ();
 sg13g2_fill_1 FILLER_28_3077 ();
 sg13g2_decap_8 FILLER_28_3086 ();
 sg13g2_decap_8 FILLER_28_3093 ();
 sg13g2_decap_8 FILLER_28_3100 ();
 sg13g2_fill_1 FILLER_28_3107 ();
 sg13g2_decap_8 FILLER_28_3116 ();
 sg13g2_decap_4 FILLER_28_3123 ();
 sg13g2_decap_4 FILLER_28_3153 ();
 sg13g2_fill_1 FILLER_28_3157 ();
 sg13g2_decap_8 FILLER_28_3184 ();
 sg13g2_decap_4 FILLER_28_3191 ();
 sg13g2_fill_2 FILLER_28_3195 ();
 sg13g2_decap_8 FILLER_28_3201 ();
 sg13g2_decap_8 FILLER_28_3208 ();
 sg13g2_decap_8 FILLER_28_3215 ();
 sg13g2_decap_8 FILLER_28_3222 ();
 sg13g2_decap_8 FILLER_28_3229 ();
 sg13g2_decap_8 FILLER_28_3236 ();
 sg13g2_decap_8 FILLER_28_3243 ();
 sg13g2_decap_8 FILLER_28_3250 ();
 sg13g2_decap_8 FILLER_28_3257 ();
 sg13g2_decap_8 FILLER_28_3264 ();
 sg13g2_decap_8 FILLER_28_3271 ();
 sg13g2_decap_8 FILLER_28_3278 ();
 sg13g2_decap_8 FILLER_28_3285 ();
 sg13g2_decap_8 FILLER_28_3292 ();
 sg13g2_decap_8 FILLER_28_3299 ();
 sg13g2_decap_8 FILLER_28_3306 ();
 sg13g2_decap_8 FILLER_28_3313 ();
 sg13g2_decap_8 FILLER_28_3320 ();
 sg13g2_decap_8 FILLER_28_3327 ();
 sg13g2_decap_8 FILLER_28_3334 ();
 sg13g2_decap_8 FILLER_28_3341 ();
 sg13g2_decap_8 FILLER_28_3348 ();
 sg13g2_decap_8 FILLER_28_3355 ();
 sg13g2_decap_8 FILLER_28_3362 ();
 sg13g2_decap_8 FILLER_28_3369 ();
 sg13g2_decap_8 FILLER_28_3376 ();
 sg13g2_decap_8 FILLER_28_3383 ();
 sg13g2_decap_8 FILLER_28_3390 ();
 sg13g2_decap_8 FILLER_28_3397 ();
 sg13g2_decap_8 FILLER_28_3404 ();
 sg13g2_decap_8 FILLER_28_3411 ();
 sg13g2_decap_8 FILLER_28_3418 ();
 sg13g2_decap_8 FILLER_28_3425 ();
 sg13g2_decap_8 FILLER_28_3432 ();
 sg13g2_decap_8 FILLER_28_3439 ();
 sg13g2_decap_8 FILLER_28_3446 ();
 sg13g2_decap_8 FILLER_28_3453 ();
 sg13g2_decap_8 FILLER_28_3460 ();
 sg13g2_decap_8 FILLER_28_3467 ();
 sg13g2_decap_8 FILLER_28_3474 ();
 sg13g2_decap_8 FILLER_28_3481 ();
 sg13g2_decap_8 FILLER_28_3488 ();
 sg13g2_decap_8 FILLER_28_3495 ();
 sg13g2_decap_8 FILLER_28_3502 ();
 sg13g2_decap_8 FILLER_28_3509 ();
 sg13g2_decap_8 FILLER_28_3516 ();
 sg13g2_decap_8 FILLER_28_3523 ();
 sg13g2_decap_8 FILLER_28_3530 ();
 sg13g2_decap_8 FILLER_28_3537 ();
 sg13g2_decap_8 FILLER_28_3544 ();
 sg13g2_decap_8 FILLER_28_3551 ();
 sg13g2_decap_8 FILLER_28_3558 ();
 sg13g2_decap_8 FILLER_28_3565 ();
 sg13g2_decap_8 FILLER_28_3572 ();
 sg13g2_fill_1 FILLER_28_3579 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_decap_4 FILLER_29_100 ();
 sg13g2_fill_1 FILLER_29_104 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_fill_2 FILLER_29_271 ();
 sg13g2_fill_1 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_333 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_344 ();
 sg13g2_decap_4 FILLER_29_362 ();
 sg13g2_fill_2 FILLER_29_366 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_fill_1 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_431 ();
 sg13g2_fill_1 FILLER_29_433 ();
 sg13g2_decap_8 FILLER_29_438 ();
 sg13g2_fill_1 FILLER_29_445 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_fill_2 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_515 ();
 sg13g2_decap_4 FILLER_29_522 ();
 sg13g2_fill_1 FILLER_29_526 ();
 sg13g2_decap_4 FILLER_29_563 ();
 sg13g2_fill_1 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_594 ();
 sg13g2_decap_4 FILLER_29_601 ();
 sg13g2_fill_1 FILLER_29_605 ();
 sg13g2_fill_1 FILLER_29_619 ();
 sg13g2_decap_8 FILLER_29_646 ();
 sg13g2_decap_8 FILLER_29_653 ();
 sg13g2_fill_1 FILLER_29_660 ();
 sg13g2_decap_8 FILLER_29_687 ();
 sg13g2_decap_8 FILLER_29_694 ();
 sg13g2_fill_2 FILLER_29_753 ();
 sg13g2_fill_2 FILLER_29_771 ();
 sg13g2_fill_2 FILLER_29_789 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_decap_8 FILLER_29_850 ();
 sg13g2_decap_8 FILLER_29_857 ();
 sg13g2_decap_4 FILLER_29_947 ();
 sg13g2_fill_2 FILLER_29_951 ();
 sg13g2_fill_1 FILLER_29_963 ();
 sg13g2_decap_8 FILLER_29_993 ();
 sg13g2_decap_8 FILLER_29_1000 ();
 sg13g2_decap_8 FILLER_29_1007 ();
 sg13g2_decap_4 FILLER_29_1014 ();
 sg13g2_fill_1 FILLER_29_1018 ();
 sg13g2_decap_8 FILLER_29_1024 ();
 sg13g2_decap_8 FILLER_29_1031 ();
 sg13g2_decap_8 FILLER_29_1038 ();
 sg13g2_decap_4 FILLER_29_1045 ();
 sg13g2_fill_2 FILLER_29_1049 ();
 sg13g2_decap_8 FILLER_29_1077 ();
 sg13g2_fill_2 FILLER_29_1084 ();
 sg13g2_fill_1 FILLER_29_1086 ();
 sg13g2_decap_8 FILLER_29_1113 ();
 sg13g2_decap_8 FILLER_29_1120 ();
 sg13g2_decap_8 FILLER_29_1127 ();
 sg13g2_decap_4 FILLER_29_1134 ();
 sg13g2_fill_2 FILLER_29_1138 ();
 sg13g2_decap_8 FILLER_29_1166 ();
 sg13g2_decap_4 FILLER_29_1173 ();
 sg13g2_fill_2 FILLER_29_1177 ();
 sg13g2_decap_8 FILLER_29_1218 ();
 sg13g2_decap_8 FILLER_29_1225 ();
 sg13g2_decap_8 FILLER_29_1232 ();
 sg13g2_decap_8 FILLER_29_1242 ();
 sg13g2_decap_8 FILLER_29_1249 ();
 sg13g2_fill_2 FILLER_29_1256 ();
 sg13g2_fill_1 FILLER_29_1258 ();
 sg13g2_decap_8 FILLER_29_1288 ();
 sg13g2_fill_1 FILLER_29_1330 ();
 sg13g2_decap_8 FILLER_29_1357 ();
 sg13g2_decap_4 FILLER_29_1364 ();
 sg13g2_fill_1 FILLER_29_1385 ();
 sg13g2_decap_8 FILLER_29_1412 ();
 sg13g2_fill_2 FILLER_29_1419 ();
 sg13g2_decap_8 FILLER_29_1466 ();
 sg13g2_fill_2 FILLER_29_1473 ();
 sg13g2_fill_2 FILLER_29_1480 ();
 sg13g2_fill_2 FILLER_29_1485 ();
 sg13g2_decap_4 FILLER_29_1544 ();
 sg13g2_fill_1 FILLER_29_1636 ();
 sg13g2_fill_2 FILLER_29_1645 ();
 sg13g2_fill_2 FILLER_29_1651 ();
 sg13g2_decap_8 FILLER_29_1696 ();
 sg13g2_decap_8 FILLER_29_1703 ();
 sg13g2_fill_2 FILLER_29_1710 ();
 sg13g2_fill_1 FILLER_29_1712 ();
 sg13g2_fill_2 FILLER_29_1717 ();
 sg13g2_fill_1 FILLER_29_1719 ();
 sg13g2_decap_8 FILLER_29_1733 ();
 sg13g2_decap_4 FILLER_29_1740 ();
 sg13g2_decap_8 FILLER_29_1770 ();
 sg13g2_decap_8 FILLER_29_1777 ();
 sg13g2_decap_8 FILLER_29_1784 ();
 sg13g2_decap_4 FILLER_29_1791 ();
 sg13g2_fill_1 FILLER_29_1795 ();
 sg13g2_fill_2 FILLER_29_1800 ();
 sg13g2_decap_4 FILLER_29_1839 ();
 sg13g2_fill_1 FILLER_29_1843 ();
 sg13g2_decap_8 FILLER_29_1887 ();
 sg13g2_decap_8 FILLER_29_1894 ();
 sg13g2_fill_1 FILLER_29_1901 ();
 sg13g2_decap_8 FILLER_29_1933 ();
 sg13g2_fill_2 FILLER_29_1940 ();
 sg13g2_fill_1 FILLER_29_1942 ();
 sg13g2_decap_8 FILLER_29_1981 ();
 sg13g2_decap_8 FILLER_29_1988 ();
 sg13g2_decap_8 FILLER_29_1995 ();
 sg13g2_fill_2 FILLER_29_2002 ();
 sg13g2_decap_4 FILLER_29_2044 ();
 sg13g2_decap_8 FILLER_29_2074 ();
 sg13g2_decap_8 FILLER_29_2081 ();
 sg13g2_decap_4 FILLER_29_2088 ();
 sg13g2_fill_2 FILLER_29_2092 ();
 sg13g2_decap_8 FILLER_29_2126 ();
 sg13g2_decap_8 FILLER_29_2133 ();
 sg13g2_decap_8 FILLER_29_2180 ();
 sg13g2_decap_8 FILLER_29_2187 ();
 sg13g2_decap_8 FILLER_29_2194 ();
 sg13g2_fill_2 FILLER_29_2201 ();
 sg13g2_decap_8 FILLER_29_2209 ();
 sg13g2_decap_8 FILLER_29_2216 ();
 sg13g2_decap_8 FILLER_29_2228 ();
 sg13g2_fill_2 FILLER_29_2235 ();
 sg13g2_fill_1 FILLER_29_2237 ();
 sg13g2_fill_2 FILLER_29_2264 ();
 sg13g2_fill_1 FILLER_29_2266 ();
 sg13g2_decap_8 FILLER_29_2293 ();
 sg13g2_decap_8 FILLER_29_2300 ();
 sg13g2_decap_4 FILLER_29_2307 ();
 sg13g2_fill_1 FILLER_29_2345 ();
 sg13g2_decap_8 FILLER_29_2403 ();
 sg13g2_fill_1 FILLER_29_2410 ();
 sg13g2_decap_8 FILLER_29_2457 ();
 sg13g2_decap_8 FILLER_29_2464 ();
 sg13g2_decap_8 FILLER_29_2471 ();
 sg13g2_fill_1 FILLER_29_2478 ();
 sg13g2_decap_8 FILLER_29_2522 ();
 sg13g2_decap_8 FILLER_29_2529 ();
 sg13g2_decap_4 FILLER_29_2536 ();
 sg13g2_fill_1 FILLER_29_2540 ();
 sg13g2_decap_8 FILLER_29_2655 ();
 sg13g2_decap_8 FILLER_29_2662 ();
 sg13g2_decap_8 FILLER_29_2669 ();
 sg13g2_decap_8 FILLER_29_2676 ();
 sg13g2_decap_8 FILLER_29_2683 ();
 sg13g2_decap_8 FILLER_29_2690 ();
 sg13g2_decap_4 FILLER_29_2697 ();
 sg13g2_decap_8 FILLER_29_2744 ();
 sg13g2_decap_8 FILLER_29_2751 ();
 sg13g2_decap_8 FILLER_29_2758 ();
 sg13g2_decap_8 FILLER_29_2765 ();
 sg13g2_decap_4 FILLER_29_2793 ();
 sg13g2_decap_8 FILLER_29_2823 ();
 sg13g2_decap_8 FILLER_29_2830 ();
 sg13g2_fill_2 FILLER_29_2837 ();
 sg13g2_fill_1 FILLER_29_2844 ();
 sg13g2_decap_4 FILLER_29_2879 ();
 sg13g2_fill_1 FILLER_29_2883 ();
 sg13g2_fill_1 FILLER_29_2936 ();
 sg13g2_decap_8 FILLER_29_2958 ();
 sg13g2_decap_8 FILLER_29_2965 ();
 sg13g2_fill_2 FILLER_29_2972 ();
 sg13g2_fill_1 FILLER_29_2974 ();
 sg13g2_fill_2 FILLER_29_3001 ();
 sg13g2_fill_1 FILLER_29_3003 ();
 sg13g2_decap_4 FILLER_29_3023 ();
 sg13g2_fill_1 FILLER_29_3027 ();
 sg13g2_fill_2 FILLER_29_3033 ();
 sg13g2_fill_2 FILLER_29_3048 ();
 sg13g2_decap_8 FILLER_29_3080 ();
 sg13g2_decap_8 FILLER_29_3087 ();
 sg13g2_fill_2 FILLER_29_3094 ();
 sg13g2_fill_1 FILLER_29_3134 ();
 sg13g2_decap_8 FILLER_29_3171 ();
 sg13g2_decap_8 FILLER_29_3182 ();
 sg13g2_fill_1 FILLER_29_3189 ();
 sg13g2_decap_8 FILLER_29_3207 ();
 sg13g2_decap_8 FILLER_29_3214 ();
 sg13g2_decap_8 FILLER_29_3221 ();
 sg13g2_decap_8 FILLER_29_3228 ();
 sg13g2_decap_8 FILLER_29_3235 ();
 sg13g2_decap_8 FILLER_29_3242 ();
 sg13g2_decap_8 FILLER_29_3249 ();
 sg13g2_decap_8 FILLER_29_3256 ();
 sg13g2_decap_8 FILLER_29_3263 ();
 sg13g2_decap_8 FILLER_29_3270 ();
 sg13g2_decap_8 FILLER_29_3277 ();
 sg13g2_decap_8 FILLER_29_3284 ();
 sg13g2_decap_8 FILLER_29_3291 ();
 sg13g2_decap_8 FILLER_29_3298 ();
 sg13g2_decap_8 FILLER_29_3305 ();
 sg13g2_decap_8 FILLER_29_3312 ();
 sg13g2_decap_8 FILLER_29_3319 ();
 sg13g2_decap_8 FILLER_29_3326 ();
 sg13g2_decap_8 FILLER_29_3333 ();
 sg13g2_decap_8 FILLER_29_3340 ();
 sg13g2_decap_8 FILLER_29_3347 ();
 sg13g2_decap_8 FILLER_29_3354 ();
 sg13g2_decap_8 FILLER_29_3361 ();
 sg13g2_decap_8 FILLER_29_3368 ();
 sg13g2_decap_8 FILLER_29_3375 ();
 sg13g2_decap_8 FILLER_29_3382 ();
 sg13g2_decap_8 FILLER_29_3389 ();
 sg13g2_decap_8 FILLER_29_3396 ();
 sg13g2_decap_8 FILLER_29_3403 ();
 sg13g2_decap_8 FILLER_29_3410 ();
 sg13g2_decap_8 FILLER_29_3417 ();
 sg13g2_decap_8 FILLER_29_3424 ();
 sg13g2_decap_8 FILLER_29_3431 ();
 sg13g2_decap_8 FILLER_29_3438 ();
 sg13g2_decap_8 FILLER_29_3445 ();
 sg13g2_decap_8 FILLER_29_3452 ();
 sg13g2_decap_8 FILLER_29_3459 ();
 sg13g2_decap_8 FILLER_29_3466 ();
 sg13g2_decap_8 FILLER_29_3473 ();
 sg13g2_decap_8 FILLER_29_3480 ();
 sg13g2_decap_8 FILLER_29_3487 ();
 sg13g2_decap_8 FILLER_29_3494 ();
 sg13g2_decap_8 FILLER_29_3501 ();
 sg13g2_decap_8 FILLER_29_3508 ();
 sg13g2_decap_8 FILLER_29_3515 ();
 sg13g2_decap_8 FILLER_29_3522 ();
 sg13g2_decap_8 FILLER_29_3529 ();
 sg13g2_decap_8 FILLER_29_3536 ();
 sg13g2_decap_8 FILLER_29_3543 ();
 sg13g2_decap_8 FILLER_29_3550 ();
 sg13g2_decap_8 FILLER_29_3557 ();
 sg13g2_decap_8 FILLER_29_3564 ();
 sg13g2_decap_8 FILLER_29_3571 ();
 sg13g2_fill_2 FILLER_29_3578 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_71 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_decap_4 FILLER_30_148 ();
 sg13g2_decap_4 FILLER_30_178 ();
 sg13g2_fill_1 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_decap_8 FILLER_30_270 ();
 sg13g2_decap_8 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_300 ();
 sg13g2_decap_4 FILLER_30_307 ();
 sg13g2_fill_2 FILLER_30_314 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_fill_2 FILLER_30_371 ();
 sg13g2_fill_1 FILLER_30_373 ();
 sg13g2_decap_4 FILLER_30_378 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_fill_2 FILLER_30_415 ();
 sg13g2_fill_1 FILLER_30_443 ();
 sg13g2_fill_2 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_478 ();
 sg13g2_decap_8 FILLER_30_485 ();
 sg13g2_decap_4 FILLER_30_492 ();
 sg13g2_decap_4 FILLER_30_500 ();
 sg13g2_decap_8 FILLER_30_508 ();
 sg13g2_decap_8 FILLER_30_515 ();
 sg13g2_decap_8 FILLER_30_522 ();
 sg13g2_decap_8 FILLER_30_529 ();
 sg13g2_fill_2 FILLER_30_536 ();
 sg13g2_fill_1 FILLER_30_538 ();
 sg13g2_decap_4 FILLER_30_565 ();
 sg13g2_fill_1 FILLER_30_569 ();
 sg13g2_fill_2 FILLER_30_601 ();
 sg13g2_fill_1 FILLER_30_603 ();
 sg13g2_fill_1 FILLER_30_608 ();
 sg13g2_decap_8 FILLER_30_640 ();
 sg13g2_fill_1 FILLER_30_647 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_fill_1 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_4 FILLER_30_782 ();
 sg13g2_decap_8 FILLER_30_846 ();
 sg13g2_decap_8 FILLER_30_853 ();
 sg13g2_decap_8 FILLER_30_860 ();
 sg13g2_fill_1 FILLER_30_867 ();
 sg13g2_decap_8 FILLER_30_897 ();
 sg13g2_decap_8 FILLER_30_904 ();
 sg13g2_decap_8 FILLER_30_911 ();
 sg13g2_fill_1 FILLER_30_918 ();
 sg13g2_fill_1 FILLER_30_922 ();
 sg13g2_decap_4 FILLER_30_954 ();
 sg13g2_fill_1 FILLER_30_958 ();
 sg13g2_decap_4 FILLER_30_993 ();
 sg13g2_fill_1 FILLER_30_997 ();
 sg13g2_fill_2 FILLER_30_1006 ();
 sg13g2_fill_1 FILLER_30_1008 ();
 sg13g2_decap_8 FILLER_30_1061 ();
 sg13g2_fill_1 FILLER_30_1068 ();
 sg13g2_decap_8 FILLER_30_1073 ();
 sg13g2_decap_8 FILLER_30_1080 ();
 sg13g2_decap_8 FILLER_30_1087 ();
 sg13g2_fill_2 FILLER_30_1094 ();
 sg13g2_decap_8 FILLER_30_1106 ();
 sg13g2_decap_4 FILLER_30_1113 ();
 sg13g2_fill_1 FILLER_30_1117 ();
 sg13g2_decap_8 FILLER_30_1144 ();
 sg13g2_fill_2 FILLER_30_1203 ();
 sg13g2_decap_4 FILLER_30_1221 ();
 sg13g2_fill_1 FILLER_30_1225 ();
 sg13g2_decap_8 FILLER_30_1252 ();
 sg13g2_fill_2 FILLER_30_1259 ();
 sg13g2_fill_1 FILLER_30_1261 ();
 sg13g2_fill_1 FILLER_30_1265 ();
 sg13g2_decap_8 FILLER_30_1273 ();
 sg13g2_fill_2 FILLER_30_1280 ();
 sg13g2_fill_1 FILLER_30_1282 ();
 sg13g2_decap_8 FILLER_30_1286 ();
 sg13g2_decap_4 FILLER_30_1293 ();
 sg13g2_fill_2 FILLER_30_1297 ();
 sg13g2_fill_1 FILLER_30_1341 ();
 sg13g2_decap_8 FILLER_30_1346 ();
 sg13g2_decap_8 FILLER_30_1353 ();
 sg13g2_decap_4 FILLER_30_1360 ();
 sg13g2_fill_1 FILLER_30_1364 ();
 sg13g2_fill_2 FILLER_30_1394 ();
 sg13g2_fill_1 FILLER_30_1396 ();
 sg13g2_fill_2 FILLER_30_1405 ();
 sg13g2_decap_8 FILLER_30_1447 ();
 sg13g2_decap_4 FILLER_30_1454 ();
 sg13g2_fill_1 FILLER_30_1458 ();
 sg13g2_fill_2 FILLER_30_1469 ();
 sg13g2_fill_2 FILLER_30_1481 ();
 sg13g2_fill_1 FILLER_30_1483 ();
 sg13g2_decap_8 FILLER_30_1546 ();
 sg13g2_decap_4 FILLER_30_1587 ();
 sg13g2_decap_8 FILLER_30_1595 ();
 sg13g2_decap_4 FILLER_30_1605 ();
 sg13g2_decap_8 FILLER_30_1625 ();
 sg13g2_decap_8 FILLER_30_1632 ();
 sg13g2_decap_4 FILLER_30_1639 ();
 sg13g2_decap_8 FILLER_30_1646 ();
 sg13g2_decap_8 FILLER_30_1653 ();
 sg13g2_decap_4 FILLER_30_1660 ();
 sg13g2_fill_2 FILLER_30_1664 ();
 sg13g2_decap_8 FILLER_30_1686 ();
 sg13g2_decap_8 FILLER_30_1693 ();
 sg13g2_decap_8 FILLER_30_1700 ();
 sg13g2_decap_8 FILLER_30_1707 ();
 sg13g2_decap_8 FILLER_30_1714 ();
 sg13g2_decap_8 FILLER_30_1721 ();
 sg13g2_fill_1 FILLER_30_1754 ();
 sg13g2_decap_8 FILLER_30_1759 ();
 sg13g2_decap_4 FILLER_30_1766 ();
 sg13g2_fill_1 FILLER_30_1770 ();
 sg13g2_decap_8 FILLER_30_1797 ();
 sg13g2_fill_2 FILLER_30_1893 ();
 sg13g2_decap_8 FILLER_30_1933 ();
 sg13g2_decap_4 FILLER_30_1940 ();
 sg13g2_fill_2 FILLER_30_1944 ();
 sg13g2_decap_8 FILLER_30_1998 ();
 sg13g2_decap_8 FILLER_30_2005 ();
 sg13g2_decap_4 FILLER_30_2012 ();
 sg13g2_decap_8 FILLER_30_2030 ();
 sg13g2_decap_8 FILLER_30_2037 ();
 sg13g2_fill_1 FILLER_30_2070 ();
 sg13g2_decap_4 FILLER_30_2083 ();
 sg13g2_decap_8 FILLER_30_2133 ();
 sg13g2_decap_4 FILLER_30_2140 ();
 sg13g2_fill_2 FILLER_30_2144 ();
 sg13g2_decap_8 FILLER_30_2178 ();
 sg13g2_decap_8 FILLER_30_2185 ();
 sg13g2_decap_4 FILLER_30_2192 ();
 sg13g2_fill_2 FILLER_30_2196 ();
 sg13g2_decap_4 FILLER_30_2250 ();
 sg13g2_fill_1 FILLER_30_2254 ();
 sg13g2_decap_8 FILLER_30_2307 ();
 sg13g2_decap_8 FILLER_30_2314 ();
 sg13g2_decap_8 FILLER_30_2321 ();
 sg13g2_decap_8 FILLER_30_2328 ();
 sg13g2_decap_8 FILLER_30_2335 ();
 sg13g2_decap_8 FILLER_30_2342 ();
 sg13g2_decap_8 FILLER_30_2392 ();
 sg13g2_decap_4 FILLER_30_2399 ();
 sg13g2_fill_1 FILLER_30_2403 ();
 sg13g2_decap_8 FILLER_30_2462 ();
 sg13g2_decap_8 FILLER_30_2469 ();
 sg13g2_decap_8 FILLER_30_2476 ();
 sg13g2_decap_8 FILLER_30_2483 ();
 sg13g2_decap_8 FILLER_30_2533 ();
 sg13g2_decap_8 FILLER_30_2540 ();
 sg13g2_decap_4 FILLER_30_2547 ();
 sg13g2_decap_8 FILLER_30_2590 ();
 sg13g2_decap_8 FILLER_30_2597 ();
 sg13g2_decap_8 FILLER_30_2604 ();
 sg13g2_decap_4 FILLER_30_2611 ();
 sg13g2_fill_2 FILLER_30_2615 ();
 sg13g2_decap_8 FILLER_30_2646 ();
 sg13g2_fill_2 FILLER_30_2653 ();
 sg13g2_fill_1 FILLER_30_2655 ();
 sg13g2_decap_8 FILLER_30_2685 ();
 sg13g2_fill_2 FILLER_30_2718 ();
 sg13g2_decap_8 FILLER_30_2742 ();
 sg13g2_decap_8 FILLER_30_2749 ();
 sg13g2_decap_8 FILLER_30_2756 ();
 sg13g2_decap_4 FILLER_30_2763 ();
 sg13g2_fill_1 FILLER_30_2767 ();
 sg13g2_decap_8 FILLER_30_2800 ();
 sg13g2_decap_8 FILLER_30_2820 ();
 sg13g2_decap_4 FILLER_30_2827 ();
 sg13g2_fill_2 FILLER_30_2831 ();
 sg13g2_fill_2 FILLER_30_2893 ();
 sg13g2_fill_1 FILLER_30_2895 ();
 sg13g2_fill_1 FILLER_30_2909 ();
 sg13g2_decap_8 FILLER_30_2962 ();
 sg13g2_fill_2 FILLER_30_2969 ();
 sg13g2_fill_2 FILLER_30_3023 ();
 sg13g2_fill_1 FILLER_30_3025 ();
 sg13g2_decap_4 FILLER_30_3031 ();
 sg13g2_fill_2 FILLER_30_3043 ();
 sg13g2_fill_1 FILLER_30_3045 ();
 sg13g2_fill_1 FILLER_30_3054 ();
 sg13g2_fill_2 FILLER_30_3094 ();
 sg13g2_decap_8 FILLER_30_3139 ();
 sg13g2_decap_4 FILLER_30_3146 ();
 sg13g2_fill_2 FILLER_30_3154 ();
 sg13g2_fill_1 FILLER_30_3156 ();
 sg13g2_decap_8 FILLER_30_3162 ();
 sg13g2_decap_4 FILLER_30_3169 ();
 sg13g2_fill_1 FILLER_30_3173 ();
 sg13g2_fill_2 FILLER_30_3179 ();
 sg13g2_fill_1 FILLER_30_3181 ();
 sg13g2_decap_8 FILLER_30_3221 ();
 sg13g2_decap_8 FILLER_30_3228 ();
 sg13g2_decap_8 FILLER_30_3235 ();
 sg13g2_decap_8 FILLER_30_3242 ();
 sg13g2_decap_8 FILLER_30_3249 ();
 sg13g2_decap_8 FILLER_30_3256 ();
 sg13g2_decap_8 FILLER_30_3263 ();
 sg13g2_decap_8 FILLER_30_3270 ();
 sg13g2_decap_8 FILLER_30_3277 ();
 sg13g2_decap_8 FILLER_30_3284 ();
 sg13g2_decap_8 FILLER_30_3291 ();
 sg13g2_decap_8 FILLER_30_3298 ();
 sg13g2_decap_8 FILLER_30_3305 ();
 sg13g2_decap_8 FILLER_30_3312 ();
 sg13g2_decap_8 FILLER_30_3319 ();
 sg13g2_decap_8 FILLER_30_3326 ();
 sg13g2_decap_8 FILLER_30_3333 ();
 sg13g2_decap_8 FILLER_30_3340 ();
 sg13g2_decap_8 FILLER_30_3347 ();
 sg13g2_decap_8 FILLER_30_3354 ();
 sg13g2_decap_8 FILLER_30_3361 ();
 sg13g2_decap_8 FILLER_30_3368 ();
 sg13g2_decap_8 FILLER_30_3375 ();
 sg13g2_decap_8 FILLER_30_3382 ();
 sg13g2_decap_8 FILLER_30_3389 ();
 sg13g2_decap_8 FILLER_30_3396 ();
 sg13g2_decap_8 FILLER_30_3403 ();
 sg13g2_decap_8 FILLER_30_3410 ();
 sg13g2_decap_8 FILLER_30_3417 ();
 sg13g2_decap_8 FILLER_30_3424 ();
 sg13g2_decap_8 FILLER_30_3431 ();
 sg13g2_decap_8 FILLER_30_3438 ();
 sg13g2_decap_8 FILLER_30_3445 ();
 sg13g2_decap_8 FILLER_30_3452 ();
 sg13g2_decap_8 FILLER_30_3459 ();
 sg13g2_decap_8 FILLER_30_3466 ();
 sg13g2_decap_8 FILLER_30_3473 ();
 sg13g2_decap_8 FILLER_30_3480 ();
 sg13g2_decap_8 FILLER_30_3487 ();
 sg13g2_decap_8 FILLER_30_3494 ();
 sg13g2_decap_8 FILLER_30_3501 ();
 sg13g2_decap_8 FILLER_30_3508 ();
 sg13g2_decap_8 FILLER_30_3515 ();
 sg13g2_decap_8 FILLER_30_3522 ();
 sg13g2_decap_8 FILLER_30_3529 ();
 sg13g2_decap_8 FILLER_30_3536 ();
 sg13g2_decap_8 FILLER_30_3543 ();
 sg13g2_decap_8 FILLER_30_3550 ();
 sg13g2_decap_8 FILLER_30_3557 ();
 sg13g2_decap_8 FILLER_30_3564 ();
 sg13g2_decap_8 FILLER_30_3571 ();
 sg13g2_fill_2 FILLER_30_3578 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_79 ();
 sg13g2_decap_8 FILLER_31_86 ();
 sg13g2_decap_4 FILLER_31_93 ();
 sg13g2_fill_2 FILLER_31_97 ();
 sg13g2_decap_8 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_152 ();
 sg13g2_decap_8 FILLER_31_159 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_fill_2 FILLER_31_180 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_255 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_decap_4 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_273 ();
 sg13g2_decap_4 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_335 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_366 ();
 sg13g2_decap_4 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_486 ();
 sg13g2_fill_2 FILLER_31_519 ();
 sg13g2_fill_2 FILLER_31_550 ();
 sg13g2_fill_1 FILLER_31_552 ();
 sg13g2_fill_2 FILLER_31_563 ();
 sg13g2_fill_1 FILLER_31_565 ();
 sg13g2_decap_8 FILLER_31_587 ();
 sg13g2_decap_8 FILLER_31_594 ();
 sg13g2_decap_8 FILLER_31_601 ();
 sg13g2_decap_8 FILLER_31_613 ();
 sg13g2_decap_8 FILLER_31_646 ();
 sg13g2_decap_8 FILLER_31_653 ();
 sg13g2_decap_4 FILLER_31_660 ();
 sg13g2_fill_2 FILLER_31_690 ();
 sg13g2_decap_8 FILLER_31_729 ();
 sg13g2_decap_8 FILLER_31_736 ();
 sg13g2_decap_8 FILLER_31_743 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_decap_8 FILLER_31_757 ();
 sg13g2_decap_8 FILLER_31_764 ();
 sg13g2_decap_8 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_778 ();
 sg13g2_fill_1 FILLER_31_785 ();
 sg13g2_fill_1 FILLER_31_789 ();
 sg13g2_fill_2 FILLER_31_794 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_849 ();
 sg13g2_decap_8 FILLER_31_856 ();
 sg13g2_decap_8 FILLER_31_863 ();
 sg13g2_decap_8 FILLER_31_870 ();
 sg13g2_decap_8 FILLER_31_887 ();
 sg13g2_decap_8 FILLER_31_894 ();
 sg13g2_decap_8 FILLER_31_901 ();
 sg13g2_decap_8 FILLER_31_908 ();
 sg13g2_fill_1 FILLER_31_915 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_fill_2 FILLER_31_945 ();
 sg13g2_fill_1 FILLER_31_947 ();
 sg13g2_decap_4 FILLER_31_953 ();
 sg13g2_decap_8 FILLER_31_972 ();
 sg13g2_decap_4 FILLER_31_979 ();
 sg13g2_fill_2 FILLER_31_983 ();
 sg13g2_decap_8 FILLER_31_1037 ();
 sg13g2_fill_2 FILLER_31_1044 ();
 sg13g2_fill_1 FILLER_31_1046 ();
 sg13g2_decap_8 FILLER_31_1076 ();
 sg13g2_fill_2 FILLER_31_1109 ();
 sg13g2_decap_8 FILLER_31_1137 ();
 sg13g2_decap_4 FILLER_31_1144 ();
 sg13g2_decap_4 FILLER_31_1184 ();
 sg13g2_fill_1 FILLER_31_1188 ();
 sg13g2_fill_2 FILLER_31_1241 ();
 sg13g2_decap_4 FILLER_31_1295 ();
 sg13g2_decap_4 FILLER_31_1302 ();
 sg13g2_fill_1 FILLER_31_1306 ();
 sg13g2_decap_8 FILLER_31_1345 ();
 sg13g2_fill_2 FILLER_31_1352 ();
 sg13g2_fill_2 FILLER_31_1406 ();
 sg13g2_fill_1 FILLER_31_1408 ();
 sg13g2_fill_1 FILLER_31_1440 ();
 sg13g2_fill_1 FILLER_31_1449 ();
 sg13g2_decap_8 FILLER_31_1455 ();
 sg13g2_fill_2 FILLER_31_1462 ();
 sg13g2_fill_2 FILLER_31_1499 ();
 sg13g2_fill_1 FILLER_31_1501 ();
 sg13g2_fill_2 FILLER_31_1522 ();
 sg13g2_fill_2 FILLER_31_1529 ();
 sg13g2_fill_1 FILLER_31_1531 ();
 sg13g2_decap_8 FILLER_31_1540 ();
 sg13g2_decap_8 FILLER_31_1547 ();
 sg13g2_decap_8 FILLER_31_1554 ();
 sg13g2_fill_2 FILLER_31_1561 ();
 sg13g2_decap_8 FILLER_31_1589 ();
 sg13g2_decap_8 FILLER_31_1596 ();
 sg13g2_decap_4 FILLER_31_1603 ();
 sg13g2_fill_1 FILLER_31_1607 ();
 sg13g2_decap_8 FILLER_31_1634 ();
 sg13g2_decap_8 FILLER_31_1641 ();
 sg13g2_decap_8 FILLER_31_1648 ();
 sg13g2_decap_8 FILLER_31_1655 ();
 sg13g2_fill_2 FILLER_31_1662 ();
 sg13g2_fill_1 FILLER_31_1664 ();
 sg13g2_decap_8 FILLER_31_1696 ();
 sg13g2_fill_1 FILLER_31_1732 ();
 sg13g2_decap_8 FILLER_31_1759 ();
 sg13g2_decap_8 FILLER_31_1766 ();
 sg13g2_fill_2 FILLER_31_1773 ();
 sg13g2_decap_8 FILLER_31_1801 ();
 sg13g2_fill_2 FILLER_31_1808 ();
 sg13g2_fill_1 FILLER_31_1810 ();
 sg13g2_decap_8 FILLER_31_1883 ();
 sg13g2_decap_8 FILLER_31_1890 ();
 sg13g2_fill_1 FILLER_31_1897 ();
 sg13g2_decap_8 FILLER_31_1924 ();
 sg13g2_decap_8 FILLER_31_1931 ();
 sg13g2_decap_4 FILLER_31_1938 ();
 sg13g2_fill_1 FILLER_31_1955 ();
 sg13g2_fill_1 FILLER_31_1982 ();
 sg13g2_decap_8 FILLER_31_2012 ();
 sg13g2_decap_8 FILLER_31_2123 ();
 sg13g2_decap_8 FILLER_31_2130 ();
 sg13g2_decap_8 FILLER_31_2137 ();
 sg13g2_fill_2 FILLER_31_2144 ();
 sg13g2_fill_1 FILLER_31_2146 ();
 sg13g2_decap_8 FILLER_31_2181 ();
 sg13g2_decap_8 FILLER_31_2248 ();
 sg13g2_decap_8 FILLER_31_2255 ();
 sg13g2_fill_2 FILLER_31_2262 ();
 sg13g2_decap_8 FILLER_31_2314 ();
 sg13g2_decap_8 FILLER_31_2321 ();
 sg13g2_decap_8 FILLER_31_2328 ();
 sg13g2_decap_4 FILLER_31_2335 ();
 sg13g2_fill_2 FILLER_31_2339 ();
 sg13g2_decap_8 FILLER_31_2381 ();
 sg13g2_decap_8 FILLER_31_2388 ();
 sg13g2_decap_8 FILLER_31_2395 ();
 sg13g2_decap_8 FILLER_31_2402 ();
 sg13g2_fill_2 FILLER_31_2409 ();
 sg13g2_fill_1 FILLER_31_2411 ();
 sg13g2_decap_4 FILLER_31_2463 ();
 sg13g2_fill_2 FILLER_31_2467 ();
 sg13g2_decap_4 FILLER_31_2521 ();
 sg13g2_fill_2 FILLER_31_2533 ();
 sg13g2_fill_1 FILLER_31_2535 ();
 sg13g2_decap_8 FILLER_31_2542 ();
 sg13g2_decap_8 FILLER_31_2549 ();
 sg13g2_fill_2 FILLER_31_2556 ();
 sg13g2_decap_8 FILLER_31_2584 ();
 sg13g2_decap_8 FILLER_31_2591 ();
 sg13g2_decap_4 FILLER_31_2598 ();
 sg13g2_fill_1 FILLER_31_2602 ();
 sg13g2_decap_8 FILLER_31_2629 ();
 sg13g2_decap_8 FILLER_31_2636 ();
 sg13g2_fill_2 FILLER_31_2643 ();
 sg13g2_fill_1 FILLER_31_2645 ();
 sg13g2_fill_1 FILLER_31_2672 ();
 sg13g2_fill_2 FILLER_31_2685 ();
 sg13g2_fill_1 FILLER_31_2687 ();
 sg13g2_fill_2 FILLER_31_2714 ();
 sg13g2_fill_1 FILLER_31_2716 ();
 sg13g2_fill_1 FILLER_31_2732 ();
 sg13g2_decap_4 FILLER_31_2759 ();
 sg13g2_decap_8 FILLER_31_2789 ();
 sg13g2_decap_8 FILLER_31_2796 ();
 sg13g2_decap_8 FILLER_31_2803 ();
 sg13g2_decap_8 FILLER_31_2810 ();
 sg13g2_decap_8 FILLER_31_2817 ();
 sg13g2_fill_1 FILLER_31_2845 ();
 sg13g2_decap_4 FILLER_31_2872 ();
 sg13g2_fill_2 FILLER_31_2876 ();
 sg13g2_decap_8 FILLER_31_2904 ();
 sg13g2_decap_4 FILLER_31_2911 ();
 sg13g2_decap_8 FILLER_31_2967 ();
 sg13g2_fill_2 FILLER_31_2974 ();
 sg13g2_fill_1 FILLER_31_2976 ();
 sg13g2_fill_1 FILLER_31_3029 ();
 sg13g2_decap_8 FILLER_31_3090 ();
 sg13g2_decap_8 FILLER_31_3097 ();
 sg13g2_decap_4 FILLER_31_3104 ();
 sg13g2_fill_1 FILLER_31_3108 ();
 sg13g2_decap_8 FILLER_31_3135 ();
 sg13g2_decap_8 FILLER_31_3147 ();
 sg13g2_fill_2 FILLER_31_3154 ();
 sg13g2_fill_2 FILLER_31_3182 ();
 sg13g2_fill_1 FILLER_31_3184 ();
 sg13g2_fill_2 FILLER_31_3198 ();
 sg13g2_decap_8 FILLER_31_3226 ();
 sg13g2_decap_8 FILLER_31_3233 ();
 sg13g2_decap_8 FILLER_31_3240 ();
 sg13g2_decap_8 FILLER_31_3247 ();
 sg13g2_decap_8 FILLER_31_3254 ();
 sg13g2_decap_8 FILLER_31_3261 ();
 sg13g2_decap_8 FILLER_31_3268 ();
 sg13g2_decap_8 FILLER_31_3275 ();
 sg13g2_decap_8 FILLER_31_3282 ();
 sg13g2_decap_8 FILLER_31_3289 ();
 sg13g2_decap_8 FILLER_31_3296 ();
 sg13g2_decap_8 FILLER_31_3303 ();
 sg13g2_decap_8 FILLER_31_3310 ();
 sg13g2_decap_8 FILLER_31_3317 ();
 sg13g2_decap_8 FILLER_31_3324 ();
 sg13g2_decap_8 FILLER_31_3331 ();
 sg13g2_decap_8 FILLER_31_3338 ();
 sg13g2_decap_8 FILLER_31_3345 ();
 sg13g2_decap_8 FILLER_31_3352 ();
 sg13g2_decap_8 FILLER_31_3359 ();
 sg13g2_decap_8 FILLER_31_3366 ();
 sg13g2_decap_8 FILLER_31_3373 ();
 sg13g2_decap_8 FILLER_31_3380 ();
 sg13g2_decap_8 FILLER_31_3387 ();
 sg13g2_decap_8 FILLER_31_3394 ();
 sg13g2_decap_8 FILLER_31_3401 ();
 sg13g2_decap_8 FILLER_31_3408 ();
 sg13g2_decap_8 FILLER_31_3415 ();
 sg13g2_decap_8 FILLER_31_3422 ();
 sg13g2_decap_8 FILLER_31_3429 ();
 sg13g2_decap_8 FILLER_31_3436 ();
 sg13g2_decap_8 FILLER_31_3443 ();
 sg13g2_decap_8 FILLER_31_3450 ();
 sg13g2_decap_8 FILLER_31_3457 ();
 sg13g2_decap_8 FILLER_31_3464 ();
 sg13g2_decap_8 FILLER_31_3471 ();
 sg13g2_decap_8 FILLER_31_3478 ();
 sg13g2_decap_8 FILLER_31_3485 ();
 sg13g2_decap_8 FILLER_31_3492 ();
 sg13g2_decap_8 FILLER_31_3499 ();
 sg13g2_decap_8 FILLER_31_3506 ();
 sg13g2_decap_8 FILLER_31_3513 ();
 sg13g2_decap_8 FILLER_31_3520 ();
 sg13g2_decap_8 FILLER_31_3527 ();
 sg13g2_decap_8 FILLER_31_3534 ();
 sg13g2_decap_8 FILLER_31_3541 ();
 sg13g2_decap_8 FILLER_31_3548 ();
 sg13g2_decap_8 FILLER_31_3555 ();
 sg13g2_decap_8 FILLER_31_3562 ();
 sg13g2_decap_8 FILLER_31_3569 ();
 sg13g2_decap_4 FILLER_31_3576 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_4 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_131 ();
 sg13g2_decap_8 FILLER_32_138 ();
 sg13g2_decap_8 FILLER_32_145 ();
 sg13g2_decap_8 FILLER_32_152 ();
 sg13g2_decap_8 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_4 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_fill_2 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_226 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_4 FILLER_32_266 ();
 sg13g2_fill_2 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_363 ();
 sg13g2_decap_8 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_32_377 ();
 sg13g2_decap_4 FILLER_32_384 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_4 FILLER_32_424 ();
 sg13g2_fill_2 FILLER_32_491 ();
 sg13g2_fill_1 FILLER_32_493 ();
 sg13g2_fill_2 FILLER_32_520 ();
 sg13g2_fill_1 FILLER_32_548 ();
 sg13g2_decap_8 FILLER_32_586 ();
 sg13g2_decap_4 FILLER_32_593 ();
 sg13g2_fill_1 FILLER_32_597 ();
 sg13g2_decap_4 FILLER_32_624 ();
 sg13g2_fill_1 FILLER_32_631 ();
 sg13g2_fill_2 FILLER_32_635 ();
 sg13g2_fill_1 FILLER_32_637 ();
 sg13g2_decap_4 FILLER_32_664 ();
 sg13g2_fill_1 FILLER_32_668 ();
 sg13g2_decap_8 FILLER_32_737 ();
 sg13g2_decap_8 FILLER_32_744 ();
 sg13g2_decap_4 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_768 ();
 sg13g2_decap_4 FILLER_32_775 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_fill_2 FILLER_32_812 ();
 sg13g2_fill_1 FILLER_32_814 ();
 sg13g2_decap_8 FILLER_32_849 ();
 sg13g2_decap_8 FILLER_32_856 ();
 sg13g2_decap_8 FILLER_32_889 ();
 sg13g2_decap_8 FILLER_32_896 ();
 sg13g2_fill_2 FILLER_32_903 ();
 sg13g2_fill_1 FILLER_32_905 ();
 sg13g2_fill_1 FILLER_32_911 ();
 sg13g2_decap_8 FILLER_32_943 ();
 sg13g2_decap_8 FILLER_32_950 ();
 sg13g2_fill_1 FILLER_32_957 ();
 sg13g2_decap_8 FILLER_32_984 ();
 sg13g2_decap_8 FILLER_32_991 ();
 sg13g2_decap_8 FILLER_32_998 ();
 sg13g2_decap_8 FILLER_32_1005 ();
 sg13g2_decap_8 FILLER_32_1038 ();
 sg13g2_fill_2 FILLER_32_1055 ();
 sg13g2_fill_2 FILLER_32_1083 ();
 sg13g2_fill_1 FILLER_32_1085 ();
 sg13g2_decap_4 FILLER_32_1138 ();
 sg13g2_decap_8 FILLER_32_1168 ();
 sg13g2_fill_1 FILLER_32_1175 ();
 sg13g2_fill_1 FILLER_32_1217 ();
 sg13g2_decap_4 FILLER_32_1310 ();
 sg13g2_fill_2 FILLER_32_1314 ();
 sg13g2_fill_2 FILLER_32_1324 ();
 sg13g2_fill_1 FILLER_32_1326 ();
 sg13g2_decap_8 FILLER_32_1353 ();
 sg13g2_decap_8 FILLER_32_1360 ();
 sg13g2_decap_8 FILLER_32_1400 ();
 sg13g2_decap_8 FILLER_32_1407 ();
 sg13g2_decap_4 FILLER_32_1414 ();
 sg13g2_fill_1 FILLER_32_1418 ();
 sg13g2_fill_1 FILLER_32_1423 ();
 sg13g2_fill_2 FILLER_32_1489 ();
 sg13g2_fill_1 FILLER_32_1491 ();
 sg13g2_fill_2 FILLER_32_1508 ();
 sg13g2_fill_1 FILLER_32_1510 ();
 sg13g2_decap_8 FILLER_32_1519 ();
 sg13g2_decap_8 FILLER_32_1526 ();
 sg13g2_decap_8 FILLER_32_1533 ();
 sg13g2_decap_8 FILLER_32_1540 ();
 sg13g2_decap_8 FILLER_32_1573 ();
 sg13g2_fill_1 FILLER_32_1580 ();
 sg13g2_decap_4 FILLER_32_1607 ();
 sg13g2_fill_2 FILLER_32_1611 ();
 sg13g2_decap_8 FILLER_32_1643 ();
 sg13g2_decap_4 FILLER_32_1706 ();
 sg13g2_fill_2 FILLER_32_1749 ();
 sg13g2_decap_8 FILLER_32_1803 ();
 sg13g2_decap_8 FILLER_32_1810 ();
 sg13g2_fill_2 FILLER_32_1817 ();
 sg13g2_decap_8 FILLER_32_1830 ();
 sg13g2_decap_8 FILLER_32_1837 ();
 sg13g2_decap_4 FILLER_32_1844 ();
 sg13g2_fill_1 FILLER_32_1848 ();
 sg13g2_decap_8 FILLER_32_1880 ();
 sg13g2_fill_2 FILLER_32_1887 ();
 sg13g2_fill_1 FILLER_32_1889 ();
 sg13g2_decap_8 FILLER_32_1922 ();
 sg13g2_decap_8 FILLER_32_1929 ();
 sg13g2_fill_2 FILLER_32_1936 ();
 sg13g2_fill_2 FILLER_32_1975 ();
 sg13g2_decap_8 FILLER_32_2003 ();
 sg13g2_decap_4 FILLER_32_2010 ();
 sg13g2_fill_1 FILLER_32_2066 ();
 sg13g2_decap_8 FILLER_32_2078 ();
 sg13g2_decap_4 FILLER_32_2085 ();
 sg13g2_decap_8 FILLER_32_2124 ();
 sg13g2_decap_8 FILLER_32_2131 ();
 sg13g2_fill_2 FILLER_32_2138 ();
 sg13g2_fill_1 FILLER_32_2140 ();
 sg13g2_decap_8 FILLER_32_2149 ();
 sg13g2_decap_8 FILLER_32_2156 ();
 sg13g2_decap_8 FILLER_32_2163 ();
 sg13g2_decap_8 FILLER_32_2170 ();
 sg13g2_decap_8 FILLER_32_2177 ();
 sg13g2_decap_8 FILLER_32_2184 ();
 sg13g2_decap_8 FILLER_32_2309 ();
 sg13g2_fill_2 FILLER_32_2316 ();
 sg13g2_decap_4 FILLER_32_2334 ();
 sg13g2_fill_1 FILLER_32_2338 ();
 sg13g2_decap_8 FILLER_32_2391 ();
 sg13g2_decap_8 FILLER_32_2398 ();
 sg13g2_decap_4 FILLER_32_2405 ();
 sg13g2_fill_2 FILLER_32_2435 ();
 sg13g2_fill_1 FILLER_32_2437 ();
 sg13g2_fill_2 FILLER_32_2470 ();
 sg13g2_fill_1 FILLER_32_2472 ();
 sg13g2_decap_8 FILLER_32_2550 ();
 sg13g2_fill_2 FILLER_32_2557 ();
 sg13g2_fill_1 FILLER_32_2559 ();
 sg13g2_decap_8 FILLER_32_2638 ();
 sg13g2_decap_4 FILLER_32_2645 ();
 sg13g2_fill_1 FILLER_32_2649 ();
 sg13g2_decap_8 FILLER_32_2685 ();
 sg13g2_decap_4 FILLER_32_2692 ();
 sg13g2_fill_2 FILLER_32_2696 ();
 sg13g2_fill_1 FILLER_32_2702 ();
 sg13g2_decap_8 FILLER_32_2707 ();
 sg13g2_fill_1 FILLER_32_2714 ();
 sg13g2_fill_2 FILLER_32_2720 ();
 sg13g2_decap_4 FILLER_32_2753 ();
 sg13g2_decap_8 FILLER_32_2783 ();
 sg13g2_decap_8 FILLER_32_2790 ();
 sg13g2_decap_8 FILLER_32_2797 ();
 sg13g2_decap_4 FILLER_32_2804 ();
 sg13g2_fill_1 FILLER_32_2808 ();
 sg13g2_fill_2 FILLER_32_2869 ();
 sg13g2_fill_1 FILLER_32_2871 ();
 sg13g2_decap_8 FILLER_32_2888 ();
 sg13g2_decap_8 FILLER_32_2895 ();
 sg13g2_decap_8 FILLER_32_2902 ();
 sg13g2_decap_4 FILLER_32_2909 ();
 sg13g2_decap_8 FILLER_32_2952 ();
 sg13g2_decap_8 FILLER_32_2959 ();
 sg13g2_decap_8 FILLER_32_2966 ();
 sg13g2_decap_8 FILLER_32_2973 ();
 sg13g2_fill_2 FILLER_32_2980 ();
 sg13g2_decap_8 FILLER_32_3018 ();
 sg13g2_decap_4 FILLER_32_3025 ();
 sg13g2_fill_2 FILLER_32_3029 ();
 sg13g2_fill_2 FILLER_32_3070 ();
 sg13g2_fill_1 FILLER_32_3072 ();
 sg13g2_decap_4 FILLER_32_3088 ();
 sg13g2_fill_2 FILLER_32_3092 ();
 sg13g2_decap_8 FILLER_32_3099 ();
 sg13g2_decap_8 FILLER_32_3106 ();
 sg13g2_decap_8 FILLER_32_3113 ();
 sg13g2_decap_8 FILLER_32_3120 ();
 sg13g2_decap_4 FILLER_32_3127 ();
 sg13g2_decap_4 FILLER_32_3154 ();
 sg13g2_fill_1 FILLER_32_3170 ();
 sg13g2_decap_8 FILLER_32_3223 ();
 sg13g2_decap_8 FILLER_32_3230 ();
 sg13g2_decap_8 FILLER_32_3237 ();
 sg13g2_decap_8 FILLER_32_3244 ();
 sg13g2_decap_8 FILLER_32_3251 ();
 sg13g2_decap_8 FILLER_32_3258 ();
 sg13g2_decap_8 FILLER_32_3265 ();
 sg13g2_decap_8 FILLER_32_3272 ();
 sg13g2_decap_8 FILLER_32_3279 ();
 sg13g2_decap_8 FILLER_32_3286 ();
 sg13g2_decap_8 FILLER_32_3293 ();
 sg13g2_decap_8 FILLER_32_3300 ();
 sg13g2_decap_8 FILLER_32_3307 ();
 sg13g2_decap_8 FILLER_32_3314 ();
 sg13g2_decap_8 FILLER_32_3321 ();
 sg13g2_decap_8 FILLER_32_3328 ();
 sg13g2_decap_8 FILLER_32_3335 ();
 sg13g2_decap_8 FILLER_32_3342 ();
 sg13g2_decap_8 FILLER_32_3349 ();
 sg13g2_decap_8 FILLER_32_3356 ();
 sg13g2_decap_8 FILLER_32_3363 ();
 sg13g2_decap_8 FILLER_32_3370 ();
 sg13g2_decap_8 FILLER_32_3377 ();
 sg13g2_decap_8 FILLER_32_3384 ();
 sg13g2_decap_8 FILLER_32_3391 ();
 sg13g2_decap_8 FILLER_32_3398 ();
 sg13g2_decap_8 FILLER_32_3405 ();
 sg13g2_decap_8 FILLER_32_3412 ();
 sg13g2_decap_8 FILLER_32_3419 ();
 sg13g2_decap_8 FILLER_32_3426 ();
 sg13g2_decap_8 FILLER_32_3433 ();
 sg13g2_decap_8 FILLER_32_3440 ();
 sg13g2_decap_8 FILLER_32_3447 ();
 sg13g2_decap_8 FILLER_32_3454 ();
 sg13g2_decap_8 FILLER_32_3461 ();
 sg13g2_decap_8 FILLER_32_3468 ();
 sg13g2_decap_8 FILLER_32_3475 ();
 sg13g2_decap_8 FILLER_32_3482 ();
 sg13g2_decap_8 FILLER_32_3489 ();
 sg13g2_decap_8 FILLER_32_3496 ();
 sg13g2_decap_8 FILLER_32_3503 ();
 sg13g2_decap_8 FILLER_32_3510 ();
 sg13g2_decap_8 FILLER_32_3517 ();
 sg13g2_decap_8 FILLER_32_3524 ();
 sg13g2_decap_8 FILLER_32_3531 ();
 sg13g2_decap_8 FILLER_32_3538 ();
 sg13g2_decap_8 FILLER_32_3545 ();
 sg13g2_decap_8 FILLER_32_3552 ();
 sg13g2_decap_8 FILLER_32_3559 ();
 sg13g2_decap_8 FILLER_32_3566 ();
 sg13g2_decap_8 FILLER_32_3573 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_78 ();
 sg13g2_decap_4 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_89 ();
 sg13g2_decap_8 FILLER_33_139 ();
 sg13g2_decap_8 FILLER_33_146 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_decap_8 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_decap_4 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_fill_2 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_fill_2 FILLER_33_422 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_fill_2 FILLER_33_441 ();
 sg13g2_decap_4 FILLER_33_451 ();
 sg13g2_fill_2 FILLER_33_455 ();
 sg13g2_fill_2 FILLER_33_465 ();
 sg13g2_fill_2 FILLER_33_480 ();
 sg13g2_decap_8 FILLER_33_512 ();
 sg13g2_decap_8 FILLER_33_519 ();
 sg13g2_decap_4 FILLER_33_591 ();
 sg13g2_decap_8 FILLER_33_736 ();
 sg13g2_decap_4 FILLER_33_743 ();
 sg13g2_fill_1 FILLER_33_747 ();
 sg13g2_decap_8 FILLER_33_774 ();
 sg13g2_fill_1 FILLER_33_781 ();
 sg13g2_decap_8 FILLER_33_850 ();
 sg13g2_decap_8 FILLER_33_857 ();
 sg13g2_decap_8 FILLER_33_864 ();
 sg13g2_decap_4 FILLER_33_871 ();
 sg13g2_fill_1 FILLER_33_875 ();
 sg13g2_fill_1 FILLER_33_880 ();
 sg13g2_decap_8 FILLER_33_886 ();
 sg13g2_fill_1 FILLER_33_893 ();
 sg13g2_decap_8 FILLER_33_946 ();
 sg13g2_decap_8 FILLER_33_953 ();
 sg13g2_fill_2 FILLER_33_960 ();
 sg13g2_fill_1 FILLER_33_962 ();
 sg13g2_decap_8 FILLER_33_989 ();
 sg13g2_decap_8 FILLER_33_996 ();
 sg13g2_decap_8 FILLER_33_1003 ();
 sg13g2_fill_2 FILLER_33_1010 ();
 sg13g2_fill_1 FILLER_33_1012 ();
 sg13g2_decap_8 FILLER_33_1077 ();
 sg13g2_fill_1 FILLER_33_1123 ();
 sg13g2_fill_1 FILLER_33_1134 ();
 sg13g2_decap_8 FILLER_33_1139 ();
 sg13g2_decap_4 FILLER_33_1146 ();
 sg13g2_fill_2 FILLER_33_1150 ();
 sg13g2_decap_8 FILLER_33_1162 ();
 sg13g2_fill_2 FILLER_33_1169 ();
 sg13g2_fill_1 FILLER_33_1171 ();
 sg13g2_decap_8 FILLER_33_1206 ();
 sg13g2_fill_2 FILLER_33_1213 ();
 sg13g2_fill_1 FILLER_33_1215 ();
 sg13g2_fill_1 FILLER_33_1248 ();
 sg13g2_fill_2 FILLER_33_1254 ();
 sg13g2_fill_1 FILLER_33_1261 ();
 sg13g2_decap_4 FILLER_33_1294 ();
 sg13g2_fill_1 FILLER_33_1298 ();
 sg13g2_decap_8 FILLER_33_1302 ();
 sg13g2_decap_8 FILLER_33_1309 ();
 sg13g2_decap_8 FILLER_33_1316 ();
 sg13g2_fill_2 FILLER_33_1341 ();
 sg13g2_fill_1 FILLER_33_1343 ();
 sg13g2_decap_8 FILLER_33_1351 ();
 sg13g2_fill_2 FILLER_33_1358 ();
 sg13g2_fill_1 FILLER_33_1360 ();
 sg13g2_decap_8 FILLER_33_1397 ();
 sg13g2_decap_8 FILLER_33_1404 ();
 sg13g2_decap_8 FILLER_33_1411 ();
 sg13g2_decap_4 FILLER_33_1418 ();
 sg13g2_fill_2 FILLER_33_1422 ();
 sg13g2_decap_8 FILLER_33_1427 ();
 sg13g2_fill_2 FILLER_33_1500 ();
 sg13g2_decap_8 FILLER_33_1528 ();
 sg13g2_decap_8 FILLER_33_1535 ();
 sg13g2_fill_1 FILLER_33_1542 ();
 sg13g2_fill_1 FILLER_33_1595 ();
 sg13g2_fill_1 FILLER_33_1705 ();
 sg13g2_decap_8 FILLER_33_1710 ();
 sg13g2_decap_4 FILLER_33_1717 ();
 sg13g2_fill_2 FILLER_33_1726 ();
 sg13g2_fill_1 FILLER_33_1728 ();
 sg13g2_decap_8 FILLER_33_1759 ();
 sg13g2_decap_8 FILLER_33_1766 ();
 sg13g2_fill_1 FILLER_33_1773 ();
 sg13g2_decap_4 FILLER_33_1816 ();
 sg13g2_decap_8 FILLER_33_1846 ();
 sg13g2_decap_8 FILLER_33_1853 ();
 sg13g2_decap_8 FILLER_33_1860 ();
 sg13g2_decap_8 FILLER_33_1867 ();
 sg13g2_decap_8 FILLER_33_1874 ();
 sg13g2_decap_8 FILLER_33_1881 ();
 sg13g2_fill_2 FILLER_33_1888 ();
 sg13g2_decap_8 FILLER_33_1916 ();
 sg13g2_decap_4 FILLER_33_1923 ();
 sg13g2_fill_1 FILLER_33_1927 ();
 sg13g2_decap_8 FILLER_33_1990 ();
 sg13g2_decap_8 FILLER_33_1997 ();
 sg13g2_decap_8 FILLER_33_2004 ();
 sg13g2_decap_8 FILLER_33_2011 ();
 sg13g2_fill_1 FILLER_33_2018 ();
 sg13g2_decap_8 FILLER_33_2028 ();
 sg13g2_decap_8 FILLER_33_2035 ();
 sg13g2_decap_8 FILLER_33_2042 ();
 sg13g2_fill_2 FILLER_33_2075 ();
 sg13g2_decap_8 FILLER_33_2085 ();
 sg13g2_decap_8 FILLER_33_2092 ();
 sg13g2_fill_2 FILLER_33_2099 ();
 sg13g2_fill_1 FILLER_33_2101 ();
 sg13g2_decap_8 FILLER_33_2128 ();
 sg13g2_decap_8 FILLER_33_2135 ();
 sg13g2_decap_8 FILLER_33_2142 ();
 sg13g2_decap_8 FILLER_33_2149 ();
 sg13g2_decap_8 FILLER_33_2156 ();
 sg13g2_fill_1 FILLER_33_2163 ();
 sg13g2_decap_8 FILLER_33_2172 ();
 sg13g2_decap_8 FILLER_33_2179 ();
 sg13g2_decap_8 FILLER_33_2186 ();
 sg13g2_decap_8 FILLER_33_2193 ();
 sg13g2_fill_2 FILLER_33_2200 ();
 sg13g2_decap_8 FILLER_33_2237 ();
 sg13g2_decap_8 FILLER_33_2244 ();
 sg13g2_decap_8 FILLER_33_2251 ();
 sg13g2_decap_8 FILLER_33_2258 ();
 sg13g2_fill_2 FILLER_33_2265 ();
 sg13g2_decap_8 FILLER_33_2298 ();
 sg13g2_decap_8 FILLER_33_2305 ();
 sg13g2_decap_8 FILLER_33_2312 ();
 sg13g2_decap_8 FILLER_33_2319 ();
 sg13g2_fill_1 FILLER_33_2326 ();
 sg13g2_decap_8 FILLER_33_2385 ();
 sg13g2_decap_8 FILLER_33_2392 ();
 sg13g2_decap_8 FILLER_33_2399 ();
 sg13g2_fill_2 FILLER_33_2406 ();
 sg13g2_fill_1 FILLER_33_2408 ();
 sg13g2_decap_8 FILLER_33_2422 ();
 sg13g2_decap_8 FILLER_33_2455 ();
 sg13g2_fill_2 FILLER_33_2462 ();
 sg13g2_decap_8 FILLER_33_2467 ();
 sg13g2_fill_2 FILLER_33_2474 ();
 sg13g2_fill_1 FILLER_33_2476 ();
 sg13g2_decap_4 FILLER_33_2552 ();
 sg13g2_fill_1 FILLER_33_2556 ();
 sg13g2_decap_4 FILLER_33_2617 ();
 sg13g2_fill_2 FILLER_33_2621 ();
 sg13g2_fill_2 FILLER_33_2649 ();
 sg13g2_fill_1 FILLER_33_2697 ();
 sg13g2_decap_8 FILLER_33_2706 ();
 sg13g2_decap_8 FILLER_33_2713 ();
 sg13g2_decap_8 FILLER_33_2720 ();
 sg13g2_decap_4 FILLER_33_2727 ();
 sg13g2_fill_2 FILLER_33_2731 ();
 sg13g2_decap_4 FILLER_33_2755 ();
 sg13g2_fill_1 FILLER_33_2759 ();
 sg13g2_fill_2 FILLER_33_2786 ();
 sg13g2_fill_1 FILLER_33_2788 ();
 sg13g2_decap_8 FILLER_33_2794 ();
 sg13g2_decap_8 FILLER_33_2801 ();
 sg13g2_decap_8 FILLER_33_2808 ();
 sg13g2_decap_8 FILLER_33_2815 ();
 sg13g2_decap_4 FILLER_33_2822 ();
 sg13g2_fill_1 FILLER_33_2826 ();
 sg13g2_fill_2 FILLER_33_2839 ();
 sg13g2_fill_1 FILLER_33_2841 ();
 sg13g2_decap_8 FILLER_33_2862 ();
 sg13g2_decap_8 FILLER_33_2869 ();
 sg13g2_decap_8 FILLER_33_2876 ();
 sg13g2_decap_8 FILLER_33_2883 ();
 sg13g2_decap_8 FILLER_33_2890 ();
 sg13g2_decap_8 FILLER_33_2897 ();
 sg13g2_decap_8 FILLER_33_2904 ();
 sg13g2_decap_4 FILLER_33_2911 ();
 sg13g2_fill_2 FILLER_33_2915 ();
 sg13g2_decap_8 FILLER_33_2959 ();
 sg13g2_fill_2 FILLER_33_2966 ();
 sg13g2_fill_1 FILLER_33_2968 ();
 sg13g2_decap_8 FILLER_33_2974 ();
 sg13g2_decap_4 FILLER_33_2981 ();
 sg13g2_fill_2 FILLER_33_2985 ();
 sg13g2_fill_1 FILLER_33_3004 ();
 sg13g2_decap_8 FILLER_33_3013 ();
 sg13g2_decap_8 FILLER_33_3020 ();
 sg13g2_decap_8 FILLER_33_3027 ();
 sg13g2_decap_4 FILLER_33_3034 ();
 sg13g2_fill_2 FILLER_33_3038 ();
 sg13g2_decap_8 FILLER_33_3045 ();
 sg13g2_fill_2 FILLER_33_3052 ();
 sg13g2_decap_4 FILLER_33_3062 ();
 sg13g2_fill_2 FILLER_33_3066 ();
 sg13g2_fill_2 FILLER_33_3094 ();
 sg13g2_decap_8 FILLER_33_3112 ();
 sg13g2_fill_2 FILLER_33_3119 ();
 sg13g2_fill_1 FILLER_33_3121 ();
 sg13g2_fill_2 FILLER_33_3130 ();
 sg13g2_decap_8 FILLER_33_3202 ();
 sg13g2_decap_8 FILLER_33_3209 ();
 sg13g2_decap_8 FILLER_33_3216 ();
 sg13g2_fill_2 FILLER_33_3223 ();
 sg13g2_fill_1 FILLER_33_3225 ();
 sg13g2_fill_2 FILLER_33_3232 ();
 sg13g2_decap_8 FILLER_33_3245 ();
 sg13g2_decap_8 FILLER_33_3252 ();
 sg13g2_decap_8 FILLER_33_3259 ();
 sg13g2_decap_8 FILLER_33_3266 ();
 sg13g2_decap_8 FILLER_33_3273 ();
 sg13g2_decap_8 FILLER_33_3280 ();
 sg13g2_decap_8 FILLER_33_3287 ();
 sg13g2_decap_8 FILLER_33_3294 ();
 sg13g2_decap_8 FILLER_33_3301 ();
 sg13g2_decap_8 FILLER_33_3308 ();
 sg13g2_decap_8 FILLER_33_3315 ();
 sg13g2_decap_8 FILLER_33_3322 ();
 sg13g2_decap_8 FILLER_33_3329 ();
 sg13g2_decap_8 FILLER_33_3336 ();
 sg13g2_decap_8 FILLER_33_3343 ();
 sg13g2_decap_8 FILLER_33_3350 ();
 sg13g2_decap_8 FILLER_33_3357 ();
 sg13g2_decap_8 FILLER_33_3364 ();
 sg13g2_decap_8 FILLER_33_3371 ();
 sg13g2_decap_8 FILLER_33_3378 ();
 sg13g2_decap_8 FILLER_33_3385 ();
 sg13g2_decap_8 FILLER_33_3392 ();
 sg13g2_decap_8 FILLER_33_3399 ();
 sg13g2_decap_8 FILLER_33_3406 ();
 sg13g2_decap_8 FILLER_33_3413 ();
 sg13g2_decap_8 FILLER_33_3420 ();
 sg13g2_decap_8 FILLER_33_3427 ();
 sg13g2_decap_8 FILLER_33_3434 ();
 sg13g2_decap_8 FILLER_33_3441 ();
 sg13g2_decap_8 FILLER_33_3448 ();
 sg13g2_decap_8 FILLER_33_3455 ();
 sg13g2_decap_8 FILLER_33_3462 ();
 sg13g2_decap_8 FILLER_33_3469 ();
 sg13g2_decap_8 FILLER_33_3476 ();
 sg13g2_decap_8 FILLER_33_3483 ();
 sg13g2_decap_8 FILLER_33_3490 ();
 sg13g2_decap_8 FILLER_33_3497 ();
 sg13g2_decap_8 FILLER_33_3504 ();
 sg13g2_decap_8 FILLER_33_3511 ();
 sg13g2_decap_8 FILLER_33_3518 ();
 sg13g2_decap_8 FILLER_33_3525 ();
 sg13g2_decap_8 FILLER_33_3532 ();
 sg13g2_decap_8 FILLER_33_3539 ();
 sg13g2_decap_8 FILLER_33_3546 ();
 sg13g2_decap_8 FILLER_33_3553 ();
 sg13g2_decap_8 FILLER_33_3560 ();
 sg13g2_decap_8 FILLER_33_3567 ();
 sg13g2_decap_4 FILLER_33_3574 ();
 sg13g2_fill_2 FILLER_33_3578 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_decap_8 FILLER_34_304 ();
 sg13g2_decap_8 FILLER_34_311 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_fill_2 FILLER_34_397 ();
 sg13g2_decap_4 FILLER_34_451 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_4 FILLER_34_483 ();
 sg13g2_fill_1 FILLER_34_487 ();
 sg13g2_decap_4 FILLER_34_518 ();
 sg13g2_fill_1 FILLER_34_522 ();
 sg13g2_decap_8 FILLER_34_526 ();
 sg13g2_decap_8 FILLER_34_533 ();
 sg13g2_fill_2 FILLER_34_540 ();
 sg13g2_fill_1 FILLER_34_542 ();
 sg13g2_fill_2 FILLER_34_549 ();
 sg13g2_fill_1 FILLER_34_551 ();
 sg13g2_decap_8 FILLER_34_598 ();
 sg13g2_decap_8 FILLER_34_605 ();
 sg13g2_decap_8 FILLER_34_612 ();
 sg13g2_decap_4 FILLER_34_619 ();
 sg13g2_fill_1 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_650 ();
 sg13g2_fill_2 FILLER_34_657 ();
 sg13g2_fill_1 FILLER_34_659 ();
 sg13g2_decap_4 FILLER_34_691 ();
 sg13g2_fill_2 FILLER_34_695 ();
 sg13g2_fill_1 FILLER_34_706 ();
 sg13g2_fill_1 FILLER_34_719 ();
 sg13g2_fill_1 FILLER_34_786 ();
 sg13g2_fill_1 FILLER_34_792 ();
 sg13g2_decap_8 FILLER_34_838 ();
 sg13g2_decap_8 FILLER_34_845 ();
 sg13g2_decap_8 FILLER_34_852 ();
 sg13g2_fill_1 FILLER_34_911 ();
 sg13g2_decap_8 FILLER_34_1000 ();
 sg13g2_decap_8 FILLER_34_1007 ();
 sg13g2_fill_1 FILLER_34_1022 ();
 sg13g2_fill_1 FILLER_34_1054 ();
 sg13g2_decap_4 FILLER_34_1063 ();
 sg13g2_fill_2 FILLER_34_1075 ();
 sg13g2_fill_2 FILLER_34_1128 ();
 sg13g2_fill_1 FILLER_34_1130 ();
 sg13g2_decap_8 FILLER_34_1148 ();
 sg13g2_fill_2 FILLER_34_1155 ();
 sg13g2_decap_8 FILLER_34_1192 ();
 sg13g2_decap_8 FILLER_34_1199 ();
 sg13g2_fill_2 FILLER_34_1206 ();
 sg13g2_fill_2 FILLER_34_1247 ();
 sg13g2_fill_2 FILLER_34_1252 ();
 sg13g2_decap_8 FILLER_34_1262 ();
 sg13g2_fill_2 FILLER_34_1269 ();
 sg13g2_decap_8 FILLER_34_1284 ();
 sg13g2_decap_8 FILLER_34_1291 ();
 sg13g2_fill_1 FILLER_34_1298 ();
 sg13g2_fill_2 FILLER_34_1328 ();
 sg13g2_decap_8 FILLER_34_1349 ();
 sg13g2_decap_8 FILLER_34_1356 ();
 sg13g2_decap_8 FILLER_34_1363 ();
 sg13g2_decap_4 FILLER_34_1370 ();
 sg13g2_fill_2 FILLER_34_1374 ();
 sg13g2_fill_1 FILLER_34_1384 ();
 sg13g2_decap_8 FILLER_34_1388 ();
 sg13g2_fill_1 FILLER_34_1395 ();
 sg13g2_decap_8 FILLER_34_1422 ();
 sg13g2_fill_1 FILLER_34_1429 ();
 sg13g2_decap_8 FILLER_34_1440 ();
 sg13g2_decap_8 FILLER_34_1447 ();
 sg13g2_decap_8 FILLER_34_1454 ();
 sg13g2_fill_2 FILLER_34_1461 ();
 sg13g2_fill_1 FILLER_34_1463 ();
 sg13g2_decap_4 FILLER_34_1472 ();
 sg13g2_fill_2 FILLER_34_1479 ();
 sg13g2_decap_4 FILLER_34_1507 ();
 sg13g2_fill_2 FILLER_34_1511 ();
 sg13g2_decap_8 FILLER_34_1543 ();
 sg13g2_decap_4 FILLER_34_1550 ();
 sg13g2_fill_2 FILLER_34_1554 ();
 sg13g2_decap_8 FILLER_34_1564 ();
 sg13g2_fill_1 FILLER_34_1571 ();
 sg13g2_decap_8 FILLER_34_1632 ();
 sg13g2_decap_8 FILLER_34_1639 ();
 sg13g2_decap_8 FILLER_34_1646 ();
 sg13g2_decap_8 FILLER_34_1653 ();
 sg13g2_decap_4 FILLER_34_1666 ();
 sg13g2_fill_1 FILLER_34_1696 ();
 sg13g2_decap_8 FILLER_34_1709 ();
 sg13g2_fill_2 FILLER_34_1727 ();
 sg13g2_fill_2 FILLER_34_1738 ();
 sg13g2_fill_1 FILLER_34_1740 ();
 sg13g2_fill_2 FILLER_34_1746 ();
 sg13g2_fill_1 FILLER_34_1748 ();
 sg13g2_fill_1 FILLER_34_1755 ();
 sg13g2_decap_8 FILLER_34_1808 ();
 sg13g2_decap_8 FILLER_34_1815 ();
 sg13g2_decap_8 FILLER_34_1822 ();
 sg13g2_decap_8 FILLER_34_1829 ();
 sg13g2_decap_4 FILLER_34_1836 ();
 sg13g2_fill_2 FILLER_34_1840 ();
 sg13g2_decap_8 FILLER_34_1847 ();
 sg13g2_decap_8 FILLER_34_1870 ();
 sg13g2_decap_8 FILLER_34_1877 ();
 sg13g2_decap_8 FILLER_34_1884 ();
 sg13g2_decap_8 FILLER_34_1891 ();
 sg13g2_fill_2 FILLER_34_1898 ();
 sg13g2_fill_2 FILLER_34_1909 ();
 sg13g2_decap_8 FILLER_34_1919 ();
 sg13g2_decap_8 FILLER_34_1926 ();
 sg13g2_fill_2 FILLER_34_1933 ();
 sg13g2_decap_4 FILLER_34_1945 ();
 sg13g2_fill_2 FILLER_34_1949 ();
 sg13g2_fill_2 FILLER_34_1980 ();
 sg13g2_fill_1 FILLER_34_1982 ();
 sg13g2_decap_8 FILLER_34_1987 ();
 sg13g2_decap_8 FILLER_34_1994 ();
 sg13g2_decap_8 FILLER_34_2001 ();
 sg13g2_fill_2 FILLER_34_2008 ();
 sg13g2_decap_4 FILLER_34_2032 ();
 sg13g2_fill_1 FILLER_34_2036 ();
 sg13g2_decap_8 FILLER_34_2042 ();
 sg13g2_decap_8 FILLER_34_2049 ();
 sg13g2_fill_1 FILLER_34_2056 ();
 sg13g2_fill_1 FILLER_34_2070 ();
 sg13g2_decap_8 FILLER_34_2076 ();
 sg13g2_fill_2 FILLER_34_2083 ();
 sg13g2_fill_1 FILLER_34_2085 ();
 sg13g2_decap_4 FILLER_34_2121 ();
 sg13g2_decap_4 FILLER_34_2203 ();
 sg13g2_fill_2 FILLER_34_2207 ();
 sg13g2_decap_8 FILLER_34_2240 ();
 sg13g2_decap_8 FILLER_34_2247 ();
 sg13g2_decap_8 FILLER_34_2254 ();
 sg13g2_decap_8 FILLER_34_2261 ();
 sg13g2_fill_2 FILLER_34_2268 ();
 sg13g2_fill_1 FILLER_34_2270 ();
 sg13g2_fill_1 FILLER_34_2289 ();
 sg13g2_decap_8 FILLER_34_2316 ();
 sg13g2_decap_8 FILLER_34_2323 ();
 sg13g2_decap_4 FILLER_34_2330 ();
 sg13g2_fill_1 FILLER_34_2334 ();
 sg13g2_decap_4 FILLER_34_2387 ();
 sg13g2_fill_2 FILLER_34_2391 ();
 sg13g2_decap_4 FILLER_34_2401 ();
 sg13g2_fill_1 FILLER_34_2405 ();
 sg13g2_decap_8 FILLER_34_2411 ();
 sg13g2_fill_1 FILLER_34_2418 ();
 sg13g2_decap_4 FILLER_34_2458 ();
 sg13g2_fill_2 FILLER_34_2462 ();
 sg13g2_decap_8 FILLER_34_2471 ();
 sg13g2_decap_4 FILLER_34_2478 ();
 sg13g2_fill_1 FILLER_34_2482 ();
 sg13g2_decap_8 FILLER_34_2553 ();
 sg13g2_fill_1 FILLER_34_2594 ();
 sg13g2_decap_8 FILLER_34_2600 ();
 sg13g2_decap_8 FILLER_34_2607 ();
 sg13g2_decap_8 FILLER_34_2614 ();
 sg13g2_fill_2 FILLER_34_2621 ();
 sg13g2_decap_8 FILLER_34_2654 ();
 sg13g2_decap_4 FILLER_34_2661 ();
 sg13g2_fill_2 FILLER_34_2682 ();
 sg13g2_decap_8 FILLER_34_2714 ();
 sg13g2_fill_2 FILLER_34_2721 ();
 sg13g2_fill_1 FILLER_34_2723 ();
 sg13g2_decap_8 FILLER_34_2732 ();
 sg13g2_decap_4 FILLER_34_2744 ();
 sg13g2_fill_1 FILLER_34_2774 ();
 sg13g2_fill_2 FILLER_34_2835 ();
 sg13g2_fill_1 FILLER_34_2837 ();
 sg13g2_decap_8 FILLER_34_2864 ();
 sg13g2_decap_4 FILLER_34_2871 ();
 sg13g2_decap_8 FILLER_34_2901 ();
 sg13g2_decap_8 FILLER_34_2908 ();
 sg13g2_fill_1 FILLER_34_2915 ();
 sg13g2_decap_4 FILLER_34_2962 ();
 sg13g2_decap_4 FILLER_34_3076 ();
 sg13g2_fill_1 FILLER_34_3106 ();
 sg13g2_decap_8 FILLER_34_3185 ();
 sg13g2_decap_8 FILLER_34_3192 ();
 sg13g2_decap_8 FILLER_34_3199 ();
 sg13g2_decap_4 FILLER_34_3206 ();
 sg13g2_fill_2 FILLER_34_3210 ();
 sg13g2_fill_1 FILLER_34_3217 ();
 sg13g2_fill_2 FILLER_34_3223 ();
 sg13g2_decap_8 FILLER_34_3251 ();
 sg13g2_decap_8 FILLER_34_3258 ();
 sg13g2_decap_8 FILLER_34_3265 ();
 sg13g2_decap_8 FILLER_34_3272 ();
 sg13g2_decap_8 FILLER_34_3279 ();
 sg13g2_decap_8 FILLER_34_3286 ();
 sg13g2_decap_8 FILLER_34_3293 ();
 sg13g2_decap_8 FILLER_34_3300 ();
 sg13g2_decap_8 FILLER_34_3307 ();
 sg13g2_decap_8 FILLER_34_3314 ();
 sg13g2_decap_8 FILLER_34_3321 ();
 sg13g2_decap_8 FILLER_34_3328 ();
 sg13g2_decap_8 FILLER_34_3335 ();
 sg13g2_decap_8 FILLER_34_3342 ();
 sg13g2_decap_8 FILLER_34_3349 ();
 sg13g2_decap_8 FILLER_34_3356 ();
 sg13g2_decap_8 FILLER_34_3363 ();
 sg13g2_decap_8 FILLER_34_3370 ();
 sg13g2_decap_8 FILLER_34_3377 ();
 sg13g2_decap_8 FILLER_34_3384 ();
 sg13g2_decap_8 FILLER_34_3391 ();
 sg13g2_decap_8 FILLER_34_3398 ();
 sg13g2_decap_8 FILLER_34_3405 ();
 sg13g2_decap_8 FILLER_34_3412 ();
 sg13g2_decap_8 FILLER_34_3419 ();
 sg13g2_decap_8 FILLER_34_3426 ();
 sg13g2_decap_8 FILLER_34_3433 ();
 sg13g2_decap_8 FILLER_34_3440 ();
 sg13g2_decap_8 FILLER_34_3447 ();
 sg13g2_decap_8 FILLER_34_3454 ();
 sg13g2_decap_8 FILLER_34_3461 ();
 sg13g2_decap_8 FILLER_34_3468 ();
 sg13g2_decap_8 FILLER_34_3475 ();
 sg13g2_decap_8 FILLER_34_3482 ();
 sg13g2_decap_8 FILLER_34_3489 ();
 sg13g2_decap_8 FILLER_34_3496 ();
 sg13g2_decap_8 FILLER_34_3503 ();
 sg13g2_decap_8 FILLER_34_3510 ();
 sg13g2_decap_8 FILLER_34_3517 ();
 sg13g2_decap_8 FILLER_34_3524 ();
 sg13g2_decap_8 FILLER_34_3531 ();
 sg13g2_decap_8 FILLER_34_3538 ();
 sg13g2_decap_8 FILLER_34_3545 ();
 sg13g2_decap_8 FILLER_34_3552 ();
 sg13g2_decap_8 FILLER_34_3559 ();
 sg13g2_decap_8 FILLER_34_3566 ();
 sg13g2_decap_8 FILLER_34_3573 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_fill_2 FILLER_35_94 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_1 FILLER_35_113 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_decap_4 FILLER_35_186 ();
 sg13g2_fill_1 FILLER_35_190 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_decap_8 FILLER_35_253 ();
 sg13g2_decap_4 FILLER_35_260 ();
 sg13g2_fill_2 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_4 FILLER_35_396 ();
 sg13g2_fill_1 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_453 ();
 sg13g2_decap_8 FILLER_35_479 ();
 sg13g2_decap_8 FILLER_35_486 ();
 sg13g2_fill_2 FILLER_35_493 ();
 sg13g2_fill_1 FILLER_35_495 ();
 sg13g2_decap_8 FILLER_35_526 ();
 sg13g2_decap_8 FILLER_35_533 ();
 sg13g2_decap_8 FILLER_35_551 ();
 sg13g2_fill_1 FILLER_35_558 ();
 sg13g2_decap_8 FILLER_35_585 ();
 sg13g2_decap_4 FILLER_35_592 ();
 sg13g2_decap_8 FILLER_35_656 ();
 sg13g2_decap_4 FILLER_35_663 ();
 sg13g2_fill_2 FILLER_35_680 ();
 sg13g2_fill_1 FILLER_35_682 ();
 sg13g2_fill_2 FILLER_35_692 ();
 sg13g2_decap_4 FILLER_35_703 ();
 sg13g2_fill_1 FILLER_35_711 ();
 sg13g2_decap_4 FILLER_35_722 ();
 sg13g2_fill_1 FILLER_35_726 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_4 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_780 ();
 sg13g2_fill_2 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_832 ();
 sg13g2_decap_8 FILLER_35_839 ();
 sg13g2_decap_8 FILLER_35_846 ();
 sg13g2_decap_8 FILLER_35_853 ();
 sg13g2_decap_8 FILLER_35_860 ();
 sg13g2_decap_4 FILLER_35_875 ();
 sg13g2_fill_1 FILLER_35_879 ();
 sg13g2_fill_2 FILLER_35_906 ();
 sg13g2_fill_1 FILLER_35_908 ();
 sg13g2_fill_1 FILLER_35_948 ();
 sg13g2_fill_2 FILLER_35_1000 ();
 sg13g2_fill_1 FILLER_35_1002 ();
 sg13g2_fill_2 FILLER_35_1008 ();
 sg13g2_fill_2 FILLER_35_1015 ();
 sg13g2_decap_4 FILLER_35_1021 ();
 sg13g2_fill_1 FILLER_35_1025 ();
 sg13g2_decap_4 FILLER_35_1029 ();
 sg13g2_fill_1 FILLER_35_1033 ();
 sg13g2_decap_4 FILLER_35_1042 ();
 sg13g2_decap_8 FILLER_35_1057 ();
 sg13g2_decap_8 FILLER_35_1064 ();
 sg13g2_decap_8 FILLER_35_1071 ();
 sg13g2_decap_8 FILLER_35_1078 ();
 sg13g2_decap_4 FILLER_35_1085 ();
 sg13g2_decap_8 FILLER_35_1120 ();
 sg13g2_decap_8 FILLER_35_1131 ();
 sg13g2_fill_2 FILLER_35_1162 ();
 sg13g2_fill_1 FILLER_35_1185 ();
 sg13g2_decap_8 FILLER_35_1202 ();
 sg13g2_decap_8 FILLER_35_1209 ();
 sg13g2_decap_8 FILLER_35_1216 ();
 sg13g2_decap_8 FILLER_35_1223 ();
 sg13g2_decap_8 FILLER_35_1230 ();
 sg13g2_decap_4 FILLER_35_1237 ();
 sg13g2_fill_1 FILLER_35_1241 ();
 sg13g2_fill_2 FILLER_35_1245 ();
 sg13g2_decap_8 FILLER_35_1252 ();
 sg13g2_decap_4 FILLER_35_1259 ();
 sg13g2_fill_1 FILLER_35_1263 ();
 sg13g2_decap_8 FILLER_35_1268 ();
 sg13g2_decap_8 FILLER_35_1275 ();
 sg13g2_decap_8 FILLER_35_1282 ();
 sg13g2_decap_8 FILLER_35_1289 ();
 sg13g2_decap_8 FILLER_35_1296 ();
 sg13g2_decap_8 FILLER_35_1303 ();
 sg13g2_fill_1 FILLER_35_1310 ();
 sg13g2_fill_1 FILLER_35_1335 ();
 sg13g2_decap_8 FILLER_35_1353 ();
 sg13g2_decap_8 FILLER_35_1360 ();
 sg13g2_fill_2 FILLER_35_1367 ();
 sg13g2_fill_1 FILLER_35_1377 ();
 sg13g2_decap_8 FILLER_35_1404 ();
 sg13g2_decap_4 FILLER_35_1411 ();
 sg13g2_fill_1 FILLER_35_1415 ();
 sg13g2_fill_2 FILLER_35_1429 ();
 sg13g2_fill_1 FILLER_35_1431 ();
 sg13g2_fill_2 FILLER_35_1437 ();
 sg13g2_decap_8 FILLER_35_1455 ();
 sg13g2_decap_8 FILLER_35_1462 ();
 sg13g2_decap_8 FILLER_35_1469 ();
 sg13g2_decap_8 FILLER_35_1476 ();
 sg13g2_decap_4 FILLER_35_1483 ();
 sg13g2_fill_1 FILLER_35_1487 ();
 sg13g2_decap_4 FILLER_35_1496 ();
 sg13g2_fill_1 FILLER_35_1500 ();
 sg13g2_decap_8 FILLER_35_1506 ();
 sg13g2_decap_4 FILLER_35_1513 ();
 sg13g2_fill_2 FILLER_35_1517 ();
 sg13g2_decap_8 FILLER_35_1548 ();
 sg13g2_decap_8 FILLER_35_1555 ();
 sg13g2_decap_8 FILLER_35_1562 ();
 sg13g2_decap_8 FILLER_35_1572 ();
 sg13g2_fill_2 FILLER_35_1579 ();
 sg13g2_fill_1 FILLER_35_1581 ();
 sg13g2_decap_8 FILLER_35_1600 ();
 sg13g2_decap_8 FILLER_35_1607 ();
 sg13g2_decap_8 FILLER_35_1614 ();
 sg13g2_fill_2 FILLER_35_1647 ();
 sg13g2_decap_8 FILLER_35_1675 ();
 sg13g2_decap_4 FILLER_35_1682 ();
 sg13g2_fill_1 FILLER_35_1686 ();
 sg13g2_fill_2 FILLER_35_1693 ();
 sg13g2_fill_1 FILLER_35_1717 ();
 sg13g2_fill_1 FILLER_35_1724 ();
 sg13g2_decap_8 FILLER_35_1743 ();
 sg13g2_fill_2 FILLER_35_1750 ();
 sg13g2_decap_8 FILLER_35_1756 ();
 sg13g2_decap_8 FILLER_35_1763 ();
 sg13g2_fill_1 FILLER_35_1770 ();
 sg13g2_fill_2 FILLER_35_1860 ();
 sg13g2_decap_8 FILLER_35_1885 ();
 sg13g2_decap_4 FILLER_35_1892 ();
 sg13g2_fill_2 FILLER_35_1896 ();
 sg13g2_decap_4 FILLER_35_1934 ();
 sg13g2_fill_1 FILLER_35_1938 ();
 sg13g2_decap_8 FILLER_35_1949 ();
 sg13g2_decap_4 FILLER_35_1956 ();
 sg13g2_fill_2 FILLER_35_1960 ();
 sg13g2_fill_2 FILLER_35_1999 ();
 sg13g2_fill_1 FILLER_35_2001 ();
 sg13g2_decap_4 FILLER_35_2010 ();
 sg13g2_fill_1 FILLER_35_2014 ();
 sg13g2_decap_8 FILLER_35_2041 ();
 sg13g2_fill_2 FILLER_35_2048 ();
 sg13g2_fill_1 FILLER_35_2055 ();
 sg13g2_fill_2 FILLER_35_2082 ();
 sg13g2_decap_8 FILLER_35_2188 ();
 sg13g2_decap_8 FILLER_35_2195 ();
 sg13g2_decap_8 FILLER_35_2202 ();
 sg13g2_decap_4 FILLER_35_2209 ();
 sg13g2_decap_4 FILLER_35_2217 ();
 sg13g2_fill_1 FILLER_35_2221 ();
 sg13g2_decap_4 FILLER_35_2248 ();
 sg13g2_fill_2 FILLER_35_2252 ();
 sg13g2_fill_2 FILLER_35_2306 ();
 sg13g2_decap_8 FILLER_35_2334 ();
 sg13g2_fill_1 FILLER_35_2400 ();
 sg13g2_fill_2 FILLER_35_2432 ();
 sg13g2_decap_4 FILLER_35_2438 ();
 sg13g2_fill_1 FILLER_35_2442 ();
 sg13g2_fill_1 FILLER_35_2448 ();
 sg13g2_fill_1 FILLER_35_2452 ();
 sg13g2_decap_4 FILLER_35_2458 ();
 sg13g2_fill_2 FILLER_35_2462 ();
 sg13g2_decap_8 FILLER_35_2467 ();
 sg13g2_decap_4 FILLER_35_2474 ();
 sg13g2_decap_8 FILLER_35_2482 ();
 sg13g2_decap_4 FILLER_35_2489 ();
 sg13g2_fill_2 FILLER_35_2506 ();
 sg13g2_fill_1 FILLER_35_2508 ();
 sg13g2_decap_8 FILLER_35_2547 ();
 sg13g2_decap_8 FILLER_35_2554 ();
 sg13g2_decap_8 FILLER_35_2561 ();
 sg13g2_decap_8 FILLER_35_2568 ();
 sg13g2_fill_1 FILLER_35_2575 ();
 sg13g2_decap_4 FILLER_35_2581 ();
 sg13g2_decap_8 FILLER_35_2590 ();
 sg13g2_decap_8 FILLER_35_2597 ();
 sg13g2_decap_8 FILLER_35_2604 ();
 sg13g2_fill_2 FILLER_35_2611 ();
 sg13g2_fill_1 FILLER_35_2613 ();
 sg13g2_decap_8 FILLER_35_2618 ();
 sg13g2_decap_4 FILLER_35_2625 ();
 sg13g2_fill_1 FILLER_35_2629 ();
 sg13g2_decap_4 FILLER_35_2661 ();
 sg13g2_fill_2 FILLER_35_2665 ();
 sg13g2_decap_8 FILLER_35_2675 ();
 sg13g2_fill_2 FILLER_35_2682 ();
 sg13g2_fill_1 FILLER_35_2684 ();
 sg13g2_decap_8 FILLER_35_2752 ();
 sg13g2_decap_4 FILLER_35_2759 ();
 sg13g2_fill_1 FILLER_35_2763 ();
 sg13g2_fill_2 FILLER_35_2798 ();
 sg13g2_fill_1 FILLER_35_2800 ();
 sg13g2_decap_8 FILLER_35_2806 ();
 sg13g2_decap_8 FILLER_35_2813 ();
 sg13g2_decap_4 FILLER_35_2820 ();
 sg13g2_fill_2 FILLER_35_2824 ();
 sg13g2_decap_8 FILLER_35_2852 ();
 sg13g2_decap_8 FILLER_35_2859 ();
 sg13g2_fill_2 FILLER_35_2866 ();
 sg13g2_fill_1 FILLER_35_2868 ();
 sg13g2_decap_8 FILLER_35_3031 ();
 sg13g2_fill_2 FILLER_35_3038 ();
 sg13g2_fill_1 FILLER_35_3040 ();
 sg13g2_decap_4 FILLER_35_3074 ();
 sg13g2_fill_2 FILLER_35_3078 ();
 sg13g2_decap_8 FILLER_35_3113 ();
 sg13g2_decap_8 FILLER_35_3120 ();
 sg13g2_fill_2 FILLER_35_3127 ();
 sg13g2_decap_8 FILLER_35_3141 ();
 sg13g2_decap_8 FILLER_35_3148 ();
 sg13g2_decap_4 FILLER_35_3155 ();
 sg13g2_decap_8 FILLER_35_3185 ();
 sg13g2_decap_4 FILLER_35_3192 ();
 sg13g2_fill_1 FILLER_35_3196 ();
 sg13g2_decap_8 FILLER_35_3275 ();
 sg13g2_decap_8 FILLER_35_3282 ();
 sg13g2_decap_8 FILLER_35_3289 ();
 sg13g2_decap_8 FILLER_35_3296 ();
 sg13g2_decap_8 FILLER_35_3303 ();
 sg13g2_decap_8 FILLER_35_3310 ();
 sg13g2_decap_8 FILLER_35_3317 ();
 sg13g2_decap_8 FILLER_35_3324 ();
 sg13g2_decap_8 FILLER_35_3331 ();
 sg13g2_decap_8 FILLER_35_3338 ();
 sg13g2_decap_8 FILLER_35_3345 ();
 sg13g2_decap_8 FILLER_35_3352 ();
 sg13g2_decap_8 FILLER_35_3359 ();
 sg13g2_decap_8 FILLER_35_3366 ();
 sg13g2_decap_8 FILLER_35_3373 ();
 sg13g2_decap_8 FILLER_35_3380 ();
 sg13g2_decap_8 FILLER_35_3387 ();
 sg13g2_decap_8 FILLER_35_3394 ();
 sg13g2_decap_8 FILLER_35_3401 ();
 sg13g2_decap_8 FILLER_35_3408 ();
 sg13g2_decap_8 FILLER_35_3415 ();
 sg13g2_decap_8 FILLER_35_3422 ();
 sg13g2_decap_8 FILLER_35_3429 ();
 sg13g2_decap_8 FILLER_35_3436 ();
 sg13g2_decap_8 FILLER_35_3443 ();
 sg13g2_decap_8 FILLER_35_3450 ();
 sg13g2_decap_8 FILLER_35_3457 ();
 sg13g2_decap_8 FILLER_35_3464 ();
 sg13g2_decap_8 FILLER_35_3471 ();
 sg13g2_decap_8 FILLER_35_3478 ();
 sg13g2_decap_8 FILLER_35_3485 ();
 sg13g2_decap_8 FILLER_35_3492 ();
 sg13g2_decap_8 FILLER_35_3499 ();
 sg13g2_decap_8 FILLER_35_3506 ();
 sg13g2_decap_8 FILLER_35_3513 ();
 sg13g2_decap_8 FILLER_35_3520 ();
 sg13g2_decap_8 FILLER_35_3527 ();
 sg13g2_decap_8 FILLER_35_3534 ();
 sg13g2_decap_8 FILLER_35_3541 ();
 sg13g2_decap_8 FILLER_35_3548 ();
 sg13g2_decap_8 FILLER_35_3555 ();
 sg13g2_decap_8 FILLER_35_3562 ();
 sg13g2_decap_8 FILLER_35_3569 ();
 sg13g2_decap_4 FILLER_35_3576 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_4 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_39 ();
 sg13g2_fill_1 FILLER_36_101 ();
 sg13g2_decap_8 FILLER_36_128 ();
 sg13g2_decap_8 FILLER_36_135 ();
 sg13g2_decap_4 FILLER_36_142 ();
 sg13g2_decap_4 FILLER_36_154 ();
 sg13g2_decap_4 FILLER_36_179 ();
 sg13g2_fill_2 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_190 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_decap_4 FILLER_36_206 ();
 sg13g2_fill_2 FILLER_36_210 ();
 sg13g2_fill_2 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_decap_4 FILLER_36_331 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_8 FILLER_36_404 ();
 sg13g2_fill_2 FILLER_36_419 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_fill_1 FILLER_36_433 ();
 sg13g2_fill_1 FILLER_36_442 ();
 sg13g2_decap_4 FILLER_36_452 ();
 sg13g2_fill_2 FILLER_36_459 ();
 sg13g2_fill_1 FILLER_36_461 ();
 sg13g2_decap_8 FILLER_36_472 ();
 sg13g2_decap_8 FILLER_36_479 ();
 sg13g2_decap_8 FILLER_36_486 ();
 sg13g2_fill_1 FILLER_36_493 ();
 sg13g2_fill_1 FILLER_36_502 ();
 sg13g2_decap_8 FILLER_36_513 ();
 sg13g2_decap_8 FILLER_36_520 ();
 sg13g2_fill_1 FILLER_36_527 ();
 sg13g2_decap_4 FILLER_36_538 ();
 sg13g2_fill_1 FILLER_36_542 ();
 sg13g2_decap_8 FILLER_36_549 ();
 sg13g2_decap_8 FILLER_36_556 ();
 sg13g2_fill_2 FILLER_36_563 ();
 sg13g2_fill_1 FILLER_36_565 ();
 sg13g2_decap_8 FILLER_36_576 ();
 sg13g2_decap_4 FILLER_36_583 ();
 sg13g2_fill_2 FILLER_36_587 ();
 sg13g2_fill_1 FILLER_36_623 ();
 sg13g2_decap_8 FILLER_36_653 ();
 sg13g2_decap_4 FILLER_36_660 ();
 sg13g2_fill_1 FILLER_36_664 ();
 sg13g2_fill_2 FILLER_36_697 ();
 sg13g2_fill_2 FILLER_36_709 ();
 sg13g2_decap_8 FILLER_36_723 ();
 sg13g2_decap_8 FILLER_36_730 ();
 sg13g2_fill_2 FILLER_36_737 ();
 sg13g2_fill_1 FILLER_36_739 ();
 sg13g2_decap_8 FILLER_36_745 ();
 sg13g2_decap_4 FILLER_36_752 ();
 sg13g2_fill_2 FILLER_36_756 ();
 sg13g2_decap_8 FILLER_36_763 ();
 sg13g2_fill_1 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_784 ();
 sg13g2_fill_2 FILLER_36_791 ();
 sg13g2_decap_8 FILLER_36_832 ();
 sg13g2_decap_8 FILLER_36_839 ();
 sg13g2_decap_8 FILLER_36_846 ();
 sg13g2_decap_4 FILLER_36_853 ();
 sg13g2_fill_1 FILLER_36_857 ();
 sg13g2_decap_8 FILLER_36_889 ();
 sg13g2_fill_2 FILLER_36_896 ();
 sg13g2_fill_1 FILLER_36_898 ();
 sg13g2_fill_2 FILLER_36_902 ();
 sg13g2_fill_2 FILLER_36_971 ();
 sg13g2_fill_1 FILLER_36_973 ();
 sg13g2_fill_2 FILLER_36_989 ();
 sg13g2_fill_2 FILLER_36_996 ();
 sg13g2_fill_1 FILLER_36_998 ();
 sg13g2_fill_2 FILLER_36_1023 ();
 sg13g2_decap_8 FILLER_36_1038 ();
 sg13g2_decap_4 FILLER_36_1045 ();
 sg13g2_decap_8 FILLER_36_1059 ();
 sg13g2_decap_8 FILLER_36_1066 ();
 sg13g2_decap_8 FILLER_36_1073 ();
 sg13g2_decap_8 FILLER_36_1080 ();
 sg13g2_decap_4 FILLER_36_1087 ();
 sg13g2_fill_2 FILLER_36_1091 ();
 sg13g2_decap_8 FILLER_36_1103 ();
 sg13g2_decap_8 FILLER_36_1110 ();
 sg13g2_decap_8 FILLER_36_1117 ();
 sg13g2_fill_2 FILLER_36_1124 ();
 sg13g2_fill_1 FILLER_36_1126 ();
 sg13g2_decap_4 FILLER_36_1135 ();
 sg13g2_fill_2 FILLER_36_1139 ();
 sg13g2_fill_1 FILLER_36_1151 ();
 sg13g2_fill_1 FILLER_36_1168 ();
 sg13g2_fill_1 FILLER_36_1206 ();
 sg13g2_fill_1 FILLER_36_1211 ();
 sg13g2_decap_8 FILLER_36_1220 ();
 sg13g2_decap_4 FILLER_36_1235 ();
 sg13g2_fill_2 FILLER_36_1239 ();
 sg13g2_fill_2 FILLER_36_1254 ();
 sg13g2_fill_1 FILLER_36_1256 ();
 sg13g2_decap_4 FILLER_36_1280 ();
 sg13g2_fill_1 FILLER_36_1284 ();
 sg13g2_fill_2 FILLER_36_1290 ();
 sg13g2_fill_1 FILLER_36_1318 ();
 sg13g2_decap_8 FILLER_36_1349 ();
 sg13g2_decap_8 FILLER_36_1395 ();
 sg13g2_decap_8 FILLER_36_1402 ();
 sg13g2_fill_1 FILLER_36_1409 ();
 sg13g2_fill_1 FILLER_36_1490 ();
 sg13g2_decap_8 FILLER_36_1495 ();
 sg13g2_decap_8 FILLER_36_1502 ();
 sg13g2_decap_8 FILLER_36_1509 ();
 sg13g2_decap_4 FILLER_36_1516 ();
 sg13g2_fill_1 FILLER_36_1520 ();
 sg13g2_fill_2 FILLER_36_1554 ();
 sg13g2_fill_1 FILLER_36_1556 ();
 sg13g2_decap_8 FILLER_36_1612 ();
 sg13g2_fill_1 FILLER_36_1619 ();
 sg13g2_fill_1 FILLER_36_1654 ();
 sg13g2_fill_2 FILLER_36_1681 ();
 sg13g2_fill_2 FILLER_36_1693 ();
 sg13g2_fill_1 FILLER_36_1708 ();
 sg13g2_decap_8 FILLER_36_1750 ();
 sg13g2_decap_8 FILLER_36_1757 ();
 sg13g2_decap_8 FILLER_36_1764 ();
 sg13g2_decap_4 FILLER_36_1771 ();
 sg13g2_fill_2 FILLER_36_1775 ();
 sg13g2_fill_2 FILLER_36_1782 ();
 sg13g2_decap_8 FILLER_36_1790 ();
 sg13g2_fill_2 FILLER_36_1797 ();
 sg13g2_decap_8 FILLER_36_1804 ();
 sg13g2_decap_8 FILLER_36_1811 ();
 sg13g2_decap_8 FILLER_36_1818 ();
 sg13g2_decap_4 FILLER_36_1825 ();
 sg13g2_fill_1 FILLER_36_1829 ();
 sg13g2_decap_8 FILLER_36_1864 ();
 sg13g2_decap_8 FILLER_36_1949 ();
 sg13g2_fill_1 FILLER_36_1956 ();
 sg13g2_fill_2 FILLER_36_1993 ();
 sg13g2_fill_1 FILLER_36_2029 ();
 sg13g2_decap_4 FILLER_36_2087 ();
 sg13g2_decap_4 FILLER_36_2153 ();
 sg13g2_decap_8 FILLER_36_2214 ();
 sg13g2_fill_2 FILLER_36_2221 ();
 sg13g2_decap_8 FILLER_36_2249 ();
 sg13g2_decap_4 FILLER_36_2256 ();
 sg13g2_decap_4 FILLER_36_2338 ();
 sg13g2_fill_2 FILLER_36_2382 ();
 sg13g2_decap_8 FILLER_36_2392 ();
 sg13g2_decap_4 FILLER_36_2399 ();
 sg13g2_fill_2 FILLER_36_2403 ();
 sg13g2_decap_8 FILLER_36_2488 ();
 sg13g2_decap_8 FILLER_36_2495 ();
 sg13g2_fill_1 FILLER_36_2502 ();
 sg13g2_decap_4 FILLER_36_2540 ();
 sg13g2_fill_2 FILLER_36_2544 ();
 sg13g2_decap_8 FILLER_36_2551 ();
 sg13g2_fill_2 FILLER_36_2558 ();
 sg13g2_fill_1 FILLER_36_2560 ();
 sg13g2_fill_1 FILLER_36_2566 ();
 sg13g2_decap_8 FILLER_36_2596 ();
 sg13g2_fill_1 FILLER_36_2629 ();
 sg13g2_fill_1 FILLER_36_2659 ();
 sg13g2_decap_8 FILLER_36_2664 ();
 sg13g2_fill_2 FILLER_36_2671 ();
 sg13g2_decap_4 FILLER_36_2725 ();
 sg13g2_decap_4 FILLER_36_2763 ();
 sg13g2_fill_2 FILLER_36_2767 ();
 sg13g2_fill_2 FILLER_36_2778 ();
 sg13g2_decap_4 FILLER_36_2800 ();
 sg13g2_fill_2 FILLER_36_2804 ();
 sg13g2_fill_2 FILLER_36_2814 ();
 sg13g2_fill_1 FILLER_36_2816 ();
 sg13g2_decap_8 FILLER_36_2857 ();
 sg13g2_fill_1 FILLER_36_2864 ();
 sg13g2_decap_8 FILLER_36_2907 ();
 sg13g2_decap_8 FILLER_36_2914 ();
 sg13g2_fill_2 FILLER_36_2921 ();
 sg13g2_fill_1 FILLER_36_2923 ();
 sg13g2_decap_8 FILLER_36_2963 ();
 sg13g2_fill_2 FILLER_36_2970 ();
 sg13g2_decap_8 FILLER_36_2980 ();
 sg13g2_decap_8 FILLER_36_3013 ();
 sg13g2_decap_4 FILLER_36_3020 ();
 sg13g2_fill_2 FILLER_36_3024 ();
 sg13g2_decap_8 FILLER_36_3033 ();
 sg13g2_fill_2 FILLER_36_3048 ();
 sg13g2_fill_1 FILLER_36_3055 ();
 sg13g2_decap_8 FILLER_36_3064 ();
 sg13g2_decap_8 FILLER_36_3071 ();
 sg13g2_decap_8 FILLER_36_3078 ();
 sg13g2_decap_8 FILLER_36_3085 ();
 sg13g2_decap_8 FILLER_36_3092 ();
 sg13g2_fill_1 FILLER_36_3099 ();
 sg13g2_decap_8 FILLER_36_3126 ();
 sg13g2_decap_8 FILLER_36_3133 ();
 sg13g2_decap_8 FILLER_36_3140 ();
 sg13g2_decap_8 FILLER_36_3147 ();
 sg13g2_decap_4 FILLER_36_3154 ();
 sg13g2_decap_8 FILLER_36_3269 ();
 sg13g2_decap_8 FILLER_36_3276 ();
 sg13g2_decap_8 FILLER_36_3283 ();
 sg13g2_decap_8 FILLER_36_3290 ();
 sg13g2_decap_8 FILLER_36_3297 ();
 sg13g2_decap_8 FILLER_36_3304 ();
 sg13g2_decap_8 FILLER_36_3311 ();
 sg13g2_decap_8 FILLER_36_3318 ();
 sg13g2_decap_8 FILLER_36_3325 ();
 sg13g2_decap_8 FILLER_36_3332 ();
 sg13g2_decap_8 FILLER_36_3339 ();
 sg13g2_decap_8 FILLER_36_3346 ();
 sg13g2_decap_8 FILLER_36_3353 ();
 sg13g2_decap_8 FILLER_36_3360 ();
 sg13g2_decap_8 FILLER_36_3367 ();
 sg13g2_decap_8 FILLER_36_3374 ();
 sg13g2_decap_8 FILLER_36_3381 ();
 sg13g2_decap_8 FILLER_36_3388 ();
 sg13g2_decap_8 FILLER_36_3395 ();
 sg13g2_decap_8 FILLER_36_3402 ();
 sg13g2_decap_8 FILLER_36_3409 ();
 sg13g2_decap_8 FILLER_36_3416 ();
 sg13g2_decap_8 FILLER_36_3423 ();
 sg13g2_decap_8 FILLER_36_3430 ();
 sg13g2_decap_8 FILLER_36_3437 ();
 sg13g2_decap_8 FILLER_36_3444 ();
 sg13g2_decap_8 FILLER_36_3451 ();
 sg13g2_decap_8 FILLER_36_3458 ();
 sg13g2_decap_8 FILLER_36_3465 ();
 sg13g2_decap_8 FILLER_36_3472 ();
 sg13g2_decap_8 FILLER_36_3479 ();
 sg13g2_decap_8 FILLER_36_3486 ();
 sg13g2_decap_8 FILLER_36_3493 ();
 sg13g2_decap_8 FILLER_36_3500 ();
 sg13g2_decap_8 FILLER_36_3507 ();
 sg13g2_decap_8 FILLER_36_3514 ();
 sg13g2_decap_8 FILLER_36_3521 ();
 sg13g2_decap_8 FILLER_36_3528 ();
 sg13g2_decap_8 FILLER_36_3535 ();
 sg13g2_decap_8 FILLER_36_3542 ();
 sg13g2_decap_8 FILLER_36_3549 ();
 sg13g2_decap_8 FILLER_36_3556 ();
 sg13g2_decap_8 FILLER_36_3563 ();
 sg13g2_decap_8 FILLER_36_3570 ();
 sg13g2_fill_2 FILLER_36_3577 ();
 sg13g2_fill_1 FILLER_36_3579 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_63 ();
 sg13g2_decap_4 FILLER_37_69 ();
 sg13g2_fill_1 FILLER_37_73 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_200 ();
 sg13g2_fill_2 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_decap_4 FILLER_37_252 ();
 sg13g2_fill_1 FILLER_37_256 ();
 sg13g2_decap_8 FILLER_37_313 ();
 sg13g2_decap_8 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_4 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_4 FILLER_37_469 ();
 sg13g2_fill_1 FILLER_37_473 ();
 sg13g2_decap_8 FILLER_37_500 ();
 sg13g2_decap_8 FILLER_37_507 ();
 sg13g2_decap_8 FILLER_37_540 ();
 sg13g2_decap_4 FILLER_37_547 ();
 sg13g2_decap_8 FILLER_37_554 ();
 sg13g2_decap_4 FILLER_37_561 ();
 sg13g2_fill_1 FILLER_37_565 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_fill_2 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_596 ();
 sg13g2_decap_8 FILLER_37_603 ();
 sg13g2_decap_8 FILLER_37_610 ();
 sg13g2_decap_8 FILLER_37_617 ();
 sg13g2_decap_4 FILLER_37_624 ();
 sg13g2_fill_1 FILLER_37_628 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_4 FILLER_37_644 ();
 sg13g2_fill_2 FILLER_37_648 ();
 sg13g2_decap_4 FILLER_37_733 ();
 sg13g2_fill_2 FILLER_37_769 ();
 sg13g2_fill_1 FILLER_37_784 ();
 sg13g2_decap_4 FILLER_37_810 ();
 sg13g2_decap_8 FILLER_37_892 ();
 sg13g2_decap_4 FILLER_37_899 ();
 sg13g2_fill_1 FILLER_37_903 ();
 sg13g2_decap_8 FILLER_37_940 ();
 sg13g2_decap_8 FILLER_37_947 ();
 sg13g2_decap_8 FILLER_37_954 ();
 sg13g2_fill_2 FILLER_37_961 ();
 sg13g2_fill_1 FILLER_37_977 ();
 sg13g2_fill_1 FILLER_37_1002 ();
 sg13g2_decap_8 FILLER_37_1025 ();
 sg13g2_fill_2 FILLER_37_1032 ();
 sg13g2_fill_1 FILLER_37_1034 ();
 sg13g2_decap_8 FILLER_37_1116 ();
 sg13g2_fill_2 FILLER_37_1123 ();
 sg13g2_fill_1 FILLER_37_1125 ();
 sg13g2_fill_1 FILLER_37_1152 ();
 sg13g2_fill_1 FILLER_37_1158 ();
 sg13g2_fill_1 FILLER_37_1167 ();
 sg13g2_fill_2 FILLER_37_1186 ();
 sg13g2_fill_1 FILLER_37_1193 ();
 sg13g2_fill_1 FILLER_37_1199 ();
 sg13g2_fill_2 FILLER_37_1208 ();
 sg13g2_fill_1 FILLER_37_1210 ();
 sg13g2_fill_1 FILLER_37_1219 ();
 sg13g2_fill_2 FILLER_37_1241 ();
 sg13g2_fill_2 FILLER_37_1277 ();
 sg13g2_decap_4 FILLER_37_1287 ();
 sg13g2_fill_2 FILLER_37_1299 ();
 sg13g2_fill_1 FILLER_37_1319 ();
 sg13g2_decap_8 FILLER_37_1334 ();
 sg13g2_fill_1 FILLER_37_1341 ();
 sg13g2_decap_4 FILLER_37_1397 ();
 sg13g2_fill_2 FILLER_37_1401 ();
 sg13g2_fill_2 FILLER_37_1411 ();
 sg13g2_fill_1 FILLER_37_1413 ();
 sg13g2_fill_2 FILLER_37_1474 ();
 sg13g2_decap_8 FILLER_37_1502 ();
 sg13g2_decap_4 FILLER_37_1509 ();
 sg13g2_decap_8 FILLER_37_1551 ();
 sg13g2_decap_8 FILLER_37_1558 ();
 sg13g2_fill_1 FILLER_37_1565 ();
 sg13g2_decap_4 FILLER_37_1628 ();
 sg13g2_fill_2 FILLER_37_1632 ();
 sg13g2_decap_4 FILLER_37_1647 ();
 sg13g2_fill_2 FILLER_37_1651 ();
 sg13g2_decap_8 FILLER_37_1684 ();
 sg13g2_decap_8 FILLER_37_1696 ();
 sg13g2_decap_4 FILLER_37_1703 ();
 sg13g2_fill_2 FILLER_37_1736 ();
 sg13g2_decap_8 FILLER_37_1756 ();
 sg13g2_decap_8 FILLER_37_1763 ();
 sg13g2_decap_4 FILLER_37_1770 ();
 sg13g2_fill_1 FILLER_37_1774 ();
 sg13g2_decap_8 FILLER_37_1801 ();
 sg13g2_decap_8 FILLER_37_1808 ();
 sg13g2_decap_8 FILLER_37_1815 ();
 sg13g2_decap_8 FILLER_37_1859 ();
 sg13g2_decap_8 FILLER_37_1866 ();
 sg13g2_decap_8 FILLER_37_1873 ();
 sg13g2_decap_4 FILLER_37_1880 ();
 sg13g2_fill_2 FILLER_37_1903 ();
 sg13g2_fill_1 FILLER_37_1920 ();
 sg13g2_decap_4 FILLER_37_1937 ();
 sg13g2_decap_8 FILLER_37_1948 ();
 sg13g2_decap_4 FILLER_37_1955 ();
 sg13g2_fill_1 FILLER_37_1959 ();
 sg13g2_decap_8 FILLER_37_2045 ();
 sg13g2_decap_8 FILLER_37_2078 ();
 sg13g2_fill_1 FILLER_37_2085 ();
 sg13g2_decap_8 FILLER_37_2090 ();
 sg13g2_decap_8 FILLER_37_2097 ();
 sg13g2_decap_8 FILLER_37_2104 ();
 sg13g2_decap_4 FILLER_37_2111 ();
 sg13g2_decap_4 FILLER_37_2119 ();
 sg13g2_decap_8 FILLER_37_2131 ();
 sg13g2_decap_8 FILLER_37_2138 ();
 sg13g2_decap_8 FILLER_37_2145 ();
 sg13g2_decap_8 FILLER_37_2152 ();
 sg13g2_fill_2 FILLER_37_2159 ();
 sg13g2_fill_1 FILLER_37_2161 ();
 sg13g2_decap_8 FILLER_37_2214 ();
 sg13g2_decap_4 FILLER_37_2221 ();
 sg13g2_decap_8 FILLER_37_2251 ();
 sg13g2_decap_4 FILLER_37_2258 ();
 sg13g2_fill_2 FILLER_37_2262 ();
 sg13g2_decap_8 FILLER_37_2316 ();
 sg13g2_decap_8 FILLER_37_2323 ();
 sg13g2_decap_8 FILLER_37_2330 ();
 sg13g2_fill_1 FILLER_37_2337 ();
 sg13g2_decap_8 FILLER_37_2370 ();
 sg13g2_decap_8 FILLER_37_2377 ();
 sg13g2_decap_8 FILLER_37_2384 ();
 sg13g2_fill_1 FILLER_37_2391 ();
 sg13g2_fill_1 FILLER_37_2397 ();
 sg13g2_fill_2 FILLER_37_2450 ();
 sg13g2_fill_1 FILLER_37_2460 ();
 sg13g2_decap_8 FILLER_37_2487 ();
 sg13g2_decap_8 FILLER_37_2494 ();
 sg13g2_decap_8 FILLER_37_2501 ();
 sg13g2_decap_4 FILLER_37_2508 ();
 sg13g2_fill_1 FILLER_37_2538 ();
 sg13g2_decap_4 FILLER_37_2551 ();
 sg13g2_fill_2 FILLER_37_2555 ();
 sg13g2_fill_2 FILLER_37_2588 ();
 sg13g2_fill_2 FILLER_37_2646 ();
 sg13g2_fill_1 FILLER_37_2648 ();
 sg13g2_decap_8 FILLER_37_2675 ();
 sg13g2_fill_2 FILLER_37_2682 ();
 sg13g2_decap_8 FILLER_37_2688 ();
 sg13g2_decap_4 FILLER_37_2695 ();
 sg13g2_decap_8 FILLER_37_2708 ();
 sg13g2_decap_4 FILLER_37_2715 ();
 sg13g2_fill_2 FILLER_37_2719 ();
 sg13g2_decap_8 FILLER_37_2759 ();
 sg13g2_decap_8 FILLER_37_2766 ();
 sg13g2_fill_1 FILLER_37_2773 ();
 sg13g2_decap_8 FILLER_37_2799 ();
 sg13g2_decap_8 FILLER_37_2806 ();
 sg13g2_fill_2 FILLER_37_2813 ();
 sg13g2_fill_2 FILLER_37_2833 ();
 sg13g2_fill_1 FILLER_37_2835 ();
 sg13g2_decap_8 FILLER_37_2843 ();
 sg13g2_fill_1 FILLER_37_2850 ();
 sg13g2_fill_2 FILLER_37_2880 ();
 sg13g2_fill_1 FILLER_37_2882 ();
 sg13g2_decap_8 FILLER_37_2896 ();
 sg13g2_fill_2 FILLER_37_2903 ();
 sg13g2_decap_8 FILLER_37_2913 ();
 sg13g2_decap_4 FILLER_37_2920 ();
 sg13g2_fill_2 FILLER_37_2924 ();
 sg13g2_decap_8 FILLER_37_2931 ();
 sg13g2_decap_8 FILLER_37_2964 ();
 sg13g2_decap_8 FILLER_37_2971 ();
 sg13g2_decap_8 FILLER_37_2978 ();
 sg13g2_decap_8 FILLER_37_2985 ();
 sg13g2_fill_2 FILLER_37_2992 ();
 sg13g2_fill_1 FILLER_37_2994 ();
 sg13g2_decap_8 FILLER_37_3000 ();
 sg13g2_decap_8 FILLER_37_3007 ();
 sg13g2_decap_8 FILLER_37_3014 ();
 sg13g2_decap_8 FILLER_37_3021 ();
 sg13g2_decap_8 FILLER_37_3028 ();
 sg13g2_decap_8 FILLER_37_3035 ();
 sg13g2_decap_8 FILLER_37_3042 ();
 sg13g2_decap_4 FILLER_37_3049 ();
 sg13g2_decap_8 FILLER_37_3079 ();
 sg13g2_decap_4 FILLER_37_3086 ();
 sg13g2_decap_8 FILLER_37_3122 ();
 sg13g2_fill_2 FILLER_37_3195 ();
 sg13g2_fill_1 FILLER_37_3197 ();
 sg13g2_fill_2 FILLER_37_3211 ();
 sg13g2_fill_2 FILLER_37_3238 ();
 sg13g2_decap_8 FILLER_37_3243 ();
 sg13g2_decap_4 FILLER_37_3250 ();
 sg13g2_decap_8 FILLER_37_3262 ();
 sg13g2_decap_8 FILLER_37_3269 ();
 sg13g2_decap_8 FILLER_37_3276 ();
 sg13g2_decap_8 FILLER_37_3283 ();
 sg13g2_decap_8 FILLER_37_3290 ();
 sg13g2_decap_8 FILLER_37_3297 ();
 sg13g2_decap_8 FILLER_37_3304 ();
 sg13g2_decap_8 FILLER_37_3311 ();
 sg13g2_decap_8 FILLER_37_3318 ();
 sg13g2_decap_8 FILLER_37_3325 ();
 sg13g2_decap_8 FILLER_37_3332 ();
 sg13g2_decap_8 FILLER_37_3339 ();
 sg13g2_decap_8 FILLER_37_3346 ();
 sg13g2_decap_8 FILLER_37_3353 ();
 sg13g2_decap_8 FILLER_37_3360 ();
 sg13g2_decap_8 FILLER_37_3367 ();
 sg13g2_decap_8 FILLER_37_3374 ();
 sg13g2_decap_8 FILLER_37_3381 ();
 sg13g2_decap_8 FILLER_37_3388 ();
 sg13g2_decap_8 FILLER_37_3395 ();
 sg13g2_decap_8 FILLER_37_3402 ();
 sg13g2_decap_8 FILLER_37_3409 ();
 sg13g2_decap_8 FILLER_37_3416 ();
 sg13g2_decap_8 FILLER_37_3423 ();
 sg13g2_decap_8 FILLER_37_3430 ();
 sg13g2_decap_8 FILLER_37_3437 ();
 sg13g2_decap_8 FILLER_37_3444 ();
 sg13g2_decap_8 FILLER_37_3451 ();
 sg13g2_decap_8 FILLER_37_3458 ();
 sg13g2_decap_8 FILLER_37_3465 ();
 sg13g2_decap_8 FILLER_37_3472 ();
 sg13g2_decap_8 FILLER_37_3479 ();
 sg13g2_decap_8 FILLER_37_3486 ();
 sg13g2_decap_8 FILLER_37_3493 ();
 sg13g2_decap_8 FILLER_37_3500 ();
 sg13g2_decap_8 FILLER_37_3507 ();
 sg13g2_decap_8 FILLER_37_3514 ();
 sg13g2_decap_8 FILLER_37_3521 ();
 sg13g2_decap_8 FILLER_37_3528 ();
 sg13g2_decap_8 FILLER_37_3535 ();
 sg13g2_decap_8 FILLER_37_3542 ();
 sg13g2_decap_8 FILLER_37_3549 ();
 sg13g2_decap_8 FILLER_37_3556 ();
 sg13g2_decap_8 FILLER_37_3563 ();
 sg13g2_decap_8 FILLER_37_3570 ();
 sg13g2_fill_2 FILLER_37_3577 ();
 sg13g2_fill_1 FILLER_37_3579 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_fill_2 FILLER_38_137 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_decap_8 FILLER_38_239 ();
 sg13g2_decap_8 FILLER_38_246 ();
 sg13g2_decap_8 FILLER_38_253 ();
 sg13g2_decap_8 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_4 FILLER_38_345 ();
 sg13g2_fill_2 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_388 ();
 sg13g2_fill_1 FILLER_38_441 ();
 sg13g2_fill_1 FILLER_38_450 ();
 sg13g2_decap_8 FILLER_38_495 ();
 sg13g2_decap_8 FILLER_38_502 ();
 sg13g2_decap_8 FILLER_38_509 ();
 sg13g2_fill_2 FILLER_38_516 ();
 sg13g2_decap_8 FILLER_38_596 ();
 sg13g2_fill_2 FILLER_38_603 ();
 sg13g2_fill_2 FILLER_38_683 ();
 sg13g2_fill_1 FILLER_38_699 ();
 sg13g2_fill_1 FILLER_38_712 ();
 sg13g2_fill_2 FILLER_38_755 ();
 sg13g2_fill_1 FILLER_38_757 ();
 sg13g2_fill_1 FILLER_38_810 ();
 sg13g2_fill_1 FILLER_38_842 ();
 sg13g2_decap_8 FILLER_38_891 ();
 sg13g2_decap_8 FILLER_38_898 ();
 sg13g2_decap_8 FILLER_38_905 ();
 sg13g2_decap_4 FILLER_38_912 ();
 sg13g2_fill_2 FILLER_38_916 ();
 sg13g2_decap_8 FILLER_38_949 ();
 sg13g2_decap_8 FILLER_38_956 ();
 sg13g2_decap_4 FILLER_38_963 ();
 sg13g2_fill_2 FILLER_38_967 ();
 sg13g2_decap_8 FILLER_38_1025 ();
 sg13g2_decap_4 FILLER_38_1032 ();
 sg13g2_fill_2 FILLER_38_1036 ();
 sg13g2_fill_2 FILLER_38_1067 ();
 sg13g2_decap_8 FILLER_38_1074 ();
 sg13g2_decap_8 FILLER_38_1081 ();
 sg13g2_decap_8 FILLER_38_1088 ();
 sg13g2_decap_8 FILLER_38_1095 ();
 sg13g2_fill_2 FILLER_38_1102 ();
 sg13g2_fill_1 FILLER_38_1104 ();
 sg13g2_decap_8 FILLER_38_1131 ();
 sg13g2_decap_8 FILLER_38_1138 ();
 sg13g2_decap_8 FILLER_38_1145 ();
 sg13g2_fill_2 FILLER_38_1152 ();
 sg13g2_decap_4 FILLER_38_1159 ();
 sg13g2_decap_8 FILLER_38_1173 ();
 sg13g2_fill_1 FILLER_38_1180 ();
 sg13g2_fill_2 FILLER_38_1186 ();
 sg13g2_fill_1 FILLER_38_1188 ();
 sg13g2_fill_2 FILLER_38_1201 ();
 sg13g2_fill_1 FILLER_38_1216 ();
 sg13g2_fill_1 FILLER_38_1256 ();
 sg13g2_fill_2 FILLER_38_1274 ();
 sg13g2_fill_1 FILLER_38_1276 ();
 sg13g2_fill_1 FILLER_38_1289 ();
 sg13g2_decap_4 FILLER_38_1298 ();
 sg13g2_decap_4 FILLER_38_1307 ();
 sg13g2_fill_1 FILLER_38_1311 ();
 sg13g2_decap_4 FILLER_38_1320 ();
 sg13g2_fill_1 FILLER_38_1324 ();
 sg13g2_fill_2 FILLER_38_1328 ();
 sg13g2_fill_1 FILLER_38_1330 ();
 sg13g2_decap_8 FILLER_38_1336 ();
 sg13g2_decap_4 FILLER_38_1343 ();
 sg13g2_fill_1 FILLER_38_1347 ();
 sg13g2_decap_4 FILLER_38_1356 ();
 sg13g2_fill_2 FILLER_38_1376 ();
 sg13g2_fill_2 FILLER_38_1394 ();
 sg13g2_decap_8 FILLER_38_1404 ();
 sg13g2_decap_4 FILLER_38_1411 ();
 sg13g2_fill_2 FILLER_38_1415 ();
 sg13g2_fill_1 FILLER_38_1430 ();
 sg13g2_fill_2 FILLER_38_1468 ();
 sg13g2_fill_1 FILLER_38_1470 ();
 sg13g2_fill_1 FILLER_38_1509 ();
 sg13g2_fill_2 FILLER_38_1554 ();
 sg13g2_fill_2 FILLER_38_1581 ();
 sg13g2_decap_4 FILLER_38_1609 ();
 sg13g2_fill_1 FILLER_38_1613 ();
 sg13g2_decap_8 FILLER_38_1627 ();
 sg13g2_decap_8 FILLER_38_1642 ();
 sg13g2_decap_8 FILLER_38_1649 ();
 sg13g2_decap_8 FILLER_38_1656 ();
 sg13g2_decap_4 FILLER_38_1663 ();
 sg13g2_decap_4 FILLER_38_1706 ();
 sg13g2_fill_1 FILLER_38_1726 ();
 sg13g2_decap_8 FILLER_38_1761 ();
 sg13g2_fill_2 FILLER_38_1768 ();
 sg13g2_fill_1 FILLER_38_1770 ();
 sg13g2_decap_8 FILLER_38_1803 ();
 sg13g2_decap_8 FILLER_38_1810 ();
 sg13g2_decap_8 FILLER_38_1817 ();
 sg13g2_fill_1 FILLER_38_1824 ();
 sg13g2_fill_2 FILLER_38_1833 ();
 sg13g2_fill_1 FILLER_38_1835 ();
 sg13g2_decap_8 FILLER_38_1865 ();
 sg13g2_fill_2 FILLER_38_1872 ();
 sg13g2_fill_1 FILLER_38_1874 ();
 sg13g2_decap_8 FILLER_38_1878 ();
 sg13g2_decap_4 FILLER_38_1885 ();
 sg13g2_fill_1 FILLER_38_1889 ();
 sg13g2_decap_4 FILLER_38_1911 ();
 sg13g2_fill_2 FILLER_38_1915 ();
 sg13g2_fill_2 FILLER_38_1920 ();
 sg13g2_decap_4 FILLER_38_1931 ();
 sg13g2_fill_1 FILLER_38_1935 ();
 sg13g2_fill_2 FILLER_38_1949 ();
 sg13g2_decap_8 FILLER_38_1959 ();
 sg13g2_fill_1 FILLER_38_1966 ();
 sg13g2_fill_2 FILLER_38_1972 ();
 sg13g2_fill_1 FILLER_38_1974 ();
 sg13g2_fill_1 FILLER_38_1988 ();
 sg13g2_fill_1 FILLER_38_2002 ();
 sg13g2_decap_8 FILLER_38_2029 ();
 sg13g2_decap_8 FILLER_38_2036 ();
 sg13g2_decap_8 FILLER_38_2043 ();
 sg13g2_decap_8 FILLER_38_2050 ();
 sg13g2_fill_2 FILLER_38_2057 ();
 sg13g2_fill_1 FILLER_38_2059 ();
 sg13g2_decap_8 FILLER_38_2065 ();
 sg13g2_decap_8 FILLER_38_2072 ();
 sg13g2_decap_4 FILLER_38_2079 ();
 sg13g2_fill_2 FILLER_38_2083 ();
 sg13g2_fill_1 FILLER_38_2089 ();
 sg13g2_fill_1 FILLER_38_2098 ();
 sg13g2_fill_2 FILLER_38_2109 ();
 sg13g2_decap_8 FILLER_38_2154 ();
 sg13g2_decap_8 FILLER_38_2161 ();
 sg13g2_decap_8 FILLER_38_2168 ();
 sg13g2_decap_8 FILLER_38_2201 ();
 sg13g2_decap_8 FILLER_38_2208 ();
 sg13g2_decap_8 FILLER_38_2215 ();
 sg13g2_fill_2 FILLER_38_2222 ();
 sg13g2_fill_2 FILLER_38_2239 ();
 sg13g2_decap_8 FILLER_38_2251 ();
 sg13g2_decap_8 FILLER_38_2258 ();
 sg13g2_decap_8 FILLER_38_2265 ();
 sg13g2_decap_8 FILLER_38_2272 ();
 sg13g2_fill_2 FILLER_38_2279 ();
 sg13g2_fill_1 FILLER_38_2300 ();
 sg13g2_decap_4 FILLER_38_2318 ();
 sg13g2_fill_2 FILLER_38_2348 ();
 sg13g2_fill_1 FILLER_38_2350 ();
 sg13g2_decap_8 FILLER_38_2377 ();
 sg13g2_decap_8 FILLER_38_2384 ();
 sg13g2_decap_8 FILLER_38_2391 ();
 sg13g2_decap_8 FILLER_38_2398 ();
 sg13g2_decap_4 FILLER_38_2405 ();
 sg13g2_fill_2 FILLER_38_2412 ();
 sg13g2_fill_1 FILLER_38_2466 ();
 sg13g2_decap_8 FILLER_38_2493 ();
 sg13g2_fill_2 FILLER_38_2500 ();
 sg13g2_fill_1 FILLER_38_2502 ();
 sg13g2_fill_2 FILLER_38_2534 ();
 sg13g2_fill_1 FILLER_38_2607 ();
 sg13g2_fill_1 FILLER_38_2634 ();
 sg13g2_decap_8 FILLER_38_2643 ();
 sg13g2_decap_4 FILLER_38_2650 ();
 sg13g2_fill_2 FILLER_38_2654 ();
 sg13g2_decap_8 FILLER_38_2664 ();
 sg13g2_decap_4 FILLER_38_2694 ();
 sg13g2_decap_8 FILLER_38_2701 ();
 sg13g2_fill_2 FILLER_38_2713 ();
 sg13g2_decap_4 FILLER_38_2723 ();
 sg13g2_fill_1 FILLER_38_2727 ();
 sg13g2_fill_2 FILLER_38_2741 ();
 sg13g2_decap_8 FILLER_38_2748 ();
 sg13g2_decap_8 FILLER_38_2755 ();
 sg13g2_decap_8 FILLER_38_2762 ();
 sg13g2_decap_8 FILLER_38_2769 ();
 sg13g2_fill_2 FILLER_38_2776 ();
 sg13g2_fill_1 FILLER_38_2778 ();
 sg13g2_decap_8 FILLER_38_2805 ();
 sg13g2_fill_1 FILLER_38_2812 ();
 sg13g2_fill_1 FILLER_38_2839 ();
 sg13g2_decap_8 FILLER_38_2869 ();
 sg13g2_decap_4 FILLER_38_2876 ();
 sg13g2_decap_4 FILLER_38_2891 ();
 sg13g2_fill_1 FILLER_38_2895 ();
 sg13g2_fill_1 FILLER_38_2922 ();
 sg13g2_fill_2 FILLER_38_2957 ();
 sg13g2_decap_8 FILLER_38_2985 ();
 sg13g2_decap_8 FILLER_38_2992 ();
 sg13g2_fill_1 FILLER_38_3030 ();
 sg13g2_decap_4 FILLER_38_3039 ();
 sg13g2_decap_8 FILLER_38_3076 ();
 sg13g2_decap_4 FILLER_38_3083 ();
 sg13g2_fill_2 FILLER_38_3099 ();
 sg13g2_decap_8 FILLER_38_3126 ();
 sg13g2_decap_8 FILLER_38_3133 ();
 sg13g2_fill_2 FILLER_38_3144 ();
 sg13g2_fill_2 FILLER_38_3200 ();
 sg13g2_decap_8 FILLER_38_3226 ();
 sg13g2_decap_8 FILLER_38_3233 ();
 sg13g2_decap_8 FILLER_38_3240 ();
 sg13g2_decap_8 FILLER_38_3247 ();
 sg13g2_decap_8 FILLER_38_3254 ();
 sg13g2_decap_8 FILLER_38_3261 ();
 sg13g2_decap_8 FILLER_38_3268 ();
 sg13g2_decap_8 FILLER_38_3275 ();
 sg13g2_decap_8 FILLER_38_3282 ();
 sg13g2_decap_8 FILLER_38_3289 ();
 sg13g2_decap_8 FILLER_38_3296 ();
 sg13g2_decap_8 FILLER_38_3303 ();
 sg13g2_decap_8 FILLER_38_3310 ();
 sg13g2_decap_8 FILLER_38_3317 ();
 sg13g2_decap_8 FILLER_38_3324 ();
 sg13g2_decap_8 FILLER_38_3331 ();
 sg13g2_decap_8 FILLER_38_3338 ();
 sg13g2_decap_8 FILLER_38_3345 ();
 sg13g2_decap_8 FILLER_38_3352 ();
 sg13g2_decap_8 FILLER_38_3359 ();
 sg13g2_decap_8 FILLER_38_3366 ();
 sg13g2_decap_8 FILLER_38_3373 ();
 sg13g2_decap_8 FILLER_38_3380 ();
 sg13g2_decap_8 FILLER_38_3387 ();
 sg13g2_decap_8 FILLER_38_3394 ();
 sg13g2_decap_8 FILLER_38_3401 ();
 sg13g2_decap_8 FILLER_38_3408 ();
 sg13g2_decap_8 FILLER_38_3415 ();
 sg13g2_decap_8 FILLER_38_3422 ();
 sg13g2_decap_8 FILLER_38_3429 ();
 sg13g2_decap_8 FILLER_38_3436 ();
 sg13g2_decap_8 FILLER_38_3443 ();
 sg13g2_decap_8 FILLER_38_3450 ();
 sg13g2_decap_8 FILLER_38_3457 ();
 sg13g2_decap_8 FILLER_38_3464 ();
 sg13g2_decap_8 FILLER_38_3471 ();
 sg13g2_decap_8 FILLER_38_3478 ();
 sg13g2_decap_8 FILLER_38_3485 ();
 sg13g2_decap_8 FILLER_38_3492 ();
 sg13g2_decap_8 FILLER_38_3499 ();
 sg13g2_decap_8 FILLER_38_3506 ();
 sg13g2_decap_8 FILLER_38_3513 ();
 sg13g2_decap_8 FILLER_38_3520 ();
 sg13g2_decap_8 FILLER_38_3527 ();
 sg13g2_decap_8 FILLER_38_3534 ();
 sg13g2_decap_8 FILLER_38_3541 ();
 sg13g2_decap_8 FILLER_38_3548 ();
 sg13g2_decap_8 FILLER_38_3555 ();
 sg13g2_decap_8 FILLER_38_3562 ();
 sg13g2_decap_8 FILLER_38_3569 ();
 sg13g2_decap_4 FILLER_38_3576 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_4 FILLER_39_84 ();
 sg13g2_fill_1 FILLER_39_88 ();
 sg13g2_decap_8 FILLER_39_93 ();
 sg13g2_decap_8 FILLER_39_100 ();
 sg13g2_decap_8 FILLER_39_107 ();
 sg13g2_decap_8 FILLER_39_114 ();
 sg13g2_decap_8 FILLER_39_121 ();
 sg13g2_decap_8 FILLER_39_128 ();
 sg13g2_decap_4 FILLER_39_135 ();
 sg13g2_fill_2 FILLER_39_139 ();
 sg13g2_fill_2 FILLER_39_171 ();
 sg13g2_decap_8 FILLER_39_176 ();
 sg13g2_decap_4 FILLER_39_183 ();
 sg13g2_fill_2 FILLER_39_216 ();
 sg13g2_decap_8 FILLER_39_251 ();
 sg13g2_decap_8 FILLER_39_258 ();
 sg13g2_decap_4 FILLER_39_265 ();
 sg13g2_fill_2 FILLER_39_298 ();
 sg13g2_decap_8 FILLER_39_303 ();
 sg13g2_decap_8 FILLER_39_310 ();
 sg13g2_decap_4 FILLER_39_317 ();
 sg13g2_fill_1 FILLER_39_321 ();
 sg13g2_fill_2 FILLER_39_325 ();
 sg13g2_fill_1 FILLER_39_327 ();
 sg13g2_decap_8 FILLER_39_338 ();
 sg13g2_decap_4 FILLER_39_345 ();
 sg13g2_decap_4 FILLER_39_388 ();
 sg13g2_fill_1 FILLER_39_392 ();
 sg13g2_fill_1 FILLER_39_445 ();
 sg13g2_fill_2 FILLER_39_492 ();
 sg13g2_fill_1 FILLER_39_494 ();
 sg13g2_decap_8 FILLER_39_499 ();
 sg13g2_decap_8 FILLER_39_587 ();
 sg13g2_decap_8 FILLER_39_594 ();
 sg13g2_fill_1 FILLER_39_601 ();
 sg13g2_decap_8 FILLER_39_605 ();
 sg13g2_decap_8 FILLER_39_612 ();
 sg13g2_decap_4 FILLER_39_619 ();
 sg13g2_fill_1 FILLER_39_623 ();
 sg13g2_decap_8 FILLER_39_650 ();
 sg13g2_decap_8 FILLER_39_657 ();
 sg13g2_fill_2 FILLER_39_664 ();
 sg13g2_decap_8 FILLER_39_770 ();
 sg13g2_decap_4 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_889 ();
 sg13g2_decap_8 FILLER_39_896 ();
 sg13g2_decap_8 FILLER_39_903 ();
 sg13g2_fill_2 FILLER_39_910 ();
 sg13g2_fill_1 FILLER_39_912 ();
 sg13g2_decap_8 FILLER_39_951 ();
 sg13g2_decap_8 FILLER_39_958 ();
 sg13g2_decap_8 FILLER_39_1025 ();
 sg13g2_decap_8 FILLER_39_1032 ();
 sg13g2_decap_8 FILLER_39_1039 ();
 sg13g2_fill_2 FILLER_39_1050 ();
 sg13g2_decap_8 FILLER_39_1057 ();
 sg13g2_decap_8 FILLER_39_1090 ();
 sg13g2_fill_2 FILLER_39_1097 ();
 sg13g2_fill_1 FILLER_39_1099 ();
 sg13g2_decap_8 FILLER_39_1152 ();
 sg13g2_fill_2 FILLER_39_1159 ();
 sg13g2_fill_1 FILLER_39_1161 ();
 sg13g2_decap_8 FILLER_39_1168 ();
 sg13g2_decap_8 FILLER_39_1175 ();
 sg13g2_decap_8 FILLER_39_1182 ();
 sg13g2_decap_8 FILLER_39_1189 ();
 sg13g2_fill_2 FILLER_39_1196 ();
 sg13g2_fill_1 FILLER_39_1198 ();
 sg13g2_fill_2 FILLER_39_1220 ();
 sg13g2_fill_1 FILLER_39_1222 ();
 sg13g2_decap_8 FILLER_39_1239 ();
 sg13g2_decap_4 FILLER_39_1246 ();
 sg13g2_fill_1 FILLER_39_1250 ();
 sg13g2_fill_2 FILLER_39_1264 ();
 sg13g2_decap_8 FILLER_39_1270 ();
 sg13g2_fill_2 FILLER_39_1277 ();
 sg13g2_fill_2 FILLER_39_1283 ();
 sg13g2_fill_2 FILLER_39_1349 ();
 sg13g2_fill_1 FILLER_39_1351 ();
 sg13g2_fill_1 FILLER_39_1360 ();
 sg13g2_decap_8 FILLER_39_1366 ();
 sg13g2_fill_2 FILLER_39_1373 ();
 sg13g2_fill_1 FILLER_39_1375 ();
 sg13g2_fill_1 FILLER_39_1389 ();
 sg13g2_decap_8 FILLER_39_1415 ();
 sg13g2_decap_8 FILLER_39_1422 ();
 sg13g2_decap_8 FILLER_39_1429 ();
 sg13g2_fill_2 FILLER_39_1436 ();
 sg13g2_decap_8 FILLER_39_1451 ();
 sg13g2_decap_8 FILLER_39_1458 ();
 sg13g2_decap_4 FILLER_39_1465 ();
 sg13g2_fill_1 FILLER_39_1506 ();
 sg13g2_decap_4 FILLER_39_1519 ();
 sg13g2_fill_2 FILLER_39_1523 ();
 sg13g2_fill_2 FILLER_39_1554 ();
 sg13g2_fill_1 FILLER_39_1556 ();
 sg13g2_decap_4 FILLER_39_1574 ();
 sg13g2_fill_1 FILLER_39_1578 ();
 sg13g2_decap_8 FILLER_39_1608 ();
 sg13g2_fill_2 FILLER_39_1615 ();
 sg13g2_fill_1 FILLER_39_1617 ();
 sg13g2_decap_8 FILLER_39_1654 ();
 sg13g2_decap_8 FILLER_39_1661 ();
 sg13g2_decap_8 FILLER_39_1668 ();
 sg13g2_decap_4 FILLER_39_1675 ();
 sg13g2_fill_1 FILLER_39_1679 ();
 sg13g2_decap_4 FILLER_39_1715 ();
 sg13g2_fill_1 FILLER_39_1719 ();
 sg13g2_fill_2 FILLER_39_1758 ();
 sg13g2_fill_1 FILLER_39_1760 ();
 sg13g2_decap_8 FILLER_39_1804 ();
 sg13g2_decap_8 FILLER_39_1811 ();
 sg13g2_fill_2 FILLER_39_1818 ();
 sg13g2_fill_1 FILLER_39_1820 ();
 sg13g2_decap_8 FILLER_39_1903 ();
 sg13g2_decap_8 FILLER_39_1910 ();
 sg13g2_fill_2 FILLER_39_1917 ();
 sg13g2_decap_8 FILLER_39_1926 ();
 sg13g2_decap_8 FILLER_39_1933 ();
 sg13g2_decap_8 FILLER_39_1940 ();
 sg13g2_decap_8 FILLER_39_1947 ();
 sg13g2_decap_4 FILLER_39_1954 ();
 sg13g2_fill_2 FILLER_39_1982 ();
 sg13g2_fill_1 FILLER_39_1984 ();
 sg13g2_decap_8 FILLER_39_2010 ();
 sg13g2_fill_1 FILLER_39_2017 ();
 sg13g2_decap_8 FILLER_39_2022 ();
 sg13g2_decap_8 FILLER_39_2029 ();
 sg13g2_decap_4 FILLER_39_2036 ();
 sg13g2_decap_8 FILLER_39_2045 ();
 sg13g2_decap_4 FILLER_39_2052 ();
 sg13g2_fill_2 FILLER_39_2056 ();
 sg13g2_decap_8 FILLER_39_2063 ();
 sg13g2_fill_1 FILLER_39_2091 ();
 sg13g2_fill_2 FILLER_39_2100 ();
 sg13g2_fill_1 FILLER_39_2102 ();
 sg13g2_fill_1 FILLER_39_2108 ();
 sg13g2_fill_1 FILLER_39_2117 ();
 sg13g2_fill_2 FILLER_39_2128 ();
 sg13g2_decap_8 FILLER_39_2156 ();
 sg13g2_fill_1 FILLER_39_2163 ();
 sg13g2_decap_8 FILLER_39_2201 ();
 sg13g2_fill_2 FILLER_39_2208 ();
 sg13g2_fill_1 FILLER_39_2210 ();
 sg13g2_fill_1 FILLER_39_2224 ();
 sg13g2_decap_8 FILLER_39_2240 ();
 sg13g2_decap_8 FILLER_39_2247 ();
 sg13g2_decap_8 FILLER_39_2332 ();
 sg13g2_decap_8 FILLER_39_2339 ();
 sg13g2_decap_4 FILLER_39_2346 ();
 sg13g2_fill_2 FILLER_39_2350 ();
 sg13g2_decap_8 FILLER_39_2383 ();
 sg13g2_decap_8 FILLER_39_2390 ();
 sg13g2_decap_8 FILLER_39_2397 ();
 sg13g2_decap_4 FILLER_39_2404 ();
 sg13g2_decap_4 FILLER_39_2448 ();
 sg13g2_fill_2 FILLER_39_2452 ();
 sg13g2_decap_8 FILLER_39_2477 ();
 sg13g2_decap_4 FILLER_39_2484 ();
 sg13g2_fill_1 FILLER_39_2488 ();
 sg13g2_decap_8 FILLER_39_2531 ();
 sg13g2_decap_8 FILLER_39_2538 ();
 sg13g2_fill_1 FILLER_39_2545 ();
 sg13g2_decap_8 FILLER_39_2551 ();
 sg13g2_decap_4 FILLER_39_2558 ();
 sg13g2_fill_2 FILLER_39_2565 ();
 sg13g2_fill_2 FILLER_39_2582 ();
 sg13g2_decap_8 FILLER_39_2587 ();
 sg13g2_decap_8 FILLER_39_2594 ();
 sg13g2_decap_8 FILLER_39_2601 ();
 sg13g2_decap_8 FILLER_39_2608 ();
 sg13g2_decap_4 FILLER_39_2615 ();
 sg13g2_decap_8 FILLER_39_2627 ();
 sg13g2_decap_8 FILLER_39_2634 ();
 sg13g2_decap_8 FILLER_39_2641 ();
 sg13g2_decap_8 FILLER_39_2648 ();
 sg13g2_decap_8 FILLER_39_2655 ();
 sg13g2_decap_8 FILLER_39_2714 ();
 sg13g2_decap_8 FILLER_39_2721 ();
 sg13g2_fill_1 FILLER_39_2728 ();
 sg13g2_fill_2 FILLER_39_2732 ();
 sg13g2_fill_1 FILLER_39_2734 ();
 sg13g2_decap_8 FILLER_39_2775 ();
 sg13g2_decap_8 FILLER_39_2782 ();
 sg13g2_decap_8 FILLER_39_2825 ();
 sg13g2_decap_4 FILLER_39_2832 ();
 sg13g2_fill_1 FILLER_39_2836 ();
 sg13g2_fill_1 FILLER_39_2861 ();
 sg13g2_decap_4 FILLER_39_2866 ();
 sg13g2_fill_1 FILLER_39_2870 ();
 sg13g2_fill_2 FILLER_39_2905 ();
 sg13g2_decap_4 FILLER_39_2911 ();
 sg13g2_fill_2 FILLER_39_2963 ();
 sg13g2_fill_1 FILLER_39_2965 ();
 sg13g2_fill_1 FILLER_39_2969 ();
 sg13g2_fill_1 FILLER_39_2974 ();
 sg13g2_fill_1 FILLER_39_3001 ();
 sg13g2_fill_2 FILLER_39_3039 ();
 sg13g2_decap_8 FILLER_39_3077 ();
 sg13g2_decap_4 FILLER_39_3084 ();
 sg13g2_fill_2 FILLER_39_3088 ();
 sg13g2_decap_8 FILLER_39_3124 ();
 sg13g2_decap_4 FILLER_39_3131 ();
 sg13g2_fill_2 FILLER_39_3135 ();
 sg13g2_decap_8 FILLER_39_3189 ();
 sg13g2_decap_8 FILLER_39_3196 ();
 sg13g2_decap_8 FILLER_39_3229 ();
 sg13g2_decap_8 FILLER_39_3236 ();
 sg13g2_decap_8 FILLER_39_3243 ();
 sg13g2_decap_8 FILLER_39_3250 ();
 sg13g2_decap_8 FILLER_39_3257 ();
 sg13g2_decap_8 FILLER_39_3264 ();
 sg13g2_decap_8 FILLER_39_3271 ();
 sg13g2_decap_8 FILLER_39_3278 ();
 sg13g2_decap_8 FILLER_39_3285 ();
 sg13g2_decap_8 FILLER_39_3292 ();
 sg13g2_decap_8 FILLER_39_3299 ();
 sg13g2_decap_8 FILLER_39_3306 ();
 sg13g2_decap_8 FILLER_39_3313 ();
 sg13g2_decap_8 FILLER_39_3320 ();
 sg13g2_decap_8 FILLER_39_3327 ();
 sg13g2_decap_8 FILLER_39_3334 ();
 sg13g2_decap_8 FILLER_39_3341 ();
 sg13g2_decap_8 FILLER_39_3348 ();
 sg13g2_decap_8 FILLER_39_3355 ();
 sg13g2_decap_8 FILLER_39_3362 ();
 sg13g2_decap_8 FILLER_39_3369 ();
 sg13g2_decap_8 FILLER_39_3376 ();
 sg13g2_decap_8 FILLER_39_3383 ();
 sg13g2_decap_8 FILLER_39_3390 ();
 sg13g2_decap_8 FILLER_39_3397 ();
 sg13g2_decap_8 FILLER_39_3404 ();
 sg13g2_decap_8 FILLER_39_3411 ();
 sg13g2_decap_8 FILLER_39_3418 ();
 sg13g2_decap_8 FILLER_39_3425 ();
 sg13g2_decap_8 FILLER_39_3432 ();
 sg13g2_decap_8 FILLER_39_3439 ();
 sg13g2_decap_8 FILLER_39_3446 ();
 sg13g2_decap_8 FILLER_39_3453 ();
 sg13g2_decap_8 FILLER_39_3460 ();
 sg13g2_decap_8 FILLER_39_3467 ();
 sg13g2_decap_8 FILLER_39_3474 ();
 sg13g2_decap_8 FILLER_39_3481 ();
 sg13g2_decap_8 FILLER_39_3488 ();
 sg13g2_decap_8 FILLER_39_3495 ();
 sg13g2_decap_8 FILLER_39_3502 ();
 sg13g2_decap_8 FILLER_39_3509 ();
 sg13g2_decap_8 FILLER_39_3516 ();
 sg13g2_decap_8 FILLER_39_3523 ();
 sg13g2_decap_8 FILLER_39_3530 ();
 sg13g2_decap_8 FILLER_39_3537 ();
 sg13g2_decap_8 FILLER_39_3544 ();
 sg13g2_decap_8 FILLER_39_3551 ();
 sg13g2_decap_8 FILLER_39_3558 ();
 sg13g2_decap_8 FILLER_39_3565 ();
 sg13g2_decap_8 FILLER_39_3572 ();
 sg13g2_fill_1 FILLER_39_3579 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_151 ();
 sg13g2_decap_8 FILLER_40_158 ();
 sg13g2_fill_2 FILLER_40_165 ();
 sg13g2_fill_1 FILLER_40_167 ();
 sg13g2_decap_8 FILLER_40_194 ();
 sg13g2_decap_8 FILLER_40_201 ();
 sg13g2_fill_2 FILLER_40_215 ();
 sg13g2_decap_8 FILLER_40_248 ();
 sg13g2_decap_8 FILLER_40_255 ();
 sg13g2_fill_2 FILLER_40_262 ();
 sg13g2_decap_4 FILLER_40_293 ();
 sg13g2_fill_1 FILLER_40_297 ();
 sg13g2_fill_1 FILLER_40_324 ();
 sg13g2_decap_8 FILLER_40_351 ();
 sg13g2_decap_4 FILLER_40_358 ();
 sg13g2_fill_2 FILLER_40_362 ();
 sg13g2_fill_2 FILLER_40_368 ();
 sg13g2_decap_4 FILLER_40_399 ();
 sg13g2_decap_4 FILLER_40_411 ();
 sg13g2_decap_4 FILLER_40_421 ();
 sg13g2_fill_1 FILLER_40_425 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_4 FILLER_40_441 ();
 sg13g2_fill_1 FILLER_40_445 ();
 sg13g2_decap_8 FILLER_40_451 ();
 sg13g2_decap_4 FILLER_40_458 ();
 sg13g2_fill_1 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_466 ();
 sg13g2_fill_2 FILLER_40_473 ();
 sg13g2_fill_1 FILLER_40_475 ();
 sg13g2_decap_8 FILLER_40_508 ();
 sg13g2_decap_8 FILLER_40_515 ();
 sg13g2_fill_2 FILLER_40_561 ();
 sg13g2_fill_1 FILLER_40_563 ();
 sg13g2_fill_1 FILLER_40_593 ();
 sg13g2_fill_2 FILLER_40_599 ();
 sg13g2_fill_1 FILLER_40_627 ();
 sg13g2_fill_1 FILLER_40_654 ();
 sg13g2_decap_8 FILLER_40_717 ();
 sg13g2_decap_4 FILLER_40_724 ();
 sg13g2_fill_2 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_733 ();
 sg13g2_decap_8 FILLER_40_766 ();
 sg13g2_decap_8 FILLER_40_773 ();
 sg13g2_decap_8 FILLER_40_780 ();
 sg13g2_decap_4 FILLER_40_787 ();
 sg13g2_fill_1 FILLER_40_791 ();
 sg13g2_decap_4 FILLER_40_828 ();
 sg13g2_fill_1 FILLER_40_832 ();
 sg13g2_fill_2 FILLER_40_838 ();
 sg13g2_fill_1 FILLER_40_891 ();
 sg13g2_fill_2 FILLER_40_897 ();
 sg13g2_fill_2 FILLER_40_904 ();
 sg13g2_decap_8 FILLER_40_943 ();
 sg13g2_decap_4 FILLER_40_950 ();
 sg13g2_fill_2 FILLER_40_954 ();
 sg13g2_decap_8 FILLER_40_960 ();
 sg13g2_decap_8 FILLER_40_1031 ();
 sg13g2_fill_2 FILLER_40_1038 ();
 sg13g2_fill_2 FILLER_40_1045 ();
 sg13g2_fill_1 FILLER_40_1047 ();
 sg13g2_decap_8 FILLER_40_1082 ();
 sg13g2_decap_8 FILLER_40_1089 ();
 sg13g2_fill_1 FILLER_40_1096 ();
 sg13g2_fill_1 FILLER_40_1155 ();
 sg13g2_decap_8 FILLER_40_1182 ();
 sg13g2_decap_8 FILLER_40_1189 ();
 sg13g2_decap_8 FILLER_40_1196 ();
 sg13g2_fill_2 FILLER_40_1203 ();
 sg13g2_fill_2 FILLER_40_1218 ();
 sg13g2_decap_8 FILLER_40_1232 ();
 sg13g2_decap_8 FILLER_40_1239 ();
 sg13g2_decap_8 FILLER_40_1246 ();
 sg13g2_decap_8 FILLER_40_1253 ();
 sg13g2_decap_8 FILLER_40_1260 ();
 sg13g2_decap_8 FILLER_40_1267 ();
 sg13g2_decap_4 FILLER_40_1274 ();
 sg13g2_fill_1 FILLER_40_1278 ();
 sg13g2_fill_2 FILLER_40_1299 ();
 sg13g2_fill_1 FILLER_40_1343 ();
 sg13g2_decap_8 FILLER_40_1352 ();
 sg13g2_decap_8 FILLER_40_1359 ();
 sg13g2_decap_8 FILLER_40_1366 ();
 sg13g2_decap_8 FILLER_40_1373 ();
 sg13g2_decap_8 FILLER_40_1380 ();
 sg13g2_decap_8 FILLER_40_1387 ();
 sg13g2_decap_4 FILLER_40_1394 ();
 sg13g2_fill_2 FILLER_40_1436 ();
 sg13g2_decap_8 FILLER_40_1447 ();
 sg13g2_decap_8 FILLER_40_1454 ();
 sg13g2_decap_4 FILLER_40_1461 ();
 sg13g2_fill_1 FILLER_40_1465 ();
 sg13g2_decap_4 FILLER_40_1474 ();
 sg13g2_fill_1 FILLER_40_1478 ();
 sg13g2_decap_4 FILLER_40_1501 ();
 sg13g2_decap_4 FILLER_40_1521 ();
 sg13g2_fill_2 FILLER_40_1525 ();
 sg13g2_fill_1 FILLER_40_1553 ();
 sg13g2_decap_8 FILLER_40_1652 ();
 sg13g2_decap_8 FILLER_40_1659 ();
 sg13g2_fill_2 FILLER_40_1666 ();
 sg13g2_fill_1 FILLER_40_1668 ();
 sg13g2_fill_2 FILLER_40_1690 ();
 sg13g2_fill_2 FILLER_40_1749 ();
 sg13g2_decap_8 FILLER_40_1803 ();
 sg13g2_decap_4 FILLER_40_1810 ();
 sg13g2_decap_8 FILLER_40_1822 ();
 sg13g2_fill_2 FILLER_40_1833 ();
 sg13g2_decap_4 FILLER_40_1844 ();
 sg13g2_fill_1 FILLER_40_1853 ();
 sg13g2_decap_8 FILLER_40_1868 ();
 sg13g2_fill_1 FILLER_40_1875 ();
 sg13g2_fill_1 FILLER_40_1982 ();
 sg13g2_decap_8 FILLER_40_1988 ();
 sg13g2_fill_2 FILLER_40_2000 ();
 sg13g2_decap_4 FILLER_40_2064 ();
 sg13g2_fill_1 FILLER_40_2095 ();
 sg13g2_fill_1 FILLER_40_2136 ();
 sg13g2_decap_8 FILLER_40_2147 ();
 sg13g2_decap_4 FILLER_40_2154 ();
 sg13g2_decap_8 FILLER_40_2196 ();
 sg13g2_fill_2 FILLER_40_2203 ();
 sg13g2_fill_1 FILLER_40_2213 ();
 sg13g2_decap_8 FILLER_40_2240 ();
 sg13g2_decap_8 FILLER_40_2247 ();
 sg13g2_fill_2 FILLER_40_2254 ();
 sg13g2_fill_1 FILLER_40_2256 ();
 sg13g2_fill_2 FILLER_40_2296 ();
 sg13g2_decap_8 FILLER_40_2324 ();
 sg13g2_decap_8 FILLER_40_2331 ();
 sg13g2_fill_2 FILLER_40_2338 ();
 sg13g2_fill_1 FILLER_40_2340 ();
 sg13g2_decap_4 FILLER_40_2349 ();
 sg13g2_decap_8 FILLER_40_2387 ();
 sg13g2_decap_8 FILLER_40_2394 ();
 sg13g2_decap_8 FILLER_40_2401 ();
 sg13g2_decap_8 FILLER_40_2408 ();
 sg13g2_decap_4 FILLER_40_2415 ();
 sg13g2_fill_1 FILLER_40_2419 ();
 sg13g2_fill_2 FILLER_40_2480 ();
 sg13g2_fill_1 FILLER_40_2482 ();
 sg13g2_fill_2 FILLER_40_2507 ();
 sg13g2_decap_8 FILLER_40_2535 ();
 sg13g2_fill_2 FILLER_40_2542 ();
 sg13g2_fill_1 FILLER_40_2544 ();
 sg13g2_decap_8 FILLER_40_2579 ();
 sg13g2_decap_8 FILLER_40_2586 ();
 sg13g2_decap_8 FILLER_40_2593 ();
 sg13g2_decap_8 FILLER_40_2600 ();
 sg13g2_decap_4 FILLER_40_2607 ();
 sg13g2_fill_1 FILLER_40_2611 ();
 sg13g2_fill_1 FILLER_40_2648 ();
 sg13g2_fill_1 FILLER_40_2701 ();
 sg13g2_fill_2 FILLER_40_2706 ();
 sg13g2_decap_8 FILLER_40_2768 ();
 sg13g2_fill_2 FILLER_40_2775 ();
 sg13g2_decap_8 FILLER_40_2782 ();
 sg13g2_fill_2 FILLER_40_2789 ();
 sg13g2_decap_8 FILLER_40_2817 ();
 sg13g2_decap_8 FILLER_40_2824 ();
 sg13g2_fill_1 FILLER_40_2831 ();
 sg13g2_decap_8 FILLER_40_2850 ();
 sg13g2_fill_2 FILLER_40_2857 ();
 sg13g2_fill_1 FILLER_40_2859 ();
 sg13g2_fill_1 FILLER_40_2868 ();
 sg13g2_fill_1 FILLER_40_2903 ();
 sg13g2_decap_8 FILLER_40_2954 ();
 sg13g2_fill_1 FILLER_40_2961 ();
 sg13g2_decap_8 FILLER_40_3077 ();
 sg13g2_fill_2 FILLER_40_3084 ();
 sg13g2_decap_8 FILLER_40_3124 ();
 sg13g2_decap_4 FILLER_40_3131 ();
 sg13g2_fill_1 FILLER_40_3135 ();
 sg13g2_decap_8 FILLER_40_3171 ();
 sg13g2_decap_8 FILLER_40_3178 ();
 sg13g2_decap_8 FILLER_40_3185 ();
 sg13g2_decap_8 FILLER_40_3192 ();
 sg13g2_fill_1 FILLER_40_3230 ();
 sg13g2_decap_8 FILLER_40_3238 ();
 sg13g2_fill_1 FILLER_40_3245 ();
 sg13g2_decap_8 FILLER_40_3250 ();
 sg13g2_decap_8 FILLER_40_3257 ();
 sg13g2_decap_8 FILLER_40_3264 ();
 sg13g2_decap_8 FILLER_40_3271 ();
 sg13g2_decap_8 FILLER_40_3278 ();
 sg13g2_decap_8 FILLER_40_3285 ();
 sg13g2_decap_8 FILLER_40_3292 ();
 sg13g2_decap_8 FILLER_40_3299 ();
 sg13g2_decap_8 FILLER_40_3306 ();
 sg13g2_decap_8 FILLER_40_3313 ();
 sg13g2_decap_8 FILLER_40_3320 ();
 sg13g2_decap_8 FILLER_40_3327 ();
 sg13g2_decap_8 FILLER_40_3334 ();
 sg13g2_decap_8 FILLER_40_3341 ();
 sg13g2_decap_8 FILLER_40_3348 ();
 sg13g2_decap_8 FILLER_40_3355 ();
 sg13g2_decap_8 FILLER_40_3362 ();
 sg13g2_decap_8 FILLER_40_3369 ();
 sg13g2_decap_8 FILLER_40_3376 ();
 sg13g2_decap_8 FILLER_40_3383 ();
 sg13g2_decap_8 FILLER_40_3390 ();
 sg13g2_decap_8 FILLER_40_3397 ();
 sg13g2_decap_8 FILLER_40_3404 ();
 sg13g2_decap_8 FILLER_40_3411 ();
 sg13g2_decap_8 FILLER_40_3418 ();
 sg13g2_decap_8 FILLER_40_3425 ();
 sg13g2_decap_8 FILLER_40_3432 ();
 sg13g2_decap_8 FILLER_40_3439 ();
 sg13g2_decap_8 FILLER_40_3446 ();
 sg13g2_decap_8 FILLER_40_3453 ();
 sg13g2_decap_8 FILLER_40_3460 ();
 sg13g2_decap_8 FILLER_40_3467 ();
 sg13g2_decap_8 FILLER_40_3474 ();
 sg13g2_decap_8 FILLER_40_3481 ();
 sg13g2_decap_8 FILLER_40_3488 ();
 sg13g2_decap_8 FILLER_40_3495 ();
 sg13g2_decap_8 FILLER_40_3502 ();
 sg13g2_decap_8 FILLER_40_3509 ();
 sg13g2_decap_8 FILLER_40_3516 ();
 sg13g2_decap_8 FILLER_40_3523 ();
 sg13g2_decap_8 FILLER_40_3530 ();
 sg13g2_decap_8 FILLER_40_3537 ();
 sg13g2_decap_8 FILLER_40_3544 ();
 sg13g2_decap_8 FILLER_40_3551 ();
 sg13g2_decap_8 FILLER_40_3558 ();
 sg13g2_decap_8 FILLER_40_3565 ();
 sg13g2_decap_8 FILLER_40_3572 ();
 sg13g2_fill_1 FILLER_40_3579 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_fill_2 FILLER_41_175 ();
 sg13g2_fill_1 FILLER_41_177 ();
 sg13g2_decap_8 FILLER_41_183 ();
 sg13g2_decap_8 FILLER_41_190 ();
 sg13g2_decap_8 FILLER_41_197 ();
 sg13g2_decap_8 FILLER_41_204 ();
 sg13g2_decap_8 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_221 ();
 sg13g2_decap_8 FILLER_41_233 ();
 sg13g2_decap_8 FILLER_41_240 ();
 sg13g2_decap_8 FILLER_41_247 ();
 sg13g2_decap_8 FILLER_41_254 ();
 sg13g2_decap_8 FILLER_41_261 ();
 sg13g2_decap_4 FILLER_41_268 ();
 sg13g2_fill_1 FILLER_41_301 ();
 sg13g2_fill_1 FILLER_41_335 ();
 sg13g2_decap_8 FILLER_41_340 ();
 sg13g2_decap_8 FILLER_41_347 ();
 sg13g2_fill_1 FILLER_41_354 ();
 sg13g2_decap_8 FILLER_41_398 ();
 sg13g2_decap_8 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_41_412 ();
 sg13g2_decap_8 FILLER_41_419 ();
 sg13g2_decap_8 FILLER_41_426 ();
 sg13g2_decap_8 FILLER_41_433 ();
 sg13g2_decap_8 FILLER_41_440 ();
 sg13g2_fill_2 FILLER_41_447 ();
 sg13g2_fill_1 FILLER_41_449 ();
 sg13g2_decap_8 FILLER_41_480 ();
 sg13g2_decap_8 FILLER_41_487 ();
 sg13g2_decap_4 FILLER_41_494 ();
 sg13g2_fill_1 FILLER_41_498 ();
 sg13g2_fill_2 FILLER_41_510 ();
 sg13g2_fill_1 FILLER_41_512 ();
 sg13g2_decap_8 FILLER_41_542 ();
 sg13g2_decap_8 FILLER_41_549 ();
 sg13g2_decap_8 FILLER_41_556 ();
 sg13g2_decap_4 FILLER_41_563 ();
 sg13g2_fill_2 FILLER_41_572 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_decap_4 FILLER_41_602 ();
 sg13g2_fill_1 FILLER_41_606 ();
 sg13g2_decap_8 FILLER_41_636 ();
 sg13g2_decap_8 FILLER_41_643 ();
 sg13g2_decap_8 FILLER_41_650 ();
 sg13g2_decap_8 FILLER_41_657 ();
 sg13g2_decap_8 FILLER_41_664 ();
 sg13g2_fill_2 FILLER_41_671 ();
 sg13g2_fill_1 FILLER_41_673 ();
 sg13g2_decap_8 FILLER_41_706 ();
 sg13g2_decap_8 FILLER_41_713 ();
 sg13g2_decap_8 FILLER_41_720 ();
 sg13g2_decap_8 FILLER_41_727 ();
 sg13g2_decap_8 FILLER_41_734 ();
 sg13g2_fill_2 FILLER_41_741 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_decap_8 FILLER_41_759 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_decap_8 FILLER_41_773 ();
 sg13g2_decap_4 FILLER_41_780 ();
 sg13g2_fill_1 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_816 ();
 sg13g2_decap_8 FILLER_41_823 ();
 sg13g2_decap_4 FILLER_41_830 ();
 sg13g2_decap_8 FILLER_41_873 ();
 sg13g2_decap_8 FILLER_41_880 ();
 sg13g2_fill_2 FILLER_41_913 ();
 sg13g2_fill_1 FILLER_41_925 ();
 sg13g2_decap_8 FILLER_41_936 ();
 sg13g2_decap_4 FILLER_41_957 ();
 sg13g2_fill_2 FILLER_41_961 ();
 sg13g2_decap_8 FILLER_41_968 ();
 sg13g2_decap_8 FILLER_41_975 ();
 sg13g2_decap_8 FILLER_41_982 ();
 sg13g2_decap_8 FILLER_41_989 ();
 sg13g2_fill_2 FILLER_41_1034 ();
 sg13g2_fill_2 FILLER_41_1062 ();
 sg13g2_fill_1 FILLER_41_1064 ();
 sg13g2_decap_4 FILLER_41_1097 ();
 sg13g2_decap_8 FILLER_41_1190 ();
 sg13g2_fill_2 FILLER_41_1205 ();
 sg13g2_fill_1 FILLER_41_1207 ();
 sg13g2_fill_1 FILLER_41_1216 ();
 sg13g2_decap_8 FILLER_41_1225 ();
 sg13g2_decap_4 FILLER_41_1232 ();
 sg13g2_fill_2 FILLER_41_1236 ();
 sg13g2_decap_4 FILLER_41_1246 ();
 sg13g2_fill_1 FILLER_41_1250 ();
 sg13g2_fill_2 FILLER_41_1277 ();
 sg13g2_decap_8 FILLER_41_1283 ();
 sg13g2_decap_8 FILLER_41_1290 ();
 sg13g2_decap_4 FILLER_41_1297 ();
 sg13g2_fill_1 FILLER_41_1301 ();
 sg13g2_fill_2 FILLER_41_1310 ();
 sg13g2_decap_8 FILLER_41_1343 ();
 sg13g2_decap_8 FILLER_41_1350 ();
 sg13g2_decap_8 FILLER_41_1357 ();
 sg13g2_decap_8 FILLER_41_1364 ();
 sg13g2_decap_4 FILLER_41_1371 ();
 sg13g2_fill_2 FILLER_41_1375 ();
 sg13g2_fill_1 FILLER_41_1403 ();
 sg13g2_fill_1 FILLER_41_1444 ();
 sg13g2_decap_8 FILLER_41_1453 ();
 sg13g2_decap_4 FILLER_41_1460 ();
 sg13g2_fill_1 FILLER_41_1464 ();
 sg13g2_decap_8 FILLER_41_1473 ();
 sg13g2_decap_8 FILLER_41_1480 ();
 sg13g2_decap_8 FILLER_41_1491 ();
 sg13g2_decap_8 FILLER_41_1498 ();
 sg13g2_decap_4 FILLER_41_1505 ();
 sg13g2_fill_1 FILLER_41_1514 ();
 sg13g2_decap_8 FILLER_41_1572 ();
 sg13g2_fill_2 FILLER_41_1579 ();
 sg13g2_decap_8 FILLER_41_1607 ();
 sg13g2_decap_8 FILLER_41_1614 ();
 sg13g2_fill_1 FILLER_41_1621 ();
 sg13g2_decap_8 FILLER_41_1651 ();
 sg13g2_decap_8 FILLER_41_1658 ();
 sg13g2_fill_2 FILLER_41_1672 ();
 sg13g2_decap_4 FILLER_41_1726 ();
 sg13g2_decap_4 FILLER_41_1750 ();
 sg13g2_decap_8 FILLER_41_1758 ();
 sg13g2_decap_8 FILLER_41_1765 ();
 sg13g2_decap_4 FILLER_41_1803 ();
 sg13g2_fill_1 FILLER_41_1807 ();
 sg13g2_decap_8 FILLER_41_1813 ();
 sg13g2_fill_2 FILLER_41_1820 ();
 sg13g2_fill_1 FILLER_41_1852 ();
 sg13g2_fill_1 FILLER_41_1904 ();
 sg13g2_decap_4 FILLER_41_1945 ();
 sg13g2_fill_1 FILLER_41_1949 ();
 sg13g2_fill_2 FILLER_41_1973 ();
 sg13g2_fill_2 FILLER_41_1988 ();
 sg13g2_fill_2 FILLER_41_2024 ();
 sg13g2_fill_1 FILLER_41_2026 ();
 sg13g2_fill_1 FILLER_41_2031 ();
 sg13g2_fill_2 FILLER_41_2036 ();
 sg13g2_fill_1 FILLER_41_2038 ();
 sg13g2_fill_1 FILLER_41_2044 ();
 sg13g2_decap_4 FILLER_41_2057 ();
 sg13g2_fill_2 FILLER_41_2061 ();
 sg13g2_fill_2 FILLER_41_2071 ();
 sg13g2_fill_1 FILLER_41_2073 ();
 sg13g2_fill_2 FILLER_41_2106 ();
 sg13g2_decap_8 FILLER_41_2137 ();
 sg13g2_decap_4 FILLER_41_2144 ();
 sg13g2_fill_1 FILLER_41_2148 ();
 sg13g2_decap_8 FILLER_41_2186 ();
 sg13g2_decap_8 FILLER_41_2193 ();
 sg13g2_decap_4 FILLER_41_2200 ();
 sg13g2_fill_1 FILLER_41_2204 ();
 sg13g2_decap_8 FILLER_41_2252 ();
 sg13g2_decap_4 FILLER_41_2274 ();
 sg13g2_decap_8 FILLER_41_2330 ();
 sg13g2_decap_8 FILLER_41_2337 ();
 sg13g2_decap_8 FILLER_41_2344 ();
 sg13g2_decap_4 FILLER_41_2351 ();
 sg13g2_decap_8 FILLER_41_2400 ();
 sg13g2_decap_8 FILLER_41_2407 ();
 sg13g2_decap_4 FILLER_41_2414 ();
 sg13g2_fill_2 FILLER_41_2418 ();
 sg13g2_decap_8 FILLER_41_2446 ();
 sg13g2_decap_8 FILLER_41_2453 ();
 sg13g2_decap_4 FILLER_41_2460 ();
 sg13g2_decap_8 FILLER_41_2477 ();
 sg13g2_decap_8 FILLER_41_2484 ();
 sg13g2_decap_8 FILLER_41_2531 ();
 sg13g2_decap_8 FILLER_41_2538 ();
 sg13g2_decap_8 FILLER_41_2579 ();
 sg13g2_decap_8 FILLER_41_2586 ();
 sg13g2_decap_8 FILLER_41_2593 ();
 sg13g2_fill_2 FILLER_41_2652 ();
 sg13g2_fill_1 FILLER_41_2654 ();
 sg13g2_fill_2 FILLER_41_2685 ();
 sg13g2_fill_1 FILLER_41_2687 ();
 sg13g2_decap_8 FILLER_41_2693 ();
 sg13g2_decap_8 FILLER_41_2700 ();
 sg13g2_fill_2 FILLER_41_2707 ();
 sg13g2_fill_1 FILLER_41_2709 ();
 sg13g2_fill_2 FILLER_41_2769 ();
 sg13g2_fill_1 FILLER_41_2771 ();
 sg13g2_decap_8 FILLER_41_2905 ();
 sg13g2_fill_1 FILLER_41_2925 ();
 sg13g2_fill_1 FILLER_41_2934 ();
 sg13g2_decap_8 FILLER_41_2948 ();
 sg13g2_decap_8 FILLER_41_2955 ();
 sg13g2_decap_8 FILLER_41_2962 ();
 sg13g2_fill_1 FILLER_41_2969 ();
 sg13g2_fill_1 FILLER_41_2977 ();
 sg13g2_fill_2 FILLER_41_3000 ();
 sg13g2_fill_2 FILLER_41_3028 ();
 sg13g2_fill_1 FILLER_41_3030 ();
 sg13g2_fill_2 FILLER_41_3052 ();
 sg13g2_decap_4 FILLER_41_3061 ();
 sg13g2_decap_4 FILLER_41_3075 ();
 sg13g2_decap_8 FILLER_41_3120 ();
 sg13g2_decap_4 FILLER_41_3127 ();
 sg13g2_decap_4 FILLER_41_3162 ();
 sg13g2_fill_2 FILLER_41_3166 ();
 sg13g2_decap_8 FILLER_41_3172 ();
 sg13g2_fill_2 FILLER_41_3179 ();
 sg13g2_fill_1 FILLER_41_3181 ();
 sg13g2_fill_2 FILLER_41_3195 ();
 sg13g2_decap_8 FILLER_41_3261 ();
 sg13g2_decap_8 FILLER_41_3268 ();
 sg13g2_decap_8 FILLER_41_3275 ();
 sg13g2_decap_8 FILLER_41_3282 ();
 sg13g2_decap_8 FILLER_41_3289 ();
 sg13g2_decap_8 FILLER_41_3296 ();
 sg13g2_decap_8 FILLER_41_3303 ();
 sg13g2_decap_8 FILLER_41_3310 ();
 sg13g2_decap_8 FILLER_41_3317 ();
 sg13g2_decap_8 FILLER_41_3324 ();
 sg13g2_decap_8 FILLER_41_3331 ();
 sg13g2_decap_8 FILLER_41_3338 ();
 sg13g2_decap_8 FILLER_41_3345 ();
 sg13g2_decap_8 FILLER_41_3352 ();
 sg13g2_decap_8 FILLER_41_3359 ();
 sg13g2_decap_8 FILLER_41_3366 ();
 sg13g2_decap_8 FILLER_41_3373 ();
 sg13g2_decap_8 FILLER_41_3380 ();
 sg13g2_decap_8 FILLER_41_3387 ();
 sg13g2_decap_8 FILLER_41_3394 ();
 sg13g2_decap_8 FILLER_41_3401 ();
 sg13g2_decap_8 FILLER_41_3408 ();
 sg13g2_decap_8 FILLER_41_3415 ();
 sg13g2_decap_8 FILLER_41_3422 ();
 sg13g2_decap_8 FILLER_41_3429 ();
 sg13g2_decap_8 FILLER_41_3436 ();
 sg13g2_decap_8 FILLER_41_3443 ();
 sg13g2_decap_8 FILLER_41_3450 ();
 sg13g2_decap_8 FILLER_41_3457 ();
 sg13g2_decap_8 FILLER_41_3464 ();
 sg13g2_decap_8 FILLER_41_3471 ();
 sg13g2_decap_8 FILLER_41_3478 ();
 sg13g2_decap_8 FILLER_41_3485 ();
 sg13g2_decap_8 FILLER_41_3492 ();
 sg13g2_decap_8 FILLER_41_3499 ();
 sg13g2_decap_8 FILLER_41_3506 ();
 sg13g2_decap_8 FILLER_41_3513 ();
 sg13g2_decap_8 FILLER_41_3520 ();
 sg13g2_decap_8 FILLER_41_3527 ();
 sg13g2_decap_8 FILLER_41_3534 ();
 sg13g2_decap_8 FILLER_41_3541 ();
 sg13g2_decap_8 FILLER_41_3548 ();
 sg13g2_decap_8 FILLER_41_3555 ();
 sg13g2_decap_8 FILLER_41_3562 ();
 sg13g2_decap_8 FILLER_41_3569 ();
 sg13g2_decap_4 FILLER_41_3576 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_4 FILLER_42_105 ();
 sg13g2_fill_1 FILLER_42_109 ();
 sg13g2_decap_8 FILLER_42_141 ();
 sg13g2_decap_8 FILLER_42_148 ();
 sg13g2_decap_8 FILLER_42_155 ();
 sg13g2_decap_4 FILLER_42_162 ();
 sg13g2_fill_1 FILLER_42_166 ();
 sg13g2_decap_8 FILLER_42_198 ();
 sg13g2_decap_8 FILLER_42_205 ();
 sg13g2_fill_2 FILLER_42_212 ();
 sg13g2_fill_1 FILLER_42_214 ();
 sg13g2_decap_8 FILLER_42_241 ();
 sg13g2_decap_8 FILLER_42_248 ();
 sg13g2_decap_8 FILLER_42_255 ();
 sg13g2_decap_8 FILLER_42_262 ();
 sg13g2_decap_4 FILLER_42_269 ();
 sg13g2_fill_1 FILLER_42_307 ();
 sg13g2_decap_8 FILLER_42_341 ();
 sg13g2_decap_8 FILLER_42_348 ();
 sg13g2_fill_2 FILLER_42_355 ();
 sg13g2_decap_8 FILLER_42_388 ();
 sg13g2_decap_8 FILLER_42_395 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_decap_4 FILLER_42_409 ();
 sg13g2_fill_1 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_443 ();
 sg13g2_decap_8 FILLER_42_450 ();
 sg13g2_fill_2 FILLER_42_457 ();
 sg13g2_fill_1 FILLER_42_459 ();
 sg13g2_decap_4 FILLER_42_492 ();
 sg13g2_decap_8 FILLER_42_500 ();
 sg13g2_fill_2 FILLER_42_507 ();
 sg13g2_fill_1 FILLER_42_509 ();
 sg13g2_decap_8 FILLER_42_543 ();
 sg13g2_fill_2 FILLER_42_550 ();
 sg13g2_fill_1 FILLER_42_552 ();
 sg13g2_fill_2 FILLER_42_556 ();
 sg13g2_fill_1 FILLER_42_558 ();
 sg13g2_decap_8 FILLER_42_563 ();
 sg13g2_decap_8 FILLER_42_578 ();
 sg13g2_decap_8 FILLER_42_585 ();
 sg13g2_decap_8 FILLER_42_592 ();
 sg13g2_fill_2 FILLER_42_599 ();
 sg13g2_fill_2 FILLER_42_604 ();
 sg13g2_decap_8 FILLER_42_636 ();
 sg13g2_decap_8 FILLER_42_643 ();
 sg13g2_decap_8 FILLER_42_650 ();
 sg13g2_decap_8 FILLER_42_657 ();
 sg13g2_decap_8 FILLER_42_664 ();
 sg13g2_decap_8 FILLER_42_671 ();
 sg13g2_decap_8 FILLER_42_678 ();
 sg13g2_fill_1 FILLER_42_685 ();
 sg13g2_decap_8 FILLER_42_692 ();
 sg13g2_decap_8 FILLER_42_699 ();
 sg13g2_decap_8 FILLER_42_706 ();
 sg13g2_decap_8 FILLER_42_713 ();
 sg13g2_decap_8 FILLER_42_720 ();
 sg13g2_decap_8 FILLER_42_727 ();
 sg13g2_decap_8 FILLER_42_734 ();
 sg13g2_fill_2 FILLER_42_741 ();
 sg13g2_decap_4 FILLER_42_769 ();
 sg13g2_decap_8 FILLER_42_799 ();
 sg13g2_decap_8 FILLER_42_806 ();
 sg13g2_decap_8 FILLER_42_813 ();
 sg13g2_decap_8 FILLER_42_820 ();
 sg13g2_decap_8 FILLER_42_827 ();
 sg13g2_decap_8 FILLER_42_834 ();
 sg13g2_fill_2 FILLER_42_841 ();
 sg13g2_fill_1 FILLER_42_843 ();
 sg13g2_decap_8 FILLER_42_870 ();
 sg13g2_decap_8 FILLER_42_877 ();
 sg13g2_decap_8 FILLER_42_884 ();
 sg13g2_decap_4 FILLER_42_891 ();
 sg13g2_fill_2 FILLER_42_895 ();
 sg13g2_decap_8 FILLER_42_923 ();
 sg13g2_decap_4 FILLER_42_930 ();
 sg13g2_fill_2 FILLER_42_934 ();
 sg13g2_decap_4 FILLER_42_951 ();
 sg13g2_fill_2 FILLER_42_965 ();
 sg13g2_decap_8 FILLER_42_975 ();
 sg13g2_decap_8 FILLER_42_982 ();
 sg13g2_decap_8 FILLER_42_989 ();
 sg13g2_decap_4 FILLER_42_996 ();
 sg13g2_fill_2 FILLER_42_1000 ();
 sg13g2_decap_8 FILLER_42_1041 ();
 sg13g2_fill_2 FILLER_42_1079 ();
 sg13g2_fill_1 FILLER_42_1081 ();
 sg13g2_fill_2 FILLER_42_1087 ();
 sg13g2_decap_4 FILLER_42_1145 ();
 sg13g2_fill_2 FILLER_42_1149 ();
 sg13g2_fill_2 FILLER_42_1189 ();
 sg13g2_fill_1 FILLER_42_1191 ();
 sg13g2_fill_2 FILLER_42_1221 ();
 sg13g2_fill_1 FILLER_42_1223 ();
 sg13g2_fill_1 FILLER_42_1236 ();
 sg13g2_decap_8 FILLER_42_1242 ();
 sg13g2_decap_8 FILLER_42_1287 ();
 sg13g2_decap_8 FILLER_42_1294 ();
 sg13g2_fill_2 FILLER_42_1301 ();
 sg13g2_fill_1 FILLER_42_1303 ();
 sg13g2_fill_1 FILLER_42_1309 ();
 sg13g2_decap_8 FILLER_42_1314 ();
 sg13g2_fill_1 FILLER_42_1321 ();
 sg13g2_fill_2 FILLER_42_1326 ();
 sg13g2_fill_1 FILLER_42_1354 ();
 sg13g2_decap_8 FILLER_42_1407 ();
 sg13g2_fill_1 FILLER_42_1414 ();
 sg13g2_decap_4 FILLER_42_1420 ();
 sg13g2_fill_2 FILLER_42_1424 ();
 sg13g2_fill_2 FILLER_42_1436 ();
 sg13g2_fill_1 FILLER_42_1438 ();
 sg13g2_fill_2 FILLER_42_1498 ();
 sg13g2_fill_1 FILLER_42_1526 ();
 sg13g2_fill_2 FILLER_42_1547 ();
 sg13g2_fill_1 FILLER_42_1552 ();
 sg13g2_fill_1 FILLER_42_1561 ();
 sg13g2_decap_8 FILLER_42_1577 ();
 sg13g2_fill_2 FILLER_42_1584 ();
 sg13g2_decap_8 FILLER_42_1612 ();
 sg13g2_decap_8 FILLER_42_1619 ();
 sg13g2_decap_4 FILLER_42_1626 ();
 sg13g2_fill_2 FILLER_42_1635 ();
 sg13g2_decap_8 FILLER_42_1645 ();
 sg13g2_decap_8 FILLER_42_1652 ();
 sg13g2_decap_8 FILLER_42_1691 ();
 sg13g2_decap_4 FILLER_42_1732 ();
 sg13g2_fill_2 FILLER_42_1736 ();
 sg13g2_decap_8 FILLER_42_1744 ();
 sg13g2_decap_8 FILLER_42_1751 ();
 sg13g2_decap_8 FILLER_42_1758 ();
 sg13g2_decap_8 FILLER_42_1816 ();
 sg13g2_decap_8 FILLER_42_1823 ();
 sg13g2_fill_1 FILLER_42_1837 ();
 sg13g2_fill_1 FILLER_42_1846 ();
 sg13g2_fill_2 FILLER_42_1860 ();
 sg13g2_fill_1 FILLER_42_1862 ();
 sg13g2_fill_1 FILLER_42_1868 ();
 sg13g2_decap_4 FILLER_42_1882 ();
 sg13g2_fill_1 FILLER_42_1886 ();
 sg13g2_decap_8 FILLER_42_1895 ();
 sg13g2_fill_2 FILLER_42_1902 ();
 sg13g2_fill_1 FILLER_42_1917 ();
 sg13g2_fill_2 FILLER_42_1949 ();
 sg13g2_fill_1 FILLER_42_1951 ();
 sg13g2_decap_8 FILLER_42_2009 ();
 sg13g2_decap_8 FILLER_42_2016 ();
 sg13g2_decap_4 FILLER_42_2062 ();
 sg13g2_fill_1 FILLER_42_2066 ();
 sg13g2_fill_2 FILLER_42_2079 ();
 sg13g2_fill_2 FILLER_42_2086 ();
 sg13g2_fill_1 FILLER_42_2088 ();
 sg13g2_fill_2 FILLER_42_2098 ();
 sg13g2_fill_1 FILLER_42_2100 ();
 sg13g2_fill_2 FILLER_42_2109 ();
 sg13g2_decap_4 FILLER_42_2128 ();
 sg13g2_decap_4 FILLER_42_2140 ();
 sg13g2_fill_1 FILLER_42_2194 ();
 sg13g2_decap_8 FILLER_42_2201 ();
 sg13g2_fill_2 FILLER_42_2208 ();
 sg13g2_decap_8 FILLER_42_2244 ();
 sg13g2_decap_8 FILLER_42_2251 ();
 sg13g2_decap_8 FILLER_42_2258 ();
 sg13g2_decap_8 FILLER_42_2306 ();
 sg13g2_decap_8 FILLER_42_2313 ();
 sg13g2_fill_1 FILLER_42_2346 ();
 sg13g2_decap_4 FILLER_42_2353 ();
 sg13g2_fill_2 FILLER_42_2386 ();
 sg13g2_fill_1 FILLER_42_2388 ();
 sg13g2_fill_2 FILLER_42_2415 ();
 sg13g2_decap_8 FILLER_42_2436 ();
 sg13g2_decap_8 FILLER_42_2443 ();
 sg13g2_decap_8 FILLER_42_2450 ();
 sg13g2_decap_8 FILLER_42_2457 ();
 sg13g2_decap_8 FILLER_42_2464 ();
 sg13g2_fill_1 FILLER_42_2471 ();
 sg13g2_decap_8 FILLER_42_2477 ();
 sg13g2_decap_8 FILLER_42_2484 ();
 sg13g2_decap_8 FILLER_42_2491 ();
 sg13g2_decap_8 FILLER_42_2498 ();
 sg13g2_decap_8 FILLER_42_2505 ();
 sg13g2_decap_8 FILLER_42_2512 ();
 sg13g2_decap_8 FILLER_42_2519 ();
 sg13g2_decap_8 FILLER_42_2526 ();
 sg13g2_decap_8 FILLER_42_2533 ();
 sg13g2_fill_2 FILLER_42_2540 ();
 sg13g2_fill_1 FILLER_42_2542 ();
 sg13g2_fill_2 FILLER_42_2595 ();
 sg13g2_decap_8 FILLER_42_2649 ();
 sg13g2_fill_2 FILLER_42_2656 ();
 sg13g2_decap_4 FILLER_42_2663 ();
 sg13g2_fill_2 FILLER_42_2667 ();
 sg13g2_decap_8 FILLER_42_2677 ();
 sg13g2_decap_8 FILLER_42_2684 ();
 sg13g2_decap_8 FILLER_42_2691 ();
 sg13g2_decap_8 FILLER_42_2698 ();
 sg13g2_decap_8 FILLER_42_2705 ();
 sg13g2_fill_1 FILLER_42_2712 ();
 sg13g2_fill_2 FILLER_42_2718 ();
 sg13g2_decap_8 FILLER_42_2760 ();
 sg13g2_decap_8 FILLER_42_2767 ();
 sg13g2_fill_2 FILLER_42_2774 ();
 sg13g2_decap_8 FILLER_42_2818 ();
 sg13g2_decap_4 FILLER_42_2825 ();
 sg13g2_fill_1 FILLER_42_2829 ();
 sg13g2_fill_2 FILLER_42_2834 ();
 sg13g2_fill_1 FILLER_42_2836 ();
 sg13g2_decap_8 FILLER_42_2867 ();
 sg13g2_decap_8 FILLER_42_2874 ();
 sg13g2_decap_8 FILLER_42_2881 ();
 sg13g2_decap_8 FILLER_42_2888 ();
 sg13g2_decap_4 FILLER_42_2895 ();
 sg13g2_fill_1 FILLER_42_2899 ();
 sg13g2_decap_8 FILLER_42_2910 ();
 sg13g2_decap_8 FILLER_42_2917 ();
 sg13g2_decap_4 FILLER_42_2924 ();
 sg13g2_fill_1 FILLER_42_2928 ();
 sg13g2_decap_8 FILLER_42_2955 ();
 sg13g2_decap_8 FILLER_42_2962 ();
 sg13g2_decap_8 FILLER_42_2969 ();
 sg13g2_decap_4 FILLER_42_2976 ();
 sg13g2_fill_1 FILLER_42_2980 ();
 sg13g2_fill_1 FILLER_42_2986 ();
 sg13g2_fill_2 FILLER_42_2992 ();
 sg13g2_fill_1 FILLER_42_2994 ();
 sg13g2_fill_2 FILLER_42_3000 ();
 sg13g2_fill_1 FILLER_42_3002 ();
 sg13g2_fill_2 FILLER_42_3011 ();
 sg13g2_decap_4 FILLER_42_3017 ();
 sg13g2_fill_2 FILLER_42_3021 ();
 sg13g2_decap_8 FILLER_42_3053 ();
 sg13g2_decap_8 FILLER_42_3060 ();
 sg13g2_decap_8 FILLER_42_3067 ();
 sg13g2_decap_4 FILLER_42_3074 ();
 sg13g2_decap_8 FILLER_42_3116 ();
 sg13g2_decap_8 FILLER_42_3123 ();
 sg13g2_fill_2 FILLER_42_3138 ();
 sg13g2_fill_2 FILLER_42_3161 ();
 sg13g2_decap_8 FILLER_42_3166 ();
 sg13g2_decap_4 FILLER_42_3199 ();
 sg13g2_fill_2 FILLER_42_3213 ();
 sg13g2_decap_8 FILLER_42_3246 ();
 sg13g2_decap_8 FILLER_42_3253 ();
 sg13g2_decap_8 FILLER_42_3260 ();
 sg13g2_decap_8 FILLER_42_3267 ();
 sg13g2_decap_8 FILLER_42_3274 ();
 sg13g2_decap_8 FILLER_42_3281 ();
 sg13g2_decap_8 FILLER_42_3288 ();
 sg13g2_decap_8 FILLER_42_3295 ();
 sg13g2_decap_8 FILLER_42_3302 ();
 sg13g2_decap_8 FILLER_42_3309 ();
 sg13g2_decap_8 FILLER_42_3316 ();
 sg13g2_decap_8 FILLER_42_3323 ();
 sg13g2_decap_8 FILLER_42_3330 ();
 sg13g2_decap_8 FILLER_42_3337 ();
 sg13g2_decap_8 FILLER_42_3344 ();
 sg13g2_decap_8 FILLER_42_3351 ();
 sg13g2_decap_8 FILLER_42_3358 ();
 sg13g2_decap_8 FILLER_42_3365 ();
 sg13g2_decap_8 FILLER_42_3372 ();
 sg13g2_decap_8 FILLER_42_3379 ();
 sg13g2_decap_8 FILLER_42_3386 ();
 sg13g2_decap_8 FILLER_42_3393 ();
 sg13g2_decap_8 FILLER_42_3400 ();
 sg13g2_decap_8 FILLER_42_3407 ();
 sg13g2_decap_8 FILLER_42_3414 ();
 sg13g2_decap_8 FILLER_42_3421 ();
 sg13g2_decap_8 FILLER_42_3428 ();
 sg13g2_decap_8 FILLER_42_3435 ();
 sg13g2_decap_8 FILLER_42_3442 ();
 sg13g2_decap_8 FILLER_42_3449 ();
 sg13g2_decap_8 FILLER_42_3456 ();
 sg13g2_decap_8 FILLER_42_3463 ();
 sg13g2_decap_8 FILLER_42_3470 ();
 sg13g2_decap_8 FILLER_42_3477 ();
 sg13g2_decap_8 FILLER_42_3484 ();
 sg13g2_decap_8 FILLER_42_3491 ();
 sg13g2_decap_8 FILLER_42_3498 ();
 sg13g2_decap_8 FILLER_42_3505 ();
 sg13g2_decap_8 FILLER_42_3512 ();
 sg13g2_decap_8 FILLER_42_3519 ();
 sg13g2_decap_8 FILLER_42_3526 ();
 sg13g2_decap_8 FILLER_42_3533 ();
 sg13g2_decap_8 FILLER_42_3540 ();
 sg13g2_decap_8 FILLER_42_3547 ();
 sg13g2_decap_8 FILLER_42_3554 ();
 sg13g2_decap_8 FILLER_42_3561 ();
 sg13g2_decap_8 FILLER_42_3568 ();
 sg13g2_decap_4 FILLER_42_3575 ();
 sg13g2_fill_1 FILLER_42_3579 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_4 FILLER_43_112 ();
 sg13g2_fill_2 FILLER_43_116 ();
 sg13g2_decap_8 FILLER_43_149 ();
 sg13g2_decap_8 FILLER_43_156 ();
 sg13g2_fill_1 FILLER_43_163 ();
 sg13g2_fill_2 FILLER_43_167 ();
 sg13g2_decap_4 FILLER_43_172 ();
 sg13g2_fill_2 FILLER_43_176 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_248 ();
 sg13g2_decap_8 FILLER_43_255 ();
 sg13g2_fill_1 FILLER_43_262 ();
 sg13g2_decap_4 FILLER_43_294 ();
 sg13g2_fill_2 FILLER_43_298 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_4 FILLER_43_350 ();
 sg13g2_fill_1 FILLER_43_354 ();
 sg13g2_decap_8 FILLER_43_447 ();
 sg13g2_fill_1 FILLER_43_454 ();
 sg13g2_fill_2 FILLER_43_511 ();
 sg13g2_fill_1 FILLER_43_513 ();
 sg13g2_fill_1 FILLER_43_527 ();
 sg13g2_decap_4 FILLER_43_540 ();
 sg13g2_fill_2 FILLER_43_544 ();
 sg13g2_decap_4 FILLER_43_572 ();
 sg13g2_fill_1 FILLER_43_576 ();
 sg13g2_decap_4 FILLER_43_647 ();
 sg13g2_fill_2 FILLER_43_651 ();
 sg13g2_fill_2 FILLER_43_661 ();
 sg13g2_decap_8 FILLER_43_689 ();
 sg13g2_decap_8 FILLER_43_696 ();
 sg13g2_decap_8 FILLER_43_703 ();
 sg13g2_fill_1 FILLER_43_710 ();
 sg13g2_fill_2 FILLER_43_737 ();
 sg13g2_fill_1 FILLER_43_739 ();
 sg13g2_fill_2 FILLER_43_771 ();
 sg13g2_fill_1 FILLER_43_802 ();
 sg13g2_decap_8 FILLER_43_821 ();
 sg13g2_decap_8 FILLER_43_828 ();
 sg13g2_decap_8 FILLER_43_835 ();
 sg13g2_fill_1 FILLER_43_842 ();
 sg13g2_decap_8 FILLER_43_869 ();
 sg13g2_decap_8 FILLER_43_876 ();
 sg13g2_fill_2 FILLER_43_883 ();
 sg13g2_fill_1 FILLER_43_885 ();
 sg13g2_fill_2 FILLER_43_918 ();
 sg13g2_fill_2 FILLER_43_952 ();
 sg13g2_fill_1 FILLER_43_954 ();
 sg13g2_decap_8 FILLER_43_984 ();
 sg13g2_decap_8 FILLER_43_991 ();
 sg13g2_decap_4 FILLER_43_998 ();
 sg13g2_fill_2 FILLER_43_1002 ();
 sg13g2_decap_4 FILLER_43_1035 ();
 sg13g2_decap_8 FILLER_43_1065 ();
 sg13g2_decap_8 FILLER_43_1072 ();
 sg13g2_decap_4 FILLER_43_1079 ();
 sg13g2_fill_2 FILLER_43_1103 ();
 sg13g2_fill_1 FILLER_43_1105 ();
 sg13g2_decap_4 FILLER_43_1112 ();
 sg13g2_decap_8 FILLER_43_1126 ();
 sg13g2_decap_8 FILLER_43_1141 ();
 sg13g2_decap_4 FILLER_43_1148 ();
 sg13g2_fill_2 FILLER_43_1152 ();
 sg13g2_decap_4 FILLER_43_1190 ();
 sg13g2_fill_2 FILLER_43_1199 ();
 sg13g2_decap_8 FILLER_43_1223 ();
 sg13g2_decap_8 FILLER_43_1230 ();
 sg13g2_decap_8 FILLER_43_1237 ();
 sg13g2_decap_4 FILLER_43_1244 ();
 sg13g2_fill_2 FILLER_43_1248 ();
 sg13g2_decap_8 FILLER_43_1286 ();
 sg13g2_decap_4 FILLER_43_1293 ();
 sg13g2_decap_8 FILLER_43_1331 ();
 sg13g2_decap_8 FILLER_43_1338 ();
 sg13g2_fill_2 FILLER_43_1345 ();
 sg13g2_fill_1 FILLER_43_1347 ();
 sg13g2_decap_8 FILLER_43_1406 ();
 sg13g2_decap_8 FILLER_43_1413 ();
 sg13g2_decap_8 FILLER_43_1420 ();
 sg13g2_decap_8 FILLER_43_1427 ();
 sg13g2_fill_2 FILLER_43_1434 ();
 sg13g2_fill_2 FILLER_43_1477 ();
 sg13g2_fill_2 FILLER_43_1495 ();
 sg13g2_fill_1 FILLER_43_1505 ();
 sg13g2_fill_1 FILLER_43_1510 ();
 sg13g2_fill_1 FILLER_43_1515 ();
 sg13g2_fill_1 FILLER_43_1526 ();
 sg13g2_fill_2 FILLER_43_1537 ();
 sg13g2_fill_2 FILLER_43_1544 ();
 sg13g2_fill_2 FILLER_43_1560 ();
 sg13g2_fill_1 FILLER_43_1569 ();
 sg13g2_decap_8 FILLER_43_1588 ();
 sg13g2_decap_8 FILLER_43_1595 ();
 sg13g2_decap_8 FILLER_43_1602 ();
 sg13g2_decap_8 FILLER_43_1609 ();
 sg13g2_decap_8 FILLER_43_1616 ();
 sg13g2_decap_8 FILLER_43_1623 ();
 sg13g2_decap_8 FILLER_43_1630 ();
 sg13g2_decap_8 FILLER_43_1637 ();
 sg13g2_decap_4 FILLER_43_1644 ();
 sg13g2_fill_2 FILLER_43_1648 ();
 sg13g2_fill_2 FILLER_43_1672 ();
 sg13g2_fill_1 FILLER_43_1674 ();
 sg13g2_decap_8 FILLER_43_1688 ();
 sg13g2_decap_8 FILLER_43_1695 ();
 sg13g2_decap_8 FILLER_43_1733 ();
 sg13g2_decap_8 FILLER_43_1740 ();
 sg13g2_decap_8 FILLER_43_1747 ();
 sg13g2_fill_2 FILLER_43_1754 ();
 sg13g2_decap_8 FILLER_43_1834 ();
 sg13g2_fill_1 FILLER_43_1841 ();
 sg13g2_decap_4 FILLER_43_1846 ();
 sg13g2_fill_2 FILLER_43_1850 ();
 sg13g2_decap_4 FILLER_43_1857 ();
 sg13g2_fill_2 FILLER_43_1861 ();
 sg13g2_fill_1 FILLER_43_1868 ();
 sg13g2_decap_8 FILLER_43_1886 ();
 sg13g2_decap_8 FILLER_43_1893 ();
 sg13g2_decap_8 FILLER_43_1900 ();
 sg13g2_decap_4 FILLER_43_1925 ();
 sg13g2_decap_8 FILLER_43_1950 ();
 sg13g2_fill_2 FILLER_43_1957 ();
 sg13g2_fill_1 FILLER_43_1959 ();
 sg13g2_fill_1 FILLER_43_1972 ();
 sg13g2_fill_2 FILLER_43_1985 ();
 sg13g2_fill_1 FILLER_43_1987 ();
 sg13g2_decap_4 FILLER_43_2019 ();
 sg13g2_fill_1 FILLER_43_2023 ();
 sg13g2_fill_2 FILLER_43_2044 ();
 sg13g2_decap_4 FILLER_43_2051 ();
 sg13g2_decap_8 FILLER_43_2059 ();
 sg13g2_decap_8 FILLER_43_2066 ();
 sg13g2_decap_8 FILLER_43_2073 ();
 sg13g2_decap_8 FILLER_43_2080 ();
 sg13g2_decap_8 FILLER_43_2091 ();
 sg13g2_decap_4 FILLER_43_2098 ();
 sg13g2_decap_4 FILLER_43_2149 ();
 sg13g2_fill_1 FILLER_43_2153 ();
 sg13g2_decap_8 FILLER_43_2186 ();
 sg13g2_decap_4 FILLER_43_2193 ();
 sg13g2_decap_4 FILLER_43_2203 ();
 sg13g2_fill_1 FILLER_43_2207 ();
 sg13g2_decap_8 FILLER_43_2242 ();
 sg13g2_decap_8 FILLER_43_2283 ();
 sg13g2_fill_2 FILLER_43_2290 ();
 sg13g2_decap_8 FILLER_43_2302 ();
 sg13g2_decap_8 FILLER_43_2309 ();
 sg13g2_decap_8 FILLER_43_2316 ();
 sg13g2_decap_8 FILLER_43_2323 ();
 sg13g2_decap_8 FILLER_43_2330 ();
 sg13g2_fill_2 FILLER_43_2337 ();
 sg13g2_fill_1 FILLER_43_2339 ();
 sg13g2_decap_8 FILLER_43_2366 ();
 sg13g2_fill_2 FILLER_43_2378 ();
 sg13g2_decap_8 FILLER_43_2442 ();
 sg13g2_fill_1 FILLER_43_2449 ();
 sg13g2_decap_8 FILLER_43_2506 ();
 sg13g2_decap_8 FILLER_43_2513 ();
 sg13g2_decap_8 FILLER_43_2520 ();
 sg13g2_decap_8 FILLER_43_2527 ();
 sg13g2_fill_2 FILLER_43_2534 ();
 sg13g2_fill_1 FILLER_43_2536 ();
 sg13g2_fill_2 FILLER_43_2569 ();
 sg13g2_fill_2 FILLER_43_2579 ();
 sg13g2_decap_4 FILLER_43_2596 ();
 sg13g2_decap_8 FILLER_43_2626 ();
 sg13g2_decap_8 FILLER_43_2633 ();
 sg13g2_fill_2 FILLER_43_2640 ();
 sg13g2_fill_1 FILLER_43_2642 ();
 sg13g2_decap_8 FILLER_43_2686 ();
 sg13g2_decap_4 FILLER_43_2693 ();
 sg13g2_fill_1 FILLER_43_2697 ();
 sg13g2_decap_8 FILLER_43_2749 ();
 sg13g2_decap_8 FILLER_43_2756 ();
 sg13g2_decap_8 FILLER_43_2771 ();
 sg13g2_decap_8 FILLER_43_2778 ();
 sg13g2_fill_1 FILLER_43_2785 ();
 sg13g2_decap_8 FILLER_43_2808 ();
 sg13g2_decap_8 FILLER_43_2815 ();
 sg13g2_decap_4 FILLER_43_2822 ();
 sg13g2_decap_8 FILLER_43_2860 ();
 sg13g2_decap_4 FILLER_43_2867 ();
 sg13g2_fill_1 FILLER_43_2871 ();
 sg13g2_decap_8 FILLER_43_2898 ();
 sg13g2_decap_8 FILLER_43_2905 ();
 sg13g2_decap_4 FILLER_43_2912 ();
 sg13g2_fill_2 FILLER_43_2916 ();
 sg13g2_decap_8 FILLER_43_2957 ();
 sg13g2_fill_1 FILLER_43_2964 ();
 sg13g2_decap_8 FILLER_43_2991 ();
 sg13g2_decap_8 FILLER_43_2998 ();
 sg13g2_decap_8 FILLER_43_3005 ();
 sg13g2_decap_8 FILLER_43_3012 ();
 sg13g2_decap_8 FILLER_43_3019 ();
 sg13g2_decap_4 FILLER_43_3026 ();
 sg13g2_fill_2 FILLER_43_3033 ();
 sg13g2_fill_2 FILLER_43_3043 ();
 sg13g2_decap_8 FILLER_43_3055 ();
 sg13g2_decap_8 FILLER_43_3062 ();
 sg13g2_decap_4 FILLER_43_3069 ();
 sg13g2_fill_1 FILLER_43_3073 ();
 sg13g2_decap_8 FILLER_43_3100 ();
 sg13g2_decap_8 FILLER_43_3107 ();
 sg13g2_decap_8 FILLER_43_3114 ();
 sg13g2_decap_8 FILLER_43_3121 ();
 sg13g2_decap_8 FILLER_43_3128 ();
 sg13g2_fill_1 FILLER_43_3135 ();
 sg13g2_fill_1 FILLER_43_3141 ();
 sg13g2_decap_4 FILLER_43_3146 ();
 sg13g2_fill_1 FILLER_43_3150 ();
 sg13g2_fill_2 FILLER_43_3155 ();
 sg13g2_fill_2 FILLER_43_3161 ();
 sg13g2_decap_8 FILLER_43_3193 ();
 sg13g2_decap_4 FILLER_43_3200 ();
 sg13g2_fill_1 FILLER_43_3243 ();
 sg13g2_decap_8 FILLER_43_3248 ();
 sg13g2_decap_8 FILLER_43_3255 ();
 sg13g2_decap_8 FILLER_43_3262 ();
 sg13g2_decap_8 FILLER_43_3269 ();
 sg13g2_decap_8 FILLER_43_3276 ();
 sg13g2_decap_8 FILLER_43_3283 ();
 sg13g2_decap_8 FILLER_43_3290 ();
 sg13g2_decap_8 FILLER_43_3297 ();
 sg13g2_decap_8 FILLER_43_3304 ();
 sg13g2_decap_8 FILLER_43_3311 ();
 sg13g2_decap_8 FILLER_43_3318 ();
 sg13g2_decap_8 FILLER_43_3325 ();
 sg13g2_decap_8 FILLER_43_3332 ();
 sg13g2_decap_8 FILLER_43_3339 ();
 sg13g2_decap_8 FILLER_43_3346 ();
 sg13g2_decap_8 FILLER_43_3353 ();
 sg13g2_decap_8 FILLER_43_3360 ();
 sg13g2_decap_8 FILLER_43_3367 ();
 sg13g2_decap_8 FILLER_43_3374 ();
 sg13g2_decap_8 FILLER_43_3381 ();
 sg13g2_decap_8 FILLER_43_3388 ();
 sg13g2_decap_8 FILLER_43_3395 ();
 sg13g2_decap_8 FILLER_43_3402 ();
 sg13g2_decap_8 FILLER_43_3409 ();
 sg13g2_decap_8 FILLER_43_3416 ();
 sg13g2_decap_8 FILLER_43_3423 ();
 sg13g2_decap_8 FILLER_43_3430 ();
 sg13g2_decap_8 FILLER_43_3437 ();
 sg13g2_decap_8 FILLER_43_3444 ();
 sg13g2_decap_8 FILLER_43_3451 ();
 sg13g2_decap_8 FILLER_43_3458 ();
 sg13g2_decap_8 FILLER_43_3465 ();
 sg13g2_decap_8 FILLER_43_3472 ();
 sg13g2_decap_8 FILLER_43_3479 ();
 sg13g2_decap_8 FILLER_43_3486 ();
 sg13g2_decap_8 FILLER_43_3493 ();
 sg13g2_decap_8 FILLER_43_3500 ();
 sg13g2_decap_8 FILLER_43_3507 ();
 sg13g2_decap_8 FILLER_43_3514 ();
 sg13g2_decap_8 FILLER_43_3521 ();
 sg13g2_decap_8 FILLER_43_3528 ();
 sg13g2_decap_8 FILLER_43_3535 ();
 sg13g2_decap_8 FILLER_43_3542 ();
 sg13g2_decap_8 FILLER_43_3549 ();
 sg13g2_decap_8 FILLER_43_3556 ();
 sg13g2_decap_8 FILLER_43_3563 ();
 sg13g2_decap_8 FILLER_43_3570 ();
 sg13g2_fill_2 FILLER_43_3577 ();
 sg13g2_fill_1 FILLER_43_3579 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_fill_2 FILLER_44_112 ();
 sg13g2_fill_1 FILLER_44_117 ();
 sg13g2_fill_1 FILLER_44_125 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_4 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_292 ();
 sg13g2_fill_1 FILLER_44_299 ();
 sg13g2_fill_1 FILLER_44_344 ();
 sg13g2_decap_4 FILLER_44_396 ();
 sg13g2_decap_8 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_fill_1 FILLER_44_469 ();
 sg13g2_fill_2 FILLER_44_478 ();
 sg13g2_fill_1 FILLER_44_480 ();
 sg13g2_decap_8 FILLER_44_489 ();
 sg13g2_decap_8 FILLER_44_496 ();
 sg13g2_decap_4 FILLER_44_503 ();
 sg13g2_fill_2 FILLER_44_507 ();
 sg13g2_fill_2 FILLER_44_787 ();
 sg13g2_decap_8 FILLER_44_864 ();
 sg13g2_decap_8 FILLER_44_871 ();
 sg13g2_decap_8 FILLER_44_878 ();
 sg13g2_decap_8 FILLER_44_885 ();
 sg13g2_decap_8 FILLER_44_892 ();
 sg13g2_decap_4 FILLER_44_899 ();
 sg13g2_fill_2 FILLER_44_903 ();
 sg13g2_decap_8 FILLER_44_993 ();
 sg13g2_decap_4 FILLER_44_1000 ();
 sg13g2_fill_1 FILLER_44_1004 ();
 sg13g2_fill_2 FILLER_44_1031 ();
 sg13g2_fill_1 FILLER_44_1033 ();
 sg13g2_decap_8 FILLER_44_1060 ();
 sg13g2_decap_8 FILLER_44_1067 ();
 sg13g2_decap_8 FILLER_44_1074 ();
 sg13g2_decap_4 FILLER_44_1081 ();
 sg13g2_decap_8 FILLER_44_1089 ();
 sg13g2_decap_8 FILLER_44_1096 ();
 sg13g2_fill_1 FILLER_44_1103 ();
 sg13g2_fill_1 FILLER_44_1108 ();
 sg13g2_decap_4 FILLER_44_1115 ();
 sg13g2_fill_1 FILLER_44_1119 ();
 sg13g2_fill_2 FILLER_44_1125 ();
 sg13g2_fill_1 FILLER_44_1127 ();
 sg13g2_decap_8 FILLER_44_1136 ();
 sg13g2_decap_8 FILLER_44_1143 ();
 sg13g2_decap_8 FILLER_44_1150 ();
 sg13g2_decap_8 FILLER_44_1157 ();
 sg13g2_decap_4 FILLER_44_1164 ();
 sg13g2_fill_2 FILLER_44_1168 ();
 sg13g2_decap_8 FILLER_44_1176 ();
 sg13g2_decap_8 FILLER_44_1183 ();
 sg13g2_decap_8 FILLER_44_1190 ();
 sg13g2_decap_4 FILLER_44_1197 ();
 sg13g2_fill_1 FILLER_44_1201 ();
 sg13g2_fill_2 FILLER_44_1206 ();
 sg13g2_fill_2 FILLER_44_1220 ();
 sg13g2_fill_1 FILLER_44_1222 ();
 sg13g2_decap_8 FILLER_44_1231 ();
 sg13g2_fill_2 FILLER_44_1238 ();
 sg13g2_fill_1 FILLER_44_1240 ();
 sg13g2_decap_4 FILLER_44_1293 ();
 sg13g2_fill_2 FILLER_44_1297 ();
 sg13g2_decap_8 FILLER_44_1335 ();
 sg13g2_decap_4 FILLER_44_1342 ();
 sg13g2_fill_2 FILLER_44_1346 ();
 sg13g2_decap_4 FILLER_44_1392 ();
 sg13g2_fill_1 FILLER_44_1396 ();
 sg13g2_decap_8 FILLER_44_1403 ();
 sg13g2_decap_8 FILLER_44_1410 ();
 sg13g2_decap_8 FILLER_44_1417 ();
 sg13g2_decap_8 FILLER_44_1424 ();
 sg13g2_fill_1 FILLER_44_1431 ();
 sg13g2_decap_4 FILLER_44_1444 ();
 sg13g2_fill_2 FILLER_44_1448 ();
 sg13g2_fill_2 FILLER_44_1490 ();
 sg13g2_fill_1 FILLER_44_1524 ();
 sg13g2_fill_1 FILLER_44_1533 ();
 sg13g2_fill_1 FILLER_44_1537 ();
 sg13g2_fill_2 FILLER_44_1602 ();
 sg13g2_decap_8 FILLER_44_1609 ();
 sg13g2_fill_2 FILLER_44_1616 ();
 sg13g2_decap_8 FILLER_44_1638 ();
 sg13g2_fill_1 FILLER_44_1645 ();
 sg13g2_fill_2 FILLER_44_1655 ();
 sg13g2_fill_1 FILLER_44_1676 ();
 sg13g2_decap_8 FILLER_44_1685 ();
 sg13g2_decap_8 FILLER_44_1692 ();
 sg13g2_decap_8 FILLER_44_1699 ();
 sg13g2_decap_4 FILLER_44_1706 ();
 sg13g2_decap_8 FILLER_44_1736 ();
 sg13g2_decap_8 FILLER_44_1743 ();
 sg13g2_decap_4 FILLER_44_1750 ();
 sg13g2_fill_1 FILLER_44_1754 ();
 sg13g2_fill_1 FILLER_44_1781 ();
 sg13g2_decap_8 FILLER_44_1814 ();
 sg13g2_decap_8 FILLER_44_1821 ();
 sg13g2_decap_8 FILLER_44_1828 ();
 sg13g2_fill_1 FILLER_44_1835 ();
 sg13g2_fill_2 FILLER_44_1862 ();
 sg13g2_fill_1 FILLER_44_1864 ();
 sg13g2_fill_2 FILLER_44_1891 ();
 sg13g2_fill_1 FILLER_44_1893 ();
 sg13g2_decap_8 FILLER_44_1898 ();
 sg13g2_decap_8 FILLER_44_1913 ();
 sg13g2_decap_8 FILLER_44_1920 ();
 sg13g2_decap_4 FILLER_44_1927 ();
 sg13g2_fill_2 FILLER_44_1931 ();
 sg13g2_decap_8 FILLER_44_1937 ();
 sg13g2_decap_8 FILLER_44_1944 ();
 sg13g2_decap_4 FILLER_44_1951 ();
 sg13g2_fill_1 FILLER_44_1955 ();
 sg13g2_decap_8 FILLER_44_1964 ();
 sg13g2_fill_2 FILLER_44_1971 ();
 sg13g2_fill_1 FILLER_44_1973 ();
 sg13g2_decap_8 FILLER_44_1985 ();
 sg13g2_decap_8 FILLER_44_1992 ();
 sg13g2_decap_8 FILLER_44_1999 ();
 sg13g2_decap_8 FILLER_44_2006 ();
 sg13g2_decap_8 FILLER_44_2013 ();
 sg13g2_decap_4 FILLER_44_2020 ();
 sg13g2_fill_1 FILLER_44_2024 ();
 sg13g2_decap_4 FILLER_44_2030 ();
 sg13g2_decap_4 FILLER_44_2038 ();
 sg13g2_fill_2 FILLER_44_2042 ();
 sg13g2_decap_8 FILLER_44_2070 ();
 sg13g2_decap_8 FILLER_44_2077 ();
 sg13g2_fill_2 FILLER_44_2084 ();
 sg13g2_decap_8 FILLER_44_2138 ();
 sg13g2_decap_8 FILLER_44_2145 ();
 sg13g2_fill_1 FILLER_44_2152 ();
 sg13g2_fill_2 FILLER_44_2163 ();
 sg13g2_decap_8 FILLER_44_2197 ();
 sg13g2_decap_8 FILLER_44_2204 ();
 sg13g2_fill_1 FILLER_44_2211 ();
 sg13g2_decap_8 FILLER_44_2264 ();
 sg13g2_decap_8 FILLER_44_2271 ();
 sg13g2_fill_2 FILLER_44_2278 ();
 sg13g2_fill_2 FILLER_44_2319 ();
 sg13g2_fill_1 FILLER_44_2321 ();
 sg13g2_decap_8 FILLER_44_2354 ();
 sg13g2_decap_8 FILLER_44_2361 ();
 sg13g2_decap_4 FILLER_44_2368 ();
 sg13g2_fill_1 FILLER_44_2372 ();
 sg13g2_decap_8 FILLER_44_2381 ();
 sg13g2_decap_8 FILLER_44_2388 ();
 sg13g2_fill_2 FILLER_44_2395 ();
 sg13g2_fill_1 FILLER_44_2397 ();
 sg13g2_fill_2 FILLER_44_2484 ();
 sg13g2_decap_4 FILLER_44_2538 ();
 sg13g2_fill_2 FILLER_44_2542 ();
 sg13g2_decap_8 FILLER_44_2604 ();
 sg13g2_decap_8 FILLER_44_2611 ();
 sg13g2_decap_8 FILLER_44_2618 ();
 sg13g2_decap_8 FILLER_44_2625 ();
 sg13g2_fill_2 FILLER_44_2632 ();
 sg13g2_fill_1 FILLER_44_2634 ();
 sg13g2_decap_8 FILLER_44_2713 ();
 sg13g2_fill_2 FILLER_44_2720 ();
 sg13g2_decap_8 FILLER_44_2748 ();
 sg13g2_decap_8 FILLER_44_2781 ();
 sg13g2_fill_2 FILLER_44_2796 ();
 sg13g2_decap_8 FILLER_44_2802 ();
 sg13g2_decap_8 FILLER_44_2809 ();
 sg13g2_decap_8 FILLER_44_2816 ();
 sg13g2_decap_4 FILLER_44_2823 ();
 sg13g2_decap_8 FILLER_44_2853 ();
 sg13g2_decap_4 FILLER_44_2860 ();
 sg13g2_decap_8 FILLER_44_2890 ();
 sg13g2_decap_8 FILLER_44_2897 ();
 sg13g2_decap_8 FILLER_44_2904 ();
 sg13g2_fill_2 FILLER_44_2942 ();
 sg13g2_decap_4 FILLER_44_2978 ();
 sg13g2_fill_2 FILLER_44_2987 ();
 sg13g2_decap_8 FILLER_44_2997 ();
 sg13g2_decap_8 FILLER_44_3004 ();
 sg13g2_decap_4 FILLER_44_3011 ();
 sg13g2_fill_1 FILLER_44_3015 ();
 sg13g2_fill_2 FILLER_44_3072 ();
 sg13g2_fill_1 FILLER_44_3074 ();
 sg13g2_fill_2 FILLER_44_3083 ();
 sg13g2_decap_4 FILLER_44_3097 ();
 sg13g2_fill_2 FILLER_44_3101 ();
 sg13g2_fill_1 FILLER_44_3107 ();
 sg13g2_decap_8 FILLER_44_3134 ();
 sg13g2_decap_4 FILLER_44_3141 ();
 sg13g2_fill_2 FILLER_44_3145 ();
 sg13g2_decap_8 FILLER_44_3186 ();
 sg13g2_decap_8 FILLER_44_3193 ();
 sg13g2_decap_8 FILLER_44_3260 ();
 sg13g2_decap_8 FILLER_44_3267 ();
 sg13g2_decap_8 FILLER_44_3274 ();
 sg13g2_decap_8 FILLER_44_3281 ();
 sg13g2_decap_8 FILLER_44_3288 ();
 sg13g2_decap_8 FILLER_44_3295 ();
 sg13g2_decap_8 FILLER_44_3302 ();
 sg13g2_decap_8 FILLER_44_3309 ();
 sg13g2_decap_8 FILLER_44_3316 ();
 sg13g2_decap_8 FILLER_44_3323 ();
 sg13g2_decap_8 FILLER_44_3330 ();
 sg13g2_decap_8 FILLER_44_3337 ();
 sg13g2_decap_8 FILLER_44_3344 ();
 sg13g2_decap_8 FILLER_44_3351 ();
 sg13g2_decap_8 FILLER_44_3358 ();
 sg13g2_decap_8 FILLER_44_3365 ();
 sg13g2_decap_8 FILLER_44_3372 ();
 sg13g2_decap_8 FILLER_44_3379 ();
 sg13g2_decap_8 FILLER_44_3386 ();
 sg13g2_decap_8 FILLER_44_3393 ();
 sg13g2_decap_8 FILLER_44_3400 ();
 sg13g2_decap_8 FILLER_44_3407 ();
 sg13g2_decap_8 FILLER_44_3414 ();
 sg13g2_decap_8 FILLER_44_3421 ();
 sg13g2_decap_8 FILLER_44_3428 ();
 sg13g2_decap_8 FILLER_44_3435 ();
 sg13g2_decap_8 FILLER_44_3442 ();
 sg13g2_decap_8 FILLER_44_3449 ();
 sg13g2_decap_8 FILLER_44_3456 ();
 sg13g2_decap_8 FILLER_44_3463 ();
 sg13g2_decap_8 FILLER_44_3470 ();
 sg13g2_decap_8 FILLER_44_3477 ();
 sg13g2_decap_8 FILLER_44_3484 ();
 sg13g2_decap_8 FILLER_44_3491 ();
 sg13g2_decap_8 FILLER_44_3498 ();
 sg13g2_decap_8 FILLER_44_3505 ();
 sg13g2_decap_8 FILLER_44_3512 ();
 sg13g2_decap_8 FILLER_44_3519 ();
 sg13g2_decap_8 FILLER_44_3526 ();
 sg13g2_decap_8 FILLER_44_3533 ();
 sg13g2_decap_8 FILLER_44_3540 ();
 sg13g2_decap_8 FILLER_44_3547 ();
 sg13g2_decap_8 FILLER_44_3554 ();
 sg13g2_decap_8 FILLER_44_3561 ();
 sg13g2_decap_8 FILLER_44_3568 ();
 sg13g2_decap_4 FILLER_44_3575 ();
 sg13g2_fill_1 FILLER_44_3579 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_fill_1 FILLER_45_105 ();
 sg13g2_decap_4 FILLER_45_135 ();
 sg13g2_fill_1 FILLER_45_139 ();
 sg13g2_decap_4 FILLER_45_147 ();
 sg13g2_fill_1 FILLER_45_151 ();
 sg13g2_fill_1 FILLER_45_193 ();
 sg13g2_fill_1 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_304 ();
 sg13g2_decap_4 FILLER_45_331 ();
 sg13g2_decap_8 FILLER_45_387 ();
 sg13g2_decap_8 FILLER_45_394 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_2 FILLER_45_468 ();
 sg13g2_decap_8 FILLER_45_496 ();
 sg13g2_decap_4 FILLER_45_503 ();
 sg13g2_decap_4 FILLER_45_538 ();
 sg13g2_fill_2 FILLER_45_542 ();
 sg13g2_fill_2 FILLER_45_586 ();
 sg13g2_fill_1 FILLER_45_588 ();
 sg13g2_fill_2 FILLER_45_593 ();
 sg13g2_fill_1 FILLER_45_599 ();
 sg13g2_decap_8 FILLER_45_608 ();
 sg13g2_fill_2 FILLER_45_632 ();
 sg13g2_decap_8 FILLER_45_639 ();
 sg13g2_fill_2 FILLER_45_646 ();
 sg13g2_decap_8 FILLER_45_686 ();
 sg13g2_fill_2 FILLER_45_693 ();
 sg13g2_fill_1 FILLER_45_695 ();
 sg13g2_decap_8 FILLER_45_731 ();
 sg13g2_decap_8 FILLER_45_738 ();
 sg13g2_fill_2 FILLER_45_745 ();
 sg13g2_decap_8 FILLER_45_774 ();
 sg13g2_fill_2 FILLER_45_807 ();
 sg13g2_fill_2 FILLER_45_814 ();
 sg13g2_fill_1 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_825 ();
 sg13g2_decap_4 FILLER_45_832 ();
 sg13g2_fill_1 FILLER_45_836 ();
 sg13g2_decap_8 FILLER_45_871 ();
 sg13g2_decap_8 FILLER_45_878 ();
 sg13g2_decap_8 FILLER_45_885 ();
 sg13g2_decap_8 FILLER_45_892 ();
 sg13g2_decap_8 FILLER_45_899 ();
 sg13g2_decap_8 FILLER_45_906 ();
 sg13g2_decap_4 FILLER_45_913 ();
 sg13g2_fill_2 FILLER_45_917 ();
 sg13g2_fill_2 FILLER_45_945 ();
 sg13g2_fill_2 FILLER_45_957 ();
 sg13g2_fill_1 FILLER_45_962 ();
 sg13g2_decap_8 FILLER_45_989 ();
 sg13g2_fill_2 FILLER_45_996 ();
 sg13g2_decap_8 FILLER_45_1006 ();
 sg13g2_decap_4 FILLER_45_1013 ();
 sg13g2_fill_1 FILLER_45_1017 ();
 sg13g2_decap_8 FILLER_45_1021 ();
 sg13g2_decap_8 FILLER_45_1028 ();
 sg13g2_decap_8 FILLER_45_1035 ();
 sg13g2_decap_8 FILLER_45_1042 ();
 sg13g2_decap_8 FILLER_45_1049 ();
 sg13g2_fill_2 FILLER_45_1056 ();
 sg13g2_fill_1 FILLER_45_1084 ();
 sg13g2_fill_2 FILLER_45_1090 ();
 sg13g2_decap_4 FILLER_45_1098 ();
 sg13g2_decap_8 FILLER_45_1136 ();
 sg13g2_decap_8 FILLER_45_1143 ();
 sg13g2_fill_1 FILLER_45_1150 ();
 sg13g2_decap_8 FILLER_45_1177 ();
 sg13g2_decap_8 FILLER_45_1184 ();
 sg13g2_decap_8 FILLER_45_1191 ();
 sg13g2_decap_8 FILLER_45_1198 ();
 sg13g2_decap_8 FILLER_45_1205 ();
 sg13g2_decap_8 FILLER_45_1237 ();
 sg13g2_decap_4 FILLER_45_1244 ();
 sg13g2_fill_1 FILLER_45_1248 ();
 sg13g2_fill_2 FILLER_45_1291 ();
 sg13g2_decap_8 FILLER_45_1383 ();
 sg13g2_decap_8 FILLER_45_1390 ();
 sg13g2_fill_2 FILLER_45_1397 ();
 sg13g2_fill_1 FILLER_45_1399 ();
 sg13g2_decap_8 FILLER_45_1426 ();
 sg13g2_fill_2 FILLER_45_1433 ();
 sg13g2_decap_8 FILLER_45_1461 ();
 sg13g2_fill_2 FILLER_45_1488 ();
 sg13g2_fill_1 FILLER_45_1542 ();
 sg13g2_fill_1 FILLER_45_1573 ();
 sg13g2_fill_2 FILLER_45_1617 ();
 sg13g2_fill_1 FILLER_45_1619 ();
 sg13g2_fill_2 FILLER_45_1624 ();
 sg13g2_fill_2 FILLER_45_1638 ();
 sg13g2_fill_1 FILLER_45_1655 ();
 sg13g2_fill_2 FILLER_45_1668 ();
 sg13g2_decap_8 FILLER_45_1676 ();
 sg13g2_decap_8 FILLER_45_1683 ();
 sg13g2_decap_8 FILLER_45_1690 ();
 sg13g2_decap_8 FILLER_45_1697 ();
 sg13g2_decap_8 FILLER_45_1704 ();
 sg13g2_decap_8 FILLER_45_1743 ();
 sg13g2_decap_8 FILLER_45_1750 ();
 sg13g2_decap_8 FILLER_45_1757 ();
 sg13g2_decap_4 FILLER_45_1764 ();
 sg13g2_fill_2 FILLER_45_1768 ();
 sg13g2_decap_8 FILLER_45_1802 ();
 sg13g2_decap_8 FILLER_45_1809 ();
 sg13g2_decap_8 FILLER_45_1816 ();
 sg13g2_decap_8 FILLER_45_1823 ();
 sg13g2_decap_8 FILLER_45_1830 ();
 sg13g2_decap_8 FILLER_45_1837 ();
 sg13g2_fill_1 FILLER_45_1844 ();
 sg13g2_fill_2 FILLER_45_1849 ();
 sg13g2_decap_8 FILLER_45_1902 ();
 sg13g2_decap_8 FILLER_45_1909 ();
 sg13g2_decap_8 FILLER_45_1916 ();
 sg13g2_decap_4 FILLER_45_1923 ();
 sg13g2_fill_2 FILLER_45_1927 ();
 sg13g2_decap_4 FILLER_45_1947 ();
 sg13g2_decap_8 FILLER_45_1994 ();
 sg13g2_decap_8 FILLER_45_2001 ();
 sg13g2_decap_4 FILLER_45_2008 ();
 sg13g2_fill_1 FILLER_45_2012 ();
 sg13g2_fill_2 FILLER_45_2025 ();
 sg13g2_fill_2 FILLER_45_2032 ();
 sg13g2_decap_8 FILLER_45_2138 ();
 sg13g2_decap_4 FILLER_45_2145 ();
 sg13g2_fill_2 FILLER_45_2163 ();
 sg13g2_fill_2 FILLER_45_2173 ();
 sg13g2_decap_8 FILLER_45_2201 ();
 sg13g2_decap_8 FILLER_45_2208 ();
 sg13g2_decap_8 FILLER_45_2215 ();
 sg13g2_fill_2 FILLER_45_2222 ();
 sg13g2_fill_1 FILLER_45_2224 ();
 sg13g2_fill_2 FILLER_45_2277 ();
 sg13g2_fill_1 FILLER_45_2279 ();
 sg13g2_fill_2 FILLER_45_2306 ();
 sg13g2_fill_1 FILLER_45_2308 ();
 sg13g2_fill_1 FILLER_45_2381 ();
 sg13g2_decap_8 FILLER_45_2390 ();
 sg13g2_fill_2 FILLER_45_2397 ();
 sg13g2_fill_1 FILLER_45_2399 ();
 sg13g2_decap_8 FILLER_45_2432 ();
 sg13g2_decap_8 FILLER_45_2439 ();
 sg13g2_decap_8 FILLER_45_2446 ();
 sg13g2_fill_1 FILLER_45_2485 ();
 sg13g2_decap_8 FILLER_45_2530 ();
 sg13g2_decap_8 FILLER_45_2537 ();
 sg13g2_decap_4 FILLER_45_2544 ();
 sg13g2_decap_8 FILLER_45_2594 ();
 sg13g2_decap_8 FILLER_45_2601 ();
 sg13g2_decap_4 FILLER_45_2608 ();
 sg13g2_fill_2 FILLER_45_2612 ();
 sg13g2_decap_4 FILLER_45_2623 ();
 sg13g2_fill_2 FILLER_45_2636 ();
 sg13g2_fill_1 FILLER_45_2638 ();
 sg13g2_decap_8 FILLER_45_2723 ();
 sg13g2_fill_2 FILLER_45_2730 ();
 sg13g2_fill_1 FILLER_45_2732 ();
 sg13g2_decap_8 FILLER_45_2737 ();
 sg13g2_decap_4 FILLER_45_2744 ();
 sg13g2_fill_1 FILLER_45_2748 ();
 sg13g2_fill_2 FILLER_45_2780 ();
 sg13g2_decap_8 FILLER_45_2812 ();
 sg13g2_fill_2 FILLER_45_2819 ();
 sg13g2_fill_1 FILLER_45_2821 ();
 sg13g2_decap_8 FILLER_45_2856 ();
 sg13g2_fill_1 FILLER_45_2863 ();
 sg13g2_fill_1 FILLER_45_2890 ();
 sg13g2_fill_1 FILLER_45_2917 ();
 sg13g2_fill_2 FILLER_45_2970 ();
 sg13g2_fill_1 FILLER_45_2972 ();
 sg13g2_decap_8 FILLER_45_3007 ();
 sg13g2_decap_8 FILLER_45_3014 ();
 sg13g2_fill_2 FILLER_45_3021 ();
 sg13g2_fill_1 FILLER_45_3023 ();
 sg13g2_fill_1 FILLER_45_3134 ();
 sg13g2_decap_4 FILLER_45_3196 ();
 sg13g2_decap_8 FILLER_45_3247 ();
 sg13g2_decap_8 FILLER_45_3254 ();
 sg13g2_decap_8 FILLER_45_3261 ();
 sg13g2_decap_8 FILLER_45_3268 ();
 sg13g2_decap_8 FILLER_45_3275 ();
 sg13g2_decap_8 FILLER_45_3282 ();
 sg13g2_decap_8 FILLER_45_3289 ();
 sg13g2_decap_8 FILLER_45_3296 ();
 sg13g2_decap_8 FILLER_45_3303 ();
 sg13g2_decap_8 FILLER_45_3310 ();
 sg13g2_decap_8 FILLER_45_3317 ();
 sg13g2_decap_8 FILLER_45_3324 ();
 sg13g2_decap_8 FILLER_45_3331 ();
 sg13g2_decap_8 FILLER_45_3338 ();
 sg13g2_decap_8 FILLER_45_3345 ();
 sg13g2_decap_8 FILLER_45_3352 ();
 sg13g2_decap_8 FILLER_45_3359 ();
 sg13g2_decap_8 FILLER_45_3366 ();
 sg13g2_decap_8 FILLER_45_3373 ();
 sg13g2_decap_8 FILLER_45_3380 ();
 sg13g2_decap_8 FILLER_45_3387 ();
 sg13g2_decap_8 FILLER_45_3394 ();
 sg13g2_decap_8 FILLER_45_3401 ();
 sg13g2_decap_8 FILLER_45_3408 ();
 sg13g2_decap_8 FILLER_45_3415 ();
 sg13g2_decap_8 FILLER_45_3422 ();
 sg13g2_decap_8 FILLER_45_3429 ();
 sg13g2_decap_8 FILLER_45_3436 ();
 sg13g2_decap_8 FILLER_45_3443 ();
 sg13g2_decap_8 FILLER_45_3450 ();
 sg13g2_decap_8 FILLER_45_3457 ();
 sg13g2_decap_8 FILLER_45_3464 ();
 sg13g2_decap_8 FILLER_45_3471 ();
 sg13g2_decap_8 FILLER_45_3478 ();
 sg13g2_decap_8 FILLER_45_3485 ();
 sg13g2_decap_8 FILLER_45_3492 ();
 sg13g2_decap_8 FILLER_45_3499 ();
 sg13g2_decap_8 FILLER_45_3506 ();
 sg13g2_decap_8 FILLER_45_3513 ();
 sg13g2_decap_8 FILLER_45_3520 ();
 sg13g2_decap_8 FILLER_45_3527 ();
 sg13g2_decap_8 FILLER_45_3534 ();
 sg13g2_decap_8 FILLER_45_3541 ();
 sg13g2_decap_8 FILLER_45_3548 ();
 sg13g2_decap_8 FILLER_45_3555 ();
 sg13g2_decap_8 FILLER_45_3562 ();
 sg13g2_decap_8 FILLER_45_3569 ();
 sg13g2_decap_4 FILLER_45_3576 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_136 ();
 sg13g2_decap_8 FILLER_46_143 ();
 sg13g2_decap_8 FILLER_46_183 ();
 sg13g2_decap_8 FILLER_46_190 ();
 sg13g2_decap_4 FILLER_46_197 ();
 sg13g2_fill_1 FILLER_46_201 ();
 sg13g2_decap_4 FILLER_46_235 ();
 sg13g2_fill_1 FILLER_46_242 ();
 sg13g2_decap_4 FILLER_46_248 ();
 sg13g2_fill_2 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_258 ();
 sg13g2_fill_2 FILLER_46_265 ();
 sg13g2_decap_8 FILLER_46_272 ();
 sg13g2_fill_1 FILLER_46_279 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_decap_8 FILLER_46_313 ();
 sg13g2_fill_1 FILLER_46_320 ();
 sg13g2_fill_1 FILLER_46_336 ();
 sg13g2_decap_4 FILLER_46_347 ();
 sg13g2_fill_2 FILLER_46_351 ();
 sg13g2_decap_8 FILLER_46_379 ();
 sg13g2_decap_8 FILLER_46_386 ();
 sg13g2_fill_2 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_fill_1 FILLER_46_438 ();
 sg13g2_fill_2 FILLER_46_462 ();
 sg13g2_fill_1 FILLER_46_464 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_4 FILLER_46_511 ();
 sg13g2_fill_1 FILLER_46_515 ();
 sg13g2_decap_8 FILLER_46_529 ();
 sg13g2_decap_8 FILLER_46_536 ();
 sg13g2_decap_8 FILLER_46_543 ();
 sg13g2_fill_2 FILLER_46_550 ();
 sg13g2_decap_8 FILLER_46_604 ();
 sg13g2_fill_1 FILLER_46_611 ();
 sg13g2_decap_4 FILLER_46_619 ();
 sg13g2_decap_8 FILLER_46_636 ();
 sg13g2_fill_2 FILLER_46_643 ();
 sg13g2_fill_2 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_689 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_fill_2 FILLER_46_721 ();
 sg13g2_fill_1 FILLER_46_731 ();
 sg13g2_fill_2 FILLER_46_740 ();
 sg13g2_fill_1 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_769 ();
 sg13g2_decap_8 FILLER_46_776 ();
 sg13g2_fill_2 FILLER_46_783 ();
 sg13g2_fill_1 FILLER_46_785 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_fill_2 FILLER_46_804 ();
 sg13g2_fill_1 FILLER_46_806 ();
 sg13g2_fill_1 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_46_831 ();
 sg13g2_decap_4 FILLER_46_838 ();
 sg13g2_decap_8 FILLER_46_881 ();
 sg13g2_decap_8 FILLER_46_888 ();
 sg13g2_decap_8 FILLER_46_895 ();
 sg13g2_decap_4 FILLER_46_902 ();
 sg13g2_fill_1 FILLER_46_906 ();
 sg13g2_decap_8 FILLER_46_933 ();
 sg13g2_decap_8 FILLER_46_940 ();
 sg13g2_decap_8 FILLER_46_947 ();
 sg13g2_decap_8 FILLER_46_957 ();
 sg13g2_decap_4 FILLER_46_964 ();
 sg13g2_decap_8 FILLER_46_989 ();
 sg13g2_decap_8 FILLER_46_996 ();
 sg13g2_decap_8 FILLER_46_1003 ();
 sg13g2_decap_4 FILLER_46_1010 ();
 sg13g2_decap_8 FILLER_46_1019 ();
 sg13g2_decap_8 FILLER_46_1026 ();
 sg13g2_decap_4 FILLER_46_1059 ();
 sg13g2_fill_1 FILLER_46_1063 ();
 sg13g2_fill_2 FILLER_46_1108 ();
 sg13g2_decap_8 FILLER_46_1144 ();
 sg13g2_decap_8 FILLER_46_1189 ();
 sg13g2_decap_4 FILLER_46_1196 ();
 sg13g2_fill_1 FILLER_46_1200 ();
 sg13g2_decap_8 FILLER_46_1251 ();
 sg13g2_decap_8 FILLER_46_1258 ();
 sg13g2_fill_2 FILLER_46_1265 ();
 sg13g2_decap_8 FILLER_46_1275 ();
 sg13g2_decap_8 FILLER_46_1282 ();
 sg13g2_decap_4 FILLER_46_1289 ();
 sg13g2_decap_4 FILLER_46_1333 ();
 sg13g2_fill_1 FILLER_46_1337 ();
 sg13g2_decap_8 FILLER_46_1376 ();
 sg13g2_decap_8 FILLER_46_1383 ();
 sg13g2_decap_8 FILLER_46_1390 ();
 sg13g2_decap_4 FILLER_46_1397 ();
 sg13g2_decap_8 FILLER_46_1443 ();
 sg13g2_decap_4 FILLER_46_1450 ();
 sg13g2_decap_8 FILLER_46_1459 ();
 sg13g2_decap_8 FILLER_46_1466 ();
 sg13g2_fill_2 FILLER_46_1473 ();
 sg13g2_fill_1 FILLER_46_1493 ();
 sg13g2_fill_2 FILLER_46_1543 ();
 sg13g2_fill_1 FILLER_46_1559 ();
 sg13g2_fill_1 FILLER_46_1578 ();
 sg13g2_fill_2 FILLER_46_1585 ();
 sg13g2_fill_1 FILLER_46_1618 ();
 sg13g2_fill_2 FILLER_46_1639 ();
 sg13g2_fill_1 FILLER_46_1667 ();
 sg13g2_decap_8 FILLER_46_1676 ();
 sg13g2_decap_8 FILLER_46_1683 ();
 sg13g2_decap_8 FILLER_46_1690 ();
 sg13g2_decap_4 FILLER_46_1697 ();
 sg13g2_fill_2 FILLER_46_1701 ();
 sg13g2_decap_8 FILLER_46_1744 ();
 sg13g2_decap_8 FILLER_46_1751 ();
 sg13g2_decap_8 FILLER_46_1758 ();
 sg13g2_fill_1 FILLER_46_1765 ();
 sg13g2_decap_8 FILLER_46_1818 ();
 sg13g2_fill_2 FILLER_46_1825 ();
 sg13g2_fill_2 FILLER_46_1835 ();
 sg13g2_fill_1 FILLER_46_1837 ();
 sg13g2_decap_8 FILLER_46_2001 ();
 sg13g2_decap_8 FILLER_46_2008 ();
 sg13g2_fill_2 FILLER_46_2015 ();
 sg13g2_fill_1 FILLER_46_2017 ();
 sg13g2_decap_8 FILLER_46_2076 ();
 sg13g2_fill_2 FILLER_46_2083 ();
 sg13g2_fill_1 FILLER_46_2085 ();
 sg13g2_fill_1 FILLER_46_2092 ();
 sg13g2_decap_8 FILLER_46_2119 ();
 sg13g2_decap_8 FILLER_46_2126 ();
 sg13g2_decap_8 FILLER_46_2133 ();
 sg13g2_fill_1 FILLER_46_2140 ();
 sg13g2_fill_1 FILLER_46_2154 ();
 sg13g2_fill_2 FILLER_46_2209 ();
 sg13g2_decap_8 FILLER_46_2237 ();
 sg13g2_fill_1 FILLER_46_2244 ();
 sg13g2_decap_8 FILLER_46_2266 ();
 sg13g2_decap_4 FILLER_46_2273 ();
 sg13g2_fill_1 FILLER_46_2277 ();
 sg13g2_fill_2 FILLER_46_2292 ();
 sg13g2_fill_1 FILLER_46_2294 ();
 sg13g2_decap_8 FILLER_46_2313 ();
 sg13g2_decap_8 FILLER_46_2320 ();
 sg13g2_decap_8 FILLER_46_2327 ();
 sg13g2_fill_2 FILLER_46_2334 ();
 sg13g2_fill_1 FILLER_46_2336 ();
 sg13g2_fill_2 FILLER_46_2389 ();
 sg13g2_decap_8 FILLER_46_2396 ();
 sg13g2_fill_1 FILLER_46_2403 ();
 sg13g2_decap_8 FILLER_46_2434 ();
 sg13g2_decap_8 FILLER_46_2441 ();
 sg13g2_decap_4 FILLER_46_2448 ();
 sg13g2_fill_1 FILLER_46_2452 ();
 sg13g2_fill_2 FILLER_46_2509 ();
 sg13g2_decap_8 FILLER_46_2542 ();
 sg13g2_decap_8 FILLER_46_2549 ();
 sg13g2_decap_8 FILLER_46_2587 ();
 sg13g2_decap_8 FILLER_46_2594 ();
 sg13g2_decap_8 FILLER_46_2601 ();
 sg13g2_decap_8 FILLER_46_2608 ();
 sg13g2_fill_1 FILLER_46_2615 ();
 sg13g2_decap_8 FILLER_46_2621 ();
 sg13g2_decap_8 FILLER_46_2628 ();
 sg13g2_fill_2 FILLER_46_2635 ();
 sg13g2_fill_2 FILLER_46_2686 ();
 sg13g2_decap_8 FILLER_46_2714 ();
 sg13g2_decap_8 FILLER_46_2721 ();
 sg13g2_decap_8 FILLER_46_2728 ();
 sg13g2_decap_8 FILLER_46_2735 ();
 sg13g2_decap_8 FILLER_46_2742 ();
 sg13g2_fill_1 FILLER_46_2749 ();
 sg13g2_decap_8 FILLER_46_2802 ();
 sg13g2_fill_2 FILLER_46_2809 ();
 sg13g2_fill_1 FILLER_46_2811 ();
 sg13g2_decap_8 FILLER_46_2852 ();
 sg13g2_decap_8 FILLER_46_2859 ();
 sg13g2_decap_8 FILLER_46_2866 ();
 sg13g2_decap_8 FILLER_46_2873 ();
 sg13g2_fill_1 FILLER_46_2880 ();
 sg13g2_decap_8 FILLER_46_2907 ();
 sg13g2_decap_8 FILLER_46_2914 ();
 sg13g2_decap_4 FILLER_46_2976 ();
 sg13g2_fill_2 FILLER_46_2980 ();
 sg13g2_decap_8 FILLER_46_3013 ();
 sg13g2_decap_8 FILLER_46_3020 ();
 sg13g2_fill_2 FILLER_46_3027 ();
 sg13g2_fill_2 FILLER_46_3075 ();
 sg13g2_fill_2 FILLER_46_3081 ();
 sg13g2_decap_8 FILLER_46_3131 ();
 sg13g2_decap_8 FILLER_46_3138 ();
 sg13g2_fill_1 FILLER_46_3145 ();
 sg13g2_fill_1 FILLER_46_3150 ();
 sg13g2_decap_8 FILLER_46_3194 ();
 sg13g2_decap_8 FILLER_46_3201 ();
 sg13g2_fill_2 FILLER_46_3208 ();
 sg13g2_decap_8 FILLER_46_3240 ();
 sg13g2_decap_8 FILLER_46_3247 ();
 sg13g2_decap_8 FILLER_46_3254 ();
 sg13g2_decap_8 FILLER_46_3261 ();
 sg13g2_decap_8 FILLER_46_3268 ();
 sg13g2_decap_8 FILLER_46_3275 ();
 sg13g2_decap_8 FILLER_46_3282 ();
 sg13g2_decap_8 FILLER_46_3289 ();
 sg13g2_decap_8 FILLER_46_3296 ();
 sg13g2_decap_8 FILLER_46_3303 ();
 sg13g2_decap_8 FILLER_46_3310 ();
 sg13g2_decap_8 FILLER_46_3317 ();
 sg13g2_decap_8 FILLER_46_3324 ();
 sg13g2_decap_8 FILLER_46_3331 ();
 sg13g2_decap_8 FILLER_46_3338 ();
 sg13g2_decap_8 FILLER_46_3345 ();
 sg13g2_decap_8 FILLER_46_3352 ();
 sg13g2_decap_8 FILLER_46_3359 ();
 sg13g2_decap_8 FILLER_46_3366 ();
 sg13g2_decap_8 FILLER_46_3373 ();
 sg13g2_decap_8 FILLER_46_3380 ();
 sg13g2_decap_8 FILLER_46_3387 ();
 sg13g2_decap_8 FILLER_46_3394 ();
 sg13g2_decap_8 FILLER_46_3401 ();
 sg13g2_decap_8 FILLER_46_3408 ();
 sg13g2_decap_8 FILLER_46_3415 ();
 sg13g2_decap_8 FILLER_46_3422 ();
 sg13g2_decap_8 FILLER_46_3429 ();
 sg13g2_decap_8 FILLER_46_3436 ();
 sg13g2_decap_8 FILLER_46_3443 ();
 sg13g2_decap_8 FILLER_46_3450 ();
 sg13g2_decap_8 FILLER_46_3457 ();
 sg13g2_decap_8 FILLER_46_3464 ();
 sg13g2_decap_8 FILLER_46_3471 ();
 sg13g2_decap_8 FILLER_46_3478 ();
 sg13g2_decap_8 FILLER_46_3485 ();
 sg13g2_decap_8 FILLER_46_3492 ();
 sg13g2_decap_8 FILLER_46_3499 ();
 sg13g2_decap_8 FILLER_46_3506 ();
 sg13g2_decap_8 FILLER_46_3513 ();
 sg13g2_decap_8 FILLER_46_3520 ();
 sg13g2_decap_8 FILLER_46_3527 ();
 sg13g2_decap_8 FILLER_46_3534 ();
 sg13g2_decap_8 FILLER_46_3541 ();
 sg13g2_decap_8 FILLER_46_3548 ();
 sg13g2_decap_8 FILLER_46_3555 ();
 sg13g2_decap_8 FILLER_46_3562 ();
 sg13g2_decap_8 FILLER_46_3569 ();
 sg13g2_decap_4 FILLER_46_3576 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_fill_1 FILLER_47_91 ();
 sg13g2_decap_4 FILLER_47_133 ();
 sg13g2_fill_1 FILLER_47_137 ();
 sg13g2_decap_8 FILLER_47_142 ();
 sg13g2_decap_8 FILLER_47_149 ();
 sg13g2_decap_8 FILLER_47_156 ();
 sg13g2_decap_8 FILLER_47_163 ();
 sg13g2_decap_4 FILLER_47_178 ();
 sg13g2_fill_2 FILLER_47_182 ();
 sg13g2_fill_1 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_247 ();
 sg13g2_decap_4 FILLER_47_254 ();
 sg13g2_fill_1 FILLER_47_292 ();
 sg13g2_decap_8 FILLER_47_303 ();
 sg13g2_fill_2 FILLER_47_310 ();
 sg13g2_decap_8 FILLER_47_338 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_fill_2 FILLER_47_385 ();
 sg13g2_fill_1 FILLER_47_387 ();
 sg13g2_decap_8 FILLER_47_393 ();
 sg13g2_decap_8 FILLER_47_400 ();
 sg13g2_fill_2 FILLER_47_433 ();
 sg13g2_fill_2 FILLER_47_443 ();
 sg13g2_fill_1 FILLER_47_445 ();
 sg13g2_fill_1 FILLER_47_472 ();
 sg13g2_decap_8 FILLER_47_507 ();
 sg13g2_decap_8 FILLER_47_514 ();
 sg13g2_decap_8 FILLER_47_521 ();
 sg13g2_decap_8 FILLER_47_528 ();
 sg13g2_decap_8 FILLER_47_535 ();
 sg13g2_fill_1 FILLER_47_542 ();
 sg13g2_decap_4 FILLER_47_548 ();
 sg13g2_fill_1 FILLER_47_552 ();
 sg13g2_decap_8 FILLER_47_566 ();
 sg13g2_decap_8 FILLER_47_573 ();
 sg13g2_decap_8 FILLER_47_580 ();
 sg13g2_fill_2 FILLER_47_587 ();
 sg13g2_decap_4 FILLER_47_593 ();
 sg13g2_fill_2 FILLER_47_597 ();
 sg13g2_decap_8 FILLER_47_628 ();
 sg13g2_decap_8 FILLER_47_635 ();
 sg13g2_decap_4 FILLER_47_746 ();
 sg13g2_decap_4 FILLER_47_784 ();
 sg13g2_fill_1 FILLER_47_788 ();
 sg13g2_decap_4 FILLER_47_815 ();
 sg13g2_decap_8 FILLER_47_829 ();
 sg13g2_decap_8 FILLER_47_836 ();
 sg13g2_fill_2 FILLER_47_843 ();
 sg13g2_fill_1 FILLER_47_845 ();
 sg13g2_decap_8 FILLER_47_872 ();
 sg13g2_decap_8 FILLER_47_879 ();
 sg13g2_fill_2 FILLER_47_886 ();
 sg13g2_fill_1 FILLER_47_888 ();
 sg13g2_fill_1 FILLER_47_928 ();
 sg13g2_decap_8 FILLER_47_981 ();
 sg13g2_decap_8 FILLER_47_988 ();
 sg13g2_decap_8 FILLER_47_995 ();
 sg13g2_decap_8 FILLER_47_1002 ();
 sg13g2_decap_4 FILLER_47_1009 ();
 sg13g2_fill_1 FILLER_47_1013 ();
 sg13g2_decap_8 FILLER_47_1019 ();
 sg13g2_decap_8 FILLER_47_1026 ();
 sg13g2_fill_1 FILLER_47_1033 ();
 sg13g2_decap_8 FILLER_47_1129 ();
 sg13g2_decap_8 FILLER_47_1251 ();
 sg13g2_decap_8 FILLER_47_1258 ();
 sg13g2_fill_1 FILLER_47_1265 ();
 sg13g2_decap_8 FILLER_47_1270 ();
 sg13g2_decap_4 FILLER_47_1277 ();
 sg13g2_fill_1 FILLER_47_1281 ();
 sg13g2_fill_1 FILLER_47_1312 ();
 sg13g2_decap_8 FILLER_47_1319 ();
 sg13g2_decap_8 FILLER_47_1326 ();
 sg13g2_decap_4 FILLER_47_1333 ();
 sg13g2_fill_2 FILLER_47_1337 ();
 sg13g2_decap_4 FILLER_47_1344 ();
 sg13g2_fill_1 FILLER_47_1348 ();
 sg13g2_decap_8 FILLER_47_1380 ();
 sg13g2_decap_8 FILLER_47_1387 ();
 sg13g2_decap_8 FILLER_47_1394 ();
 sg13g2_decap_8 FILLER_47_1427 ();
 sg13g2_decap_8 FILLER_47_1434 ();
 sg13g2_decap_8 FILLER_47_1441 ();
 sg13g2_decap_4 FILLER_47_1448 ();
 sg13g2_fill_1 FILLER_47_1452 ();
 sg13g2_decap_8 FILLER_47_1474 ();
 sg13g2_fill_2 FILLER_47_1481 ();
 sg13g2_fill_1 FILLER_47_1483 ();
 sg13g2_fill_2 FILLER_47_1499 ();
 sg13g2_fill_2 FILLER_47_1533 ();
 sg13g2_fill_1 FILLER_47_1540 ();
 sg13g2_fill_2 FILLER_47_1587 ();
 sg13g2_fill_1 FILLER_47_1669 ();
 sg13g2_decap_8 FILLER_47_1682 ();
 sg13g2_decap_4 FILLER_47_1689 ();
 sg13g2_fill_2 FILLER_47_1794 ();
 sg13g2_fill_2 FILLER_47_1874 ();
 sg13g2_decap_8 FILLER_47_1902 ();
 sg13g2_decap_8 FILLER_47_1909 ();
 sg13g2_fill_2 FILLER_47_1928 ();
 sg13g2_fill_1 FILLER_47_1930 ();
 sg13g2_fill_1 FILLER_47_1963 ();
 sg13g2_decap_8 FILLER_47_1990 ();
 sg13g2_decap_4 FILLER_47_1997 ();
 sg13g2_fill_2 FILLER_47_2053 ();
 sg13g2_fill_1 FILLER_47_2055 ();
 sg13g2_fill_2 FILLER_47_2082 ();
 sg13g2_decap_8 FILLER_47_2089 ();
 sg13g2_decap_4 FILLER_47_2096 ();
 sg13g2_fill_2 FILLER_47_2100 ();
 sg13g2_fill_1 FILLER_47_2128 ();
 sg13g2_fill_2 FILLER_47_2149 ();
 sg13g2_decap_4 FILLER_47_2155 ();
 sg13g2_fill_2 FILLER_47_2159 ();
 sg13g2_decap_8 FILLER_47_2250 ();
 sg13g2_decap_8 FILLER_47_2257 ();
 sg13g2_decap_8 FILLER_47_2264 ();
 sg13g2_decap_4 FILLER_47_2271 ();
 sg13g2_fill_2 FILLER_47_2275 ();
 sg13g2_decap_8 FILLER_47_2303 ();
 sg13g2_decap_8 FILLER_47_2310 ();
 sg13g2_decap_8 FILLER_47_2317 ();
 sg13g2_decap_8 FILLER_47_2324 ();
 sg13g2_decap_4 FILLER_47_2331 ();
 sg13g2_fill_1 FILLER_47_2335 ();
 sg13g2_fill_2 FILLER_47_2362 ();
 sg13g2_fill_1 FILLER_47_2367 ();
 sg13g2_decap_4 FILLER_47_2382 ();
 sg13g2_fill_1 FILLER_47_2398 ();
 sg13g2_fill_1 FILLER_47_2416 ();
 sg13g2_fill_1 FILLER_47_2422 ();
 sg13g2_fill_2 FILLER_47_2431 ();
 sg13g2_decap_4 FILLER_47_2438 ();
 sg13g2_fill_1 FILLER_47_2442 ();
 sg13g2_fill_2 FILLER_47_2495 ();
 sg13g2_fill_1 FILLER_47_2497 ();
 sg13g2_decap_8 FILLER_47_2536 ();
 sg13g2_decap_8 FILLER_47_2543 ();
 sg13g2_decap_8 FILLER_47_2550 ();
 sg13g2_decap_8 FILLER_47_2557 ();
 sg13g2_fill_1 FILLER_47_2564 ();
 sg13g2_decap_4 FILLER_47_2568 ();
 sg13g2_fill_1 FILLER_47_2572 ();
 sg13g2_decap_4 FILLER_47_2599 ();
 sg13g2_fill_1 FILLER_47_2603 ();
 sg13g2_fill_2 FILLER_47_2609 ();
 sg13g2_fill_1 FILLER_47_2611 ();
 sg13g2_decap_4 FILLER_47_2643 ();
 sg13g2_fill_2 FILLER_47_2678 ();
 sg13g2_decap_8 FILLER_47_2732 ();
 sg13g2_decap_4 FILLER_47_2739 ();
 sg13g2_decap_8 FILLER_47_2795 ();
 sg13g2_decap_8 FILLER_47_2802 ();
 sg13g2_decap_8 FILLER_47_2809 ();
 sg13g2_fill_2 FILLER_47_2816 ();
 sg13g2_fill_1 FILLER_47_2818 ();
 sg13g2_decap_8 FILLER_47_2849 ();
 sg13g2_decap_8 FILLER_47_2856 ();
 sg13g2_decap_8 FILLER_47_2863 ();
 sg13g2_fill_2 FILLER_47_2870 ();
 sg13g2_decap_8 FILLER_47_2915 ();
 sg13g2_decap_4 FILLER_47_2922 ();
 sg13g2_fill_2 FILLER_47_2926 ();
 sg13g2_fill_2 FILLER_47_2938 ();
 sg13g2_fill_1 FILLER_47_2940 ();
 sg13g2_fill_2 FILLER_47_2949 ();
 sg13g2_fill_1 FILLER_47_2951 ();
 sg13g2_decap_8 FILLER_47_2970 ();
 sg13g2_decap_8 FILLER_47_2977 ();
 sg13g2_decap_8 FILLER_47_2984 ();
 sg13g2_decap_4 FILLER_47_2991 ();
 sg13g2_fill_2 FILLER_47_2995 ();
 sg13g2_decap_8 FILLER_47_3023 ();
 sg13g2_decap_8 FILLER_47_3030 ();
 sg13g2_fill_1 FILLER_47_3037 ();
 sg13g2_fill_2 FILLER_47_3055 ();
 sg13g2_fill_1 FILLER_47_3057 ();
 sg13g2_decap_8 FILLER_47_3076 ();
 sg13g2_decap_8 FILLER_47_3083 ();
 sg13g2_decap_4 FILLER_47_3090 ();
 sg13g2_decap_8 FILLER_47_3098 ();
 sg13g2_fill_2 FILLER_47_3105 ();
 sg13g2_fill_1 FILLER_47_3107 ();
 sg13g2_decap_8 FILLER_47_3113 ();
 sg13g2_decap_8 FILLER_47_3120 ();
 sg13g2_decap_8 FILLER_47_3127 ();
 sg13g2_decap_8 FILLER_47_3134 ();
 sg13g2_decap_8 FILLER_47_3141 ();
 sg13g2_decap_8 FILLER_47_3148 ();
 sg13g2_fill_2 FILLER_47_3155 ();
 sg13g2_decap_8 FILLER_47_3183 ();
 sg13g2_decap_8 FILLER_47_3190 ();
 sg13g2_decap_8 FILLER_47_3197 ();
 sg13g2_decap_8 FILLER_47_3204 ();
 sg13g2_decap_8 FILLER_47_3211 ();
 sg13g2_decap_4 FILLER_47_3218 ();
 sg13g2_fill_1 FILLER_47_3222 ();
 sg13g2_decap_8 FILLER_47_3226 ();
 sg13g2_decap_8 FILLER_47_3233 ();
 sg13g2_decap_8 FILLER_47_3240 ();
 sg13g2_decap_8 FILLER_47_3247 ();
 sg13g2_decap_8 FILLER_47_3254 ();
 sg13g2_decap_8 FILLER_47_3261 ();
 sg13g2_decap_8 FILLER_47_3268 ();
 sg13g2_decap_8 FILLER_47_3275 ();
 sg13g2_decap_8 FILLER_47_3282 ();
 sg13g2_decap_8 FILLER_47_3289 ();
 sg13g2_decap_8 FILLER_47_3296 ();
 sg13g2_decap_8 FILLER_47_3303 ();
 sg13g2_decap_8 FILLER_47_3310 ();
 sg13g2_decap_8 FILLER_47_3317 ();
 sg13g2_decap_8 FILLER_47_3324 ();
 sg13g2_decap_8 FILLER_47_3331 ();
 sg13g2_decap_8 FILLER_47_3338 ();
 sg13g2_decap_8 FILLER_47_3345 ();
 sg13g2_decap_8 FILLER_47_3352 ();
 sg13g2_decap_8 FILLER_47_3359 ();
 sg13g2_decap_8 FILLER_47_3366 ();
 sg13g2_decap_8 FILLER_47_3373 ();
 sg13g2_decap_8 FILLER_47_3380 ();
 sg13g2_decap_8 FILLER_47_3387 ();
 sg13g2_decap_8 FILLER_47_3394 ();
 sg13g2_decap_8 FILLER_47_3401 ();
 sg13g2_decap_8 FILLER_47_3408 ();
 sg13g2_decap_8 FILLER_47_3415 ();
 sg13g2_decap_8 FILLER_47_3422 ();
 sg13g2_decap_8 FILLER_47_3429 ();
 sg13g2_decap_8 FILLER_47_3436 ();
 sg13g2_decap_8 FILLER_47_3443 ();
 sg13g2_decap_8 FILLER_47_3450 ();
 sg13g2_decap_8 FILLER_47_3457 ();
 sg13g2_decap_8 FILLER_47_3464 ();
 sg13g2_decap_8 FILLER_47_3471 ();
 sg13g2_decap_8 FILLER_47_3478 ();
 sg13g2_decap_8 FILLER_47_3485 ();
 sg13g2_decap_8 FILLER_47_3492 ();
 sg13g2_decap_8 FILLER_47_3499 ();
 sg13g2_decap_8 FILLER_47_3506 ();
 sg13g2_decap_8 FILLER_47_3513 ();
 sg13g2_decap_8 FILLER_47_3520 ();
 sg13g2_decap_8 FILLER_47_3527 ();
 sg13g2_decap_8 FILLER_47_3534 ();
 sg13g2_decap_8 FILLER_47_3541 ();
 sg13g2_decap_8 FILLER_47_3548 ();
 sg13g2_decap_8 FILLER_47_3555 ();
 sg13g2_decap_8 FILLER_47_3562 ();
 sg13g2_decap_8 FILLER_47_3569 ();
 sg13g2_decap_4 FILLER_47_3576 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_4 FILLER_48_143 ();
 sg13g2_fill_2 FILLER_48_147 ();
 sg13g2_fill_1 FILLER_48_152 ();
 sg13g2_fill_2 FILLER_48_241 ();
 sg13g2_fill_1 FILLER_48_254 ();
 sg13g2_decap_8 FILLER_48_307 ();
 sg13g2_decap_4 FILLER_48_314 ();
 sg13g2_fill_2 FILLER_48_318 ();
 sg13g2_decap_8 FILLER_48_328 ();
 sg13g2_decap_4 FILLER_48_335 ();
 sg13g2_fill_2 FILLER_48_339 ();
 sg13g2_decap_8 FILLER_48_367 ();
 sg13g2_decap_8 FILLER_48_374 ();
 sg13g2_fill_2 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_48_417 ();
 sg13g2_fill_1 FILLER_48_424 ();
 sg13g2_fill_2 FILLER_48_430 ();
 sg13g2_fill_1 FILLER_48_432 ();
 sg13g2_decap_4 FILLER_48_438 ();
 sg13g2_fill_1 FILLER_48_442 ();
 sg13g2_decap_8 FILLER_48_459 ();
 sg13g2_fill_1 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_520 ();
 sg13g2_decap_4 FILLER_48_527 ();
 sg13g2_fill_2 FILLER_48_557 ();
 sg13g2_fill_1 FILLER_48_559 ();
 sg13g2_decap_8 FILLER_48_576 ();
 sg13g2_decap_8 FILLER_48_583 ();
 sg13g2_fill_2 FILLER_48_668 ();
 sg13g2_decap_8 FILLER_48_684 ();
 sg13g2_decap_8 FILLER_48_691 ();
 sg13g2_decap_4 FILLER_48_698 ();
 sg13g2_fill_2 FILLER_48_702 ();
 sg13g2_decap_8 FILLER_48_737 ();
 sg13g2_decap_8 FILLER_48_744 ();
 sg13g2_fill_2 FILLER_48_751 ();
 sg13g2_fill_1 FILLER_48_753 ();
 sg13g2_fill_2 FILLER_48_758 ();
 sg13g2_fill_1 FILLER_48_760 ();
 sg13g2_fill_2 FILLER_48_817 ();
 sg13g2_decap_4 FILLER_48_832 ();
 sg13g2_decap_8 FILLER_48_870 ();
 sg13g2_decap_4 FILLER_48_877 ();
 sg13g2_fill_2 FILLER_48_881 ();
 sg13g2_decap_4 FILLER_48_922 ();
 sg13g2_decap_8 FILLER_48_971 ();
 sg13g2_decap_4 FILLER_48_1104 ();
 sg13g2_decap_4 FILLER_48_1112 ();
 sg13g2_fill_1 FILLER_48_1116 ();
 sg13g2_fill_2 FILLER_48_1178 ();
 sg13g2_fill_1 FILLER_48_1180 ();
 sg13g2_fill_1 FILLER_48_1241 ();
 sg13g2_fill_2 FILLER_48_1247 ();
 sg13g2_decap_8 FILLER_48_1261 ();
 sg13g2_decap_4 FILLER_48_1330 ();
 sg13g2_fill_1 FILLER_48_1334 ();
 sg13g2_decap_8 FILLER_48_1379 ();
 sg13g2_fill_2 FILLER_48_1386 ();
 sg13g2_fill_1 FILLER_48_1388 ();
 sg13g2_decap_8 FILLER_48_1434 ();
 sg13g2_fill_1 FILLER_48_1441 ();
 sg13g2_fill_2 FILLER_48_1480 ();
 sg13g2_fill_1 FILLER_48_1482 ();
 sg13g2_fill_2 FILLER_48_1527 ();
 sg13g2_fill_1 FILLER_48_1621 ();
 sg13g2_fill_2 FILLER_48_1656 ();
 sg13g2_fill_1 FILLER_48_1658 ();
 sg13g2_fill_2 FILLER_48_1664 ();
 sg13g2_fill_1 FILLER_48_1666 ();
 sg13g2_decap_4 FILLER_48_1687 ();
 sg13g2_fill_1 FILLER_48_1691 ();
 sg13g2_fill_2 FILLER_48_1704 ();
 sg13g2_fill_1 FILLER_48_1706 ();
 sg13g2_decap_8 FILLER_48_1744 ();
 sg13g2_decap_8 FILLER_48_1751 ();
 sg13g2_fill_1 FILLER_48_1758 ();
 sg13g2_decap_4 FILLER_48_1797 ();
 sg13g2_decap_8 FILLER_48_1807 ();
 sg13g2_decap_8 FILLER_48_1814 ();
 sg13g2_decap_8 FILLER_48_1821 ();
 sg13g2_decap_8 FILLER_48_1833 ();
 sg13g2_fill_1 FILLER_48_1882 ();
 sg13g2_decap_8 FILLER_48_1889 ();
 sg13g2_fill_2 FILLER_48_1896 ();
 sg13g2_fill_1 FILLER_48_1898 ();
 sg13g2_fill_2 FILLER_48_1907 ();
 sg13g2_decap_8 FILLER_48_1961 ();
 sg13g2_decap_4 FILLER_48_1968 ();
 sg13g2_fill_2 FILLER_48_1972 ();
 sg13g2_decap_4 FILLER_48_1980 ();
 sg13g2_fill_1 FILLER_48_2028 ();
 sg13g2_fill_2 FILLER_48_2035 ();
 sg13g2_fill_1 FILLER_48_2037 ();
 sg13g2_decap_8 FILLER_48_2095 ();
 sg13g2_decap_8 FILLER_48_2102 ();
 sg13g2_decap_8 FILLER_48_2109 ();
 sg13g2_decap_4 FILLER_48_2116 ();
 sg13g2_fill_2 FILLER_48_2120 ();
 sg13g2_fill_1 FILLER_48_2177 ();
 sg13g2_decap_4 FILLER_48_2184 ();
 sg13g2_decap_8 FILLER_48_2240 ();
 sg13g2_decap_8 FILLER_48_2247 ();
 sg13g2_decap_4 FILLER_48_2254 ();
 sg13g2_fill_1 FILLER_48_2258 ();
 sg13g2_decap_8 FILLER_48_2264 ();
 sg13g2_decap_8 FILLER_48_2271 ();
 sg13g2_fill_2 FILLER_48_2278 ();
 sg13g2_fill_1 FILLER_48_2280 ();
 sg13g2_fill_2 FILLER_48_2290 ();
 sg13g2_fill_1 FILLER_48_2292 ();
 sg13g2_decap_8 FILLER_48_2319 ();
 sg13g2_decap_8 FILLER_48_2326 ();
 sg13g2_decap_8 FILLER_48_2333 ();
 sg13g2_decap_8 FILLER_48_2340 ();
 sg13g2_fill_1 FILLER_48_2347 ();
 sg13g2_decap_8 FILLER_48_2360 ();
 sg13g2_decap_4 FILLER_48_2367 ();
 sg13g2_fill_1 FILLER_48_2371 ();
 sg13g2_fill_2 FILLER_48_2383 ();
 sg13g2_fill_2 FILLER_48_2417 ();
 sg13g2_fill_2 FILLER_48_2435 ();
 sg13g2_fill_1 FILLER_48_2437 ();
 sg13g2_decap_4 FILLER_48_2469 ();
 sg13g2_fill_1 FILLER_48_2473 ();
 sg13g2_fill_2 FILLER_48_2479 ();
 sg13g2_decap_8 FILLER_48_2489 ();
 sg13g2_decap_4 FILLER_48_2496 ();
 sg13g2_fill_2 FILLER_48_2500 ();
 sg13g2_decap_4 FILLER_48_2598 ();
 sg13g2_fill_1 FILLER_48_2602 ();
 sg13g2_decap_4 FILLER_48_2642 ();
 sg13g2_fill_1 FILLER_48_2646 ();
 sg13g2_decap_8 FILLER_48_2699 ();
 sg13g2_decap_4 FILLER_48_2706 ();
 sg13g2_fill_1 FILLER_48_2710 ();
 sg13g2_decap_8 FILLER_48_2721 ();
 sg13g2_decap_8 FILLER_48_2728 ();
 sg13g2_decap_8 FILLER_48_2735 ();
 sg13g2_decap_8 FILLER_48_2742 ();
 sg13g2_fill_2 FILLER_48_2749 ();
 sg13g2_fill_1 FILLER_48_2751 ();
 sg13g2_decap_8 FILLER_48_2783 ();
 sg13g2_decap_8 FILLER_48_2790 ();
 sg13g2_decap_8 FILLER_48_2797 ();
 sg13g2_fill_2 FILLER_48_2804 ();
 sg13g2_fill_1 FILLER_48_2806 ();
 sg13g2_decap_8 FILLER_48_2923 ();
 sg13g2_decap_8 FILLER_48_2930 ();
 sg13g2_decap_8 FILLER_48_2937 ();
 sg13g2_decap_4 FILLER_48_2944 ();
 sg13g2_fill_1 FILLER_48_2948 ();
 sg13g2_decap_8 FILLER_48_2975 ();
 sg13g2_decap_8 FILLER_48_2982 ();
 sg13g2_decap_8 FILLER_48_2994 ();
 sg13g2_fill_2 FILLER_48_3001 ();
 sg13g2_decap_8 FILLER_48_3029 ();
 sg13g2_decap_8 FILLER_48_3036 ();
 sg13g2_fill_2 FILLER_48_3043 ();
 sg13g2_fill_1 FILLER_48_3045 ();
 sg13g2_decap_8 FILLER_48_3072 ();
 sg13g2_decap_8 FILLER_48_3079 ();
 sg13g2_decap_8 FILLER_48_3086 ();
 sg13g2_decap_8 FILLER_48_3093 ();
 sg13g2_decap_8 FILLER_48_3100 ();
 sg13g2_decap_8 FILLER_48_3107 ();
 sg13g2_decap_8 FILLER_48_3114 ();
 sg13g2_decap_8 FILLER_48_3121 ();
 sg13g2_decap_8 FILLER_48_3128 ();
 sg13g2_decap_8 FILLER_48_3135 ();
 sg13g2_decap_8 FILLER_48_3142 ();
 sg13g2_decap_8 FILLER_48_3149 ();
 sg13g2_decap_4 FILLER_48_3156 ();
 sg13g2_fill_2 FILLER_48_3160 ();
 sg13g2_fill_2 FILLER_48_3166 ();
 sg13g2_decap_8 FILLER_48_3172 ();
 sg13g2_decap_8 FILLER_48_3179 ();
 sg13g2_decap_8 FILLER_48_3186 ();
 sg13g2_decap_8 FILLER_48_3193 ();
 sg13g2_decap_8 FILLER_48_3200 ();
 sg13g2_decap_8 FILLER_48_3207 ();
 sg13g2_decap_8 FILLER_48_3214 ();
 sg13g2_decap_8 FILLER_48_3221 ();
 sg13g2_decap_8 FILLER_48_3228 ();
 sg13g2_decap_8 FILLER_48_3235 ();
 sg13g2_decap_8 FILLER_48_3242 ();
 sg13g2_decap_8 FILLER_48_3249 ();
 sg13g2_decap_8 FILLER_48_3256 ();
 sg13g2_decap_8 FILLER_48_3263 ();
 sg13g2_decap_8 FILLER_48_3270 ();
 sg13g2_decap_8 FILLER_48_3277 ();
 sg13g2_decap_8 FILLER_48_3284 ();
 sg13g2_decap_8 FILLER_48_3291 ();
 sg13g2_decap_8 FILLER_48_3298 ();
 sg13g2_decap_8 FILLER_48_3305 ();
 sg13g2_decap_8 FILLER_48_3312 ();
 sg13g2_decap_8 FILLER_48_3319 ();
 sg13g2_decap_8 FILLER_48_3326 ();
 sg13g2_decap_8 FILLER_48_3333 ();
 sg13g2_decap_8 FILLER_48_3340 ();
 sg13g2_decap_8 FILLER_48_3347 ();
 sg13g2_decap_8 FILLER_48_3354 ();
 sg13g2_decap_8 FILLER_48_3361 ();
 sg13g2_decap_8 FILLER_48_3368 ();
 sg13g2_decap_8 FILLER_48_3375 ();
 sg13g2_decap_8 FILLER_48_3382 ();
 sg13g2_decap_8 FILLER_48_3389 ();
 sg13g2_decap_8 FILLER_48_3396 ();
 sg13g2_decap_8 FILLER_48_3403 ();
 sg13g2_decap_8 FILLER_48_3410 ();
 sg13g2_decap_8 FILLER_48_3417 ();
 sg13g2_decap_8 FILLER_48_3424 ();
 sg13g2_decap_8 FILLER_48_3431 ();
 sg13g2_decap_8 FILLER_48_3438 ();
 sg13g2_decap_8 FILLER_48_3445 ();
 sg13g2_decap_8 FILLER_48_3452 ();
 sg13g2_decap_8 FILLER_48_3459 ();
 sg13g2_decap_8 FILLER_48_3466 ();
 sg13g2_decap_8 FILLER_48_3473 ();
 sg13g2_decap_8 FILLER_48_3480 ();
 sg13g2_decap_8 FILLER_48_3487 ();
 sg13g2_decap_8 FILLER_48_3494 ();
 sg13g2_decap_8 FILLER_48_3501 ();
 sg13g2_decap_8 FILLER_48_3508 ();
 sg13g2_decap_8 FILLER_48_3515 ();
 sg13g2_decap_8 FILLER_48_3522 ();
 sg13g2_decap_8 FILLER_48_3529 ();
 sg13g2_decap_8 FILLER_48_3536 ();
 sg13g2_decap_8 FILLER_48_3543 ();
 sg13g2_decap_8 FILLER_48_3550 ();
 sg13g2_decap_8 FILLER_48_3557 ();
 sg13g2_decap_8 FILLER_48_3564 ();
 sg13g2_decap_8 FILLER_48_3571 ();
 sg13g2_fill_2 FILLER_48_3578 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_4 FILLER_49_84 ();
 sg13g2_fill_1 FILLER_49_88 ();
 sg13g2_fill_2 FILLER_49_118 ();
 sg13g2_decap_8 FILLER_49_188 ();
 sg13g2_decap_8 FILLER_49_195 ();
 sg13g2_fill_2 FILLER_49_202 ();
 sg13g2_fill_2 FILLER_49_230 ();
 sg13g2_fill_1 FILLER_49_232 ();
 sg13g2_decap_8 FILLER_49_267 ();
 sg13g2_decap_8 FILLER_49_274 ();
 sg13g2_fill_2 FILLER_49_281 ();
 sg13g2_decap_4 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_362 ();
 sg13g2_fill_1 FILLER_49_376 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_4 FILLER_49_455 ();
 sg13g2_fill_2 FILLER_49_459 ();
 sg13g2_fill_2 FILLER_49_487 ();
 sg13g2_fill_2 FILLER_49_494 ();
 sg13g2_fill_1 FILLER_49_496 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_decap_4 FILLER_49_543 ();
 sg13g2_fill_2 FILLER_49_547 ();
 sg13g2_decap_8 FILLER_49_580 ();
 sg13g2_decap_8 FILLER_49_587 ();
 sg13g2_decap_4 FILLER_49_594 ();
 sg13g2_fill_1 FILLER_49_598 ();
 sg13g2_decap_4 FILLER_49_641 ();
 sg13g2_fill_2 FILLER_49_645 ();
 sg13g2_fill_2 FILLER_49_650 ();
 sg13g2_decap_8 FILLER_49_656 ();
 sg13g2_fill_2 FILLER_49_663 ();
 sg13g2_fill_1 FILLER_49_665 ();
 sg13g2_decap_4 FILLER_49_676 ();
 sg13g2_fill_1 FILLER_49_680 ();
 sg13g2_decap_8 FILLER_49_689 ();
 sg13g2_decap_8 FILLER_49_696 ();
 sg13g2_decap_4 FILLER_49_703 ();
 sg13g2_decap_8 FILLER_49_737 ();
 sg13g2_decap_8 FILLER_49_744 ();
 sg13g2_decap_8 FILLER_49_751 ();
 sg13g2_decap_8 FILLER_49_758 ();
 sg13g2_decap_8 FILLER_49_765 ();
 sg13g2_decap_8 FILLER_49_780 ();
 sg13g2_decap_8 FILLER_49_787 ();
 sg13g2_fill_2 FILLER_49_794 ();
 sg13g2_fill_1 FILLER_49_796 ();
 sg13g2_decap_8 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_831 ();
 sg13g2_decap_4 FILLER_49_838 ();
 sg13g2_fill_2 FILLER_49_842 ();
 sg13g2_decap_8 FILLER_49_874 ();
 sg13g2_decap_8 FILLER_49_881 ();
 sg13g2_fill_2 FILLER_49_932 ();
 sg13g2_decap_8 FILLER_49_963 ();
 sg13g2_decap_4 FILLER_49_970 ();
 sg13g2_fill_2 FILLER_49_974 ();
 sg13g2_fill_2 FILLER_49_1033 ();
 sg13g2_decap_4 FILLER_49_1061 ();
 sg13g2_fill_2 FILLER_49_1065 ();
 sg13g2_decap_8 FILLER_49_1125 ();
 sg13g2_fill_2 FILLER_49_1132 ();
 sg13g2_fill_2 FILLER_49_1160 ();
 sg13g2_fill_1 FILLER_49_1176 ();
 sg13g2_decap_8 FILLER_49_1183 ();
 sg13g2_decap_8 FILLER_49_1190 ();
 sg13g2_fill_2 FILLER_49_1197 ();
 sg13g2_fill_1 FILLER_49_1199 ();
 sg13g2_fill_1 FILLER_49_1268 ();
 sg13g2_decap_8 FILLER_49_1321 ();
 sg13g2_decap_8 FILLER_49_1328 ();
 sg13g2_fill_1 FILLER_49_1369 ();
 sg13g2_decap_8 FILLER_49_1428 ();
 sg13g2_decap_4 FILLER_49_1435 ();
 sg13g2_fill_1 FILLER_49_1439 ();
 sg13g2_fill_1 FILLER_49_1492 ();
 sg13g2_fill_1 FILLER_49_1504 ();
 sg13g2_fill_2 FILLER_49_1515 ();
 sg13g2_fill_1 FILLER_49_1530 ();
 sg13g2_fill_1 FILLER_49_1541 ();
 sg13g2_fill_1 FILLER_49_1620 ();
 sg13g2_fill_1 FILLER_49_1631 ();
 sg13g2_fill_1 FILLER_49_1642 ();
 sg13g2_fill_2 FILLER_49_1654 ();
 sg13g2_decap_4 FILLER_49_1688 ();
 sg13g2_fill_1 FILLER_49_1692 ();
 sg13g2_fill_2 FILLER_49_1703 ();
 sg13g2_fill_2 FILLER_49_1710 ();
 sg13g2_decap_8 FILLER_49_1738 ();
 sg13g2_decap_4 FILLER_49_1777 ();
 sg13g2_decap_8 FILLER_49_1800 ();
 sg13g2_decap_8 FILLER_49_1807 ();
 sg13g2_decap_4 FILLER_49_1814 ();
 sg13g2_fill_1 FILLER_49_1818 ();
 sg13g2_decap_8 FILLER_49_1831 ();
 sg13g2_fill_2 FILLER_49_1838 ();
 sg13g2_fill_1 FILLER_49_1866 ();
 sg13g2_decap_8 FILLER_49_1872 ();
 sg13g2_decap_8 FILLER_49_1879 ();
 sg13g2_decap_4 FILLER_49_1886 ();
 sg13g2_decap_4 FILLER_49_1924 ();
 sg13g2_fill_2 FILLER_49_1928 ();
 sg13g2_decap_4 FILLER_49_1964 ();
 sg13g2_fill_1 FILLER_49_1968 ();
 sg13g2_decap_4 FILLER_49_1984 ();
 sg13g2_fill_1 FILLER_49_1988 ();
 sg13g2_decap_8 FILLER_49_2022 ();
 sg13g2_decap_8 FILLER_49_2029 ();
 sg13g2_decap_8 FILLER_49_2036 ();
 sg13g2_decap_8 FILLER_49_2043 ();
 sg13g2_decap_8 FILLER_49_2050 ();
 sg13g2_fill_2 FILLER_49_2057 ();
 sg13g2_fill_2 FILLER_49_2085 ();
 sg13g2_fill_1 FILLER_49_2087 ();
 sg13g2_decap_4 FILLER_49_2127 ();
 sg13g2_decap_8 FILLER_49_2162 ();
 sg13g2_fill_2 FILLER_49_2169 ();
 sg13g2_fill_1 FILLER_49_2171 ();
 sg13g2_fill_1 FILLER_49_2198 ();
 sg13g2_decap_8 FILLER_49_2205 ();
 sg13g2_fill_2 FILLER_49_2212 ();
 sg13g2_decap_8 FILLER_49_2240 ();
 sg13g2_fill_2 FILLER_49_2247 ();
 sg13g2_fill_1 FILLER_49_2249 ();
 sg13g2_decap_4 FILLER_49_2254 ();
 sg13g2_fill_2 FILLER_49_2258 ();
 sg13g2_decap_8 FILLER_49_2265 ();
 sg13g2_fill_1 FILLER_49_2272 ();
 sg13g2_decap_8 FILLER_49_2299 ();
 sg13g2_decap_8 FILLER_49_2306 ();
 sg13g2_decap_8 FILLER_49_2313 ();
 sg13g2_fill_2 FILLER_49_2320 ();
 sg13g2_fill_1 FILLER_49_2322 ();
 sg13g2_fill_2 FILLER_49_2354 ();
 sg13g2_fill_1 FILLER_49_2356 ();
 sg13g2_fill_1 FILLER_49_2379 ();
 sg13g2_fill_1 FILLER_49_2399 ();
 sg13g2_decap_4 FILLER_49_2409 ();
 sg13g2_fill_2 FILLER_49_2413 ();
 sg13g2_decap_4 FILLER_49_2431 ();
 sg13g2_fill_1 FILLER_49_2440 ();
 sg13g2_decap_8 FILLER_49_2457 ();
 sg13g2_decap_8 FILLER_49_2464 ();
 sg13g2_decap_8 FILLER_49_2497 ();
 sg13g2_decap_8 FILLER_49_2504 ();
 sg13g2_decap_8 FILLER_49_2537 ();
 sg13g2_decap_8 FILLER_49_2544 ();
 sg13g2_fill_1 FILLER_49_2608 ();
 sg13g2_decap_4 FILLER_49_2648 ();
 sg13g2_fill_2 FILLER_49_2652 ();
 sg13g2_decap_8 FILLER_49_2693 ();
 sg13g2_decap_4 FILLER_49_2726 ();
 sg13g2_fill_1 FILLER_49_2740 ();
 sg13g2_decap_8 FILLER_49_2747 ();
 sg13g2_fill_2 FILLER_49_2754 ();
 sg13g2_fill_1 FILLER_49_2756 ();
 sg13g2_decap_4 FILLER_49_2762 ();
 sg13g2_fill_1 FILLER_49_2766 ();
 sg13g2_fill_1 FILLER_49_2772 ();
 sg13g2_decap_8 FILLER_49_2799 ();
 sg13g2_decap_4 FILLER_49_2806 ();
 sg13g2_fill_2 FILLER_49_2810 ();
 sg13g2_decap_4 FILLER_49_2851 ();
 sg13g2_fill_2 FILLER_49_2855 ();
 sg13g2_fill_1 FILLER_49_2872 ();
 sg13g2_decap_4 FILLER_49_2931 ();
 sg13g2_fill_2 FILLER_49_2935 ();
 sg13g2_fill_2 FILLER_49_2978 ();
 sg13g2_fill_1 FILLER_49_2980 ();
 sg13g2_decap_8 FILLER_49_3033 ();
 sg13g2_decap_8 FILLER_49_3040 ();
 sg13g2_fill_2 FILLER_49_3047 ();
 sg13g2_fill_1 FILLER_49_3049 ();
 sg13g2_decap_8 FILLER_49_3076 ();
 sg13g2_decap_8 FILLER_49_3083 ();
 sg13g2_decap_8 FILLER_49_3090 ();
 sg13g2_decap_8 FILLER_49_3097 ();
 sg13g2_decap_8 FILLER_49_3104 ();
 sg13g2_decap_8 FILLER_49_3111 ();
 sg13g2_decap_8 FILLER_49_3118 ();
 sg13g2_decap_8 FILLER_49_3125 ();
 sg13g2_decap_8 FILLER_49_3132 ();
 sg13g2_decap_8 FILLER_49_3139 ();
 sg13g2_decap_8 FILLER_49_3146 ();
 sg13g2_decap_8 FILLER_49_3153 ();
 sg13g2_decap_8 FILLER_49_3160 ();
 sg13g2_decap_8 FILLER_49_3167 ();
 sg13g2_decap_8 FILLER_49_3174 ();
 sg13g2_decap_8 FILLER_49_3181 ();
 sg13g2_decap_8 FILLER_49_3188 ();
 sg13g2_decap_8 FILLER_49_3195 ();
 sg13g2_decap_8 FILLER_49_3202 ();
 sg13g2_decap_8 FILLER_49_3209 ();
 sg13g2_decap_8 FILLER_49_3216 ();
 sg13g2_decap_8 FILLER_49_3223 ();
 sg13g2_decap_8 FILLER_49_3230 ();
 sg13g2_decap_8 FILLER_49_3237 ();
 sg13g2_decap_8 FILLER_49_3244 ();
 sg13g2_decap_8 FILLER_49_3251 ();
 sg13g2_decap_8 FILLER_49_3258 ();
 sg13g2_decap_8 FILLER_49_3265 ();
 sg13g2_decap_8 FILLER_49_3272 ();
 sg13g2_decap_8 FILLER_49_3279 ();
 sg13g2_decap_8 FILLER_49_3286 ();
 sg13g2_decap_8 FILLER_49_3293 ();
 sg13g2_decap_8 FILLER_49_3300 ();
 sg13g2_decap_8 FILLER_49_3307 ();
 sg13g2_decap_8 FILLER_49_3314 ();
 sg13g2_decap_8 FILLER_49_3321 ();
 sg13g2_decap_8 FILLER_49_3328 ();
 sg13g2_decap_8 FILLER_49_3335 ();
 sg13g2_decap_8 FILLER_49_3342 ();
 sg13g2_decap_8 FILLER_49_3349 ();
 sg13g2_decap_8 FILLER_49_3356 ();
 sg13g2_decap_8 FILLER_49_3363 ();
 sg13g2_decap_8 FILLER_49_3370 ();
 sg13g2_decap_8 FILLER_49_3377 ();
 sg13g2_decap_8 FILLER_49_3384 ();
 sg13g2_decap_8 FILLER_49_3391 ();
 sg13g2_decap_8 FILLER_49_3398 ();
 sg13g2_decap_8 FILLER_49_3405 ();
 sg13g2_decap_8 FILLER_49_3412 ();
 sg13g2_decap_8 FILLER_49_3419 ();
 sg13g2_decap_8 FILLER_49_3426 ();
 sg13g2_decap_8 FILLER_49_3433 ();
 sg13g2_decap_8 FILLER_49_3440 ();
 sg13g2_decap_8 FILLER_49_3447 ();
 sg13g2_decap_8 FILLER_49_3454 ();
 sg13g2_decap_8 FILLER_49_3461 ();
 sg13g2_decap_8 FILLER_49_3468 ();
 sg13g2_decap_8 FILLER_49_3475 ();
 sg13g2_decap_8 FILLER_49_3482 ();
 sg13g2_decap_8 FILLER_49_3489 ();
 sg13g2_decap_8 FILLER_49_3496 ();
 sg13g2_decap_8 FILLER_49_3503 ();
 sg13g2_decap_8 FILLER_49_3510 ();
 sg13g2_decap_8 FILLER_49_3517 ();
 sg13g2_decap_8 FILLER_49_3524 ();
 sg13g2_decap_8 FILLER_49_3531 ();
 sg13g2_decap_8 FILLER_49_3538 ();
 sg13g2_decap_8 FILLER_49_3545 ();
 sg13g2_decap_8 FILLER_49_3552 ();
 sg13g2_decap_8 FILLER_49_3559 ();
 sg13g2_decap_8 FILLER_49_3566 ();
 sg13g2_decap_8 FILLER_49_3573 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_4 FILLER_50_77 ();
 sg13g2_fill_2 FILLER_50_81 ();
 sg13g2_decap_4 FILLER_50_142 ();
 sg13g2_fill_2 FILLER_50_146 ();
 sg13g2_decap_8 FILLER_50_238 ();
 sg13g2_decap_8 FILLER_50_245 ();
 sg13g2_decap_4 FILLER_50_281 ();
 sg13g2_fill_1 FILLER_50_285 ();
 sg13g2_decap_8 FILLER_50_303 ();
 sg13g2_decap_8 FILLER_50_310 ();
 sg13g2_decap_4 FILLER_50_317 ();
 sg13g2_fill_1 FILLER_50_321 ();
 sg13g2_decap_4 FILLER_50_329 ();
 sg13g2_fill_1 FILLER_50_349 ();
 sg13g2_decap_4 FILLER_50_358 ();
 sg13g2_decap_8 FILLER_50_443 ();
 sg13g2_decap_8 FILLER_50_450 ();
 sg13g2_decap_8 FILLER_50_457 ();
 sg13g2_decap_8 FILLER_50_464 ();
 sg13g2_fill_1 FILLER_50_471 ();
 sg13g2_fill_2 FILLER_50_498 ();
 sg13g2_fill_1 FILLER_50_500 ();
 sg13g2_fill_1 FILLER_50_536 ();
 sg13g2_fill_1 FILLER_50_544 ();
 sg13g2_fill_2 FILLER_50_554 ();
 sg13g2_decap_8 FILLER_50_582 ();
 sg13g2_decap_8 FILLER_50_589 ();
 sg13g2_decap_8 FILLER_50_596 ();
 sg13g2_decap_8 FILLER_50_603 ();
 sg13g2_decap_8 FILLER_50_639 ();
 sg13g2_fill_2 FILLER_50_646 ();
 sg13g2_fill_1 FILLER_50_648 ();
 sg13g2_decap_8 FILLER_50_652 ();
 sg13g2_decap_4 FILLER_50_695 ();
 sg13g2_fill_2 FILLER_50_699 ();
 sg13g2_decap_8 FILLER_50_731 ();
 sg13g2_fill_2 FILLER_50_764 ();
 sg13g2_fill_2 FILLER_50_792 ();
 sg13g2_fill_1 FILLER_50_794 ();
 sg13g2_decap_4 FILLER_50_805 ();
 sg13g2_fill_1 FILLER_50_819 ();
 sg13g2_decap_8 FILLER_50_836 ();
 sg13g2_decap_4 FILLER_50_843 ();
 sg13g2_fill_2 FILLER_50_847 ();
 sg13g2_decap_4 FILLER_50_879 ();
 sg13g2_fill_1 FILLER_50_883 ();
 sg13g2_fill_1 FILLER_50_915 ();
 sg13g2_fill_1 FILLER_50_919 ();
 sg13g2_decap_4 FILLER_50_924 ();
 sg13g2_decap_4 FILLER_50_933 ();
 sg13g2_decap_8 FILLER_50_963 ();
 sg13g2_decap_8 FILLER_50_970 ();
 sg13g2_decap_8 FILLER_50_977 ();
 sg13g2_decap_8 FILLER_50_984 ();
 sg13g2_decap_8 FILLER_50_996 ();
 sg13g2_decap_4 FILLER_50_1003 ();
 sg13g2_fill_2 FILLER_50_1007 ();
 sg13g2_decap_8 FILLER_50_1052 ();
 sg13g2_decap_8 FILLER_50_1059 ();
 sg13g2_decap_8 FILLER_50_1066 ();
 sg13g2_decap_8 FILLER_50_1082 ();
 sg13g2_decap_8 FILLER_50_1089 ();
 sg13g2_decap_4 FILLER_50_1096 ();
 sg13g2_fill_1 FILLER_50_1100 ();
 sg13g2_decap_8 FILLER_50_1136 ();
 sg13g2_decap_8 FILLER_50_1143 ();
 sg13g2_decap_8 FILLER_50_1150 ();
 sg13g2_fill_1 FILLER_50_1157 ();
 sg13g2_decap_4 FILLER_50_1190 ();
 sg13g2_decap_8 FILLER_50_1202 ();
 sg13g2_decap_8 FILLER_50_1209 ();
 sg13g2_decap_4 FILLER_50_1216 ();
 sg13g2_fill_2 FILLER_50_1224 ();
 sg13g2_fill_1 FILLER_50_1226 ();
 sg13g2_decap_8 FILLER_50_1253 ();
 sg13g2_decap_8 FILLER_50_1260 ();
 sg13g2_fill_2 FILLER_50_1267 ();
 sg13g2_fill_1 FILLER_50_1269 ();
 sg13g2_decap_8 FILLER_50_1309 ();
 sg13g2_decap_8 FILLER_50_1316 ();
 sg13g2_decap_8 FILLER_50_1323 ();
 sg13g2_fill_1 FILLER_50_1330 ();
 sg13g2_fill_1 FILLER_50_1367 ();
 sg13g2_decap_8 FILLER_50_1417 ();
 sg13g2_decap_8 FILLER_50_1424 ();
 sg13g2_decap_8 FILLER_50_1431 ();
 sg13g2_fill_2 FILLER_50_1438 ();
 sg13g2_decap_8 FILLER_50_1481 ();
 sg13g2_decap_8 FILLER_50_1488 ();
 sg13g2_decap_8 FILLER_50_1495 ();
 sg13g2_decap_4 FILLER_50_1502 ();
 sg13g2_fill_2 FILLER_50_1506 ();
 sg13g2_fill_2 FILLER_50_1511 ();
 sg13g2_fill_1 FILLER_50_1544 ();
 sg13g2_fill_1 FILLER_50_1560 ();
 sg13g2_fill_2 FILLER_50_1608 ();
 sg13g2_fill_1 FILLER_50_1610 ();
 sg13g2_decap_4 FILLER_50_1620 ();
 sg13g2_fill_2 FILLER_50_1628 ();
 sg13g2_decap_4 FILLER_50_1642 ();
 sg13g2_fill_1 FILLER_50_1646 ();
 sg13g2_fill_2 FILLER_50_1651 ();
 sg13g2_fill_1 FILLER_50_1653 ();
 sg13g2_decap_8 FILLER_50_1680 ();
 sg13g2_fill_2 FILLER_50_1692 ();
 sg13g2_decap_8 FILLER_50_1735 ();
 sg13g2_decap_8 FILLER_50_1742 ();
 sg13g2_decap_4 FILLER_50_1749 ();
 sg13g2_decap_8 FILLER_50_1777 ();
 sg13g2_decap_8 FILLER_50_1795 ();
 sg13g2_decap_8 FILLER_50_1802 ();
 sg13g2_fill_2 FILLER_50_1809 ();
 sg13g2_fill_1 FILLER_50_1811 ();
 sg13g2_fill_1 FILLER_50_1817 ();
 sg13g2_fill_1 FILLER_50_1823 ();
 sg13g2_decap_8 FILLER_50_1833 ();
 sg13g2_fill_1 FILLER_50_1840 ();
 sg13g2_decap_4 FILLER_50_1849 ();
 sg13g2_fill_2 FILLER_50_1853 ();
 sg13g2_decap_8 FILLER_50_1866 ();
 sg13g2_decap_8 FILLER_50_1873 ();
 sg13g2_decap_4 FILLER_50_1932 ();
 sg13g2_decap_8 FILLER_50_1942 ();
 sg13g2_fill_1 FILLER_50_1949 ();
 sg13g2_fill_1 FILLER_50_1971 ();
 sg13g2_fill_2 FILLER_50_1998 ();
 sg13g2_decap_8 FILLER_50_2005 ();
 sg13g2_fill_2 FILLER_50_2012 ();
 sg13g2_fill_1 FILLER_50_2014 ();
 sg13g2_fill_1 FILLER_50_2028 ();
 sg13g2_decap_8 FILLER_50_2040 ();
 sg13g2_decap_8 FILLER_50_2047 ();
 sg13g2_decap_8 FILLER_50_2054 ();
 sg13g2_decap_8 FILLER_50_2067 ();
 sg13g2_fill_1 FILLER_50_2082 ();
 sg13g2_decap_8 FILLER_50_2109 ();
 sg13g2_decap_4 FILLER_50_2116 ();
 sg13g2_fill_1 FILLER_50_2120 ();
 sg13g2_fill_2 FILLER_50_2137 ();
 sg13g2_decap_8 FILLER_50_2144 ();
 sg13g2_decap_8 FILLER_50_2151 ();
 sg13g2_decap_8 FILLER_50_2162 ();
 sg13g2_decap_8 FILLER_50_2169 ();
 sg13g2_decap_8 FILLER_50_2176 ();
 sg13g2_decap_4 FILLER_50_2183 ();
 sg13g2_fill_1 FILLER_50_2187 ();
 sg13g2_decap_8 FILLER_50_2192 ();
 sg13g2_decap_4 FILLER_50_2199 ();
 sg13g2_fill_1 FILLER_50_2203 ();
 sg13g2_decap_8 FILLER_50_2230 ();
 sg13g2_decap_8 FILLER_50_2237 ();
 sg13g2_decap_4 FILLER_50_2244 ();
 sg13g2_fill_1 FILLER_50_2248 ();
 sg13g2_decap_8 FILLER_50_2257 ();
 sg13g2_decap_8 FILLER_50_2264 ();
 sg13g2_decap_8 FILLER_50_2389 ();
 sg13g2_decap_4 FILLER_50_2396 ();
 sg13g2_decap_8 FILLER_50_2408 ();
 sg13g2_decap_8 FILLER_50_2415 ();
 sg13g2_decap_8 FILLER_50_2422 ();
 sg13g2_decap_8 FILLER_50_2429 ();
 sg13g2_decap_4 FILLER_50_2436 ();
 sg13g2_fill_2 FILLER_50_2440 ();
 sg13g2_fill_1 FILLER_50_2450 ();
 sg13g2_decap_8 FILLER_50_2496 ();
 sg13g2_decap_8 FILLER_50_2503 ();
 sg13g2_fill_1 FILLER_50_2510 ();
 sg13g2_decap_8 FILLER_50_2537 ();
 sg13g2_decap_4 FILLER_50_2544 ();
 sg13g2_fill_1 FILLER_50_2548 ();
 sg13g2_decap_4 FILLER_50_2595 ();
 sg13g2_fill_2 FILLER_50_2609 ();
 sg13g2_decap_8 FILLER_50_2640 ();
 sg13g2_decap_8 FILLER_50_2647 ();
 sg13g2_decap_8 FILLER_50_2654 ();
 sg13g2_decap_8 FILLER_50_2661 ();
 sg13g2_fill_1 FILLER_50_2668 ();
 sg13g2_decap_8 FILLER_50_2680 ();
 sg13g2_decap_8 FILLER_50_2687 ();
 sg13g2_fill_2 FILLER_50_2694 ();
 sg13g2_decap_4 FILLER_50_2722 ();
 sg13g2_fill_1 FILLER_50_2726 ();
 sg13g2_fill_2 FILLER_50_2753 ();
 sg13g2_fill_1 FILLER_50_2755 ();
 sg13g2_decap_8 FILLER_50_2799 ();
 sg13g2_decap_8 FILLER_50_2806 ();
 sg13g2_fill_1 FILLER_50_2813 ();
 sg13g2_fill_1 FILLER_50_2819 ();
 sg13g2_fill_1 FILLER_50_2852 ();
 sg13g2_fill_2 FILLER_50_2931 ();
 sg13g2_decap_8 FILLER_50_3025 ();
 sg13g2_decap_8 FILLER_50_3032 ();
 sg13g2_decap_8 FILLER_50_3039 ();
 sg13g2_decap_8 FILLER_50_3046 ();
 sg13g2_decap_4 FILLER_50_3053 ();
 sg13g2_decap_8 FILLER_50_3065 ();
 sg13g2_decap_8 FILLER_50_3072 ();
 sg13g2_decap_8 FILLER_50_3079 ();
 sg13g2_decap_8 FILLER_50_3086 ();
 sg13g2_decap_8 FILLER_50_3093 ();
 sg13g2_decap_8 FILLER_50_3100 ();
 sg13g2_decap_8 FILLER_50_3107 ();
 sg13g2_decap_8 FILLER_50_3114 ();
 sg13g2_decap_8 FILLER_50_3121 ();
 sg13g2_decap_8 FILLER_50_3128 ();
 sg13g2_decap_8 FILLER_50_3135 ();
 sg13g2_decap_8 FILLER_50_3142 ();
 sg13g2_decap_8 FILLER_50_3149 ();
 sg13g2_decap_8 FILLER_50_3156 ();
 sg13g2_decap_8 FILLER_50_3163 ();
 sg13g2_decap_8 FILLER_50_3170 ();
 sg13g2_decap_8 FILLER_50_3177 ();
 sg13g2_decap_8 FILLER_50_3184 ();
 sg13g2_decap_8 FILLER_50_3191 ();
 sg13g2_decap_8 FILLER_50_3198 ();
 sg13g2_decap_8 FILLER_50_3205 ();
 sg13g2_decap_8 FILLER_50_3212 ();
 sg13g2_decap_8 FILLER_50_3219 ();
 sg13g2_decap_8 FILLER_50_3226 ();
 sg13g2_decap_8 FILLER_50_3233 ();
 sg13g2_decap_8 FILLER_50_3240 ();
 sg13g2_decap_8 FILLER_50_3247 ();
 sg13g2_decap_8 FILLER_50_3254 ();
 sg13g2_decap_8 FILLER_50_3261 ();
 sg13g2_decap_8 FILLER_50_3268 ();
 sg13g2_decap_8 FILLER_50_3275 ();
 sg13g2_decap_8 FILLER_50_3282 ();
 sg13g2_decap_8 FILLER_50_3289 ();
 sg13g2_decap_8 FILLER_50_3296 ();
 sg13g2_decap_8 FILLER_50_3303 ();
 sg13g2_decap_8 FILLER_50_3310 ();
 sg13g2_decap_8 FILLER_50_3317 ();
 sg13g2_decap_8 FILLER_50_3324 ();
 sg13g2_decap_8 FILLER_50_3331 ();
 sg13g2_decap_8 FILLER_50_3338 ();
 sg13g2_decap_8 FILLER_50_3345 ();
 sg13g2_decap_8 FILLER_50_3352 ();
 sg13g2_decap_8 FILLER_50_3359 ();
 sg13g2_decap_8 FILLER_50_3366 ();
 sg13g2_decap_8 FILLER_50_3373 ();
 sg13g2_decap_8 FILLER_50_3380 ();
 sg13g2_decap_8 FILLER_50_3387 ();
 sg13g2_decap_8 FILLER_50_3394 ();
 sg13g2_decap_8 FILLER_50_3401 ();
 sg13g2_decap_8 FILLER_50_3408 ();
 sg13g2_decap_8 FILLER_50_3415 ();
 sg13g2_decap_8 FILLER_50_3422 ();
 sg13g2_decap_8 FILLER_50_3429 ();
 sg13g2_decap_8 FILLER_50_3436 ();
 sg13g2_decap_8 FILLER_50_3443 ();
 sg13g2_decap_8 FILLER_50_3450 ();
 sg13g2_decap_8 FILLER_50_3457 ();
 sg13g2_decap_8 FILLER_50_3464 ();
 sg13g2_decap_8 FILLER_50_3471 ();
 sg13g2_decap_8 FILLER_50_3478 ();
 sg13g2_decap_8 FILLER_50_3485 ();
 sg13g2_decap_8 FILLER_50_3492 ();
 sg13g2_decap_8 FILLER_50_3499 ();
 sg13g2_decap_8 FILLER_50_3506 ();
 sg13g2_decap_8 FILLER_50_3513 ();
 sg13g2_decap_8 FILLER_50_3520 ();
 sg13g2_decap_8 FILLER_50_3527 ();
 sg13g2_decap_8 FILLER_50_3534 ();
 sg13g2_decap_8 FILLER_50_3541 ();
 sg13g2_decap_8 FILLER_50_3548 ();
 sg13g2_decap_8 FILLER_50_3555 ();
 sg13g2_decap_8 FILLER_50_3562 ();
 sg13g2_decap_8 FILLER_50_3569 ();
 sg13g2_decap_4 FILLER_50_3576 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_132 ();
 sg13g2_decap_8 FILLER_51_139 ();
 sg13g2_decap_8 FILLER_51_146 ();
 sg13g2_fill_2 FILLER_51_153 ();
 sg13g2_decap_8 FILLER_51_158 ();
 sg13g2_decap_8 FILLER_51_165 ();
 sg13g2_fill_1 FILLER_51_172 ();
 sg13g2_decap_8 FILLER_51_177 ();
 sg13g2_decap_8 FILLER_51_184 ();
 sg13g2_decap_8 FILLER_51_191 ();
 sg13g2_decap_8 FILLER_51_198 ();
 sg13g2_fill_1 FILLER_51_205 ();
 sg13g2_decap_8 FILLER_51_235 ();
 sg13g2_decap_8 FILLER_51_242 ();
 sg13g2_decap_4 FILLER_51_249 ();
 sg13g2_fill_2 FILLER_51_253 ();
 sg13g2_decap_8 FILLER_51_310 ();
 sg13g2_decap_8 FILLER_51_356 ();
 sg13g2_decap_8 FILLER_51_363 ();
 sg13g2_decap_8 FILLER_51_370 ();
 sg13g2_decap_4 FILLER_51_377 ();
 sg13g2_fill_1 FILLER_51_381 ();
 sg13g2_fill_1 FILLER_51_399 ();
 sg13g2_fill_2 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_51_431 ();
 sg13g2_decap_8 FILLER_51_438 ();
 sg13g2_decap_8 FILLER_51_445 ();
 sg13g2_decap_8 FILLER_51_452 ();
 sg13g2_decap_4 FILLER_51_459 ();
 sg13g2_fill_2 FILLER_51_468 ();
 sg13g2_fill_1 FILLER_51_470 ();
 sg13g2_decap_8 FILLER_51_497 ();
 sg13g2_decap_4 FILLER_51_504 ();
 sg13g2_fill_1 FILLER_51_508 ();
 sg13g2_decap_8 FILLER_51_586 ();
 sg13g2_fill_2 FILLER_51_671 ();
 sg13g2_fill_1 FILLER_51_673 ();
 sg13g2_fill_2 FILLER_51_679 ();
 sg13g2_decap_8 FILLER_51_694 ();
 sg13g2_decap_4 FILLER_51_701 ();
 sg13g2_fill_2 FILLER_51_705 ();
 sg13g2_fill_2 FILLER_51_733 ();
 sg13g2_fill_1 FILLER_51_735 ();
 sg13g2_decap_4 FILLER_51_762 ();
 sg13g2_decap_4 FILLER_51_799 ();
 sg13g2_fill_2 FILLER_51_813 ();
 sg13g2_fill_2 FILLER_51_820 ();
 sg13g2_decap_8 FILLER_51_830 ();
 sg13g2_decap_8 FILLER_51_837 ();
 sg13g2_decap_8 FILLER_51_844 ();
 sg13g2_fill_2 FILLER_51_851 ();
 sg13g2_decap_8 FILLER_51_883 ();
 sg13g2_fill_1 FILLER_51_890 ();
 sg13g2_fill_1 FILLER_51_917 ();
 sg13g2_decap_8 FILLER_51_947 ();
 sg13g2_fill_2 FILLER_51_954 ();
 sg13g2_fill_1 FILLER_51_956 ();
 sg13g2_decap_4 FILLER_51_960 ();
 sg13g2_fill_1 FILLER_51_964 ();
 sg13g2_fill_2 FILLER_51_973 ();
 sg13g2_fill_1 FILLER_51_975 ();
 sg13g2_fill_2 FILLER_51_1028 ();
 sg13g2_decap_4 FILLER_51_1056 ();
 sg13g2_fill_1 FILLER_51_1072 ();
 sg13g2_decap_8 FILLER_51_1088 ();
 sg13g2_fill_2 FILLER_51_1095 ();
 sg13g2_fill_2 FILLER_51_1113 ();
 sg13g2_fill_1 FILLER_51_1115 ();
 sg13g2_decap_4 FILLER_51_1137 ();
 sg13g2_fill_1 FILLER_51_1141 ();
 sg13g2_decap_8 FILLER_51_1147 ();
 sg13g2_decap_4 FILLER_51_1154 ();
 sg13g2_fill_2 FILLER_51_1158 ();
 sg13g2_decap_8 FILLER_51_1198 ();
 sg13g2_decap_8 FILLER_51_1205 ();
 sg13g2_decap_8 FILLER_51_1212 ();
 sg13g2_decap_4 FILLER_51_1219 ();
 sg13g2_fill_2 FILLER_51_1223 ();
 sg13g2_decap_8 FILLER_51_1261 ();
 sg13g2_decap_4 FILLER_51_1268 ();
 sg13g2_fill_1 FILLER_51_1272 ();
 sg13g2_fill_2 FILLER_51_1310 ();
 sg13g2_fill_1 FILLER_51_1312 ();
 sg13g2_decap_4 FILLER_51_1389 ();
 sg13g2_fill_1 FILLER_51_1399 ();
 sg13g2_fill_1 FILLER_51_1417 ();
 sg13g2_decap_8 FILLER_51_1423 ();
 sg13g2_decap_8 FILLER_51_1430 ();
 sg13g2_fill_1 FILLER_51_1437 ();
 sg13g2_fill_2 FILLER_51_1451 ();
 sg13g2_fill_1 FILLER_51_1453 ();
 sg13g2_decap_8 FILLER_51_1470 ();
 sg13g2_decap_8 FILLER_51_1477 ();
 sg13g2_decap_8 FILLER_51_1484 ();
 sg13g2_decap_8 FILLER_51_1491 ();
 sg13g2_decap_8 FILLER_51_1498 ();
 sg13g2_decap_4 FILLER_51_1505 ();
 sg13g2_fill_2 FILLER_51_1509 ();
 sg13g2_fill_1 FILLER_51_1567 ();
 sg13g2_fill_2 FILLER_51_1580 ();
 sg13g2_fill_1 FILLER_51_1582 ();
 sg13g2_fill_1 FILLER_51_1587 ();
 sg13g2_fill_1 FILLER_51_1592 ();
 sg13g2_fill_1 FILLER_51_1601 ();
 sg13g2_decap_8 FILLER_51_1607 ();
 sg13g2_decap_8 FILLER_51_1614 ();
 sg13g2_decap_8 FILLER_51_1621 ();
 sg13g2_fill_2 FILLER_51_1628 ();
 sg13g2_fill_1 FILLER_51_1630 ();
 sg13g2_decap_8 FILLER_51_1635 ();
 sg13g2_decap_8 FILLER_51_1642 ();
 sg13g2_decap_8 FILLER_51_1649 ();
 sg13g2_decap_4 FILLER_51_1656 ();
 sg13g2_fill_1 FILLER_51_1660 ();
 sg13g2_fill_2 FILLER_51_1687 ();
 sg13g2_decap_8 FILLER_51_1736 ();
 sg13g2_fill_1 FILLER_51_1743 ();
 sg13g2_fill_2 FILLER_51_1796 ();
 sg13g2_decap_4 FILLER_51_1806 ();
 sg13g2_fill_2 FILLER_51_1823 ();
 sg13g2_fill_2 FILLER_51_1833 ();
 sg13g2_decap_8 FILLER_51_1843 ();
 sg13g2_decap_4 FILLER_51_1850 ();
 sg13g2_fill_2 FILLER_51_1854 ();
 sg13g2_fill_2 FILLER_51_1882 ();
 sg13g2_fill_2 FILLER_51_1888 ();
 sg13g2_fill_2 FILLER_51_1895 ();
 sg13g2_decap_8 FILLER_51_1928 ();
 sg13g2_decap_8 FILLER_51_1935 ();
 sg13g2_decap_8 FILLER_51_1942 ();
 sg13g2_fill_2 FILLER_51_1949 ();
 sg13g2_fill_1 FILLER_51_1951 ();
 sg13g2_fill_1 FILLER_51_1964 ();
 sg13g2_fill_2 FILLER_51_2000 ();
 sg13g2_fill_1 FILLER_51_2002 ();
 sg13g2_fill_2 FILLER_51_2008 ();
 sg13g2_fill_1 FILLER_51_2024 ();
 sg13g2_decap_8 FILLER_51_2051 ();
 sg13g2_decap_8 FILLER_51_2058 ();
 sg13g2_fill_2 FILLER_51_2065 ();
 sg13g2_fill_1 FILLER_51_2067 ();
 sg13g2_decap_4 FILLER_51_2112 ();
 sg13g2_fill_2 FILLER_51_2129 ();
 sg13g2_decap_4 FILLER_51_2157 ();
 sg13g2_decap_4 FILLER_51_2169 ();
 sg13g2_fill_1 FILLER_51_2173 ();
 sg13g2_decap_4 FILLER_51_2179 ();
 sg13g2_fill_1 FILLER_51_2183 ();
 sg13g2_fill_2 FILLER_51_2195 ();
 sg13g2_fill_1 FILLER_51_2197 ();
 sg13g2_decap_8 FILLER_51_2392 ();
 sg13g2_decap_8 FILLER_51_2399 ();
 sg13g2_decap_8 FILLER_51_2414 ();
 sg13g2_fill_2 FILLER_51_2421 ();
 sg13g2_decap_8 FILLER_51_2428 ();
 sg13g2_decap_8 FILLER_51_2435 ();
 sg13g2_decap_4 FILLER_51_2442 ();
 sg13g2_fill_2 FILLER_51_2446 ();
 sg13g2_decap_4 FILLER_51_2506 ();
 sg13g2_fill_1 FILLER_51_2510 ();
 sg13g2_decap_8 FILLER_51_2519 ();
 sg13g2_decap_8 FILLER_51_2526 ();
 sg13g2_decap_8 FILLER_51_2533 ();
 sg13g2_decap_8 FILLER_51_2540 ();
 sg13g2_decap_8 FILLER_51_2547 ();
 sg13g2_decap_8 FILLER_51_2554 ();
 sg13g2_fill_1 FILLER_51_2561 ();
 sg13g2_decap_8 FILLER_51_2588 ();
 sg13g2_decap_8 FILLER_51_2595 ();
 sg13g2_decap_8 FILLER_51_2602 ();
 sg13g2_fill_2 FILLER_51_2609 ();
 sg13g2_fill_1 FILLER_51_2611 ();
 sg13g2_decap_8 FILLER_51_2646 ();
 sg13g2_decap_8 FILLER_51_2653 ();
 sg13g2_decap_8 FILLER_51_2660 ();
 sg13g2_decap_8 FILLER_51_2667 ();
 sg13g2_decap_8 FILLER_51_2674 ();
 sg13g2_decap_8 FILLER_51_2681 ();
 sg13g2_fill_2 FILLER_51_2688 ();
 sg13g2_fill_1 FILLER_51_2690 ();
 sg13g2_decap_8 FILLER_51_2695 ();
 sg13g2_fill_1 FILLER_51_2702 ();
 sg13g2_fill_2 FILLER_51_2706 ();
 sg13g2_fill_1 FILLER_51_2708 ();
 sg13g2_decap_4 FILLER_51_2829 ();
 sg13g2_fill_2 FILLER_51_2833 ();
 sg13g2_decap_8 FILLER_51_2861 ();
 sg13g2_decap_8 FILLER_51_2868 ();
 sg13g2_decap_8 FILLER_51_2915 ();
 sg13g2_decap_8 FILLER_51_2922 ();
 sg13g2_decap_8 FILLER_51_2929 ();
 sg13g2_decap_8 FILLER_51_2936 ();
 sg13g2_decap_8 FILLER_51_2975 ();
 sg13g2_decap_4 FILLER_51_2982 ();
 sg13g2_fill_1 FILLER_51_2986 ();
 sg13g2_decap_8 FILLER_51_3021 ();
 sg13g2_decap_8 FILLER_51_3028 ();
 sg13g2_decap_8 FILLER_51_3035 ();
 sg13g2_decap_8 FILLER_51_3042 ();
 sg13g2_decap_8 FILLER_51_3049 ();
 sg13g2_decap_8 FILLER_51_3056 ();
 sg13g2_decap_8 FILLER_51_3063 ();
 sg13g2_decap_8 FILLER_51_3070 ();
 sg13g2_decap_8 FILLER_51_3077 ();
 sg13g2_decap_8 FILLER_51_3084 ();
 sg13g2_decap_8 FILLER_51_3091 ();
 sg13g2_decap_8 FILLER_51_3098 ();
 sg13g2_decap_8 FILLER_51_3105 ();
 sg13g2_decap_8 FILLER_51_3112 ();
 sg13g2_decap_8 FILLER_51_3119 ();
 sg13g2_decap_8 FILLER_51_3126 ();
 sg13g2_decap_8 FILLER_51_3133 ();
 sg13g2_decap_8 FILLER_51_3140 ();
 sg13g2_decap_8 FILLER_51_3147 ();
 sg13g2_decap_8 FILLER_51_3154 ();
 sg13g2_decap_8 FILLER_51_3161 ();
 sg13g2_decap_8 FILLER_51_3168 ();
 sg13g2_decap_8 FILLER_51_3175 ();
 sg13g2_decap_8 FILLER_51_3182 ();
 sg13g2_decap_8 FILLER_51_3189 ();
 sg13g2_decap_8 FILLER_51_3196 ();
 sg13g2_decap_8 FILLER_51_3203 ();
 sg13g2_decap_8 FILLER_51_3210 ();
 sg13g2_decap_8 FILLER_51_3217 ();
 sg13g2_decap_8 FILLER_51_3224 ();
 sg13g2_decap_8 FILLER_51_3231 ();
 sg13g2_decap_8 FILLER_51_3238 ();
 sg13g2_decap_8 FILLER_51_3245 ();
 sg13g2_decap_8 FILLER_51_3252 ();
 sg13g2_decap_8 FILLER_51_3259 ();
 sg13g2_decap_8 FILLER_51_3266 ();
 sg13g2_decap_8 FILLER_51_3273 ();
 sg13g2_decap_8 FILLER_51_3280 ();
 sg13g2_decap_8 FILLER_51_3287 ();
 sg13g2_decap_8 FILLER_51_3294 ();
 sg13g2_decap_8 FILLER_51_3301 ();
 sg13g2_decap_8 FILLER_51_3308 ();
 sg13g2_decap_8 FILLER_51_3315 ();
 sg13g2_decap_8 FILLER_51_3322 ();
 sg13g2_decap_8 FILLER_51_3329 ();
 sg13g2_decap_8 FILLER_51_3336 ();
 sg13g2_decap_8 FILLER_51_3343 ();
 sg13g2_decap_8 FILLER_51_3350 ();
 sg13g2_decap_8 FILLER_51_3357 ();
 sg13g2_decap_8 FILLER_51_3364 ();
 sg13g2_decap_8 FILLER_51_3371 ();
 sg13g2_decap_8 FILLER_51_3378 ();
 sg13g2_decap_8 FILLER_51_3385 ();
 sg13g2_decap_8 FILLER_51_3392 ();
 sg13g2_decap_8 FILLER_51_3399 ();
 sg13g2_decap_8 FILLER_51_3406 ();
 sg13g2_decap_8 FILLER_51_3413 ();
 sg13g2_decap_8 FILLER_51_3420 ();
 sg13g2_decap_8 FILLER_51_3427 ();
 sg13g2_decap_8 FILLER_51_3434 ();
 sg13g2_decap_8 FILLER_51_3441 ();
 sg13g2_decap_8 FILLER_51_3448 ();
 sg13g2_decap_8 FILLER_51_3455 ();
 sg13g2_decap_8 FILLER_51_3462 ();
 sg13g2_decap_8 FILLER_51_3469 ();
 sg13g2_decap_8 FILLER_51_3476 ();
 sg13g2_decap_8 FILLER_51_3483 ();
 sg13g2_decap_8 FILLER_51_3490 ();
 sg13g2_decap_8 FILLER_51_3497 ();
 sg13g2_decap_8 FILLER_51_3504 ();
 sg13g2_decap_8 FILLER_51_3511 ();
 sg13g2_decap_8 FILLER_51_3518 ();
 sg13g2_decap_8 FILLER_51_3525 ();
 sg13g2_decap_8 FILLER_51_3532 ();
 sg13g2_decap_8 FILLER_51_3539 ();
 sg13g2_decap_8 FILLER_51_3546 ();
 sg13g2_decap_8 FILLER_51_3553 ();
 sg13g2_decap_8 FILLER_51_3560 ();
 sg13g2_decap_8 FILLER_51_3567 ();
 sg13g2_decap_4 FILLER_51_3574 ();
 sg13g2_fill_2 FILLER_51_3578 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_4 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_150 ();
 sg13g2_decap_8 FILLER_52_157 ();
 sg13g2_decap_8 FILLER_52_164 ();
 sg13g2_decap_8 FILLER_52_171 ();
 sg13g2_decap_8 FILLER_52_178 ();
 sg13g2_decap_8 FILLER_52_185 ();
 sg13g2_decap_8 FILLER_52_192 ();
 sg13g2_decap_8 FILLER_52_199 ();
 sg13g2_decap_8 FILLER_52_206 ();
 sg13g2_fill_1 FILLER_52_213 ();
 sg13g2_decap_8 FILLER_52_217 ();
 sg13g2_decap_8 FILLER_52_224 ();
 sg13g2_decap_8 FILLER_52_231 ();
 sg13g2_decap_8 FILLER_52_238 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_decap_8 FILLER_52_252 ();
 sg13g2_decap_8 FILLER_52_259 ();
 sg13g2_decap_4 FILLER_52_266 ();
 sg13g2_decap_4 FILLER_52_273 ();
 sg13g2_fill_1 FILLER_52_277 ();
 sg13g2_fill_1 FILLER_52_283 ();
 sg13g2_decap_8 FILLER_52_310 ();
 sg13g2_fill_2 FILLER_52_317 ();
 sg13g2_decap_8 FILLER_52_363 ();
 sg13g2_fill_2 FILLER_52_370 ();
 sg13g2_fill_1 FILLER_52_372 ();
 sg13g2_fill_1 FILLER_52_395 ();
 sg13g2_decap_8 FILLER_52_401 ();
 sg13g2_decap_8 FILLER_52_408 ();
 sg13g2_fill_2 FILLER_52_415 ();
 sg13g2_fill_1 FILLER_52_417 ();
 sg13g2_decap_8 FILLER_52_425 ();
 sg13g2_decap_4 FILLER_52_432 ();
 sg13g2_fill_1 FILLER_52_436 ();
 sg13g2_fill_2 FILLER_52_440 ();
 sg13g2_decap_4 FILLER_52_455 ();
 sg13g2_decap_8 FILLER_52_492 ();
 sg13g2_decap_4 FILLER_52_499 ();
 sg13g2_fill_2 FILLER_52_503 ();
 sg13g2_decap_8 FILLER_52_581 ();
 sg13g2_decap_8 FILLER_52_588 ();
 sg13g2_decap_8 FILLER_52_595 ();
 sg13g2_decap_8 FILLER_52_602 ();
 sg13g2_fill_2 FILLER_52_643 ();
 sg13g2_fill_1 FILLER_52_645 ();
 sg13g2_fill_2 FILLER_52_649 ();
 sg13g2_fill_1 FILLER_52_651 ();
 sg13g2_decap_4 FILLER_52_665 ();
 sg13g2_fill_1 FILLER_52_693 ();
 sg13g2_decap_8 FILLER_52_699 ();
 sg13g2_fill_2 FILLER_52_706 ();
 sg13g2_fill_1 FILLER_52_717 ();
 sg13g2_fill_1 FILLER_52_722 ();
 sg13g2_fill_2 FILLER_52_757 ();
 sg13g2_fill_2 FILLER_52_814 ();
 sg13g2_fill_1 FILLER_52_829 ();
 sg13g2_decap_8 FILLER_52_843 ();
 sg13g2_decap_8 FILLER_52_850 ();
 sg13g2_decap_4 FILLER_52_887 ();
 sg13g2_fill_1 FILLER_52_891 ();
 sg13g2_fill_1 FILLER_52_902 ();
 sg13g2_decap_8 FILLER_52_942 ();
 sg13g2_fill_2 FILLER_52_949 ();
 sg13g2_fill_1 FILLER_52_1087 ();
 sg13g2_decap_8 FILLER_52_1136 ();
 sg13g2_fill_2 FILLER_52_1143 ();
 sg13g2_fill_1 FILLER_52_1145 ();
 sg13g2_decap_4 FILLER_52_1209 ();
 sg13g2_fill_1 FILLER_52_1213 ();
 sg13g2_decap_8 FILLER_52_1274 ();
 sg13g2_decap_8 FILLER_52_1281 ();
 sg13g2_fill_2 FILLER_52_1288 ();
 sg13g2_decap_8 FILLER_52_1298 ();
 sg13g2_decap_8 FILLER_52_1305 ();
 sg13g2_fill_1 FILLER_52_1312 ();
 sg13g2_decap_8 FILLER_52_1369 ();
 sg13g2_decap_8 FILLER_52_1376 ();
 sg13g2_decap_4 FILLER_52_1383 ();
 sg13g2_fill_2 FILLER_52_1431 ();
 sg13g2_fill_1 FILLER_52_1433 ();
 sg13g2_fill_2 FILLER_52_1458 ();
 sg13g2_fill_1 FILLER_52_1460 ();
 sg13g2_decap_8 FILLER_52_1499 ();
 sg13g2_fill_1 FILLER_52_1515 ();
 sg13g2_fill_2 FILLER_52_1550 ();
 sg13g2_decap_8 FILLER_52_1570 ();
 sg13g2_decap_8 FILLER_52_1587 ();
 sg13g2_fill_2 FILLER_52_1594 ();
 sg13g2_decap_8 FILLER_52_1630 ();
 sg13g2_decap_8 FILLER_52_1637 ();
 sg13g2_fill_2 FILLER_52_1644 ();
 sg13g2_fill_1 FILLER_52_1646 ();
 sg13g2_decap_8 FILLER_52_1725 ();
 sg13g2_decap_8 FILLER_52_1732 ();
 sg13g2_fill_1 FILLER_52_1739 ();
 sg13g2_fill_2 FILLER_52_1808 ();
 sg13g2_fill_2 FILLER_52_1844 ();
 sg13g2_fill_1 FILLER_52_1846 ();
 sg13g2_decap_8 FILLER_52_1873 ();
 sg13g2_decap_8 FILLER_52_1880 ();
 sg13g2_decap_8 FILLER_52_1887 ();
 sg13g2_decap_8 FILLER_52_1894 ();
 sg13g2_fill_2 FILLER_52_1906 ();
 sg13g2_decap_8 FILLER_52_1934 ();
 sg13g2_decap_8 FILLER_52_1941 ();
 sg13g2_fill_2 FILLER_52_1948 ();
 sg13g2_fill_1 FILLER_52_1950 ();
 sg13g2_fill_1 FILLER_52_1957 ();
 sg13g2_fill_1 FILLER_52_1963 ();
 sg13g2_decap_4 FILLER_52_1976 ();
 sg13g2_fill_2 FILLER_52_1980 ();
 sg13g2_decap_8 FILLER_52_1988 ();
 sg13g2_decap_4 FILLER_52_1995 ();
 sg13g2_decap_8 FILLER_52_2057 ();
 sg13g2_decap_4 FILLER_52_2064 ();
 sg13g2_fill_2 FILLER_52_2068 ();
 sg13g2_fill_2 FILLER_52_2090 ();
 sg13g2_fill_2 FILLER_52_2108 ();
 sg13g2_fill_1 FILLER_52_2110 ();
 sg13g2_fill_1 FILLER_52_2122 ();
 sg13g2_decap_8 FILLER_52_2165 ();
 sg13g2_decap_8 FILLER_52_2172 ();
 sg13g2_decap_8 FILLER_52_2179 ();
 sg13g2_fill_2 FILLER_52_2186 ();
 sg13g2_fill_1 FILLER_52_2188 ();
 sg13g2_fill_1 FILLER_52_2195 ();
 sg13g2_fill_2 FILLER_52_2202 ();
 sg13g2_decap_8 FILLER_52_2282 ();
 sg13g2_decap_8 FILLER_52_2289 ();
 sg13g2_decap_8 FILLER_52_2296 ();
 sg13g2_decap_8 FILLER_52_2303 ();
 sg13g2_decap_8 FILLER_52_2310 ();
 sg13g2_fill_2 FILLER_52_2317 ();
 sg13g2_fill_1 FILLER_52_2319 ();
 sg13g2_decap_4 FILLER_52_2398 ();
 sg13g2_fill_1 FILLER_52_2402 ();
 sg13g2_decap_4 FILLER_52_2419 ();
 sg13g2_fill_2 FILLER_52_2423 ();
 sg13g2_fill_1 FILLER_52_2430 ();
 sg13g2_decap_8 FILLER_52_2439 ();
 sg13g2_decap_8 FILLER_52_2446 ();
 sg13g2_decap_8 FILLER_52_2453 ();
 sg13g2_fill_1 FILLER_52_2460 ();
 sg13g2_decap_8 FILLER_52_2499 ();
 sg13g2_decap_8 FILLER_52_2506 ();
 sg13g2_decap_8 FILLER_52_2513 ();
 sg13g2_decap_4 FILLER_52_2520 ();
 sg13g2_decap_8 FILLER_52_2564 ();
 sg13g2_decap_8 FILLER_52_2571 ();
 sg13g2_decap_8 FILLER_52_2578 ();
 sg13g2_fill_2 FILLER_52_2585 ();
 sg13g2_fill_1 FILLER_52_2587 ();
 sg13g2_fill_2 FILLER_52_2604 ();
 sg13g2_fill_1 FILLER_52_2606 ();
 sg13g2_fill_2 FILLER_52_2633 ();
 sg13g2_fill_1 FILLER_52_2635 ();
 sg13g2_decap_8 FILLER_52_2662 ();
 sg13g2_fill_1 FILLER_52_2695 ();
 sg13g2_decap_8 FILLER_52_2701 ();
 sg13g2_decap_8 FILLER_52_2708 ();
 sg13g2_fill_1 FILLER_52_2715 ();
 sg13g2_fill_1 FILLER_52_2720 ();
 sg13g2_fill_1 FILLER_52_2726 ();
 sg13g2_decap_4 FILLER_52_2758 ();
 sg13g2_decap_8 FILLER_52_2801 ();
 sg13g2_decap_8 FILLER_52_2808 ();
 sg13g2_fill_1 FILLER_52_2815 ();
 sg13g2_decap_8 FILLER_52_2842 ();
 sg13g2_decap_8 FILLER_52_2849 ();
 sg13g2_decap_8 FILLER_52_2856 ();
 sg13g2_decap_8 FILLER_52_2863 ();
 sg13g2_decap_4 FILLER_52_2870 ();
 sg13g2_fill_1 FILLER_52_2874 ();
 sg13g2_decap_8 FILLER_52_2909 ();
 sg13g2_decap_8 FILLER_52_2916 ();
 sg13g2_decap_8 FILLER_52_2923 ();
 sg13g2_decap_4 FILLER_52_2930 ();
 sg13g2_fill_1 FILLER_52_2934 ();
 sg13g2_decap_4 FILLER_52_2948 ();
 sg13g2_fill_1 FILLER_52_2952 ();
 sg13g2_decap_8 FILLER_52_2979 ();
 sg13g2_decap_8 FILLER_52_2986 ();
 sg13g2_decap_8 FILLER_52_2993 ();
 sg13g2_fill_1 FILLER_52_3000 ();
 sg13g2_decap_8 FILLER_52_3027 ();
 sg13g2_decap_8 FILLER_52_3034 ();
 sg13g2_decap_8 FILLER_52_3041 ();
 sg13g2_decap_8 FILLER_52_3048 ();
 sg13g2_decap_8 FILLER_52_3055 ();
 sg13g2_decap_8 FILLER_52_3062 ();
 sg13g2_decap_8 FILLER_52_3069 ();
 sg13g2_decap_8 FILLER_52_3076 ();
 sg13g2_decap_8 FILLER_52_3083 ();
 sg13g2_decap_8 FILLER_52_3090 ();
 sg13g2_decap_8 FILLER_52_3097 ();
 sg13g2_decap_8 FILLER_52_3104 ();
 sg13g2_decap_8 FILLER_52_3111 ();
 sg13g2_decap_8 FILLER_52_3118 ();
 sg13g2_decap_8 FILLER_52_3125 ();
 sg13g2_decap_8 FILLER_52_3132 ();
 sg13g2_decap_8 FILLER_52_3139 ();
 sg13g2_decap_8 FILLER_52_3146 ();
 sg13g2_decap_8 FILLER_52_3153 ();
 sg13g2_decap_8 FILLER_52_3160 ();
 sg13g2_decap_8 FILLER_52_3167 ();
 sg13g2_decap_8 FILLER_52_3174 ();
 sg13g2_decap_8 FILLER_52_3181 ();
 sg13g2_decap_8 FILLER_52_3188 ();
 sg13g2_decap_8 FILLER_52_3195 ();
 sg13g2_decap_8 FILLER_52_3202 ();
 sg13g2_decap_8 FILLER_52_3209 ();
 sg13g2_decap_8 FILLER_52_3216 ();
 sg13g2_decap_8 FILLER_52_3223 ();
 sg13g2_decap_8 FILLER_52_3230 ();
 sg13g2_decap_8 FILLER_52_3237 ();
 sg13g2_decap_8 FILLER_52_3244 ();
 sg13g2_decap_8 FILLER_52_3251 ();
 sg13g2_decap_8 FILLER_52_3258 ();
 sg13g2_decap_8 FILLER_52_3265 ();
 sg13g2_decap_8 FILLER_52_3272 ();
 sg13g2_decap_8 FILLER_52_3279 ();
 sg13g2_decap_8 FILLER_52_3286 ();
 sg13g2_decap_8 FILLER_52_3293 ();
 sg13g2_decap_8 FILLER_52_3300 ();
 sg13g2_decap_8 FILLER_52_3307 ();
 sg13g2_decap_8 FILLER_52_3314 ();
 sg13g2_decap_8 FILLER_52_3321 ();
 sg13g2_decap_8 FILLER_52_3328 ();
 sg13g2_decap_8 FILLER_52_3335 ();
 sg13g2_decap_8 FILLER_52_3342 ();
 sg13g2_decap_8 FILLER_52_3349 ();
 sg13g2_decap_8 FILLER_52_3356 ();
 sg13g2_decap_8 FILLER_52_3363 ();
 sg13g2_decap_8 FILLER_52_3370 ();
 sg13g2_decap_8 FILLER_52_3377 ();
 sg13g2_decap_8 FILLER_52_3384 ();
 sg13g2_decap_8 FILLER_52_3391 ();
 sg13g2_decap_8 FILLER_52_3398 ();
 sg13g2_decap_8 FILLER_52_3405 ();
 sg13g2_decap_8 FILLER_52_3412 ();
 sg13g2_decap_8 FILLER_52_3419 ();
 sg13g2_decap_8 FILLER_52_3426 ();
 sg13g2_decap_8 FILLER_52_3433 ();
 sg13g2_decap_8 FILLER_52_3440 ();
 sg13g2_decap_8 FILLER_52_3447 ();
 sg13g2_decap_8 FILLER_52_3454 ();
 sg13g2_decap_8 FILLER_52_3461 ();
 sg13g2_decap_8 FILLER_52_3468 ();
 sg13g2_decap_8 FILLER_52_3475 ();
 sg13g2_decap_8 FILLER_52_3482 ();
 sg13g2_decap_8 FILLER_52_3489 ();
 sg13g2_decap_8 FILLER_52_3496 ();
 sg13g2_decap_8 FILLER_52_3503 ();
 sg13g2_decap_8 FILLER_52_3510 ();
 sg13g2_decap_8 FILLER_52_3517 ();
 sg13g2_decap_8 FILLER_52_3524 ();
 sg13g2_decap_8 FILLER_52_3531 ();
 sg13g2_decap_8 FILLER_52_3538 ();
 sg13g2_decap_8 FILLER_52_3545 ();
 sg13g2_decap_8 FILLER_52_3552 ();
 sg13g2_decap_8 FILLER_52_3559 ();
 sg13g2_decap_8 FILLER_52_3566 ();
 sg13g2_decap_8 FILLER_52_3573 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_4 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_134 ();
 sg13g2_decap_8 FILLER_53_141 ();
 sg13g2_decap_8 FILLER_53_148 ();
 sg13g2_decap_8 FILLER_53_155 ();
 sg13g2_decap_8 FILLER_53_162 ();
 sg13g2_decap_8 FILLER_53_169 ();
 sg13g2_decap_8 FILLER_53_176 ();
 sg13g2_decap_8 FILLER_53_183 ();
 sg13g2_decap_8 FILLER_53_190 ();
 sg13g2_decap_8 FILLER_53_197 ();
 sg13g2_decap_8 FILLER_53_204 ();
 sg13g2_decap_8 FILLER_53_211 ();
 sg13g2_decap_8 FILLER_53_218 ();
 sg13g2_decap_8 FILLER_53_225 ();
 sg13g2_decap_8 FILLER_53_232 ();
 sg13g2_decap_8 FILLER_53_239 ();
 sg13g2_decap_8 FILLER_53_246 ();
 sg13g2_decap_8 FILLER_53_253 ();
 sg13g2_decap_8 FILLER_53_260 ();
 sg13g2_fill_2 FILLER_53_267 ();
 sg13g2_decap_8 FILLER_53_300 ();
 sg13g2_decap_8 FILLER_53_307 ();
 sg13g2_decap_8 FILLER_53_314 ();
 sg13g2_decap_8 FILLER_53_321 ();
 sg13g2_fill_1 FILLER_53_328 ();
 sg13g2_fill_1 FILLER_53_342 ();
 sg13g2_decap_4 FILLER_53_363 ();
 sg13g2_fill_2 FILLER_53_367 ();
 sg13g2_fill_2 FILLER_53_411 ();
 sg13g2_decap_8 FILLER_53_416 ();
 sg13g2_decap_4 FILLER_53_423 ();
 sg13g2_decap_8 FILLER_53_500 ();
 sg13g2_fill_1 FILLER_53_507 ();
 sg13g2_decap_8 FILLER_53_572 ();
 sg13g2_decap_8 FILLER_53_579 ();
 sg13g2_decap_8 FILLER_53_586 ();
 sg13g2_fill_2 FILLER_53_593 ();
 sg13g2_fill_1 FILLER_53_595 ();
 sg13g2_decap_8 FILLER_53_601 ();
 sg13g2_fill_2 FILLER_53_608 ();
 sg13g2_fill_1 FILLER_53_610 ();
 sg13g2_decap_4 FILLER_53_616 ();
 sg13g2_fill_1 FILLER_53_620 ();
 sg13g2_decap_8 FILLER_53_629 ();
 sg13g2_decap_4 FILLER_53_636 ();
 sg13g2_fill_1 FILLER_53_640 ();
 sg13g2_decap_4 FILLER_53_667 ();
 sg13g2_fill_2 FILLER_53_710 ();
 sg13g2_decap_8 FILLER_53_720 ();
 sg13g2_fill_1 FILLER_53_727 ();
 sg13g2_decap_8 FILLER_53_758 ();
 sg13g2_fill_2 FILLER_53_765 ();
 sg13g2_fill_2 FILLER_53_797 ();
 sg13g2_fill_1 FILLER_53_799 ();
 sg13g2_fill_2 FILLER_53_837 ();
 sg13g2_decap_8 FILLER_53_852 ();
 sg13g2_fill_1 FILLER_53_859 ();
 sg13g2_decap_8 FILLER_53_938 ();
 sg13g2_decap_4 FILLER_53_945 ();
 sg13g2_fill_1 FILLER_53_949 ();
 sg13g2_decap_8 FILLER_53_976 ();
 sg13g2_decap_8 FILLER_53_983 ();
 sg13g2_decap_8 FILLER_53_990 ();
 sg13g2_decap_4 FILLER_53_997 ();
 sg13g2_decap_8 FILLER_53_1007 ();
 sg13g2_decap_8 FILLER_53_1014 ();
 sg13g2_decap_8 FILLER_53_1047 ();
 sg13g2_decap_4 FILLER_53_1054 ();
 sg13g2_fill_2 FILLER_53_1090 ();
 sg13g2_fill_1 FILLER_53_1092 ();
 sg13g2_fill_2 FILLER_53_1221 ();
 sg13g2_decap_4 FILLER_53_1255 ();
 sg13g2_decap_8 FILLER_53_1283 ();
 sg13g2_decap_8 FILLER_53_1290 ();
 sg13g2_decap_4 FILLER_53_1301 ();
 sg13g2_fill_1 FILLER_53_1305 ();
 sg13g2_decap_8 FILLER_53_1336 ();
 sg13g2_fill_2 FILLER_53_1343 ();
 sg13g2_fill_1 FILLER_53_1345 ();
 sg13g2_decap_8 FILLER_53_1360 ();
 sg13g2_decap_8 FILLER_53_1367 ();
 sg13g2_decap_8 FILLER_53_1374 ();
 sg13g2_fill_2 FILLER_53_1381 ();
 sg13g2_decap_4 FILLER_53_1387 ();
 sg13g2_fill_2 FILLER_53_1400 ();
 sg13g2_fill_2 FILLER_53_1411 ();
 sg13g2_fill_1 FILLER_53_1413 ();
 sg13g2_fill_2 FILLER_53_1419 ();
 sg13g2_fill_1 FILLER_53_1421 ();
 sg13g2_fill_2 FILLER_53_1440 ();
 sg13g2_fill_1 FILLER_53_1447 ();
 sg13g2_fill_1 FILLER_53_1463 ();
 sg13g2_fill_2 FILLER_53_1469 ();
 sg13g2_fill_2 FILLER_53_1476 ();
 sg13g2_fill_1 FILLER_53_1504 ();
 sg13g2_fill_2 FILLER_53_1531 ();
 sg13g2_fill_2 FILLER_53_1541 ();
 sg13g2_decap_8 FILLER_53_1569 ();
 sg13g2_decap_8 FILLER_53_1576 ();
 sg13g2_decap_8 FILLER_53_1583 ();
 sg13g2_decap_4 FILLER_53_1590 ();
 sg13g2_fill_1 FILLER_53_1594 ();
 sg13g2_decap_8 FILLER_53_1636 ();
 sg13g2_decap_8 FILLER_53_1695 ();
 sg13g2_fill_1 FILLER_53_1702 ();
 sg13g2_decap_8 FILLER_53_1729 ();
 sg13g2_decap_8 FILLER_53_1736 ();
 sg13g2_decap_4 FILLER_53_1743 ();
 sg13g2_fill_2 FILLER_53_1747 ();
 sg13g2_fill_2 FILLER_53_1797 ();
 sg13g2_fill_1 FILLER_53_1799 ();
 sg13g2_fill_2 FILLER_53_1816 ();
 sg13g2_decap_4 FILLER_53_1842 ();
 sg13g2_fill_2 FILLER_53_1846 ();
 sg13g2_decap_8 FILLER_53_1892 ();
 sg13g2_decap_8 FILLER_53_1899 ();
 sg13g2_decap_4 FILLER_53_1906 ();
 sg13g2_fill_2 FILLER_53_1910 ();
 sg13g2_decap_8 FILLER_53_1915 ();
 sg13g2_decap_8 FILLER_53_1922 ();
 sg13g2_decap_8 FILLER_53_1929 ();
 sg13g2_decap_8 FILLER_53_1936 ();
 sg13g2_fill_2 FILLER_53_1943 ();
 sg13g2_decap_8 FILLER_53_1997 ();
 sg13g2_fill_2 FILLER_53_2004 ();
 sg13g2_fill_1 FILLER_53_2006 ();
 sg13g2_decap_8 FILLER_53_2065 ();
 sg13g2_fill_2 FILLER_53_2072 ();
 sg13g2_fill_1 FILLER_53_2074 ();
 sg13g2_decap_8 FILLER_53_2083 ();
 sg13g2_decap_8 FILLER_53_2090 ();
 sg13g2_fill_2 FILLER_53_2097 ();
 sg13g2_fill_1 FILLER_53_2099 ();
 sg13g2_fill_2 FILLER_53_2137 ();
 sg13g2_fill_1 FILLER_53_2139 ();
 sg13g2_decap_4 FILLER_53_2192 ();
 sg13g2_fill_2 FILLER_53_2196 ();
 sg13g2_fill_1 FILLER_53_2204 ();
 sg13g2_decap_4 FILLER_53_2231 ();
 sg13g2_fill_2 FILLER_53_2235 ();
 sg13g2_decap_8 FILLER_53_2268 ();
 sg13g2_decap_8 FILLER_53_2275 ();
 sg13g2_decap_8 FILLER_53_2282 ();
 sg13g2_decap_8 FILLER_53_2289 ();
 sg13g2_decap_8 FILLER_53_2296 ();
 sg13g2_decap_8 FILLER_53_2303 ();
 sg13g2_decap_8 FILLER_53_2310 ();
 sg13g2_decap_8 FILLER_53_2317 ();
 sg13g2_fill_2 FILLER_53_2324 ();
 sg13g2_decap_8 FILLER_53_2334 ();
 sg13g2_decap_8 FILLER_53_2341 ();
 sg13g2_fill_2 FILLER_53_2348 ();
 sg13g2_fill_1 FILLER_53_2350 ();
 sg13g2_decap_8 FILLER_53_2391 ();
 sg13g2_decap_4 FILLER_53_2398 ();
 sg13g2_fill_2 FILLER_53_2402 ();
 sg13g2_fill_1 FILLER_53_2417 ();
 sg13g2_decap_4 FILLER_53_2424 ();
 sg13g2_decap_4 FILLER_53_2436 ();
 sg13g2_decap_4 FILLER_53_2518 ();
 sg13g2_fill_2 FILLER_53_2522 ();
 sg13g2_decap_4 FILLER_53_2576 ();
 sg13g2_fill_2 FILLER_53_2580 ();
 sg13g2_decap_4 FILLER_53_2606 ();
 sg13g2_decap_8 FILLER_53_2706 ();
 sg13g2_decap_8 FILLER_53_2713 ();
 sg13g2_decap_4 FILLER_53_2720 ();
 sg13g2_decap_8 FILLER_53_2755 ();
 sg13g2_decap_8 FILLER_53_2762 ();
 sg13g2_decap_8 FILLER_53_2769 ();
 sg13g2_decap_4 FILLER_53_2776 ();
 sg13g2_decap_8 FILLER_53_2806 ();
 sg13g2_decap_8 FILLER_53_2813 ();
 sg13g2_decap_8 FILLER_53_2820 ();
 sg13g2_decap_8 FILLER_53_2827 ();
 sg13g2_decap_8 FILLER_53_2866 ();
 sg13g2_decap_8 FILLER_53_2873 ();
 sg13g2_decap_8 FILLER_53_2880 ();
 sg13g2_decap_8 FILLER_53_2887 ();
 sg13g2_decap_4 FILLER_53_2894 ();
 sg13g2_decap_8 FILLER_53_2990 ();
 sg13g2_decap_8 FILLER_53_2997 ();
 sg13g2_decap_8 FILLER_53_3004 ();
 sg13g2_decap_8 FILLER_53_3011 ();
 sg13g2_decap_8 FILLER_53_3018 ();
 sg13g2_decap_8 FILLER_53_3025 ();
 sg13g2_decap_8 FILLER_53_3032 ();
 sg13g2_decap_8 FILLER_53_3039 ();
 sg13g2_decap_8 FILLER_53_3046 ();
 sg13g2_decap_8 FILLER_53_3053 ();
 sg13g2_decap_8 FILLER_53_3060 ();
 sg13g2_decap_8 FILLER_53_3067 ();
 sg13g2_decap_8 FILLER_53_3074 ();
 sg13g2_decap_8 FILLER_53_3081 ();
 sg13g2_decap_8 FILLER_53_3088 ();
 sg13g2_decap_8 FILLER_53_3095 ();
 sg13g2_decap_8 FILLER_53_3102 ();
 sg13g2_decap_8 FILLER_53_3109 ();
 sg13g2_decap_8 FILLER_53_3116 ();
 sg13g2_decap_8 FILLER_53_3123 ();
 sg13g2_decap_8 FILLER_53_3130 ();
 sg13g2_decap_8 FILLER_53_3137 ();
 sg13g2_decap_8 FILLER_53_3144 ();
 sg13g2_decap_8 FILLER_53_3151 ();
 sg13g2_decap_8 FILLER_53_3158 ();
 sg13g2_decap_8 FILLER_53_3165 ();
 sg13g2_decap_8 FILLER_53_3172 ();
 sg13g2_decap_8 FILLER_53_3179 ();
 sg13g2_decap_8 FILLER_53_3186 ();
 sg13g2_decap_8 FILLER_53_3193 ();
 sg13g2_decap_8 FILLER_53_3200 ();
 sg13g2_decap_8 FILLER_53_3207 ();
 sg13g2_decap_8 FILLER_53_3214 ();
 sg13g2_decap_8 FILLER_53_3221 ();
 sg13g2_decap_8 FILLER_53_3228 ();
 sg13g2_decap_8 FILLER_53_3235 ();
 sg13g2_decap_8 FILLER_53_3242 ();
 sg13g2_decap_8 FILLER_53_3249 ();
 sg13g2_decap_8 FILLER_53_3256 ();
 sg13g2_decap_8 FILLER_53_3263 ();
 sg13g2_decap_8 FILLER_53_3270 ();
 sg13g2_decap_8 FILLER_53_3277 ();
 sg13g2_decap_8 FILLER_53_3284 ();
 sg13g2_decap_8 FILLER_53_3291 ();
 sg13g2_decap_8 FILLER_53_3298 ();
 sg13g2_decap_8 FILLER_53_3305 ();
 sg13g2_decap_8 FILLER_53_3312 ();
 sg13g2_decap_8 FILLER_53_3319 ();
 sg13g2_decap_8 FILLER_53_3326 ();
 sg13g2_decap_8 FILLER_53_3333 ();
 sg13g2_decap_8 FILLER_53_3340 ();
 sg13g2_decap_8 FILLER_53_3347 ();
 sg13g2_decap_8 FILLER_53_3354 ();
 sg13g2_decap_8 FILLER_53_3361 ();
 sg13g2_decap_8 FILLER_53_3368 ();
 sg13g2_decap_8 FILLER_53_3375 ();
 sg13g2_decap_8 FILLER_53_3382 ();
 sg13g2_decap_8 FILLER_53_3389 ();
 sg13g2_decap_8 FILLER_53_3396 ();
 sg13g2_decap_8 FILLER_53_3403 ();
 sg13g2_decap_8 FILLER_53_3410 ();
 sg13g2_decap_8 FILLER_53_3417 ();
 sg13g2_decap_8 FILLER_53_3424 ();
 sg13g2_decap_8 FILLER_53_3431 ();
 sg13g2_decap_8 FILLER_53_3438 ();
 sg13g2_decap_8 FILLER_53_3445 ();
 sg13g2_decap_8 FILLER_53_3452 ();
 sg13g2_decap_8 FILLER_53_3459 ();
 sg13g2_decap_8 FILLER_53_3466 ();
 sg13g2_decap_8 FILLER_53_3473 ();
 sg13g2_decap_8 FILLER_53_3480 ();
 sg13g2_decap_8 FILLER_53_3487 ();
 sg13g2_decap_8 FILLER_53_3494 ();
 sg13g2_decap_8 FILLER_53_3501 ();
 sg13g2_decap_8 FILLER_53_3508 ();
 sg13g2_decap_8 FILLER_53_3515 ();
 sg13g2_decap_8 FILLER_53_3522 ();
 sg13g2_decap_8 FILLER_53_3529 ();
 sg13g2_decap_8 FILLER_53_3536 ();
 sg13g2_decap_8 FILLER_53_3543 ();
 sg13g2_decap_8 FILLER_53_3550 ();
 sg13g2_decap_8 FILLER_53_3557 ();
 sg13g2_decap_8 FILLER_53_3564 ();
 sg13g2_decap_8 FILLER_53_3571 ();
 sg13g2_fill_2 FILLER_53_3578 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_decap_8 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_182 ();
 sg13g2_decap_8 FILLER_54_189 ();
 sg13g2_decap_8 FILLER_54_196 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_decap_8 FILLER_54_210 ();
 sg13g2_decap_8 FILLER_54_217 ();
 sg13g2_decap_8 FILLER_54_224 ();
 sg13g2_decap_8 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_238 ();
 sg13g2_decap_8 FILLER_54_245 ();
 sg13g2_decap_8 FILLER_54_252 ();
 sg13g2_decap_8 FILLER_54_259 ();
 sg13g2_decap_8 FILLER_54_266 ();
 sg13g2_decap_4 FILLER_54_273 ();
 sg13g2_fill_2 FILLER_54_277 ();
 sg13g2_decap_8 FILLER_54_283 ();
 sg13g2_decap_8 FILLER_54_290 ();
 sg13g2_decap_8 FILLER_54_297 ();
 sg13g2_decap_8 FILLER_54_304 ();
 sg13g2_decap_8 FILLER_54_311 ();
 sg13g2_decap_8 FILLER_54_318 ();
 sg13g2_fill_1 FILLER_54_385 ();
 sg13g2_fill_2 FILLER_54_421 ();
 sg13g2_decap_4 FILLER_54_436 ();
 sg13g2_fill_1 FILLER_54_440 ();
 sg13g2_fill_2 FILLER_54_467 ();
 sg13g2_fill_1 FILLER_54_469 ();
 sg13g2_decap_8 FILLER_54_499 ();
 sg13g2_decap_8 FILLER_54_506 ();
 sg13g2_decap_8 FILLER_54_513 ();
 sg13g2_decap_8 FILLER_54_525 ();
 sg13g2_decap_8 FILLER_54_532 ();
 sg13g2_decap_4 FILLER_54_539 ();
 sg13g2_fill_1 FILLER_54_543 ();
 sg13g2_decap_8 FILLER_54_573 ();
 sg13g2_fill_2 FILLER_54_580 ();
 sg13g2_fill_1 FILLER_54_582 ();
 sg13g2_decap_8 FILLER_54_609 ();
 sg13g2_decap_8 FILLER_54_616 ();
 sg13g2_decap_8 FILLER_54_623 ();
 sg13g2_decap_8 FILLER_54_630 ();
 sg13g2_fill_2 FILLER_54_637 ();
 sg13g2_fill_2 FILLER_54_670 ();
 sg13g2_fill_2 FILLER_54_677 ();
 sg13g2_fill_1 FILLER_54_679 ();
 sg13g2_fill_2 FILLER_54_700 ();
 sg13g2_fill_2 FILLER_54_715 ();
 sg13g2_decap_8 FILLER_54_725 ();
 sg13g2_decap_8 FILLER_54_732 ();
 sg13g2_decap_4 FILLER_54_739 ();
 sg13g2_decap_8 FILLER_54_747 ();
 sg13g2_decap_8 FILLER_54_754 ();
 sg13g2_decap_8 FILLER_54_761 ();
 sg13g2_decap_8 FILLER_54_768 ();
 sg13g2_decap_4 FILLER_54_775 ();
 sg13g2_fill_1 FILLER_54_779 ();
 sg13g2_decap_8 FILLER_54_791 ();
 sg13g2_fill_2 FILLER_54_805 ();
 sg13g2_fill_1 FILLER_54_810 ();
 sg13g2_decap_8 FILLER_54_815 ();
 sg13g2_fill_2 FILLER_54_822 ();
 sg13g2_fill_1 FILLER_54_835 ();
 sg13g2_decap_4 FILLER_54_841 ();
 sg13g2_decap_8 FILLER_54_853 ();
 sg13g2_decap_8 FILLER_54_860 ();
 sg13g2_fill_1 FILLER_54_867 ();
 sg13g2_decap_8 FILLER_54_876 ();
 sg13g2_decap_8 FILLER_54_883 ();
 sg13g2_decap_8 FILLER_54_890 ();
 sg13g2_decap_4 FILLER_54_907 ();
 sg13g2_fill_2 FILLER_54_911 ();
 sg13g2_decap_8 FILLER_54_939 ();
 sg13g2_decap_8 FILLER_54_982 ();
 sg13g2_decap_8 FILLER_54_989 ();
 sg13g2_decap_4 FILLER_54_996 ();
 sg13g2_fill_1 FILLER_54_1000 ();
 sg13g2_decap_8 FILLER_54_1027 ();
 sg13g2_decap_8 FILLER_54_1034 ();
 sg13g2_decap_8 FILLER_54_1041 ();
 sg13g2_fill_2 FILLER_54_1048 ();
 sg13g2_decap_8 FILLER_54_1134 ();
 sg13g2_fill_1 FILLER_54_1141 ();
 sg13g2_decap_4 FILLER_54_1172 ();
 sg13g2_fill_1 FILLER_54_1176 ();
 sg13g2_decap_8 FILLER_54_1203 ();
 sg13g2_fill_2 FILLER_54_1210 ();
 sg13g2_decap_8 FILLER_54_1249 ();
 sg13g2_fill_2 FILLER_54_1256 ();
 sg13g2_decap_4 FILLER_54_1288 ();
 sg13g2_decap_8 FILLER_54_1318 ();
 sg13g2_decap_8 FILLER_54_1325 ();
 sg13g2_decap_4 FILLER_54_1332 ();
 sg13g2_decap_4 FILLER_54_1360 ();
 sg13g2_fill_2 FILLER_54_1364 ();
 sg13g2_fill_2 FILLER_54_1374 ();
 sg13g2_fill_1 FILLER_54_1376 ();
 sg13g2_decap_8 FILLER_54_1398 ();
 sg13g2_fill_2 FILLER_54_1405 ();
 sg13g2_fill_1 FILLER_54_1407 ();
 sg13g2_decap_8 FILLER_54_1501 ();
 sg13g2_decap_8 FILLER_54_1508 ();
 sg13g2_decap_4 FILLER_54_1515 ();
 sg13g2_decap_8 FILLER_54_1571 ();
 sg13g2_decap_8 FILLER_54_1578 ();
 sg13g2_fill_1 FILLER_54_1585 ();
 sg13g2_fill_1 FILLER_54_1615 ();
 sg13g2_fill_2 FILLER_54_1620 ();
 sg13g2_decap_8 FILLER_54_1674 ();
 sg13g2_decap_8 FILLER_54_1681 ();
 sg13g2_fill_2 FILLER_54_1688 ();
 sg13g2_decap_8 FILLER_54_1716 ();
 sg13g2_decap_8 FILLER_54_1723 ();
 sg13g2_decap_8 FILLER_54_1730 ();
 sg13g2_decap_8 FILLER_54_1737 ();
 sg13g2_decap_8 FILLER_54_1744 ();
 sg13g2_decap_4 FILLER_54_1751 ();
 sg13g2_decap_8 FILLER_54_1781 ();
 sg13g2_decap_8 FILLER_54_1788 ();
 sg13g2_decap_8 FILLER_54_1795 ();
 sg13g2_decap_8 FILLER_54_1802 ();
 sg13g2_fill_2 FILLER_54_1809 ();
 sg13g2_decap_8 FILLER_54_1837 ();
 sg13g2_decap_8 FILLER_54_1844 ();
 sg13g2_fill_1 FILLER_54_1851 ();
 sg13g2_fill_2 FILLER_54_1878 ();
 sg13g2_decap_8 FILLER_54_1906 ();
 sg13g2_decap_8 FILLER_54_1913 ();
 sg13g2_decap_8 FILLER_54_1920 ();
 sg13g2_decap_4 FILLER_54_1927 ();
 sg13g2_fill_2 FILLER_54_1931 ();
 sg13g2_fill_2 FILLER_54_2011 ();
 sg13g2_fill_1 FILLER_54_2013 ();
 sg13g2_decap_8 FILLER_54_2066 ();
 sg13g2_decap_8 FILLER_54_2073 ();
 sg13g2_decap_8 FILLER_54_2080 ();
 sg13g2_decap_8 FILLER_54_2087 ();
 sg13g2_fill_1 FILLER_54_2094 ();
 sg13g2_decap_8 FILLER_54_2147 ();
 sg13g2_decap_8 FILLER_54_2154 ();
 sg13g2_decap_8 FILLER_54_2161 ();
 sg13g2_fill_2 FILLER_54_2168 ();
 sg13g2_decap_4 FILLER_54_2202 ();
 sg13g2_fill_1 FILLER_54_2232 ();
 sg13g2_decap_8 FILLER_54_2259 ();
 sg13g2_decap_8 FILLER_54_2266 ();
 sg13g2_decap_8 FILLER_54_2273 ();
 sg13g2_decap_8 FILLER_54_2280 ();
 sg13g2_decap_8 FILLER_54_2287 ();
 sg13g2_decap_8 FILLER_54_2294 ();
 sg13g2_decap_8 FILLER_54_2301 ();
 sg13g2_decap_8 FILLER_54_2308 ();
 sg13g2_fill_2 FILLER_54_2315 ();
 sg13g2_fill_1 FILLER_54_2317 ();
 sg13g2_decap_8 FILLER_54_2344 ();
 sg13g2_decap_4 FILLER_54_2351 ();
 sg13g2_fill_1 FILLER_54_2355 ();
 sg13g2_decap_8 FILLER_54_2450 ();
 sg13g2_decap_4 FILLER_54_2457 ();
 sg13g2_fill_1 FILLER_54_2461 ();
 sg13g2_decap_8 FILLER_54_2501 ();
 sg13g2_decap_4 FILLER_54_2508 ();
 sg13g2_decap_4 FILLER_54_2588 ();
 sg13g2_fill_1 FILLER_54_2592 ();
 sg13g2_decap_8 FILLER_54_2601 ();
 sg13g2_decap_4 FILLER_54_2608 ();
 sg13g2_fill_2 FILLER_54_2612 ();
 sg13g2_fill_2 FILLER_54_2653 ();
 sg13g2_decap_8 FILLER_54_2712 ();
 sg13g2_decap_8 FILLER_54_2719 ();
 sg13g2_decap_8 FILLER_54_2726 ();
 sg13g2_fill_2 FILLER_54_2733 ();
 sg13g2_fill_1 FILLER_54_2735 ();
 sg13g2_decap_8 FILLER_54_2762 ();
 sg13g2_fill_2 FILLER_54_2803 ();
 sg13g2_fill_2 FILLER_54_2810 ();
 sg13g2_decap_8 FILLER_54_2817 ();
 sg13g2_decap_4 FILLER_54_2824 ();
 sg13g2_fill_2 FILLER_54_2828 ();
 sg13g2_fill_2 FILLER_54_2882 ();
 sg13g2_fill_1 FILLER_54_2916 ();
 sg13g2_decap_8 FILLER_54_2925 ();
 sg13g2_decap_8 FILLER_54_2932 ();
 sg13g2_decap_8 FILLER_54_2939 ();
 sg13g2_decap_8 FILLER_54_3004 ();
 sg13g2_decap_8 FILLER_54_3011 ();
 sg13g2_decap_8 FILLER_54_3018 ();
 sg13g2_decap_8 FILLER_54_3025 ();
 sg13g2_decap_8 FILLER_54_3032 ();
 sg13g2_decap_8 FILLER_54_3039 ();
 sg13g2_decap_8 FILLER_54_3046 ();
 sg13g2_decap_8 FILLER_54_3053 ();
 sg13g2_decap_8 FILLER_54_3060 ();
 sg13g2_decap_8 FILLER_54_3067 ();
 sg13g2_decap_8 FILLER_54_3074 ();
 sg13g2_decap_8 FILLER_54_3081 ();
 sg13g2_decap_8 FILLER_54_3088 ();
 sg13g2_decap_8 FILLER_54_3095 ();
 sg13g2_decap_8 FILLER_54_3102 ();
 sg13g2_decap_8 FILLER_54_3109 ();
 sg13g2_decap_8 FILLER_54_3116 ();
 sg13g2_decap_8 FILLER_54_3123 ();
 sg13g2_decap_8 FILLER_54_3130 ();
 sg13g2_decap_8 FILLER_54_3137 ();
 sg13g2_decap_8 FILLER_54_3144 ();
 sg13g2_decap_8 FILLER_54_3151 ();
 sg13g2_decap_8 FILLER_54_3158 ();
 sg13g2_decap_8 FILLER_54_3165 ();
 sg13g2_decap_8 FILLER_54_3172 ();
 sg13g2_decap_8 FILLER_54_3179 ();
 sg13g2_decap_8 FILLER_54_3186 ();
 sg13g2_decap_8 FILLER_54_3193 ();
 sg13g2_decap_8 FILLER_54_3200 ();
 sg13g2_decap_8 FILLER_54_3207 ();
 sg13g2_decap_8 FILLER_54_3214 ();
 sg13g2_decap_8 FILLER_54_3221 ();
 sg13g2_decap_8 FILLER_54_3228 ();
 sg13g2_decap_8 FILLER_54_3235 ();
 sg13g2_decap_8 FILLER_54_3242 ();
 sg13g2_decap_8 FILLER_54_3249 ();
 sg13g2_decap_8 FILLER_54_3256 ();
 sg13g2_decap_8 FILLER_54_3263 ();
 sg13g2_decap_8 FILLER_54_3270 ();
 sg13g2_decap_8 FILLER_54_3277 ();
 sg13g2_decap_8 FILLER_54_3284 ();
 sg13g2_decap_8 FILLER_54_3291 ();
 sg13g2_decap_8 FILLER_54_3298 ();
 sg13g2_decap_8 FILLER_54_3305 ();
 sg13g2_decap_8 FILLER_54_3312 ();
 sg13g2_decap_8 FILLER_54_3319 ();
 sg13g2_decap_8 FILLER_54_3326 ();
 sg13g2_decap_8 FILLER_54_3333 ();
 sg13g2_decap_8 FILLER_54_3340 ();
 sg13g2_decap_8 FILLER_54_3347 ();
 sg13g2_decap_8 FILLER_54_3354 ();
 sg13g2_decap_8 FILLER_54_3361 ();
 sg13g2_decap_8 FILLER_54_3368 ();
 sg13g2_decap_8 FILLER_54_3375 ();
 sg13g2_decap_8 FILLER_54_3382 ();
 sg13g2_decap_8 FILLER_54_3389 ();
 sg13g2_decap_8 FILLER_54_3396 ();
 sg13g2_decap_8 FILLER_54_3403 ();
 sg13g2_decap_8 FILLER_54_3410 ();
 sg13g2_decap_8 FILLER_54_3417 ();
 sg13g2_decap_8 FILLER_54_3424 ();
 sg13g2_decap_8 FILLER_54_3431 ();
 sg13g2_decap_8 FILLER_54_3438 ();
 sg13g2_decap_8 FILLER_54_3445 ();
 sg13g2_decap_8 FILLER_54_3452 ();
 sg13g2_decap_8 FILLER_54_3459 ();
 sg13g2_decap_8 FILLER_54_3466 ();
 sg13g2_decap_8 FILLER_54_3473 ();
 sg13g2_decap_8 FILLER_54_3480 ();
 sg13g2_decap_8 FILLER_54_3487 ();
 sg13g2_decap_8 FILLER_54_3494 ();
 sg13g2_decap_8 FILLER_54_3501 ();
 sg13g2_decap_8 FILLER_54_3508 ();
 sg13g2_decap_8 FILLER_54_3515 ();
 sg13g2_decap_8 FILLER_54_3522 ();
 sg13g2_decap_8 FILLER_54_3529 ();
 sg13g2_decap_8 FILLER_54_3536 ();
 sg13g2_decap_8 FILLER_54_3543 ();
 sg13g2_decap_8 FILLER_54_3550 ();
 sg13g2_decap_8 FILLER_54_3557 ();
 sg13g2_decap_8 FILLER_54_3564 ();
 sg13g2_decap_8 FILLER_54_3571 ();
 sg13g2_fill_2 FILLER_54_3578 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_decap_8 FILLER_55_189 ();
 sg13g2_decap_8 FILLER_55_196 ();
 sg13g2_decap_8 FILLER_55_203 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_8 FILLER_55_224 ();
 sg13g2_decap_8 FILLER_55_231 ();
 sg13g2_decap_8 FILLER_55_238 ();
 sg13g2_decap_8 FILLER_55_245 ();
 sg13g2_decap_8 FILLER_55_252 ();
 sg13g2_decap_8 FILLER_55_259 ();
 sg13g2_decap_8 FILLER_55_266 ();
 sg13g2_decap_8 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_8 FILLER_55_287 ();
 sg13g2_decap_8 FILLER_55_294 ();
 sg13g2_decap_8 FILLER_55_301 ();
 sg13g2_decap_8 FILLER_55_308 ();
 sg13g2_decap_8 FILLER_55_315 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_1 FILLER_55_324 ();
 sg13g2_decap_8 FILLER_55_354 ();
 sg13g2_fill_2 FILLER_55_361 ();
 sg13g2_fill_1 FILLER_55_389 ();
 sg13g2_fill_1 FILLER_55_398 ();
 sg13g2_fill_2 FILLER_55_466 ();
 sg13g2_fill_1 FILLER_55_468 ();
 sg13g2_decap_8 FILLER_55_493 ();
 sg13g2_fill_1 FILLER_55_500 ();
 sg13g2_decap_8 FILLER_55_505 ();
 sg13g2_decap_8 FILLER_55_512 ();
 sg13g2_decap_8 FILLER_55_519 ();
 sg13g2_decap_8 FILLER_55_526 ();
 sg13g2_decap_8 FILLER_55_533 ();
 sg13g2_decap_8 FILLER_55_540 ();
 sg13g2_fill_1 FILLER_55_547 ();
 sg13g2_decap_8 FILLER_55_622 ();
 sg13g2_decap_8 FILLER_55_681 ();
 sg13g2_decap_8 FILLER_55_688 ();
 sg13g2_decap_4 FILLER_55_695 ();
 sg13g2_fill_1 FILLER_55_699 ();
 sg13g2_decap_8 FILLER_55_703 ();
 sg13g2_decap_8 FILLER_55_710 ();
 sg13g2_fill_2 FILLER_55_717 ();
 sg13g2_fill_2 FILLER_55_728 ();
 sg13g2_decap_8 FILLER_55_738 ();
 sg13g2_decap_8 FILLER_55_745 ();
 sg13g2_fill_2 FILLER_55_752 ();
 sg13g2_fill_1 FILLER_55_754 ();
 sg13g2_fill_2 FILLER_55_781 ();
 sg13g2_fill_1 FILLER_55_848 ();
 sg13g2_fill_2 FILLER_55_865 ();
 sg13g2_fill_2 FILLER_55_872 ();
 sg13g2_decap_8 FILLER_55_903 ();
 sg13g2_decap_4 FILLER_55_936 ();
 sg13g2_fill_2 FILLER_55_940 ();
 sg13g2_decap_4 FILLER_55_994 ();
 sg13g2_fill_2 FILLER_55_998 ();
 sg13g2_decap_8 FILLER_55_1010 ();
 sg13g2_fill_2 FILLER_55_1017 ();
 sg13g2_fill_1 FILLER_55_1019 ();
 sg13g2_decap_8 FILLER_55_1046 ();
 sg13g2_decap_8 FILLER_55_1053 ();
 sg13g2_decap_4 FILLER_55_1060 ();
 sg13g2_decap_8 FILLER_55_1072 ();
 sg13g2_decap_8 FILLER_55_1079 ();
 sg13g2_decap_8 FILLER_55_1086 ();
 sg13g2_decap_4 FILLER_55_1093 ();
 sg13g2_fill_1 FILLER_55_1097 ();
 sg13g2_decap_8 FILLER_55_1129 ();
 sg13g2_decap_8 FILLER_55_1136 ();
 sg13g2_decap_8 FILLER_55_1143 ();
 sg13g2_decap_8 FILLER_55_1150 ();
 sg13g2_decap_4 FILLER_55_1157 ();
 sg13g2_fill_2 FILLER_55_1161 ();
 sg13g2_fill_2 FILLER_55_1169 ();
 sg13g2_decap_8 FILLER_55_1177 ();
 sg13g2_decap_8 FILLER_55_1184 ();
 sg13g2_decap_4 FILLER_55_1191 ();
 sg13g2_fill_2 FILLER_55_1195 ();
 sg13g2_decap_8 FILLER_55_1202 ();
 sg13g2_decap_8 FILLER_55_1209 ();
 sg13g2_decap_8 FILLER_55_1216 ();
 sg13g2_decap_4 FILLER_55_1223 ();
 sg13g2_fill_1 FILLER_55_1227 ();
 sg13g2_fill_1 FILLER_55_1233 ();
 sg13g2_decap_8 FILLER_55_1244 ();
 sg13g2_decap_8 FILLER_55_1251 ();
 sg13g2_fill_2 FILLER_55_1258 ();
 sg13g2_fill_1 FILLER_55_1260 ();
 sg13g2_decap_8 FILLER_55_1339 ();
 sg13g2_decap_8 FILLER_55_1350 ();
 sg13g2_fill_2 FILLER_55_1357 ();
 sg13g2_fill_1 FILLER_55_1359 ();
 sg13g2_decap_8 FILLER_55_1389 ();
 sg13g2_fill_1 FILLER_55_1396 ();
 sg13g2_decap_8 FILLER_55_1501 ();
 sg13g2_decap_8 FILLER_55_1508 ();
 sg13g2_decap_8 FILLER_55_1515 ();
 sg13g2_decap_8 FILLER_55_1568 ();
 sg13g2_decap_8 FILLER_55_1575 ();
 sg13g2_decap_8 FILLER_55_1582 ();
 sg13g2_decap_4 FILLER_55_1589 ();
 sg13g2_decap_8 FILLER_55_1631 ();
 sg13g2_fill_2 FILLER_55_1638 ();
 sg13g2_decap_8 FILLER_55_1648 ();
 sg13g2_decap_8 FILLER_55_1655 ();
 sg13g2_fill_1 FILLER_55_1662 ();
 sg13g2_decap_8 FILLER_55_1668 ();
 sg13g2_decap_8 FILLER_55_1675 ();
 sg13g2_decap_4 FILLER_55_1682 ();
 sg13g2_fill_2 FILLER_55_1686 ();
 sg13g2_fill_1 FILLER_55_1693 ();
 sg13g2_decap_8 FILLER_55_1732 ();
 sg13g2_decap_8 FILLER_55_1739 ();
 sg13g2_decap_8 FILLER_55_1746 ();
 sg13g2_decap_8 FILLER_55_1753 ();
 sg13g2_decap_8 FILLER_55_1760 ();
 sg13g2_fill_1 FILLER_55_1767 ();
 sg13g2_fill_2 FILLER_55_1803 ();
 sg13g2_decap_8 FILLER_55_1844 ();
 sg13g2_decap_8 FILLER_55_1851 ();
 sg13g2_fill_1 FILLER_55_1858 ();
 sg13g2_decap_4 FILLER_55_1863 ();
 sg13g2_decap_8 FILLER_55_1940 ();
 sg13g2_fill_2 FILLER_55_1947 ();
 sg13g2_decap_8 FILLER_55_2001 ();
 sg13g2_decap_8 FILLER_55_2008 ();
 sg13g2_decap_8 FILLER_55_2015 ();
 sg13g2_decap_4 FILLER_55_2022 ();
 sg13g2_decap_8 FILLER_55_2052 ();
 sg13g2_decap_8 FILLER_55_2059 ();
 sg13g2_decap_8 FILLER_55_2066 ();
 sg13g2_decap_8 FILLER_55_2073 ();
 sg13g2_fill_2 FILLER_55_2080 ();
 sg13g2_fill_1 FILLER_55_2082 ();
 sg13g2_decap_8 FILLER_55_2135 ();
 sg13g2_decap_8 FILLER_55_2142 ();
 sg13g2_decap_8 FILLER_55_2149 ();
 sg13g2_decap_8 FILLER_55_2156 ();
 sg13g2_decap_8 FILLER_55_2163 ();
 sg13g2_decap_4 FILLER_55_2170 ();
 sg13g2_fill_1 FILLER_55_2174 ();
 sg13g2_decap_8 FILLER_55_2227 ();
 sg13g2_decap_8 FILLER_55_2234 ();
 sg13g2_decap_4 FILLER_55_2241 ();
 sg13g2_fill_1 FILLER_55_2245 ();
 sg13g2_decap_8 FILLER_55_2272 ();
 sg13g2_decap_8 FILLER_55_2279 ();
 sg13g2_decap_8 FILLER_55_2286 ();
 sg13g2_decap_8 FILLER_55_2293 ();
 sg13g2_decap_8 FILLER_55_2300 ();
 sg13g2_decap_4 FILLER_55_2307 ();
 sg13g2_fill_1 FILLER_55_2311 ();
 sg13g2_decap_8 FILLER_55_2442 ();
 sg13g2_fill_2 FILLER_55_2449 ();
 sg13g2_fill_1 FILLER_55_2451 ();
 sg13g2_decap_8 FILLER_55_2495 ();
 sg13g2_decap_8 FILLER_55_2502 ();
 sg13g2_decap_8 FILLER_55_2509 ();
 sg13g2_decap_4 FILLER_55_2516 ();
 sg13g2_fill_1 FILLER_55_2552 ();
 sg13g2_decap_8 FILLER_55_2584 ();
 sg13g2_decap_8 FILLER_55_2591 ();
 sg13g2_decap_8 FILLER_55_2598 ();
 sg13g2_decap_8 FILLER_55_2605 ();
 sg13g2_decap_8 FILLER_55_2612 ();
 sg13g2_fill_2 FILLER_55_2619 ();
 sg13g2_fill_1 FILLER_55_2673 ();
 sg13g2_decap_8 FILLER_55_2717 ();
 sg13g2_decap_8 FILLER_55_2724 ();
 sg13g2_decap_8 FILLER_55_2731 ();
 sg13g2_decap_8 FILLER_55_2809 ();
 sg13g2_decap_8 FILLER_55_2816 ();
 sg13g2_decap_8 FILLER_55_2823 ();
 sg13g2_fill_1 FILLER_55_2830 ();
 sg13g2_decap_8 FILLER_55_2869 ();
 sg13g2_decap_8 FILLER_55_2876 ();
 sg13g2_decap_8 FILLER_55_2883 ();
 sg13g2_fill_2 FILLER_55_2890 ();
 sg13g2_decap_8 FILLER_55_2929 ();
 sg13g2_decap_8 FILLER_55_2936 ();
 sg13g2_decap_8 FILLER_55_2943 ();
 sg13g2_fill_2 FILLER_55_2950 ();
 sg13g2_fill_1 FILLER_55_2952 ();
 sg13g2_decap_8 FILLER_55_2991 ();
 sg13g2_decap_8 FILLER_55_2998 ();
 sg13g2_decap_8 FILLER_55_3005 ();
 sg13g2_decap_8 FILLER_55_3012 ();
 sg13g2_decap_8 FILLER_55_3019 ();
 sg13g2_decap_8 FILLER_55_3026 ();
 sg13g2_decap_8 FILLER_55_3033 ();
 sg13g2_decap_8 FILLER_55_3040 ();
 sg13g2_decap_8 FILLER_55_3047 ();
 sg13g2_decap_8 FILLER_55_3054 ();
 sg13g2_decap_8 FILLER_55_3061 ();
 sg13g2_decap_8 FILLER_55_3068 ();
 sg13g2_decap_8 FILLER_55_3075 ();
 sg13g2_decap_8 FILLER_55_3082 ();
 sg13g2_decap_8 FILLER_55_3089 ();
 sg13g2_decap_8 FILLER_55_3096 ();
 sg13g2_decap_8 FILLER_55_3103 ();
 sg13g2_decap_8 FILLER_55_3110 ();
 sg13g2_decap_8 FILLER_55_3117 ();
 sg13g2_decap_8 FILLER_55_3124 ();
 sg13g2_decap_8 FILLER_55_3131 ();
 sg13g2_decap_8 FILLER_55_3138 ();
 sg13g2_decap_8 FILLER_55_3145 ();
 sg13g2_decap_8 FILLER_55_3152 ();
 sg13g2_decap_8 FILLER_55_3159 ();
 sg13g2_decap_8 FILLER_55_3166 ();
 sg13g2_decap_8 FILLER_55_3173 ();
 sg13g2_decap_8 FILLER_55_3180 ();
 sg13g2_decap_8 FILLER_55_3187 ();
 sg13g2_decap_8 FILLER_55_3194 ();
 sg13g2_decap_8 FILLER_55_3201 ();
 sg13g2_decap_8 FILLER_55_3208 ();
 sg13g2_decap_8 FILLER_55_3215 ();
 sg13g2_decap_8 FILLER_55_3222 ();
 sg13g2_decap_8 FILLER_55_3229 ();
 sg13g2_decap_8 FILLER_55_3236 ();
 sg13g2_decap_8 FILLER_55_3243 ();
 sg13g2_decap_8 FILLER_55_3250 ();
 sg13g2_decap_8 FILLER_55_3257 ();
 sg13g2_decap_8 FILLER_55_3264 ();
 sg13g2_decap_8 FILLER_55_3271 ();
 sg13g2_decap_8 FILLER_55_3278 ();
 sg13g2_decap_8 FILLER_55_3285 ();
 sg13g2_decap_8 FILLER_55_3292 ();
 sg13g2_decap_8 FILLER_55_3299 ();
 sg13g2_decap_8 FILLER_55_3306 ();
 sg13g2_decap_8 FILLER_55_3313 ();
 sg13g2_decap_8 FILLER_55_3320 ();
 sg13g2_decap_8 FILLER_55_3327 ();
 sg13g2_decap_8 FILLER_55_3334 ();
 sg13g2_decap_8 FILLER_55_3341 ();
 sg13g2_decap_8 FILLER_55_3348 ();
 sg13g2_decap_8 FILLER_55_3355 ();
 sg13g2_decap_8 FILLER_55_3362 ();
 sg13g2_decap_8 FILLER_55_3369 ();
 sg13g2_decap_8 FILLER_55_3376 ();
 sg13g2_decap_8 FILLER_55_3383 ();
 sg13g2_decap_8 FILLER_55_3390 ();
 sg13g2_decap_8 FILLER_55_3397 ();
 sg13g2_decap_8 FILLER_55_3404 ();
 sg13g2_decap_8 FILLER_55_3411 ();
 sg13g2_decap_8 FILLER_55_3418 ();
 sg13g2_decap_8 FILLER_55_3425 ();
 sg13g2_decap_8 FILLER_55_3432 ();
 sg13g2_decap_8 FILLER_55_3439 ();
 sg13g2_decap_8 FILLER_55_3446 ();
 sg13g2_decap_8 FILLER_55_3453 ();
 sg13g2_decap_8 FILLER_55_3460 ();
 sg13g2_decap_8 FILLER_55_3467 ();
 sg13g2_decap_8 FILLER_55_3474 ();
 sg13g2_decap_8 FILLER_55_3481 ();
 sg13g2_decap_8 FILLER_55_3488 ();
 sg13g2_decap_8 FILLER_55_3495 ();
 sg13g2_decap_8 FILLER_55_3502 ();
 sg13g2_decap_8 FILLER_55_3509 ();
 sg13g2_decap_8 FILLER_55_3516 ();
 sg13g2_decap_8 FILLER_55_3523 ();
 sg13g2_decap_8 FILLER_55_3530 ();
 sg13g2_decap_8 FILLER_55_3537 ();
 sg13g2_decap_8 FILLER_55_3544 ();
 sg13g2_decap_8 FILLER_55_3551 ();
 sg13g2_decap_8 FILLER_55_3558 ();
 sg13g2_decap_8 FILLER_55_3565 ();
 sg13g2_decap_8 FILLER_55_3572 ();
 sg13g2_fill_1 FILLER_55_3579 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_decap_8 FILLER_56_182 ();
 sg13g2_decap_8 FILLER_56_189 ();
 sg13g2_decap_8 FILLER_56_196 ();
 sg13g2_decap_8 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_decap_8 FILLER_56_224 ();
 sg13g2_decap_8 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_238 ();
 sg13g2_decap_8 FILLER_56_245 ();
 sg13g2_decap_8 FILLER_56_252 ();
 sg13g2_decap_8 FILLER_56_259 ();
 sg13g2_decap_8 FILLER_56_266 ();
 sg13g2_decap_8 FILLER_56_273 ();
 sg13g2_decap_8 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_287 ();
 sg13g2_decap_8 FILLER_56_294 ();
 sg13g2_decap_8 FILLER_56_301 ();
 sg13g2_decap_8 FILLER_56_308 ();
 sg13g2_decap_8 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_322 ();
 sg13g2_fill_1 FILLER_56_329 ();
 sg13g2_decap_8 FILLER_56_356 ();
 sg13g2_fill_2 FILLER_56_363 ();
 sg13g2_fill_2 FILLER_56_381 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_56_446 ();
 sg13g2_decap_8 FILLER_56_453 ();
 sg13g2_decap_8 FILLER_56_460 ();
 sg13g2_fill_1 FILLER_56_506 ();
 sg13g2_fill_2 FILLER_56_512 ();
 sg13g2_fill_1 FILLER_56_514 ();
 sg13g2_decap_4 FILLER_56_546 ();
 sg13g2_decap_8 FILLER_56_615 ();
 sg13g2_fill_2 FILLER_56_622 ();
 sg13g2_fill_1 FILLER_56_624 ();
 sg13g2_decap_8 FILLER_56_638 ();
 sg13g2_fill_1 FILLER_56_645 ();
 sg13g2_decap_4 FILLER_56_662 ();
 sg13g2_fill_2 FILLER_56_670 ();
 sg13g2_decap_8 FILLER_56_751 ();
 sg13g2_fill_1 FILLER_56_758 ();
 sg13g2_decap_8 FILLER_56_789 ();
 sg13g2_fill_1 FILLER_56_804 ();
 sg13g2_fill_1 FILLER_56_835 ();
 sg13g2_fill_2 FILLER_56_849 ();
 sg13g2_fill_2 FILLER_56_880 ();
 sg13g2_fill_1 FILLER_56_882 ();
 sg13g2_decap_4 FILLER_56_909 ();
 sg13g2_fill_1 FILLER_56_913 ();
 sg13g2_decap_4 FILLER_56_944 ();
 sg13g2_fill_2 FILLER_56_948 ();
 sg13g2_decap_4 FILLER_56_976 ();
 sg13g2_fill_1 FILLER_56_980 ();
 sg13g2_fill_1 FILLER_56_1010 ();
 sg13g2_decap_8 FILLER_56_1053 ();
 sg13g2_decap_8 FILLER_56_1060 ();
 sg13g2_decap_8 FILLER_56_1067 ();
 sg13g2_decap_8 FILLER_56_1074 ();
 sg13g2_decap_8 FILLER_56_1081 ();
 sg13g2_decap_8 FILLER_56_1088 ();
 sg13g2_decap_8 FILLER_56_1121 ();
 sg13g2_decap_8 FILLER_56_1128 ();
 sg13g2_decap_8 FILLER_56_1135 ();
 sg13g2_decap_8 FILLER_56_1142 ();
 sg13g2_decap_8 FILLER_56_1149 ();
 sg13g2_decap_8 FILLER_56_1156 ();
 sg13g2_decap_8 FILLER_56_1163 ();
 sg13g2_decap_8 FILLER_56_1170 ();
 sg13g2_decap_8 FILLER_56_1177 ();
 sg13g2_fill_2 FILLER_56_1184 ();
 sg13g2_decap_8 FILLER_56_1212 ();
 sg13g2_decap_8 FILLER_56_1219 ();
 sg13g2_decap_4 FILLER_56_1226 ();
 sg13g2_fill_2 FILLER_56_1230 ();
 sg13g2_fill_2 FILLER_56_1258 ();
 sg13g2_decap_8 FILLER_56_1299 ();
 sg13g2_fill_2 FILLER_56_1306 ();
 sg13g2_decap_8 FILLER_56_1339 ();
 sg13g2_decap_8 FILLER_56_1346 ();
 sg13g2_decap_8 FILLER_56_1353 ();
 sg13g2_fill_2 FILLER_56_1360 ();
 sg13g2_fill_2 FILLER_56_1371 ();
 sg13g2_decap_8 FILLER_56_1404 ();
 sg13g2_decap_8 FILLER_56_1411 ();
 sg13g2_fill_2 FILLER_56_1418 ();
 sg13g2_decap_8 FILLER_56_1446 ();
 sg13g2_decap_4 FILLER_56_1453 ();
 sg13g2_decap_8 FILLER_56_1488 ();
 sg13g2_decap_8 FILLER_56_1495 ();
 sg13g2_decap_8 FILLER_56_1502 ();
 sg13g2_decap_8 FILLER_56_1509 ();
 sg13g2_decap_8 FILLER_56_1516 ();
 sg13g2_decap_4 FILLER_56_1523 ();
 sg13g2_fill_2 FILLER_56_1527 ();
 sg13g2_decap_8 FILLER_56_1558 ();
 sg13g2_decap_8 FILLER_56_1565 ();
 sg13g2_decap_8 FILLER_56_1572 ();
 sg13g2_decap_4 FILLER_56_1579 ();
 sg13g2_fill_2 FILLER_56_1662 ();
 sg13g2_fill_1 FILLER_56_1664 ();
 sg13g2_fill_2 FILLER_56_1691 ();
 sg13g2_decap_8 FILLER_56_1732 ();
 sg13g2_decap_8 FILLER_56_1739 ();
 sg13g2_decap_4 FILLER_56_1746 ();
 sg13g2_fill_1 FILLER_56_1750 ();
 sg13g2_decap_8 FILLER_56_1818 ();
 sg13g2_decap_8 FILLER_56_1825 ();
 sg13g2_fill_1 FILLER_56_1832 ();
 sg13g2_decap_8 FILLER_56_1862 ();
 sg13g2_fill_1 FILLER_56_1869 ();
 sg13g2_fill_2 FILLER_56_1922 ();
 sg13g2_decap_8 FILLER_56_1934 ();
 sg13g2_decap_8 FILLER_56_1941 ();
 sg13g2_fill_1 FILLER_56_1948 ();
 sg13g2_decap_4 FILLER_56_1954 ();
 sg13g2_decap_8 FILLER_56_1966 ();
 sg13g2_decap_8 FILLER_56_1973 ();
 sg13g2_decap_8 FILLER_56_1980 ();
 sg13g2_decap_8 FILLER_56_1987 ();
 sg13g2_decap_8 FILLER_56_1994 ();
 sg13g2_decap_8 FILLER_56_2001 ();
 sg13g2_decap_8 FILLER_56_2008 ();
 sg13g2_decap_8 FILLER_56_2015 ();
 sg13g2_decap_8 FILLER_56_2022 ();
 sg13g2_decap_8 FILLER_56_2029 ();
 sg13g2_decap_4 FILLER_56_2088 ();
 sg13g2_fill_1 FILLER_56_2092 ();
 sg13g2_decap_8 FILLER_56_2145 ();
 sg13g2_decap_8 FILLER_56_2152 ();
 sg13g2_decap_8 FILLER_56_2159 ();
 sg13g2_decap_8 FILLER_56_2166 ();
 sg13g2_fill_2 FILLER_56_2173 ();
 sg13g2_fill_1 FILLER_56_2175 ();
 sg13g2_decap_8 FILLER_56_2202 ();
 sg13g2_decap_4 FILLER_56_2209 ();
 sg13g2_fill_2 FILLER_56_2213 ();
 sg13g2_decap_8 FILLER_56_2241 ();
 sg13g2_decap_8 FILLER_56_2248 ();
 sg13g2_decap_8 FILLER_56_2255 ();
 sg13g2_decap_8 FILLER_56_2262 ();
 sg13g2_decap_8 FILLER_56_2269 ();
 sg13g2_decap_8 FILLER_56_2276 ();
 sg13g2_decap_8 FILLER_56_2283 ();
 sg13g2_decap_8 FILLER_56_2290 ();
 sg13g2_decap_8 FILLER_56_2297 ();
 sg13g2_decap_8 FILLER_56_2304 ();
 sg13g2_decap_8 FILLER_56_2311 ();
 sg13g2_decap_8 FILLER_56_2318 ();
 sg13g2_decap_8 FILLER_56_2325 ();
 sg13g2_decap_8 FILLER_56_2332 ();
 sg13g2_fill_2 FILLER_56_2339 ();
 sg13g2_fill_1 FILLER_56_2341 ();
 sg13g2_fill_1 FILLER_56_2394 ();
 sg13g2_decap_8 FILLER_56_2447 ();
 sg13g2_decap_4 FILLER_56_2454 ();
 sg13g2_fill_2 FILLER_56_2458 ();
 sg13g2_fill_2 FILLER_56_2512 ();
 sg13g2_fill_1 FILLER_56_2514 ();
 sg13g2_fill_2 FILLER_56_2541 ();
 sg13g2_fill_1 FILLER_56_2543 ();
 sg13g2_fill_1 FILLER_56_2557 ();
 sg13g2_decap_8 FILLER_56_2584 ();
 sg13g2_decap_8 FILLER_56_2591 ();
 sg13g2_decap_8 FILLER_56_2598 ();
 sg13g2_decap_8 FILLER_56_2605 ();
 sg13g2_decap_4 FILLER_56_2612 ();
 sg13g2_fill_2 FILLER_56_2616 ();
 sg13g2_decap_8 FILLER_56_2649 ();
 sg13g2_decap_8 FILLER_56_2656 ();
 sg13g2_decap_8 FILLER_56_2663 ();
 sg13g2_decap_4 FILLER_56_2670 ();
 sg13g2_fill_2 FILLER_56_2674 ();
 sg13g2_fill_2 FILLER_56_2681 ();
 sg13g2_fill_1 FILLER_56_2683 ();
 sg13g2_fill_2 FILLER_56_2724 ();
 sg13g2_fill_1 FILLER_56_2726 ();
 sg13g2_decap_8 FILLER_56_2735 ();
 sg13g2_fill_1 FILLER_56_2742 ();
 sg13g2_decap_8 FILLER_56_2805 ();
 sg13g2_decap_8 FILLER_56_2812 ();
 sg13g2_decap_4 FILLER_56_2819 ();
 sg13g2_fill_1 FILLER_56_2823 ();
 sg13g2_decap_8 FILLER_56_2871 ();
 sg13g2_decap_8 FILLER_56_2878 ();
 sg13g2_decap_8 FILLER_56_2937 ();
 sg13g2_fill_2 FILLER_56_3007 ();
 sg13g2_fill_1 FILLER_56_3009 ();
 sg13g2_decap_8 FILLER_56_3036 ();
 sg13g2_decap_8 FILLER_56_3043 ();
 sg13g2_decap_8 FILLER_56_3050 ();
 sg13g2_decap_8 FILLER_56_3057 ();
 sg13g2_decap_8 FILLER_56_3064 ();
 sg13g2_decap_8 FILLER_56_3071 ();
 sg13g2_decap_8 FILLER_56_3078 ();
 sg13g2_decap_8 FILLER_56_3085 ();
 sg13g2_decap_8 FILLER_56_3092 ();
 sg13g2_decap_8 FILLER_56_3099 ();
 sg13g2_decap_8 FILLER_56_3106 ();
 sg13g2_decap_8 FILLER_56_3113 ();
 sg13g2_decap_8 FILLER_56_3120 ();
 sg13g2_decap_8 FILLER_56_3127 ();
 sg13g2_decap_8 FILLER_56_3134 ();
 sg13g2_decap_8 FILLER_56_3141 ();
 sg13g2_decap_8 FILLER_56_3148 ();
 sg13g2_decap_8 FILLER_56_3155 ();
 sg13g2_decap_8 FILLER_56_3162 ();
 sg13g2_decap_8 FILLER_56_3169 ();
 sg13g2_decap_8 FILLER_56_3176 ();
 sg13g2_decap_8 FILLER_56_3183 ();
 sg13g2_decap_8 FILLER_56_3190 ();
 sg13g2_decap_8 FILLER_56_3197 ();
 sg13g2_decap_8 FILLER_56_3204 ();
 sg13g2_decap_8 FILLER_56_3211 ();
 sg13g2_decap_8 FILLER_56_3218 ();
 sg13g2_decap_8 FILLER_56_3225 ();
 sg13g2_decap_8 FILLER_56_3232 ();
 sg13g2_decap_8 FILLER_56_3239 ();
 sg13g2_decap_8 FILLER_56_3246 ();
 sg13g2_decap_8 FILLER_56_3253 ();
 sg13g2_decap_8 FILLER_56_3260 ();
 sg13g2_decap_8 FILLER_56_3267 ();
 sg13g2_decap_8 FILLER_56_3274 ();
 sg13g2_decap_8 FILLER_56_3281 ();
 sg13g2_decap_8 FILLER_56_3288 ();
 sg13g2_decap_8 FILLER_56_3295 ();
 sg13g2_decap_8 FILLER_56_3302 ();
 sg13g2_decap_8 FILLER_56_3309 ();
 sg13g2_decap_8 FILLER_56_3316 ();
 sg13g2_decap_8 FILLER_56_3323 ();
 sg13g2_decap_8 FILLER_56_3330 ();
 sg13g2_decap_8 FILLER_56_3337 ();
 sg13g2_decap_8 FILLER_56_3344 ();
 sg13g2_decap_8 FILLER_56_3351 ();
 sg13g2_decap_8 FILLER_56_3358 ();
 sg13g2_decap_8 FILLER_56_3365 ();
 sg13g2_decap_8 FILLER_56_3372 ();
 sg13g2_decap_8 FILLER_56_3379 ();
 sg13g2_decap_8 FILLER_56_3386 ();
 sg13g2_decap_8 FILLER_56_3393 ();
 sg13g2_decap_8 FILLER_56_3400 ();
 sg13g2_decap_8 FILLER_56_3407 ();
 sg13g2_decap_8 FILLER_56_3414 ();
 sg13g2_decap_8 FILLER_56_3421 ();
 sg13g2_decap_8 FILLER_56_3428 ();
 sg13g2_decap_8 FILLER_56_3435 ();
 sg13g2_decap_8 FILLER_56_3442 ();
 sg13g2_decap_8 FILLER_56_3449 ();
 sg13g2_decap_8 FILLER_56_3456 ();
 sg13g2_decap_8 FILLER_56_3463 ();
 sg13g2_decap_8 FILLER_56_3470 ();
 sg13g2_decap_8 FILLER_56_3477 ();
 sg13g2_decap_8 FILLER_56_3484 ();
 sg13g2_decap_8 FILLER_56_3491 ();
 sg13g2_decap_8 FILLER_56_3498 ();
 sg13g2_decap_8 FILLER_56_3505 ();
 sg13g2_decap_8 FILLER_56_3512 ();
 sg13g2_decap_8 FILLER_56_3519 ();
 sg13g2_decap_8 FILLER_56_3526 ();
 sg13g2_decap_8 FILLER_56_3533 ();
 sg13g2_decap_8 FILLER_56_3540 ();
 sg13g2_decap_8 FILLER_56_3547 ();
 sg13g2_decap_8 FILLER_56_3554 ();
 sg13g2_decap_8 FILLER_56_3561 ();
 sg13g2_decap_8 FILLER_56_3568 ();
 sg13g2_decap_4 FILLER_56_3575 ();
 sg13g2_fill_1 FILLER_56_3579 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_decap_8 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_231 ();
 sg13g2_decap_8 FILLER_57_238 ();
 sg13g2_decap_8 FILLER_57_245 ();
 sg13g2_decap_8 FILLER_57_252 ();
 sg13g2_decap_8 FILLER_57_259 ();
 sg13g2_decap_8 FILLER_57_266 ();
 sg13g2_decap_8 FILLER_57_273 ();
 sg13g2_decap_8 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_287 ();
 sg13g2_decap_8 FILLER_57_294 ();
 sg13g2_decap_8 FILLER_57_301 ();
 sg13g2_decap_8 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_decap_8 FILLER_57_322 ();
 sg13g2_decap_8 FILLER_57_329 ();
 sg13g2_decap_8 FILLER_57_336 ();
 sg13g2_decap_8 FILLER_57_343 ();
 sg13g2_decap_8 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_364 ();
 sg13g2_decap_8 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_4 FILLER_57_385 ();
 sg13g2_fill_1 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_57_452 ();
 sg13g2_fill_2 FILLER_57_459 ();
 sg13g2_decap_4 FILLER_57_549 ();
 sg13g2_fill_2 FILLER_57_553 ();
 sg13g2_fill_2 FILLER_57_584 ();
 sg13g2_decap_8 FILLER_57_643 ();
 sg13g2_decap_8 FILLER_57_650 ();
 sg13g2_fill_2 FILLER_57_657 ();
 sg13g2_fill_1 FILLER_57_659 ();
 sg13g2_decap_8 FILLER_57_665 ();
 sg13g2_decap_4 FILLER_57_672 ();
 sg13g2_fill_1 FILLER_57_676 ();
 sg13g2_fill_2 FILLER_57_711 ();
 sg13g2_decap_8 FILLER_57_750 ();
 sg13g2_fill_2 FILLER_57_881 ();
 sg13g2_fill_1 FILLER_57_883 ();
 sg13g2_fill_1 FILLER_57_905 ();
 sg13g2_decap_8 FILLER_57_914 ();
 sg13g2_decap_8 FILLER_57_921 ();
 sg13g2_fill_1 FILLER_57_928 ();
 sg13g2_decap_8 FILLER_57_933 ();
 sg13g2_decap_8 FILLER_57_940 ();
 sg13g2_decap_8 FILLER_57_947 ();
 sg13g2_fill_1 FILLER_57_954 ();
 sg13g2_fill_1 FILLER_57_958 ();
 sg13g2_fill_1 FILLER_57_988 ();
 sg13g2_decap_8 FILLER_57_1054 ();
 sg13g2_decap_8 FILLER_57_1061 ();
 sg13g2_decap_8 FILLER_57_1068 ();
 sg13g2_decap_8 FILLER_57_1075 ();
 sg13g2_decap_8 FILLER_57_1134 ();
 sg13g2_decap_8 FILLER_57_1141 ();
 sg13g2_decap_8 FILLER_57_1174 ();
 sg13g2_decap_4 FILLER_57_1181 ();
 sg13g2_fill_1 FILLER_57_1185 ();
 sg13g2_decap_4 FILLER_57_1295 ();
 sg13g2_fill_1 FILLER_57_1299 ();
 sg13g2_decap_8 FILLER_57_1305 ();
 sg13g2_decap_8 FILLER_57_1312 ();
 sg13g2_decap_8 FILLER_57_1319 ();
 sg13g2_fill_2 FILLER_57_1326 ();
 sg13g2_fill_1 FILLER_57_1328 ();
 sg13g2_decap_8 FILLER_57_1355 ();
 sg13g2_decap_8 FILLER_57_1362 ();
 sg13g2_fill_1 FILLER_57_1407 ();
 sg13g2_decap_8 FILLER_57_1439 ();
 sg13g2_decap_8 FILLER_57_1446 ();
 sg13g2_decap_8 FILLER_57_1453 ();
 sg13g2_decap_8 FILLER_57_1460 ();
 sg13g2_decap_4 FILLER_57_1467 ();
 sg13g2_decap_8 FILLER_57_1497 ();
 sg13g2_decap_8 FILLER_57_1504 ();
 sg13g2_decap_8 FILLER_57_1511 ();
 sg13g2_decap_8 FILLER_57_1518 ();
 sg13g2_fill_1 FILLER_57_1525 ();
 sg13g2_fill_2 FILLER_57_1558 ();
 sg13g2_decap_8 FILLER_57_1567 ();
 sg13g2_fill_1 FILLER_57_1574 ();
 sg13g2_decap_8 FILLER_57_1618 ();
 sg13g2_decap_8 FILLER_57_1625 ();
 sg13g2_fill_2 FILLER_57_1632 ();
 sg13g2_decap_8 FILLER_57_1639 ();
 sg13g2_fill_1 FILLER_57_1672 ();
 sg13g2_decap_8 FILLER_57_1732 ();
 sg13g2_decap_8 FILLER_57_1748 ();
 sg13g2_fill_2 FILLER_57_1755 ();
 sg13g2_fill_1 FILLER_57_1757 ();
 sg13g2_decap_4 FILLER_57_1822 ();
 sg13g2_decap_8 FILLER_57_1862 ();
 sg13g2_decap_8 FILLER_57_1869 ();
 sg13g2_decap_8 FILLER_57_1876 ();
 sg13g2_decap_8 FILLER_57_1912 ();
 sg13g2_decap_8 FILLER_57_1919 ();
 sg13g2_decap_8 FILLER_57_1926 ();
 sg13g2_decap_8 FILLER_57_1933 ();
 sg13g2_decap_4 FILLER_57_1940 ();
 sg13g2_fill_2 FILLER_57_1944 ();
 sg13g2_fill_1 FILLER_57_1972 ();
 sg13g2_fill_2 FILLER_57_2025 ();
 sg13g2_fill_2 FILLER_57_2035 ();
 sg13g2_decap_8 FILLER_57_2089 ();
 sg13g2_fill_2 FILLER_57_2096 ();
 sg13g2_fill_1 FILLER_57_2098 ();
 sg13g2_decap_8 FILLER_57_2104 ();
 sg13g2_decap_8 FILLER_57_2111 ();
 sg13g2_decap_8 FILLER_57_2155 ();
 sg13g2_decap_8 FILLER_57_2162 ();
 sg13g2_decap_8 FILLER_57_2169 ();
 sg13g2_decap_8 FILLER_57_2176 ();
 sg13g2_fill_2 FILLER_57_2183 ();
 sg13g2_fill_1 FILLER_57_2185 ();
 sg13g2_decap_8 FILLER_57_2212 ();
 sg13g2_decap_8 FILLER_57_2227 ();
 sg13g2_decap_8 FILLER_57_2234 ();
 sg13g2_decap_8 FILLER_57_2241 ();
 sg13g2_decap_8 FILLER_57_2248 ();
 sg13g2_decap_8 FILLER_57_2255 ();
 sg13g2_decap_8 FILLER_57_2262 ();
 sg13g2_decap_8 FILLER_57_2269 ();
 sg13g2_decap_8 FILLER_57_2276 ();
 sg13g2_decap_8 FILLER_57_2283 ();
 sg13g2_decap_8 FILLER_57_2290 ();
 sg13g2_decap_8 FILLER_57_2297 ();
 sg13g2_decap_8 FILLER_57_2304 ();
 sg13g2_decap_8 FILLER_57_2311 ();
 sg13g2_decap_8 FILLER_57_2318 ();
 sg13g2_decap_8 FILLER_57_2325 ();
 sg13g2_decap_8 FILLER_57_2332 ();
 sg13g2_decap_8 FILLER_57_2339 ();
 sg13g2_decap_8 FILLER_57_2346 ();
 sg13g2_decap_8 FILLER_57_2353 ();
 sg13g2_decap_8 FILLER_57_2360 ();
 sg13g2_decap_4 FILLER_57_2367 ();
 sg13g2_fill_2 FILLER_57_2371 ();
 sg13g2_decap_8 FILLER_57_2399 ();
 sg13g2_fill_2 FILLER_57_2406 ();
 sg13g2_fill_1 FILLER_57_2408 ();
 sg13g2_decap_4 FILLER_57_2461 ();
 sg13g2_fill_1 FILLER_57_2465 ();
 sg13g2_decap_8 FILLER_57_2492 ();
 sg13g2_decap_8 FILLER_57_2499 ();
 sg13g2_decap_8 FILLER_57_2506 ();
 sg13g2_decap_8 FILLER_57_2513 ();
 sg13g2_decap_8 FILLER_57_2582 ();
 sg13g2_fill_1 FILLER_57_2589 ();
 sg13g2_decap_4 FILLER_57_2616 ();
 sg13g2_fill_2 FILLER_57_2626 ();
 sg13g2_fill_1 FILLER_57_2628 ();
 sg13g2_decap_8 FILLER_57_2643 ();
 sg13g2_decap_8 FILLER_57_2650 ();
 sg13g2_decap_8 FILLER_57_2657 ();
 sg13g2_decap_8 FILLER_57_2664 ();
 sg13g2_decap_4 FILLER_57_2671 ();
 sg13g2_fill_1 FILLER_57_2675 ();
 sg13g2_fill_1 FILLER_57_2702 ();
 sg13g2_decap_4 FILLER_57_2709 ();
 sg13g2_decap_8 FILLER_57_2729 ();
 sg13g2_fill_2 FILLER_57_2736 ();
 sg13g2_fill_2 FILLER_57_2776 ();
 sg13g2_decap_8 FILLER_57_2814 ();
 sg13g2_decap_4 FILLER_57_2821 ();
 sg13g2_fill_2 FILLER_57_2836 ();
 sg13g2_fill_1 FILLER_57_2838 ();
 sg13g2_decap_8 FILLER_57_2870 ();
 sg13g2_decap_8 FILLER_57_2877 ();
 sg13g2_decap_8 FILLER_57_2884 ();
 sg13g2_fill_2 FILLER_57_2891 ();
 sg13g2_fill_2 FILLER_57_2950 ();
 sg13g2_fill_1 FILLER_57_2952 ();
 sg13g2_decap_8 FILLER_57_2987 ();
 sg13g2_decap_4 FILLER_57_2994 ();
 sg13g2_fill_2 FILLER_57_2998 ();
 sg13g2_decap_8 FILLER_57_3026 ();
 sg13g2_decap_8 FILLER_57_3033 ();
 sg13g2_decap_8 FILLER_57_3040 ();
 sg13g2_decap_8 FILLER_57_3047 ();
 sg13g2_decap_8 FILLER_57_3054 ();
 sg13g2_decap_8 FILLER_57_3061 ();
 sg13g2_decap_8 FILLER_57_3068 ();
 sg13g2_decap_8 FILLER_57_3075 ();
 sg13g2_decap_8 FILLER_57_3082 ();
 sg13g2_decap_8 FILLER_57_3089 ();
 sg13g2_decap_8 FILLER_57_3096 ();
 sg13g2_decap_8 FILLER_57_3103 ();
 sg13g2_decap_8 FILLER_57_3110 ();
 sg13g2_decap_8 FILLER_57_3117 ();
 sg13g2_decap_8 FILLER_57_3124 ();
 sg13g2_decap_8 FILLER_57_3131 ();
 sg13g2_decap_8 FILLER_57_3138 ();
 sg13g2_decap_8 FILLER_57_3145 ();
 sg13g2_decap_8 FILLER_57_3152 ();
 sg13g2_decap_8 FILLER_57_3159 ();
 sg13g2_decap_8 FILLER_57_3166 ();
 sg13g2_decap_8 FILLER_57_3173 ();
 sg13g2_decap_8 FILLER_57_3180 ();
 sg13g2_decap_8 FILLER_57_3187 ();
 sg13g2_decap_8 FILLER_57_3194 ();
 sg13g2_decap_8 FILLER_57_3201 ();
 sg13g2_decap_8 FILLER_57_3208 ();
 sg13g2_decap_8 FILLER_57_3215 ();
 sg13g2_decap_8 FILLER_57_3222 ();
 sg13g2_decap_8 FILLER_57_3229 ();
 sg13g2_decap_8 FILLER_57_3236 ();
 sg13g2_decap_8 FILLER_57_3243 ();
 sg13g2_decap_8 FILLER_57_3250 ();
 sg13g2_decap_8 FILLER_57_3257 ();
 sg13g2_decap_8 FILLER_57_3264 ();
 sg13g2_decap_8 FILLER_57_3271 ();
 sg13g2_decap_8 FILLER_57_3278 ();
 sg13g2_decap_8 FILLER_57_3285 ();
 sg13g2_decap_8 FILLER_57_3292 ();
 sg13g2_decap_8 FILLER_57_3299 ();
 sg13g2_decap_8 FILLER_57_3306 ();
 sg13g2_decap_8 FILLER_57_3313 ();
 sg13g2_decap_8 FILLER_57_3320 ();
 sg13g2_decap_8 FILLER_57_3327 ();
 sg13g2_decap_8 FILLER_57_3334 ();
 sg13g2_decap_8 FILLER_57_3341 ();
 sg13g2_decap_8 FILLER_57_3348 ();
 sg13g2_decap_8 FILLER_57_3355 ();
 sg13g2_decap_8 FILLER_57_3362 ();
 sg13g2_decap_8 FILLER_57_3369 ();
 sg13g2_decap_8 FILLER_57_3376 ();
 sg13g2_decap_8 FILLER_57_3383 ();
 sg13g2_decap_8 FILLER_57_3390 ();
 sg13g2_decap_8 FILLER_57_3397 ();
 sg13g2_decap_8 FILLER_57_3404 ();
 sg13g2_decap_8 FILLER_57_3411 ();
 sg13g2_decap_8 FILLER_57_3418 ();
 sg13g2_decap_8 FILLER_57_3425 ();
 sg13g2_decap_8 FILLER_57_3432 ();
 sg13g2_decap_8 FILLER_57_3439 ();
 sg13g2_decap_8 FILLER_57_3446 ();
 sg13g2_decap_8 FILLER_57_3453 ();
 sg13g2_decap_8 FILLER_57_3460 ();
 sg13g2_decap_8 FILLER_57_3467 ();
 sg13g2_decap_8 FILLER_57_3474 ();
 sg13g2_decap_8 FILLER_57_3481 ();
 sg13g2_decap_8 FILLER_57_3488 ();
 sg13g2_decap_8 FILLER_57_3495 ();
 sg13g2_decap_8 FILLER_57_3502 ();
 sg13g2_decap_8 FILLER_57_3509 ();
 sg13g2_decap_8 FILLER_57_3516 ();
 sg13g2_decap_8 FILLER_57_3523 ();
 sg13g2_decap_8 FILLER_57_3530 ();
 sg13g2_decap_8 FILLER_57_3537 ();
 sg13g2_decap_8 FILLER_57_3544 ();
 sg13g2_decap_8 FILLER_57_3551 ();
 sg13g2_decap_8 FILLER_57_3558 ();
 sg13g2_decap_8 FILLER_57_3565 ();
 sg13g2_decap_8 FILLER_57_3572 ();
 sg13g2_fill_1 FILLER_57_3579 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_210 ();
 sg13g2_decap_8 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_224 ();
 sg13g2_decap_8 FILLER_58_231 ();
 sg13g2_decap_8 FILLER_58_238 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_decap_8 FILLER_58_252 ();
 sg13g2_decap_8 FILLER_58_259 ();
 sg13g2_decap_8 FILLER_58_266 ();
 sg13g2_decap_8 FILLER_58_273 ();
 sg13g2_decap_8 FILLER_58_280 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_8 FILLER_58_301 ();
 sg13g2_decap_8 FILLER_58_308 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_decap_8 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_343 ();
 sg13g2_decap_8 FILLER_58_350 ();
 sg13g2_decap_8 FILLER_58_357 ();
 sg13g2_decap_8 FILLER_58_364 ();
 sg13g2_decap_8 FILLER_58_371 ();
 sg13g2_decap_8 FILLER_58_378 ();
 sg13g2_decap_8 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_392 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_decap_8 FILLER_58_458 ();
 sg13g2_decap_4 FILLER_58_465 ();
 sg13g2_decap_4 FILLER_58_553 ();
 sg13g2_fill_1 FILLER_58_557 ();
 sg13g2_fill_1 FILLER_58_584 ();
 sg13g2_fill_2 FILLER_58_603 ();
 sg13g2_fill_1 FILLER_58_605 ();
 sg13g2_fill_2 FILLER_58_616 ();
 sg13g2_decap_8 FILLER_58_644 ();
 sg13g2_fill_2 FILLER_58_651 ();
 sg13g2_fill_1 FILLER_58_653 ();
 sg13g2_fill_2 FILLER_58_715 ();
 sg13g2_decap_8 FILLER_58_746 ();
 sg13g2_decap_8 FILLER_58_753 ();
 sg13g2_fill_2 FILLER_58_760 ();
 sg13g2_fill_1 FILLER_58_762 ();
 sg13g2_decap_8 FILLER_58_798 ();
 sg13g2_decap_4 FILLER_58_805 ();
 sg13g2_fill_1 FILLER_58_809 ();
 sg13g2_fill_2 FILLER_58_813 ();
 sg13g2_fill_1 FILLER_58_815 ();
 sg13g2_decap_4 FILLER_58_820 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_4 FILLER_58_835 ();
 sg13g2_fill_1 FILLER_58_842 ();
 sg13g2_fill_1 FILLER_58_852 ();
 sg13g2_decap_4 FILLER_58_858 ();
 sg13g2_decap_8 FILLER_58_867 ();
 sg13g2_fill_1 FILLER_58_874 ();
 sg13g2_decap_8 FILLER_58_878 ();
 sg13g2_decap_4 FILLER_58_885 ();
 sg13g2_fill_1 FILLER_58_889 ();
 sg13g2_fill_1 FILLER_58_895 ();
 sg13g2_decap_8 FILLER_58_899 ();
 sg13g2_fill_1 FILLER_58_919 ();
 sg13g2_decap_8 FILLER_58_946 ();
 sg13g2_decap_8 FILLER_58_953 ();
 sg13g2_decap_8 FILLER_58_960 ();
 sg13g2_fill_1 FILLER_58_967 ();
 sg13g2_decap_8 FILLER_58_973 ();
 sg13g2_fill_2 FILLER_58_980 ();
 sg13g2_fill_1 FILLER_58_982 ();
 sg13g2_fill_2 FILLER_58_1017 ();
 sg13g2_fill_1 FILLER_58_1019 ();
 sg13g2_decap_8 FILLER_58_1030 ();
 sg13g2_decap_8 FILLER_58_1037 ();
 sg13g2_fill_2 FILLER_58_1044 ();
 sg13g2_fill_1 FILLER_58_1046 ();
 sg13g2_fill_1 FILLER_58_1076 ();
 sg13g2_decap_8 FILLER_58_1129 ();
 sg13g2_fill_2 FILLER_58_1222 ();
 sg13g2_fill_1 FILLER_58_1224 ();
 sg13g2_fill_2 FILLER_58_1257 ();
 sg13g2_decap_8 FILLER_58_1291 ();
 sg13g2_decap_4 FILLER_58_1298 ();
 sg13g2_fill_1 FILLER_58_1302 ();
 sg13g2_fill_1 FILLER_58_1311 ();
 sg13g2_decap_8 FILLER_58_1317 ();
 sg13g2_decap_4 FILLER_58_1324 ();
 sg13g2_decap_8 FILLER_58_1354 ();
 sg13g2_decap_8 FILLER_58_1361 ();
 sg13g2_decap_8 FILLER_58_1368 ();
 sg13g2_fill_2 FILLER_58_1375 ();
 sg13g2_fill_1 FILLER_58_1377 ();
 sg13g2_fill_1 FILLER_58_1387 ();
 sg13g2_decap_8 FILLER_58_1445 ();
 sg13g2_decap_8 FILLER_58_1452 ();
 sg13g2_decap_8 FILLER_58_1459 ();
 sg13g2_decap_4 FILLER_58_1466 ();
 sg13g2_fill_2 FILLER_58_1470 ();
 sg13g2_decap_8 FILLER_58_1498 ();
 sg13g2_decap_8 FILLER_58_1505 ();
 sg13g2_decap_4 FILLER_58_1512 ();
 sg13g2_fill_2 FILLER_58_1516 ();
 sg13g2_fill_2 FILLER_58_1557 ();
 sg13g2_fill_1 FILLER_58_1572 ();
 sg13g2_decap_8 FILLER_58_1599 ();
 sg13g2_fill_1 FILLER_58_1606 ();
 sg13g2_fill_2 FILLER_58_1633 ();
 sg13g2_fill_1 FILLER_58_1635 ();
 sg13g2_decap_4 FILLER_58_1728 ();
 sg13g2_decap_8 FILLER_58_1808 ();
 sg13g2_decap_4 FILLER_58_1815 ();
 sg13g2_fill_1 FILLER_58_1819 ();
 sg13g2_decap_8 FILLER_58_1877 ();
 sg13g2_decap_8 FILLER_58_1884 ();
 sg13g2_decap_8 FILLER_58_1917 ();
 sg13g2_decap_8 FILLER_58_1924 ();
 sg13g2_fill_2 FILLER_58_1931 ();
 sg13g2_decap_4 FILLER_58_2037 ();
 sg13g2_fill_2 FILLER_58_2041 ();
 sg13g2_decap_4 FILLER_58_2048 ();
 sg13g2_decap_8 FILLER_58_2078 ();
 sg13g2_decap_4 FILLER_58_2085 ();
 sg13g2_fill_1 FILLER_58_2089 ();
 sg13g2_fill_2 FILLER_58_2121 ();
 sg13g2_fill_1 FILLER_58_2123 ();
 sg13g2_decap_4 FILLER_58_2132 ();
 sg13g2_fill_1 FILLER_58_2136 ();
 sg13g2_decap_8 FILLER_58_2168 ();
 sg13g2_fill_2 FILLER_58_2175 ();
 sg13g2_decap_8 FILLER_58_2242 ();
 sg13g2_decap_8 FILLER_58_2249 ();
 sg13g2_decap_8 FILLER_58_2256 ();
 sg13g2_decap_8 FILLER_58_2263 ();
 sg13g2_decap_8 FILLER_58_2270 ();
 sg13g2_decap_8 FILLER_58_2277 ();
 sg13g2_decap_8 FILLER_58_2284 ();
 sg13g2_decap_8 FILLER_58_2291 ();
 sg13g2_decap_8 FILLER_58_2298 ();
 sg13g2_decap_8 FILLER_58_2305 ();
 sg13g2_decap_8 FILLER_58_2312 ();
 sg13g2_decap_8 FILLER_58_2319 ();
 sg13g2_decap_8 FILLER_58_2326 ();
 sg13g2_decap_8 FILLER_58_2333 ();
 sg13g2_decap_8 FILLER_58_2340 ();
 sg13g2_decap_8 FILLER_58_2347 ();
 sg13g2_decap_8 FILLER_58_2354 ();
 sg13g2_decap_8 FILLER_58_2361 ();
 sg13g2_decap_8 FILLER_58_2368 ();
 sg13g2_decap_8 FILLER_58_2375 ();
 sg13g2_decap_8 FILLER_58_2382 ();
 sg13g2_decap_8 FILLER_58_2389 ();
 sg13g2_fill_1 FILLER_58_2396 ();
 sg13g2_decap_8 FILLER_58_2449 ();
 sg13g2_decap_8 FILLER_58_2456 ();
 sg13g2_decap_4 FILLER_58_2463 ();
 sg13g2_fill_2 FILLER_58_2467 ();
 sg13g2_decap_8 FILLER_58_2495 ();
 sg13g2_decap_8 FILLER_58_2502 ();
 sg13g2_decap_4 FILLER_58_2509 ();
 sg13g2_fill_2 FILLER_58_2539 ();
 sg13g2_fill_1 FILLER_58_2541 ();
 sg13g2_fill_2 FILLER_58_2568 ();
 sg13g2_fill_2 FILLER_58_2575 ();
 sg13g2_decap_4 FILLER_58_2660 ();
 sg13g2_fill_2 FILLER_58_2664 ();
 sg13g2_decap_8 FILLER_58_2674 ();
 sg13g2_decap_4 FILLER_58_2681 ();
 sg13g2_fill_1 FILLER_58_2685 ();
 sg13g2_decap_8 FILLER_58_2733 ();
 sg13g2_fill_2 FILLER_58_2740 ();
 sg13g2_fill_1 FILLER_58_2742 ();
 sg13g2_decap_8 FILLER_58_2775 ();
 sg13g2_fill_2 FILLER_58_2782 ();
 sg13g2_decap_8 FILLER_58_2810 ();
 sg13g2_decap_8 FILLER_58_2817 ();
 sg13g2_decap_8 FILLER_58_2824 ();
 sg13g2_fill_2 FILLER_58_2831 ();
 sg13g2_fill_1 FILLER_58_2833 ();
 sg13g2_decap_4 FILLER_58_2877 ();
 sg13g2_fill_2 FILLER_58_2881 ();
 sg13g2_fill_2 FILLER_58_2888 ();
 sg13g2_fill_1 FILLER_58_2890 ();
 sg13g2_decap_4 FILLER_58_2899 ();
 sg13g2_fill_1 FILLER_58_2903 ();
 sg13g2_decap_8 FILLER_58_2936 ();
 sg13g2_fill_2 FILLER_58_2943 ();
 sg13g2_fill_2 FILLER_58_2953 ();
 sg13g2_decap_8 FILLER_58_3033 ();
 sg13g2_decap_8 FILLER_58_3040 ();
 sg13g2_decap_8 FILLER_58_3047 ();
 sg13g2_decap_8 FILLER_58_3054 ();
 sg13g2_decap_8 FILLER_58_3061 ();
 sg13g2_decap_8 FILLER_58_3068 ();
 sg13g2_decap_8 FILLER_58_3075 ();
 sg13g2_decap_8 FILLER_58_3082 ();
 sg13g2_decap_8 FILLER_58_3089 ();
 sg13g2_decap_8 FILLER_58_3096 ();
 sg13g2_decap_8 FILLER_58_3103 ();
 sg13g2_decap_8 FILLER_58_3110 ();
 sg13g2_decap_8 FILLER_58_3117 ();
 sg13g2_decap_8 FILLER_58_3124 ();
 sg13g2_decap_8 FILLER_58_3131 ();
 sg13g2_decap_8 FILLER_58_3138 ();
 sg13g2_decap_8 FILLER_58_3145 ();
 sg13g2_decap_8 FILLER_58_3152 ();
 sg13g2_decap_8 FILLER_58_3159 ();
 sg13g2_decap_8 FILLER_58_3166 ();
 sg13g2_decap_8 FILLER_58_3173 ();
 sg13g2_decap_8 FILLER_58_3180 ();
 sg13g2_decap_8 FILLER_58_3187 ();
 sg13g2_decap_8 FILLER_58_3194 ();
 sg13g2_decap_8 FILLER_58_3201 ();
 sg13g2_decap_8 FILLER_58_3208 ();
 sg13g2_decap_8 FILLER_58_3215 ();
 sg13g2_decap_8 FILLER_58_3222 ();
 sg13g2_decap_8 FILLER_58_3229 ();
 sg13g2_decap_8 FILLER_58_3236 ();
 sg13g2_decap_8 FILLER_58_3243 ();
 sg13g2_decap_8 FILLER_58_3250 ();
 sg13g2_decap_8 FILLER_58_3257 ();
 sg13g2_decap_8 FILLER_58_3264 ();
 sg13g2_decap_8 FILLER_58_3271 ();
 sg13g2_decap_8 FILLER_58_3278 ();
 sg13g2_decap_8 FILLER_58_3285 ();
 sg13g2_decap_8 FILLER_58_3292 ();
 sg13g2_decap_8 FILLER_58_3299 ();
 sg13g2_decap_8 FILLER_58_3306 ();
 sg13g2_decap_8 FILLER_58_3313 ();
 sg13g2_decap_8 FILLER_58_3320 ();
 sg13g2_decap_8 FILLER_58_3327 ();
 sg13g2_decap_8 FILLER_58_3334 ();
 sg13g2_decap_8 FILLER_58_3341 ();
 sg13g2_decap_8 FILLER_58_3348 ();
 sg13g2_decap_8 FILLER_58_3355 ();
 sg13g2_decap_8 FILLER_58_3362 ();
 sg13g2_decap_8 FILLER_58_3369 ();
 sg13g2_decap_8 FILLER_58_3376 ();
 sg13g2_decap_8 FILLER_58_3383 ();
 sg13g2_decap_8 FILLER_58_3390 ();
 sg13g2_decap_8 FILLER_58_3397 ();
 sg13g2_decap_8 FILLER_58_3404 ();
 sg13g2_decap_8 FILLER_58_3411 ();
 sg13g2_decap_8 FILLER_58_3418 ();
 sg13g2_decap_8 FILLER_58_3425 ();
 sg13g2_decap_8 FILLER_58_3432 ();
 sg13g2_decap_8 FILLER_58_3439 ();
 sg13g2_decap_8 FILLER_58_3446 ();
 sg13g2_decap_8 FILLER_58_3453 ();
 sg13g2_decap_8 FILLER_58_3460 ();
 sg13g2_decap_8 FILLER_58_3467 ();
 sg13g2_decap_8 FILLER_58_3474 ();
 sg13g2_decap_8 FILLER_58_3481 ();
 sg13g2_decap_8 FILLER_58_3488 ();
 sg13g2_decap_8 FILLER_58_3495 ();
 sg13g2_decap_8 FILLER_58_3502 ();
 sg13g2_decap_8 FILLER_58_3509 ();
 sg13g2_decap_8 FILLER_58_3516 ();
 sg13g2_decap_8 FILLER_58_3523 ();
 sg13g2_decap_8 FILLER_58_3530 ();
 sg13g2_decap_8 FILLER_58_3537 ();
 sg13g2_decap_8 FILLER_58_3544 ();
 sg13g2_decap_8 FILLER_58_3551 ();
 sg13g2_decap_8 FILLER_58_3558 ();
 sg13g2_decap_8 FILLER_58_3565 ();
 sg13g2_decap_8 FILLER_58_3572 ();
 sg13g2_fill_1 FILLER_58_3579 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_decap_8 FILLER_59_210 ();
 sg13g2_decap_8 FILLER_59_217 ();
 sg13g2_decap_8 FILLER_59_224 ();
 sg13g2_decap_8 FILLER_59_231 ();
 sg13g2_decap_8 FILLER_59_238 ();
 sg13g2_decap_8 FILLER_59_245 ();
 sg13g2_decap_8 FILLER_59_252 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_decap_8 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_decap_8 FILLER_59_287 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_301 ();
 sg13g2_decap_8 FILLER_59_308 ();
 sg13g2_decap_8 FILLER_59_315 ();
 sg13g2_decap_8 FILLER_59_322 ();
 sg13g2_decap_8 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_336 ();
 sg13g2_decap_8 FILLER_59_343 ();
 sg13g2_decap_8 FILLER_59_350 ();
 sg13g2_decap_8 FILLER_59_357 ();
 sg13g2_decap_8 FILLER_59_364 ();
 sg13g2_decap_8 FILLER_59_371 ();
 sg13g2_decap_8 FILLER_59_378 ();
 sg13g2_decap_8 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_406 ();
 sg13g2_fill_2 FILLER_59_413 ();
 sg13g2_decap_8 FILLER_59_440 ();
 sg13g2_decap_8 FILLER_59_447 ();
 sg13g2_decap_8 FILLER_59_454 ();
 sg13g2_decap_8 FILLER_59_461 ();
 sg13g2_decap_8 FILLER_59_468 ();
 sg13g2_decap_4 FILLER_59_475 ();
 sg13g2_decap_8 FILLER_59_550 ();
 sg13g2_decap_8 FILLER_59_557 ();
 sg13g2_decap_4 FILLER_59_564 ();
 sg13g2_fill_1 FILLER_59_568 ();
 sg13g2_fill_1 FILLER_59_608 ();
 sg13g2_fill_2 FILLER_59_614 ();
 sg13g2_fill_1 FILLER_59_616 ();
 sg13g2_decap_8 FILLER_59_643 ();
 sg13g2_decap_8 FILLER_59_650 ();
 sg13g2_decap_8 FILLER_59_657 ();
 sg13g2_fill_1 FILLER_59_664 ();
 sg13g2_decap_8 FILLER_59_669 ();
 sg13g2_fill_1 FILLER_59_680 ();
 sg13g2_decap_4 FILLER_59_684 ();
 sg13g2_fill_2 FILLER_59_688 ();
 sg13g2_decap_8 FILLER_59_694 ();
 sg13g2_decap_8 FILLER_59_701 ();
 sg13g2_decap_8 FILLER_59_708 ();
 sg13g2_decap_4 FILLER_59_715 ();
 sg13g2_fill_2 FILLER_59_719 ();
 sg13g2_fill_1 FILLER_59_731 ();
 sg13g2_decap_8 FILLER_59_737 ();
 sg13g2_decap_8 FILLER_59_749 ();
 sg13g2_decap_8 FILLER_59_756 ();
 sg13g2_decap_8 FILLER_59_763 ();
 sg13g2_decap_4 FILLER_59_774 ();
 sg13g2_fill_1 FILLER_59_778 ();
 sg13g2_fill_1 FILLER_59_783 ();
 sg13g2_decap_8 FILLER_59_793 ();
 sg13g2_decap_8 FILLER_59_800 ();
 sg13g2_decap_8 FILLER_59_807 ();
 sg13g2_decap_8 FILLER_59_814 ();
 sg13g2_decap_8 FILLER_59_821 ();
 sg13g2_decap_8 FILLER_59_828 ();
 sg13g2_decap_8 FILLER_59_835 ();
 sg13g2_fill_2 FILLER_59_842 ();
 sg13g2_fill_1 FILLER_59_844 ();
 sg13g2_decap_8 FILLER_59_848 ();
 sg13g2_decap_8 FILLER_59_855 ();
 sg13g2_fill_2 FILLER_59_862 ();
 sg13g2_fill_1 FILLER_59_864 ();
 sg13g2_fill_2 FILLER_59_891 ();
 sg13g2_decap_8 FILLER_59_936 ();
 sg13g2_decap_4 FILLER_59_943 ();
 sg13g2_decap_8 FILLER_59_973 ();
 sg13g2_decap_8 FILLER_59_980 ();
 sg13g2_decap_4 FILLER_59_987 ();
 sg13g2_fill_1 FILLER_59_991 ();
 sg13g2_fill_1 FILLER_59_1017 ();
 sg13g2_decap_8 FILLER_59_1023 ();
 sg13g2_decap_8 FILLER_59_1030 ();
 sg13g2_fill_2 FILLER_59_1177 ();
 sg13g2_fill_1 FILLER_59_1179 ();
 sg13g2_decap_8 FILLER_59_1224 ();
 sg13g2_fill_2 FILLER_59_1231 ();
 sg13g2_decap_8 FILLER_59_1247 ();
 sg13g2_decap_8 FILLER_59_1254 ();
 sg13g2_fill_2 FILLER_59_1272 ();
 sg13g2_fill_1 FILLER_59_1274 ();
 sg13g2_fill_2 FILLER_59_1301 ();
 sg13g2_fill_1 FILLER_59_1355 ();
 sg13g2_decap_8 FILLER_59_1382 ();
 sg13g2_decap_8 FILLER_59_1389 ();
 sg13g2_decap_4 FILLER_59_1396 ();
 sg13g2_fill_2 FILLER_59_1400 ();
 sg13g2_decap_8 FILLER_59_1454 ();
 sg13g2_fill_1 FILLER_59_1461 ();
 sg13g2_decap_8 FILLER_59_1502 ();
 sg13g2_fill_2 FILLER_59_1509 ();
 sg13g2_fill_1 FILLER_59_1511 ();
 sg13g2_decap_8 FILLER_59_1604 ();
 sg13g2_decap_8 FILLER_59_1611 ();
 sg13g2_decap_8 FILLER_59_1622 ();
 sg13g2_decap_4 FILLER_59_1629 ();
 sg13g2_fill_2 FILLER_59_1633 ();
 sg13g2_fill_1 FILLER_59_1644 ();
 sg13g2_decap_8 FILLER_59_1658 ();
 sg13g2_decap_8 FILLER_59_1665 ();
 sg13g2_decap_8 FILLER_59_1672 ();
 sg13g2_decap_8 FILLER_59_1679 ();
 sg13g2_decap_8 FILLER_59_1686 ();
 sg13g2_decap_4 FILLER_59_1693 ();
 sg13g2_decap_4 FILLER_59_1703 ();
 sg13g2_decap_8 FILLER_59_1721 ();
 sg13g2_decap_4 FILLER_59_1728 ();
 sg13g2_fill_2 FILLER_59_1732 ();
 sg13g2_decap_8 FILLER_59_1750 ();
 sg13g2_decap_8 FILLER_59_1757 ();
 sg13g2_decap_8 FILLER_59_1764 ();
 sg13g2_fill_2 FILLER_59_1771 ();
 sg13g2_fill_1 FILLER_59_1773 ();
 sg13g2_fill_1 FILLER_59_1787 ();
 sg13g2_decap_8 FILLER_59_1812 ();
 sg13g2_decap_8 FILLER_59_1819 ();
 sg13g2_decap_8 FILLER_59_1826 ();
 sg13g2_fill_2 FILLER_59_1833 ();
 sg13g2_fill_1 FILLER_59_1835 ();
 sg13g2_decap_8 FILLER_59_1852 ();
 sg13g2_decap_4 FILLER_59_1859 ();
 sg13g2_fill_2 FILLER_59_1863 ();
 sg13g2_fill_2 FILLER_59_1894 ();
 sg13g2_decap_4 FILLER_59_1904 ();
 sg13g2_fill_1 FILLER_59_1970 ();
 sg13g2_decap_8 FILLER_59_1981 ();
 sg13g2_fill_2 FILLER_59_1988 ();
 sg13g2_decap_8 FILLER_59_2038 ();
 sg13g2_decap_4 FILLER_59_2045 ();
 sg13g2_decap_4 FILLER_59_2064 ();
 sg13g2_fill_1 FILLER_59_2068 ();
 sg13g2_decap_8 FILLER_59_2119 ();
 sg13g2_fill_1 FILLER_59_2126 ();
 sg13g2_fill_1 FILLER_59_2167 ();
 sg13g2_decap_8 FILLER_59_2175 ();
 sg13g2_decap_8 FILLER_59_2182 ();
 sg13g2_fill_1 FILLER_59_2189 ();
 sg13g2_decap_8 FILLER_59_2242 ();
 sg13g2_decap_8 FILLER_59_2249 ();
 sg13g2_decap_8 FILLER_59_2256 ();
 sg13g2_decap_8 FILLER_59_2263 ();
 sg13g2_decap_8 FILLER_59_2270 ();
 sg13g2_decap_8 FILLER_59_2277 ();
 sg13g2_decap_8 FILLER_59_2284 ();
 sg13g2_decap_8 FILLER_59_2291 ();
 sg13g2_decap_8 FILLER_59_2298 ();
 sg13g2_decap_8 FILLER_59_2305 ();
 sg13g2_decap_8 FILLER_59_2312 ();
 sg13g2_decap_8 FILLER_59_2319 ();
 sg13g2_decap_8 FILLER_59_2326 ();
 sg13g2_decap_8 FILLER_59_2333 ();
 sg13g2_decap_8 FILLER_59_2340 ();
 sg13g2_decap_8 FILLER_59_2347 ();
 sg13g2_decap_8 FILLER_59_2354 ();
 sg13g2_decap_8 FILLER_59_2361 ();
 sg13g2_decap_8 FILLER_59_2368 ();
 sg13g2_decap_8 FILLER_59_2375 ();
 sg13g2_decap_8 FILLER_59_2382 ();
 sg13g2_decap_8 FILLER_59_2389 ();
 sg13g2_decap_8 FILLER_59_2396 ();
 sg13g2_decap_8 FILLER_59_2403 ();
 sg13g2_decap_8 FILLER_59_2410 ();
 sg13g2_decap_8 FILLER_59_2417 ();
 sg13g2_decap_8 FILLER_59_2450 ();
 sg13g2_decap_8 FILLER_59_2457 ();
 sg13g2_decap_8 FILLER_59_2464 ();
 sg13g2_decap_8 FILLER_59_2471 ();
 sg13g2_decap_8 FILLER_59_2478 ();
 sg13g2_decap_8 FILLER_59_2485 ();
 sg13g2_decap_8 FILLER_59_2492 ();
 sg13g2_decap_8 FILLER_59_2499 ();
 sg13g2_decap_8 FILLER_59_2506 ();
 sg13g2_decap_8 FILLER_59_2513 ();
 sg13g2_fill_2 FILLER_59_2520 ();
 sg13g2_fill_1 FILLER_59_2522 ();
 sg13g2_fill_2 FILLER_59_2549 ();
 sg13g2_fill_1 FILLER_59_2603 ();
 sg13g2_decap_8 FILLER_59_2662 ();
 sg13g2_decap_8 FILLER_59_2669 ();
 sg13g2_decap_8 FILLER_59_2676 ();
 sg13g2_decap_4 FILLER_59_2683 ();
 sg13g2_fill_2 FILLER_59_2687 ();
 sg13g2_decap_8 FILLER_59_2741 ();
 sg13g2_decap_8 FILLER_59_2748 ();
 sg13g2_fill_1 FILLER_59_2760 ();
 sg13g2_decap_8 FILLER_59_2771 ();
 sg13g2_decap_8 FILLER_59_2778 ();
 sg13g2_fill_2 FILLER_59_2785 ();
 sg13g2_decap_8 FILLER_59_2821 ();
 sg13g2_decap_8 FILLER_59_2828 ();
 sg13g2_decap_8 FILLER_59_2835 ();
 sg13g2_fill_2 FILLER_59_2842 ();
 sg13g2_decap_4 FILLER_59_2896 ();
 sg13g2_fill_2 FILLER_59_2958 ();
 sg13g2_fill_1 FILLER_59_2960 ();
 sg13g2_fill_2 FILLER_59_2966 ();
 sg13g2_fill_1 FILLER_59_2968 ();
 sg13g2_decap_8 FILLER_59_3029 ();
 sg13g2_decap_8 FILLER_59_3036 ();
 sg13g2_decap_8 FILLER_59_3043 ();
 sg13g2_decap_8 FILLER_59_3050 ();
 sg13g2_decap_8 FILLER_59_3057 ();
 sg13g2_decap_8 FILLER_59_3064 ();
 sg13g2_decap_8 FILLER_59_3071 ();
 sg13g2_decap_8 FILLER_59_3078 ();
 sg13g2_decap_8 FILLER_59_3085 ();
 sg13g2_decap_8 FILLER_59_3092 ();
 sg13g2_decap_8 FILLER_59_3099 ();
 sg13g2_decap_8 FILLER_59_3106 ();
 sg13g2_decap_8 FILLER_59_3113 ();
 sg13g2_decap_8 FILLER_59_3120 ();
 sg13g2_decap_8 FILLER_59_3127 ();
 sg13g2_decap_8 FILLER_59_3134 ();
 sg13g2_decap_8 FILLER_59_3141 ();
 sg13g2_decap_8 FILLER_59_3148 ();
 sg13g2_decap_8 FILLER_59_3155 ();
 sg13g2_decap_8 FILLER_59_3162 ();
 sg13g2_decap_8 FILLER_59_3169 ();
 sg13g2_decap_8 FILLER_59_3176 ();
 sg13g2_decap_8 FILLER_59_3183 ();
 sg13g2_decap_8 FILLER_59_3190 ();
 sg13g2_decap_8 FILLER_59_3197 ();
 sg13g2_decap_8 FILLER_59_3204 ();
 sg13g2_decap_8 FILLER_59_3211 ();
 sg13g2_decap_8 FILLER_59_3218 ();
 sg13g2_decap_8 FILLER_59_3225 ();
 sg13g2_decap_8 FILLER_59_3232 ();
 sg13g2_decap_8 FILLER_59_3239 ();
 sg13g2_decap_8 FILLER_59_3246 ();
 sg13g2_decap_8 FILLER_59_3253 ();
 sg13g2_decap_8 FILLER_59_3260 ();
 sg13g2_decap_8 FILLER_59_3267 ();
 sg13g2_decap_8 FILLER_59_3274 ();
 sg13g2_decap_8 FILLER_59_3281 ();
 sg13g2_decap_8 FILLER_59_3288 ();
 sg13g2_decap_8 FILLER_59_3295 ();
 sg13g2_decap_8 FILLER_59_3302 ();
 sg13g2_decap_8 FILLER_59_3309 ();
 sg13g2_decap_8 FILLER_59_3316 ();
 sg13g2_decap_8 FILLER_59_3323 ();
 sg13g2_decap_8 FILLER_59_3330 ();
 sg13g2_decap_8 FILLER_59_3337 ();
 sg13g2_decap_8 FILLER_59_3344 ();
 sg13g2_decap_8 FILLER_59_3351 ();
 sg13g2_decap_8 FILLER_59_3358 ();
 sg13g2_decap_8 FILLER_59_3365 ();
 sg13g2_decap_8 FILLER_59_3372 ();
 sg13g2_decap_8 FILLER_59_3379 ();
 sg13g2_decap_8 FILLER_59_3386 ();
 sg13g2_decap_8 FILLER_59_3393 ();
 sg13g2_decap_8 FILLER_59_3400 ();
 sg13g2_decap_8 FILLER_59_3407 ();
 sg13g2_decap_8 FILLER_59_3414 ();
 sg13g2_decap_8 FILLER_59_3421 ();
 sg13g2_decap_8 FILLER_59_3428 ();
 sg13g2_decap_8 FILLER_59_3435 ();
 sg13g2_decap_8 FILLER_59_3442 ();
 sg13g2_decap_8 FILLER_59_3449 ();
 sg13g2_decap_8 FILLER_59_3456 ();
 sg13g2_decap_8 FILLER_59_3463 ();
 sg13g2_decap_8 FILLER_59_3470 ();
 sg13g2_decap_8 FILLER_59_3477 ();
 sg13g2_decap_8 FILLER_59_3484 ();
 sg13g2_decap_8 FILLER_59_3491 ();
 sg13g2_decap_8 FILLER_59_3498 ();
 sg13g2_decap_8 FILLER_59_3505 ();
 sg13g2_decap_8 FILLER_59_3512 ();
 sg13g2_decap_8 FILLER_59_3519 ();
 sg13g2_decap_8 FILLER_59_3526 ();
 sg13g2_decap_8 FILLER_59_3533 ();
 sg13g2_decap_8 FILLER_59_3540 ();
 sg13g2_decap_8 FILLER_59_3547 ();
 sg13g2_decap_8 FILLER_59_3554 ();
 sg13g2_decap_8 FILLER_59_3561 ();
 sg13g2_decap_8 FILLER_59_3568 ();
 sg13g2_decap_4 FILLER_59_3575 ();
 sg13g2_fill_1 FILLER_59_3579 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_196 ();
 sg13g2_decap_8 FILLER_60_203 ();
 sg13g2_decap_8 FILLER_60_210 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_decap_8 FILLER_60_245 ();
 sg13g2_decap_8 FILLER_60_252 ();
 sg13g2_decap_8 FILLER_60_259 ();
 sg13g2_decap_8 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_decap_8 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_294 ();
 sg13g2_decap_8 FILLER_60_301 ();
 sg13g2_decap_8 FILLER_60_308 ();
 sg13g2_decap_8 FILLER_60_315 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_343 ();
 sg13g2_decap_8 FILLER_60_350 ();
 sg13g2_decap_8 FILLER_60_357 ();
 sg13g2_decap_8 FILLER_60_364 ();
 sg13g2_decap_8 FILLER_60_371 ();
 sg13g2_decap_8 FILLER_60_378 ();
 sg13g2_decap_8 FILLER_60_385 ();
 sg13g2_decap_8 FILLER_60_392 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_decap_8 FILLER_60_406 ();
 sg13g2_decap_8 FILLER_60_413 ();
 sg13g2_fill_1 FILLER_60_440 ();
 sg13g2_decap_8 FILLER_60_467 ();
 sg13g2_fill_2 FILLER_60_474 ();
 sg13g2_fill_1 FILLER_60_476 ();
 sg13g2_decap_8 FILLER_60_516 ();
 sg13g2_decap_8 FILLER_60_523 ();
 sg13g2_decap_8 FILLER_60_530 ();
 sg13g2_decap_8 FILLER_60_537 ();
 sg13g2_decap_8 FILLER_60_544 ();
 sg13g2_decap_8 FILLER_60_551 ();
 sg13g2_fill_2 FILLER_60_584 ();
 sg13g2_decap_8 FILLER_60_637 ();
 sg13g2_decap_8 FILLER_60_644 ();
 sg13g2_decap_8 FILLER_60_651 ();
 sg13g2_decap_8 FILLER_60_658 ();
 sg13g2_fill_2 FILLER_60_694 ();
 sg13g2_fill_1 FILLER_60_696 ();
 sg13g2_decap_8 FILLER_60_704 ();
 sg13g2_decap_4 FILLER_60_711 ();
 sg13g2_fill_2 FILLER_60_715 ();
 sg13g2_fill_1 FILLER_60_748 ();
 sg13g2_decap_8 FILLER_60_757 ();
 sg13g2_decap_4 FILLER_60_764 ();
 sg13g2_fill_1 FILLER_60_768 ();
 sg13g2_decap_8 FILLER_60_799 ();
 sg13g2_decap_4 FILLER_60_806 ();
 sg13g2_fill_2 FILLER_60_810 ();
 sg13g2_decap_4 FILLER_60_838 ();
 sg13g2_fill_1 FILLER_60_868 ();
 sg13g2_fill_1 FILLER_60_899 ();
 sg13g2_decap_8 FILLER_60_929 ();
 sg13g2_decap_8 FILLER_60_936 ();
 sg13g2_decap_4 FILLER_60_943 ();
 sg13g2_fill_2 FILLER_60_947 ();
 sg13g2_decap_8 FILLER_60_979 ();
 sg13g2_decap_4 FILLER_60_986 ();
 sg13g2_fill_2 FILLER_60_1027 ();
 sg13g2_fill_1 FILLER_60_1029 ();
 sg13g2_fill_1 FILLER_60_1077 ();
 sg13g2_decap_8 FILLER_60_1083 ();
 sg13g2_fill_1 FILLER_60_1090 ();
 sg13g2_fill_1 FILLER_60_1121 ();
 sg13g2_fill_1 FILLER_60_1127 ();
 sg13g2_decap_8 FILLER_60_1162 ();
 sg13g2_decap_4 FILLER_60_1195 ();
 sg13g2_decap_8 FILLER_60_1213 ();
 sg13g2_decap_8 FILLER_60_1220 ();
 sg13g2_decap_8 FILLER_60_1227 ();
 sg13g2_decap_8 FILLER_60_1234 ();
 sg13g2_decap_8 FILLER_60_1241 ();
 sg13g2_decap_8 FILLER_60_1248 ();
 sg13g2_decap_8 FILLER_60_1255 ();
 sg13g2_decap_8 FILLER_60_1262 ();
 sg13g2_decap_8 FILLER_60_1269 ();
 sg13g2_decap_4 FILLER_60_1276 ();
 sg13g2_fill_2 FILLER_60_1280 ();
 sg13g2_decap_8 FILLER_60_1383 ();
 sg13g2_decap_4 FILLER_60_1390 ();
 sg13g2_fill_2 FILLER_60_1394 ();
 sg13g2_decap_8 FILLER_60_1454 ();
 sg13g2_decap_8 FILLER_60_1461 ();
 sg13g2_fill_1 FILLER_60_1468 ();
 sg13g2_decap_8 FILLER_60_1501 ();
 sg13g2_decap_8 FILLER_60_1516 ();
 sg13g2_decap_8 FILLER_60_1594 ();
 sg13g2_decap_8 FILLER_60_1601 ();
 sg13g2_decap_8 FILLER_60_1608 ();
 sg13g2_decap_8 FILLER_60_1615 ();
 sg13g2_decap_4 FILLER_60_1622 ();
 sg13g2_fill_1 FILLER_60_1626 ();
 sg13g2_decap_8 FILLER_60_1653 ();
 sg13g2_decap_8 FILLER_60_1660 ();
 sg13g2_decap_4 FILLER_60_1667 ();
 sg13g2_fill_1 FILLER_60_1671 ();
 sg13g2_fill_2 FILLER_60_1698 ();
 sg13g2_fill_1 FILLER_60_1700 ();
 sg13g2_decap_4 FILLER_60_1731 ();
 sg13g2_decap_8 FILLER_60_1749 ();
 sg13g2_decap_8 FILLER_60_1756 ();
 sg13g2_decap_8 FILLER_60_1763 ();
 sg13g2_decap_8 FILLER_60_1770 ();
 sg13g2_fill_2 FILLER_60_1777 ();
 sg13g2_fill_1 FILLER_60_1779 ();
 sg13g2_decap_8 FILLER_60_1819 ();
 sg13g2_fill_1 FILLER_60_1826 ();
 sg13g2_decap_4 FILLER_60_1853 ();
 sg13g2_fill_1 FILLER_60_1857 ();
 sg13g2_decap_4 FILLER_60_1902 ();
 sg13g2_fill_1 FILLER_60_1932 ();
 sg13g2_fill_2 FILLER_60_1941 ();
 sg13g2_fill_1 FILLER_60_1966 ();
 sg13g2_decap_8 FILLER_60_1972 ();
 sg13g2_decap_8 FILLER_60_1979 ();
 sg13g2_decap_8 FILLER_60_1986 ();
 sg13g2_decap_8 FILLER_60_1993 ();
 sg13g2_decap_8 FILLER_60_2000 ();
 sg13g2_decap_4 FILLER_60_2007 ();
 sg13g2_decap_8 FILLER_60_2053 ();
 sg13g2_decap_8 FILLER_60_2060 ();
 sg13g2_decap_4 FILLER_60_2067 ();
 sg13g2_fill_2 FILLER_60_2118 ();
 sg13g2_fill_1 FILLER_60_2176 ();
 sg13g2_decap_8 FILLER_60_2255 ();
 sg13g2_decap_8 FILLER_60_2262 ();
 sg13g2_decap_8 FILLER_60_2269 ();
 sg13g2_decap_8 FILLER_60_2276 ();
 sg13g2_decap_8 FILLER_60_2283 ();
 sg13g2_decap_8 FILLER_60_2290 ();
 sg13g2_decap_8 FILLER_60_2297 ();
 sg13g2_decap_8 FILLER_60_2304 ();
 sg13g2_decap_8 FILLER_60_2311 ();
 sg13g2_decap_8 FILLER_60_2318 ();
 sg13g2_decap_8 FILLER_60_2325 ();
 sg13g2_decap_8 FILLER_60_2332 ();
 sg13g2_decap_8 FILLER_60_2339 ();
 sg13g2_decap_8 FILLER_60_2346 ();
 sg13g2_decap_8 FILLER_60_2353 ();
 sg13g2_decap_8 FILLER_60_2360 ();
 sg13g2_decap_8 FILLER_60_2367 ();
 sg13g2_decap_8 FILLER_60_2374 ();
 sg13g2_decap_8 FILLER_60_2381 ();
 sg13g2_decap_8 FILLER_60_2388 ();
 sg13g2_decap_8 FILLER_60_2395 ();
 sg13g2_decap_8 FILLER_60_2402 ();
 sg13g2_decap_8 FILLER_60_2409 ();
 sg13g2_decap_8 FILLER_60_2416 ();
 sg13g2_decap_8 FILLER_60_2423 ();
 sg13g2_decap_8 FILLER_60_2430 ();
 sg13g2_decap_8 FILLER_60_2437 ();
 sg13g2_decap_8 FILLER_60_2444 ();
 sg13g2_decap_8 FILLER_60_2451 ();
 sg13g2_decap_8 FILLER_60_2458 ();
 sg13g2_decap_8 FILLER_60_2465 ();
 sg13g2_decap_8 FILLER_60_2472 ();
 sg13g2_decap_8 FILLER_60_2479 ();
 sg13g2_decap_8 FILLER_60_2486 ();
 sg13g2_decap_8 FILLER_60_2493 ();
 sg13g2_decap_8 FILLER_60_2500 ();
 sg13g2_decap_8 FILLER_60_2507 ();
 sg13g2_decap_8 FILLER_60_2514 ();
 sg13g2_decap_8 FILLER_60_2521 ();
 sg13g2_decap_8 FILLER_60_2528 ();
 sg13g2_decap_8 FILLER_60_2535 ();
 sg13g2_decap_8 FILLER_60_2542 ();
 sg13g2_fill_2 FILLER_60_2549 ();
 sg13g2_decap_4 FILLER_60_2555 ();
 sg13g2_decap_8 FILLER_60_2563 ();
 sg13g2_decap_8 FILLER_60_2570 ();
 sg13g2_decap_4 FILLER_60_2577 ();
 sg13g2_fill_1 FILLER_60_2581 ();
 sg13g2_fill_1 FILLER_60_2613 ();
 sg13g2_fill_2 FILLER_60_2640 ();
 sg13g2_decap_8 FILLER_60_2668 ();
 sg13g2_decap_8 FILLER_60_2675 ();
 sg13g2_decap_4 FILLER_60_2682 ();
 sg13g2_decap_4 FILLER_60_2712 ();
 sg13g2_decap_4 FILLER_60_2742 ();
 sg13g2_fill_2 FILLER_60_2746 ();
 sg13g2_fill_2 FILLER_60_2774 ();
 sg13g2_fill_2 FILLER_60_2781 ();
 sg13g2_fill_2 FILLER_60_2791 ();
 sg13g2_decap_8 FILLER_60_2828 ();
 sg13g2_fill_1 FILLER_60_2843 ();
 sg13g2_decap_8 FILLER_60_2870 ();
 sg13g2_decap_4 FILLER_60_2877 ();
 sg13g2_fill_1 FILLER_60_2881 ();
 sg13g2_decap_8 FILLER_60_2947 ();
 sg13g2_decap_8 FILLER_60_2954 ();
 sg13g2_decap_8 FILLER_60_2961 ();
 sg13g2_decap_8 FILLER_60_2973 ();
 sg13g2_decap_8 FILLER_60_2980 ();
 sg13g2_decap_8 FILLER_60_2987 ();
 sg13g2_decap_8 FILLER_60_2994 ();
 sg13g2_decap_8 FILLER_60_3001 ();
 sg13g2_decap_8 FILLER_60_3034 ();
 sg13g2_decap_8 FILLER_60_3041 ();
 sg13g2_decap_8 FILLER_60_3048 ();
 sg13g2_decap_8 FILLER_60_3055 ();
 sg13g2_decap_8 FILLER_60_3062 ();
 sg13g2_decap_8 FILLER_60_3069 ();
 sg13g2_decap_8 FILLER_60_3076 ();
 sg13g2_decap_8 FILLER_60_3083 ();
 sg13g2_decap_8 FILLER_60_3090 ();
 sg13g2_decap_8 FILLER_60_3097 ();
 sg13g2_decap_8 FILLER_60_3104 ();
 sg13g2_decap_8 FILLER_60_3111 ();
 sg13g2_decap_8 FILLER_60_3118 ();
 sg13g2_decap_8 FILLER_60_3125 ();
 sg13g2_decap_8 FILLER_60_3132 ();
 sg13g2_decap_8 FILLER_60_3139 ();
 sg13g2_decap_8 FILLER_60_3146 ();
 sg13g2_decap_8 FILLER_60_3153 ();
 sg13g2_decap_8 FILLER_60_3160 ();
 sg13g2_decap_8 FILLER_60_3167 ();
 sg13g2_decap_8 FILLER_60_3174 ();
 sg13g2_decap_8 FILLER_60_3181 ();
 sg13g2_decap_8 FILLER_60_3188 ();
 sg13g2_decap_8 FILLER_60_3195 ();
 sg13g2_decap_8 FILLER_60_3202 ();
 sg13g2_decap_8 FILLER_60_3209 ();
 sg13g2_decap_8 FILLER_60_3216 ();
 sg13g2_decap_8 FILLER_60_3223 ();
 sg13g2_decap_8 FILLER_60_3230 ();
 sg13g2_decap_8 FILLER_60_3237 ();
 sg13g2_decap_8 FILLER_60_3244 ();
 sg13g2_decap_8 FILLER_60_3251 ();
 sg13g2_decap_8 FILLER_60_3258 ();
 sg13g2_decap_8 FILLER_60_3265 ();
 sg13g2_decap_8 FILLER_60_3272 ();
 sg13g2_decap_8 FILLER_60_3279 ();
 sg13g2_decap_8 FILLER_60_3286 ();
 sg13g2_decap_8 FILLER_60_3293 ();
 sg13g2_decap_8 FILLER_60_3300 ();
 sg13g2_decap_8 FILLER_60_3307 ();
 sg13g2_decap_8 FILLER_60_3314 ();
 sg13g2_decap_8 FILLER_60_3321 ();
 sg13g2_decap_8 FILLER_60_3328 ();
 sg13g2_decap_8 FILLER_60_3335 ();
 sg13g2_decap_8 FILLER_60_3342 ();
 sg13g2_decap_8 FILLER_60_3349 ();
 sg13g2_decap_8 FILLER_60_3356 ();
 sg13g2_decap_8 FILLER_60_3363 ();
 sg13g2_decap_8 FILLER_60_3370 ();
 sg13g2_decap_8 FILLER_60_3377 ();
 sg13g2_decap_8 FILLER_60_3384 ();
 sg13g2_decap_8 FILLER_60_3391 ();
 sg13g2_decap_8 FILLER_60_3398 ();
 sg13g2_decap_8 FILLER_60_3405 ();
 sg13g2_decap_8 FILLER_60_3412 ();
 sg13g2_decap_8 FILLER_60_3419 ();
 sg13g2_decap_8 FILLER_60_3426 ();
 sg13g2_decap_8 FILLER_60_3433 ();
 sg13g2_decap_8 FILLER_60_3440 ();
 sg13g2_decap_8 FILLER_60_3447 ();
 sg13g2_decap_8 FILLER_60_3454 ();
 sg13g2_decap_8 FILLER_60_3461 ();
 sg13g2_decap_8 FILLER_60_3468 ();
 sg13g2_decap_8 FILLER_60_3475 ();
 sg13g2_decap_8 FILLER_60_3482 ();
 sg13g2_decap_8 FILLER_60_3489 ();
 sg13g2_decap_8 FILLER_60_3496 ();
 sg13g2_decap_8 FILLER_60_3503 ();
 sg13g2_decap_8 FILLER_60_3510 ();
 sg13g2_decap_8 FILLER_60_3517 ();
 sg13g2_decap_8 FILLER_60_3524 ();
 sg13g2_decap_8 FILLER_60_3531 ();
 sg13g2_decap_8 FILLER_60_3538 ();
 sg13g2_decap_8 FILLER_60_3545 ();
 sg13g2_decap_8 FILLER_60_3552 ();
 sg13g2_decap_8 FILLER_60_3559 ();
 sg13g2_decap_8 FILLER_60_3566 ();
 sg13g2_decap_8 FILLER_60_3573 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_decap_8 FILLER_61_189 ();
 sg13g2_decap_8 FILLER_61_196 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_217 ();
 sg13g2_decap_8 FILLER_61_224 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_decap_8 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_decap_8 FILLER_61_252 ();
 sg13g2_decap_8 FILLER_61_259 ();
 sg13g2_decap_8 FILLER_61_266 ();
 sg13g2_decap_8 FILLER_61_273 ();
 sg13g2_decap_8 FILLER_61_280 ();
 sg13g2_decap_8 FILLER_61_287 ();
 sg13g2_decap_8 FILLER_61_294 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_decap_8 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_322 ();
 sg13g2_decap_8 FILLER_61_329 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_61_357 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_441 ();
 sg13g2_decap_8 FILLER_61_468 ();
 sg13g2_fill_1 FILLER_61_475 ();
 sg13g2_decap_8 FILLER_61_517 ();
 sg13g2_decap_8 FILLER_61_524 ();
 sg13g2_decap_4 FILLER_61_531 ();
 sg13g2_fill_1 FILLER_61_535 ();
 sg13g2_decap_8 FILLER_61_543 ();
 sg13g2_decap_8 FILLER_61_550 ();
 sg13g2_fill_2 FILLER_61_557 ();
 sg13g2_decap_8 FILLER_61_566 ();
 sg13g2_decap_8 FILLER_61_573 ();
 sg13g2_decap_8 FILLER_61_580 ();
 sg13g2_decap_8 FILLER_61_608 ();
 sg13g2_decap_4 FILLER_61_615 ();
 sg13g2_fill_2 FILLER_61_619 ();
 sg13g2_decap_8 FILLER_61_625 ();
 sg13g2_fill_2 FILLER_61_632 ();
 sg13g2_fill_1 FILLER_61_634 ();
 sg13g2_fill_2 FILLER_61_661 ();
 sg13g2_fill_2 FILLER_61_715 ();
 sg13g2_fill_2 FILLER_61_746 ();
 sg13g2_fill_1 FILLER_61_764 ();
 sg13g2_fill_1 FILLER_61_843 ();
 sg13g2_fill_1 FILLER_61_875 ();
 sg13g2_fill_1 FILLER_61_905 ();
 sg13g2_decap_8 FILLER_61_919 ();
 sg13g2_decap_8 FILLER_61_926 ();
 sg13g2_decap_4 FILLER_61_933 ();
 sg13g2_fill_2 FILLER_61_937 ();
 sg13g2_decap_8 FILLER_61_973 ();
 sg13g2_decap_8 FILLER_61_980 ();
 sg13g2_fill_1 FILLER_61_987 ();
 sg13g2_decap_8 FILLER_61_1071 ();
 sg13g2_decap_8 FILLER_61_1078 ();
 sg13g2_decap_8 FILLER_61_1093 ();
 sg13g2_decap_8 FILLER_61_1100 ();
 sg13g2_decap_8 FILLER_61_1107 ();
 sg13g2_decap_4 FILLER_61_1114 ();
 sg13g2_fill_2 FILLER_61_1118 ();
 sg13g2_decap_8 FILLER_61_1151 ();
 sg13g2_decap_4 FILLER_61_1158 ();
 sg13g2_fill_1 FILLER_61_1162 ();
 sg13g2_decap_8 FILLER_61_1201 ();
 sg13g2_decap_4 FILLER_61_1208 ();
 sg13g2_fill_1 FILLER_61_1212 ();
 sg13g2_decap_4 FILLER_61_1218 ();
 sg13g2_decap_8 FILLER_61_1260 ();
 sg13g2_decap_8 FILLER_61_1267 ();
 sg13g2_decap_8 FILLER_61_1274 ();
 sg13g2_fill_2 FILLER_61_1281 ();
 sg13g2_fill_1 FILLER_61_1283 ();
 sg13g2_decap_8 FILLER_61_1316 ();
 sg13g2_fill_2 FILLER_61_1323 ();
 sg13g2_decap_4 FILLER_61_1357 ();
 sg13g2_decap_8 FILLER_61_1369 ();
 sg13g2_decap_8 FILLER_61_1376 ();
 sg13g2_decap_8 FILLER_61_1383 ();
 sg13g2_decap_8 FILLER_61_1390 ();
 sg13g2_fill_2 FILLER_61_1397 ();
 sg13g2_fill_1 FILLER_61_1399 ();
 sg13g2_decap_8 FILLER_61_1406 ();
 sg13g2_fill_2 FILLER_61_1413 ();
 sg13g2_decap_8 FILLER_61_1447 ();
 sg13g2_decap_8 FILLER_61_1454 ();
 sg13g2_fill_2 FILLER_61_1461 ();
 sg13g2_fill_2 FILLER_61_1471 ();
 sg13g2_fill_1 FILLER_61_1473 ();
 sg13g2_decap_4 FILLER_61_1513 ();
 sg13g2_decap_4 FILLER_61_1523 ();
 sg13g2_fill_2 FILLER_61_1549 ();
 sg13g2_decap_8 FILLER_61_1556 ();
 sg13g2_decap_8 FILLER_61_1563 ();
 sg13g2_fill_1 FILLER_61_1570 ();
 sg13g2_decap_8 FILLER_61_1597 ();
 sg13g2_decap_8 FILLER_61_1604 ();
 sg13g2_decap_8 FILLER_61_1611 ();
 sg13g2_fill_2 FILLER_61_1618 ();
 sg13g2_fill_1 FILLER_61_1620 ();
 sg13g2_decap_8 FILLER_61_1736 ();
 sg13g2_fill_2 FILLER_61_1743 ();
 sg13g2_decap_8 FILLER_61_1829 ();
 sg13g2_decap_8 FILLER_61_1836 ();
 sg13g2_fill_2 FILLER_61_1843 ();
 sg13g2_fill_1 FILLER_61_1845 ();
 sg13g2_fill_2 FILLER_61_1872 ();
 sg13g2_fill_1 FILLER_61_1874 ();
 sg13g2_fill_2 FILLER_61_1883 ();
 sg13g2_fill_1 FILLER_61_1885 ();
 sg13g2_decap_4 FILLER_61_1899 ();
 sg13g2_fill_2 FILLER_61_1903 ();
 sg13g2_decap_8 FILLER_61_1924 ();
 sg13g2_fill_2 FILLER_61_1931 ();
 sg13g2_fill_1 FILLER_61_1936 ();
 sg13g2_fill_2 FILLER_61_1953 ();
 sg13g2_decap_8 FILLER_61_1959 ();
 sg13g2_decap_8 FILLER_61_1966 ();
 sg13g2_decap_8 FILLER_61_1973 ();
 sg13g2_decap_8 FILLER_61_1980 ();
 sg13g2_decap_4 FILLER_61_1987 ();
 sg13g2_fill_1 FILLER_61_1991 ();
 sg13g2_decap_8 FILLER_61_1997 ();
 sg13g2_fill_1 FILLER_61_2004 ();
 sg13g2_decap_8 FILLER_61_2057 ();
 sg13g2_decap_8 FILLER_61_2064 ();
 sg13g2_decap_4 FILLER_61_2071 ();
 sg13g2_fill_1 FILLER_61_2075 ();
 sg13g2_decap_4 FILLER_61_2121 ();
 sg13g2_fill_2 FILLER_61_2125 ();
 sg13g2_fill_2 FILLER_61_2179 ();
 sg13g2_fill_1 FILLER_61_2181 ();
 sg13g2_fill_2 FILLER_61_2213 ();
 sg13g2_decap_8 FILLER_61_2241 ();
 sg13g2_decap_8 FILLER_61_2248 ();
 sg13g2_decap_8 FILLER_61_2255 ();
 sg13g2_decap_8 FILLER_61_2262 ();
 sg13g2_decap_8 FILLER_61_2269 ();
 sg13g2_decap_8 FILLER_61_2276 ();
 sg13g2_decap_8 FILLER_61_2283 ();
 sg13g2_decap_8 FILLER_61_2290 ();
 sg13g2_decap_8 FILLER_61_2297 ();
 sg13g2_decap_8 FILLER_61_2304 ();
 sg13g2_decap_8 FILLER_61_2311 ();
 sg13g2_decap_8 FILLER_61_2318 ();
 sg13g2_decap_8 FILLER_61_2325 ();
 sg13g2_decap_8 FILLER_61_2332 ();
 sg13g2_decap_8 FILLER_61_2339 ();
 sg13g2_decap_8 FILLER_61_2346 ();
 sg13g2_decap_8 FILLER_61_2353 ();
 sg13g2_decap_8 FILLER_61_2360 ();
 sg13g2_decap_8 FILLER_61_2367 ();
 sg13g2_decap_8 FILLER_61_2374 ();
 sg13g2_decap_8 FILLER_61_2381 ();
 sg13g2_decap_8 FILLER_61_2388 ();
 sg13g2_decap_8 FILLER_61_2395 ();
 sg13g2_decap_8 FILLER_61_2402 ();
 sg13g2_decap_8 FILLER_61_2409 ();
 sg13g2_decap_8 FILLER_61_2416 ();
 sg13g2_decap_8 FILLER_61_2423 ();
 sg13g2_decap_8 FILLER_61_2430 ();
 sg13g2_decap_8 FILLER_61_2437 ();
 sg13g2_decap_8 FILLER_61_2444 ();
 sg13g2_decap_8 FILLER_61_2451 ();
 sg13g2_decap_8 FILLER_61_2458 ();
 sg13g2_decap_8 FILLER_61_2465 ();
 sg13g2_decap_8 FILLER_61_2472 ();
 sg13g2_decap_8 FILLER_61_2479 ();
 sg13g2_decap_8 FILLER_61_2486 ();
 sg13g2_decap_8 FILLER_61_2493 ();
 sg13g2_decap_8 FILLER_61_2500 ();
 sg13g2_decap_8 FILLER_61_2507 ();
 sg13g2_decap_8 FILLER_61_2514 ();
 sg13g2_decap_8 FILLER_61_2521 ();
 sg13g2_decap_8 FILLER_61_2528 ();
 sg13g2_decap_8 FILLER_61_2535 ();
 sg13g2_decap_8 FILLER_61_2542 ();
 sg13g2_decap_8 FILLER_61_2549 ();
 sg13g2_decap_8 FILLER_61_2556 ();
 sg13g2_decap_8 FILLER_61_2563 ();
 sg13g2_decap_8 FILLER_61_2570 ();
 sg13g2_decap_8 FILLER_61_2577 ();
 sg13g2_decap_8 FILLER_61_2584 ();
 sg13g2_decap_8 FILLER_61_2591 ();
 sg13g2_decap_8 FILLER_61_2598 ();
 sg13g2_decap_8 FILLER_61_2665 ();
 sg13g2_decap_8 FILLER_61_2672 ();
 sg13g2_decap_8 FILLER_61_2679 ();
 sg13g2_decap_4 FILLER_61_2686 ();
 sg13g2_fill_2 FILLER_61_2742 ();
 sg13g2_fill_1 FILLER_61_2744 ();
 sg13g2_decap_8 FILLER_61_2823 ();
 sg13g2_fill_2 FILLER_61_2830 ();
 sg13g2_fill_1 FILLER_61_2832 ();
 sg13g2_decap_8 FILLER_61_2859 ();
 sg13g2_decap_8 FILLER_61_2866 ();
 sg13g2_decap_8 FILLER_61_2873 ();
 sg13g2_decap_8 FILLER_61_2880 ();
 sg13g2_decap_4 FILLER_61_2887 ();
 sg13g2_fill_1 FILLER_61_2891 ();
 sg13g2_decap_8 FILLER_61_2944 ();
 sg13g2_decap_8 FILLER_61_2951 ();
 sg13g2_decap_8 FILLER_61_2958 ();
 sg13g2_decap_8 FILLER_61_2965 ();
 sg13g2_decap_8 FILLER_61_2972 ();
 sg13g2_decap_8 FILLER_61_2979 ();
 sg13g2_decap_8 FILLER_61_2986 ();
 sg13g2_decap_8 FILLER_61_2993 ();
 sg13g2_decap_8 FILLER_61_3000 ();
 sg13g2_decap_8 FILLER_61_3007 ();
 sg13g2_decap_8 FILLER_61_3014 ();
 sg13g2_decap_8 FILLER_61_3021 ();
 sg13g2_decap_8 FILLER_61_3028 ();
 sg13g2_decap_8 FILLER_61_3035 ();
 sg13g2_decap_8 FILLER_61_3042 ();
 sg13g2_decap_8 FILLER_61_3049 ();
 sg13g2_decap_8 FILLER_61_3056 ();
 sg13g2_decap_8 FILLER_61_3063 ();
 sg13g2_decap_8 FILLER_61_3070 ();
 sg13g2_decap_8 FILLER_61_3077 ();
 sg13g2_decap_8 FILLER_61_3084 ();
 sg13g2_decap_8 FILLER_61_3091 ();
 sg13g2_decap_8 FILLER_61_3098 ();
 sg13g2_decap_8 FILLER_61_3105 ();
 sg13g2_decap_8 FILLER_61_3112 ();
 sg13g2_decap_8 FILLER_61_3119 ();
 sg13g2_decap_8 FILLER_61_3126 ();
 sg13g2_decap_8 FILLER_61_3133 ();
 sg13g2_decap_8 FILLER_61_3140 ();
 sg13g2_decap_8 FILLER_61_3147 ();
 sg13g2_decap_8 FILLER_61_3154 ();
 sg13g2_decap_8 FILLER_61_3161 ();
 sg13g2_decap_8 FILLER_61_3168 ();
 sg13g2_decap_8 FILLER_61_3175 ();
 sg13g2_decap_8 FILLER_61_3182 ();
 sg13g2_decap_8 FILLER_61_3189 ();
 sg13g2_decap_8 FILLER_61_3196 ();
 sg13g2_decap_8 FILLER_61_3203 ();
 sg13g2_decap_8 FILLER_61_3210 ();
 sg13g2_decap_8 FILLER_61_3217 ();
 sg13g2_decap_8 FILLER_61_3224 ();
 sg13g2_decap_8 FILLER_61_3231 ();
 sg13g2_decap_8 FILLER_61_3238 ();
 sg13g2_decap_8 FILLER_61_3245 ();
 sg13g2_decap_8 FILLER_61_3252 ();
 sg13g2_decap_8 FILLER_61_3259 ();
 sg13g2_decap_8 FILLER_61_3266 ();
 sg13g2_decap_8 FILLER_61_3273 ();
 sg13g2_decap_8 FILLER_61_3280 ();
 sg13g2_decap_8 FILLER_61_3287 ();
 sg13g2_decap_8 FILLER_61_3294 ();
 sg13g2_decap_8 FILLER_61_3301 ();
 sg13g2_decap_8 FILLER_61_3308 ();
 sg13g2_decap_8 FILLER_61_3315 ();
 sg13g2_decap_8 FILLER_61_3322 ();
 sg13g2_decap_8 FILLER_61_3329 ();
 sg13g2_decap_8 FILLER_61_3336 ();
 sg13g2_decap_8 FILLER_61_3343 ();
 sg13g2_decap_8 FILLER_61_3350 ();
 sg13g2_decap_8 FILLER_61_3357 ();
 sg13g2_decap_8 FILLER_61_3364 ();
 sg13g2_decap_8 FILLER_61_3371 ();
 sg13g2_decap_8 FILLER_61_3378 ();
 sg13g2_decap_8 FILLER_61_3385 ();
 sg13g2_decap_8 FILLER_61_3392 ();
 sg13g2_decap_8 FILLER_61_3399 ();
 sg13g2_decap_8 FILLER_61_3406 ();
 sg13g2_decap_8 FILLER_61_3413 ();
 sg13g2_decap_8 FILLER_61_3420 ();
 sg13g2_decap_8 FILLER_61_3427 ();
 sg13g2_decap_8 FILLER_61_3434 ();
 sg13g2_decap_8 FILLER_61_3441 ();
 sg13g2_decap_8 FILLER_61_3448 ();
 sg13g2_decap_8 FILLER_61_3455 ();
 sg13g2_decap_8 FILLER_61_3462 ();
 sg13g2_decap_8 FILLER_61_3469 ();
 sg13g2_decap_8 FILLER_61_3476 ();
 sg13g2_decap_8 FILLER_61_3483 ();
 sg13g2_decap_8 FILLER_61_3490 ();
 sg13g2_decap_8 FILLER_61_3497 ();
 sg13g2_decap_8 FILLER_61_3504 ();
 sg13g2_decap_8 FILLER_61_3511 ();
 sg13g2_decap_8 FILLER_61_3518 ();
 sg13g2_decap_8 FILLER_61_3525 ();
 sg13g2_decap_8 FILLER_61_3532 ();
 sg13g2_decap_8 FILLER_61_3539 ();
 sg13g2_decap_8 FILLER_61_3546 ();
 sg13g2_decap_8 FILLER_61_3553 ();
 sg13g2_decap_8 FILLER_61_3560 ();
 sg13g2_decap_8 FILLER_61_3567 ();
 sg13g2_decap_4 FILLER_61_3574 ();
 sg13g2_fill_2 FILLER_61_3578 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_decap_8 FILLER_62_245 ();
 sg13g2_decap_8 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_decap_8 FILLER_62_273 ();
 sg13g2_decap_8 FILLER_62_280 ();
 sg13g2_decap_8 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_294 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_decap_4 FILLER_62_406 ();
 sg13g2_decap_8 FILLER_62_467 ();
 sg13g2_decap_4 FILLER_62_474 ();
 sg13g2_decap_8 FILLER_62_524 ();
 sg13g2_decap_8 FILLER_62_531 ();
 sg13g2_fill_1 FILLER_62_538 ();
 sg13g2_decap_8 FILLER_62_577 ();
 sg13g2_decap_4 FILLER_62_584 ();
 sg13g2_fill_2 FILLER_62_588 ();
 sg13g2_fill_2 FILLER_62_605 ();
 sg13g2_decap_4 FILLER_62_659 ();
 sg13g2_fill_1 FILLER_62_663 ();
 sg13g2_decap_8 FILLER_62_755 ();
 sg13g2_fill_2 FILLER_62_762 ();
 sg13g2_fill_1 FILLER_62_764 ();
 sg13g2_decap_8 FILLER_62_800 ();
 sg13g2_fill_2 FILLER_62_807 ();
 sg13g2_fill_2 FILLER_62_813 ();
 sg13g2_decap_8 FILLER_62_845 ();
 sg13g2_fill_1 FILLER_62_852 ();
 sg13g2_fill_2 FILLER_62_857 ();
 sg13g2_fill_1 FILLER_62_859 ();
 sg13g2_decap_8 FILLER_62_864 ();
 sg13g2_fill_1 FILLER_62_871 ();
 sg13g2_decap_8 FILLER_62_877 ();
 sg13g2_fill_1 FILLER_62_888 ();
 sg13g2_fill_2 FILLER_62_902 ();
 sg13g2_decap_8 FILLER_62_908 ();
 sg13g2_decap_8 FILLER_62_915 ();
 sg13g2_decap_8 FILLER_62_922 ();
 sg13g2_decap_4 FILLER_62_929 ();
 sg13g2_decap_8 FILLER_62_968 ();
 sg13g2_decap_4 FILLER_62_975 ();
 sg13g2_fill_2 FILLER_62_979 ();
 sg13g2_decap_8 FILLER_62_1015 ();
 sg13g2_decap_8 FILLER_62_1022 ();
 sg13g2_fill_2 FILLER_62_1029 ();
 sg13g2_fill_1 FILLER_62_1044 ();
 sg13g2_decap_8 FILLER_62_1074 ();
 sg13g2_decap_8 FILLER_62_1081 ();
 sg13g2_decap_8 FILLER_62_1088 ();
 sg13g2_decap_8 FILLER_62_1095 ();
 sg13g2_decap_8 FILLER_62_1102 ();
 sg13g2_decap_8 FILLER_62_1109 ();
 sg13g2_decap_8 FILLER_62_1116 ();
 sg13g2_decap_8 FILLER_62_1123 ();
 sg13g2_decap_8 FILLER_62_1130 ();
 sg13g2_decap_8 FILLER_62_1137 ();
 sg13g2_decap_8 FILLER_62_1144 ();
 sg13g2_decap_8 FILLER_62_1151 ();
 sg13g2_decap_8 FILLER_62_1158 ();
 sg13g2_decap_4 FILLER_62_1165 ();
 sg13g2_fill_2 FILLER_62_1169 ();
 sg13g2_fill_2 FILLER_62_1211 ();
 sg13g2_decap_8 FILLER_62_1265 ();
 sg13g2_decap_8 FILLER_62_1272 ();
 sg13g2_decap_8 FILLER_62_1279 ();
 sg13g2_decap_8 FILLER_62_1317 ();
 sg13g2_decap_4 FILLER_62_1324 ();
 sg13g2_fill_1 FILLER_62_1328 ();
 sg13g2_decap_8 FILLER_62_1360 ();
 sg13g2_fill_2 FILLER_62_1367 ();
 sg13g2_decap_8 FILLER_62_1440 ();
 sg13g2_decap_8 FILLER_62_1447 ();
 sg13g2_decap_8 FILLER_62_1454 ();
 sg13g2_fill_2 FILLER_62_1461 ();
 sg13g2_fill_1 FILLER_62_1463 ();
 sg13g2_decap_8 FILLER_62_1532 ();
 sg13g2_decap_8 FILLER_62_1539 ();
 sg13g2_decap_4 FILLER_62_1546 ();
 sg13g2_fill_2 FILLER_62_1576 ();
 sg13g2_decap_8 FILLER_62_1604 ();
 sg13g2_decap_8 FILLER_62_1611 ();
 sg13g2_fill_1 FILLER_62_1618 ();
 sg13g2_decap_4 FILLER_62_1676 ();
 sg13g2_decap_4 FILLER_62_1734 ();
 sg13g2_fill_1 FILLER_62_1738 ();
 sg13g2_fill_2 FILLER_62_1791 ();
 sg13g2_fill_1 FILLER_62_1793 ();
 sg13g2_decap_4 FILLER_62_1828 ();
 sg13g2_fill_2 FILLER_62_1832 ();
 sg13g2_fill_1 FILLER_62_1838 ();
 sg13g2_decap_8 FILLER_62_1870 ();
 sg13g2_fill_2 FILLER_62_1877 ();
 sg13g2_fill_1 FILLER_62_1879 ();
 sg13g2_decap_8 FILLER_62_1888 ();
 sg13g2_decap_8 FILLER_62_1895 ();
 sg13g2_decap_8 FILLER_62_1902 ();
 sg13g2_fill_1 FILLER_62_1909 ();
 sg13g2_decap_4 FILLER_62_1918 ();
 sg13g2_fill_2 FILLER_62_1922 ();
 sg13g2_fill_1 FILLER_62_1930 ();
 sg13g2_fill_1 FILLER_62_1940 ();
 sg13g2_decap_8 FILLER_62_1954 ();
 sg13g2_fill_2 FILLER_62_1971 ();
 sg13g2_decap_8 FILLER_62_2064 ();
 sg13g2_decap_8 FILLER_62_2071 ();
 sg13g2_fill_1 FILLER_62_2078 ();
 sg13g2_decap_8 FILLER_62_2119 ();
 sg13g2_decap_8 FILLER_62_2126 ();
 sg13g2_fill_2 FILLER_62_2133 ();
 sg13g2_decap_8 FILLER_62_2185 ();
 sg13g2_decap_8 FILLER_62_2192 ();
 sg13g2_decap_8 FILLER_62_2199 ();
 sg13g2_decap_8 FILLER_62_2206 ();
 sg13g2_fill_2 FILLER_62_2213 ();
 sg13g2_fill_1 FILLER_62_2215 ();
 sg13g2_decap_8 FILLER_62_2242 ();
 sg13g2_decap_8 FILLER_62_2249 ();
 sg13g2_decap_8 FILLER_62_2256 ();
 sg13g2_decap_8 FILLER_62_2263 ();
 sg13g2_decap_8 FILLER_62_2270 ();
 sg13g2_decap_8 FILLER_62_2277 ();
 sg13g2_decap_8 FILLER_62_2284 ();
 sg13g2_decap_8 FILLER_62_2291 ();
 sg13g2_decap_8 FILLER_62_2298 ();
 sg13g2_decap_8 FILLER_62_2305 ();
 sg13g2_decap_8 FILLER_62_2312 ();
 sg13g2_decap_8 FILLER_62_2319 ();
 sg13g2_decap_8 FILLER_62_2326 ();
 sg13g2_decap_8 FILLER_62_2333 ();
 sg13g2_decap_8 FILLER_62_2340 ();
 sg13g2_decap_8 FILLER_62_2347 ();
 sg13g2_decap_8 FILLER_62_2354 ();
 sg13g2_decap_8 FILLER_62_2361 ();
 sg13g2_decap_8 FILLER_62_2368 ();
 sg13g2_decap_8 FILLER_62_2375 ();
 sg13g2_decap_8 FILLER_62_2382 ();
 sg13g2_decap_8 FILLER_62_2389 ();
 sg13g2_decap_8 FILLER_62_2396 ();
 sg13g2_decap_8 FILLER_62_2403 ();
 sg13g2_decap_8 FILLER_62_2410 ();
 sg13g2_decap_8 FILLER_62_2417 ();
 sg13g2_decap_8 FILLER_62_2424 ();
 sg13g2_decap_8 FILLER_62_2431 ();
 sg13g2_decap_8 FILLER_62_2438 ();
 sg13g2_decap_8 FILLER_62_2445 ();
 sg13g2_decap_8 FILLER_62_2452 ();
 sg13g2_decap_8 FILLER_62_2459 ();
 sg13g2_decap_8 FILLER_62_2466 ();
 sg13g2_decap_8 FILLER_62_2473 ();
 sg13g2_decap_8 FILLER_62_2480 ();
 sg13g2_decap_8 FILLER_62_2487 ();
 sg13g2_decap_8 FILLER_62_2494 ();
 sg13g2_decap_8 FILLER_62_2501 ();
 sg13g2_decap_8 FILLER_62_2508 ();
 sg13g2_decap_8 FILLER_62_2515 ();
 sg13g2_decap_8 FILLER_62_2522 ();
 sg13g2_decap_8 FILLER_62_2529 ();
 sg13g2_decap_8 FILLER_62_2536 ();
 sg13g2_decap_8 FILLER_62_2543 ();
 sg13g2_decap_8 FILLER_62_2550 ();
 sg13g2_decap_8 FILLER_62_2557 ();
 sg13g2_decap_8 FILLER_62_2564 ();
 sg13g2_decap_8 FILLER_62_2571 ();
 sg13g2_decap_8 FILLER_62_2578 ();
 sg13g2_decap_8 FILLER_62_2585 ();
 sg13g2_decap_8 FILLER_62_2592 ();
 sg13g2_fill_2 FILLER_62_2599 ();
 sg13g2_fill_1 FILLER_62_2601 ();
 sg13g2_decap_4 FILLER_62_2680 ();
 sg13g2_fill_2 FILLER_62_2710 ();
 sg13g2_fill_1 FILLER_62_2738 ();
 sg13g2_decap_4 FILLER_62_2791 ();
 sg13g2_fill_1 FILLER_62_2795 ();
 sg13g2_decap_8 FILLER_62_2874 ();
 sg13g2_decap_8 FILLER_62_2881 ();
 sg13g2_decap_8 FILLER_62_2888 ();
 sg13g2_fill_2 FILLER_62_2895 ();
 sg13g2_decap_8 FILLER_62_2923 ();
 sg13g2_decap_8 FILLER_62_2930 ();
 sg13g2_decap_8 FILLER_62_2937 ();
 sg13g2_decap_8 FILLER_62_2944 ();
 sg13g2_decap_8 FILLER_62_2951 ();
 sg13g2_decap_8 FILLER_62_2958 ();
 sg13g2_decap_8 FILLER_62_2965 ();
 sg13g2_decap_8 FILLER_62_2972 ();
 sg13g2_decap_8 FILLER_62_2979 ();
 sg13g2_decap_8 FILLER_62_2986 ();
 sg13g2_decap_8 FILLER_62_2993 ();
 sg13g2_decap_8 FILLER_62_3000 ();
 sg13g2_decap_8 FILLER_62_3007 ();
 sg13g2_decap_8 FILLER_62_3014 ();
 sg13g2_decap_8 FILLER_62_3021 ();
 sg13g2_decap_8 FILLER_62_3028 ();
 sg13g2_decap_8 FILLER_62_3035 ();
 sg13g2_decap_8 FILLER_62_3042 ();
 sg13g2_decap_8 FILLER_62_3049 ();
 sg13g2_decap_8 FILLER_62_3056 ();
 sg13g2_decap_8 FILLER_62_3063 ();
 sg13g2_decap_8 FILLER_62_3070 ();
 sg13g2_decap_8 FILLER_62_3077 ();
 sg13g2_decap_8 FILLER_62_3084 ();
 sg13g2_decap_8 FILLER_62_3091 ();
 sg13g2_decap_8 FILLER_62_3098 ();
 sg13g2_decap_8 FILLER_62_3105 ();
 sg13g2_decap_8 FILLER_62_3112 ();
 sg13g2_decap_8 FILLER_62_3119 ();
 sg13g2_decap_8 FILLER_62_3126 ();
 sg13g2_decap_8 FILLER_62_3133 ();
 sg13g2_decap_8 FILLER_62_3140 ();
 sg13g2_decap_8 FILLER_62_3147 ();
 sg13g2_decap_8 FILLER_62_3154 ();
 sg13g2_decap_8 FILLER_62_3161 ();
 sg13g2_decap_8 FILLER_62_3168 ();
 sg13g2_decap_8 FILLER_62_3175 ();
 sg13g2_decap_8 FILLER_62_3182 ();
 sg13g2_decap_8 FILLER_62_3189 ();
 sg13g2_decap_8 FILLER_62_3196 ();
 sg13g2_decap_8 FILLER_62_3203 ();
 sg13g2_decap_8 FILLER_62_3210 ();
 sg13g2_decap_8 FILLER_62_3217 ();
 sg13g2_decap_8 FILLER_62_3224 ();
 sg13g2_decap_8 FILLER_62_3231 ();
 sg13g2_decap_8 FILLER_62_3238 ();
 sg13g2_decap_8 FILLER_62_3245 ();
 sg13g2_decap_8 FILLER_62_3252 ();
 sg13g2_decap_8 FILLER_62_3259 ();
 sg13g2_decap_8 FILLER_62_3266 ();
 sg13g2_decap_8 FILLER_62_3273 ();
 sg13g2_decap_8 FILLER_62_3280 ();
 sg13g2_decap_8 FILLER_62_3287 ();
 sg13g2_decap_8 FILLER_62_3294 ();
 sg13g2_decap_8 FILLER_62_3301 ();
 sg13g2_decap_8 FILLER_62_3308 ();
 sg13g2_decap_8 FILLER_62_3315 ();
 sg13g2_decap_8 FILLER_62_3322 ();
 sg13g2_decap_8 FILLER_62_3329 ();
 sg13g2_decap_8 FILLER_62_3336 ();
 sg13g2_decap_8 FILLER_62_3343 ();
 sg13g2_decap_8 FILLER_62_3350 ();
 sg13g2_decap_8 FILLER_62_3357 ();
 sg13g2_decap_8 FILLER_62_3364 ();
 sg13g2_decap_8 FILLER_62_3371 ();
 sg13g2_decap_8 FILLER_62_3378 ();
 sg13g2_decap_8 FILLER_62_3385 ();
 sg13g2_decap_8 FILLER_62_3392 ();
 sg13g2_decap_8 FILLER_62_3399 ();
 sg13g2_decap_8 FILLER_62_3406 ();
 sg13g2_decap_8 FILLER_62_3413 ();
 sg13g2_decap_8 FILLER_62_3420 ();
 sg13g2_decap_8 FILLER_62_3427 ();
 sg13g2_decap_8 FILLER_62_3434 ();
 sg13g2_decap_8 FILLER_62_3441 ();
 sg13g2_decap_8 FILLER_62_3448 ();
 sg13g2_decap_8 FILLER_62_3455 ();
 sg13g2_decap_8 FILLER_62_3462 ();
 sg13g2_decap_8 FILLER_62_3469 ();
 sg13g2_decap_8 FILLER_62_3476 ();
 sg13g2_decap_8 FILLER_62_3483 ();
 sg13g2_decap_8 FILLER_62_3490 ();
 sg13g2_decap_8 FILLER_62_3497 ();
 sg13g2_decap_8 FILLER_62_3504 ();
 sg13g2_decap_8 FILLER_62_3511 ();
 sg13g2_decap_8 FILLER_62_3518 ();
 sg13g2_decap_8 FILLER_62_3525 ();
 sg13g2_decap_8 FILLER_62_3532 ();
 sg13g2_decap_8 FILLER_62_3539 ();
 sg13g2_decap_8 FILLER_62_3546 ();
 sg13g2_decap_8 FILLER_62_3553 ();
 sg13g2_decap_8 FILLER_62_3560 ();
 sg13g2_decap_8 FILLER_62_3567 ();
 sg13g2_decap_4 FILLER_62_3574 ();
 sg13g2_fill_2 FILLER_62_3578 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_217 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_252 ();
 sg13g2_decap_8 FILLER_63_259 ();
 sg13g2_decap_8 FILLER_63_266 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_decap_8 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_301 ();
 sg13g2_decap_8 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_315 ();
 sg13g2_decap_8 FILLER_63_322 ();
 sg13g2_decap_8 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_371 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_decap_4 FILLER_63_413 ();
 sg13g2_fill_2 FILLER_63_417 ();
 sg13g2_decap_8 FILLER_63_473 ();
 sg13g2_decap_4 FILLER_63_480 ();
 sg13g2_fill_1 FILLER_63_484 ();
 sg13g2_decap_4 FILLER_63_518 ();
 sg13g2_fill_2 FILLER_63_522 ();
 sg13g2_fill_2 FILLER_63_553 ();
 sg13g2_decap_4 FILLER_63_581 ();
 sg13g2_fill_2 FILLER_63_630 ();
 sg13g2_decap_8 FILLER_63_663 ();
 sg13g2_decap_4 FILLER_63_670 ();
 sg13g2_decap_4 FILLER_63_678 ();
 sg13g2_fill_2 FILLER_63_716 ();
 sg13g2_decap_4 FILLER_63_738 ();
 sg13g2_decap_8 FILLER_63_747 ();
 sg13g2_decap_4 FILLER_63_754 ();
 sg13g2_fill_1 FILLER_63_758 ();
 sg13g2_decap_4 FILLER_63_762 ();
 sg13g2_decap_8 FILLER_63_792 ();
 sg13g2_decap_8 FILLER_63_799 ();
 sg13g2_decap_8 FILLER_63_806 ();
 sg13g2_fill_2 FILLER_63_821 ();
 sg13g2_decap_8 FILLER_63_832 ();
 sg13g2_decap_8 FILLER_63_839 ();
 sg13g2_fill_2 FILLER_63_846 ();
 sg13g2_fill_1 FILLER_63_848 ();
 sg13g2_decap_8 FILLER_63_857 ();
 sg13g2_fill_2 FILLER_63_864 ();
 sg13g2_decap_8 FILLER_63_916 ();
 sg13g2_decap_4 FILLER_63_923 ();
 sg13g2_fill_1 FILLER_63_927 ();
 sg13g2_fill_2 FILLER_63_939 ();
 sg13g2_fill_1 FILLER_63_941 ();
 sg13g2_fill_2 FILLER_63_952 ();
 sg13g2_fill_1 FILLER_63_954 ();
 sg13g2_fill_2 FILLER_63_963 ();
 sg13g2_decap_4 FILLER_63_973 ();
 sg13g2_decap_8 FILLER_63_982 ();
 sg13g2_fill_1 FILLER_63_989 ();
 sg13g2_decap_8 FILLER_63_1020 ();
 sg13g2_decap_4 FILLER_63_1027 ();
 sg13g2_fill_1 FILLER_63_1031 ();
 sg13g2_fill_1 FILLER_63_1042 ();
 sg13g2_decap_4 FILLER_63_1121 ();
 sg13g2_fill_2 FILLER_63_1125 ();
 sg13g2_decap_8 FILLER_63_1270 ();
 sg13g2_decap_8 FILLER_63_1277 ();
 sg13g2_fill_1 FILLER_63_1288 ();
 sg13g2_decap_4 FILLER_63_1294 ();
 sg13g2_fill_1 FILLER_63_1298 ();
 sg13g2_fill_2 FILLER_63_1304 ();
 sg13g2_fill_1 FILLER_63_1306 ();
 sg13g2_fill_2 FILLER_63_1320 ();
 sg13g2_fill_1 FILLER_63_1322 ();
 sg13g2_fill_2 FILLER_63_1349 ();
 sg13g2_fill_2 FILLER_63_1357 ();
 sg13g2_fill_1 FILLER_63_1364 ();
 sg13g2_decap_8 FILLER_63_1371 ();
 sg13g2_decap_8 FILLER_63_1378 ();
 sg13g2_fill_2 FILLER_63_1385 ();
 sg13g2_fill_1 FILLER_63_1387 ();
 sg13g2_decap_8 FILLER_63_1458 ();
 sg13g2_fill_1 FILLER_63_1465 ();
 sg13g2_fill_2 FILLER_63_1492 ();
 sg13g2_fill_1 FILLER_63_1494 ();
 sg13g2_decap_8 FILLER_63_1521 ();
 sg13g2_decap_8 FILLER_63_1528 ();
 sg13g2_decap_8 FILLER_63_1535 ();
 sg13g2_decap_4 FILLER_63_1542 ();
 sg13g2_fill_1 FILLER_63_1546 ();
 sg13g2_decap_8 FILLER_63_1555 ();
 sg13g2_fill_2 FILLER_63_1562 ();
 sg13g2_decap_8 FILLER_63_1601 ();
 sg13g2_decap_8 FILLER_63_1608 ();
 sg13g2_decap_8 FILLER_63_1615 ();
 sg13g2_decap_8 FILLER_63_1622 ();
 sg13g2_decap_4 FILLER_63_1629 ();
 sg13g2_decap_8 FILLER_63_1667 ();
 sg13g2_decap_8 FILLER_63_1674 ();
 sg13g2_decap_8 FILLER_63_1681 ();
 sg13g2_decap_8 FILLER_63_1688 ();
 sg13g2_fill_2 FILLER_63_1695 ();
 sg13g2_decap_4 FILLER_63_1703 ();
 sg13g2_fill_1 FILLER_63_1707 ();
 sg13g2_decap_8 FILLER_63_1722 ();
 sg13g2_decap_8 FILLER_63_1729 ();
 sg13g2_decap_8 FILLER_63_1736 ();
 sg13g2_decap_8 FILLER_63_1743 ();
 sg13g2_decap_4 FILLER_63_1750 ();
 sg13g2_fill_2 FILLER_63_1754 ();
 sg13g2_decap_4 FILLER_63_1788 ();
 sg13g2_decap_8 FILLER_63_1823 ();
 sg13g2_decap_8 FILLER_63_1830 ();
 sg13g2_decap_8 FILLER_63_1837 ();
 sg13g2_decap_4 FILLER_63_1882 ();
 sg13g2_decap_8 FILLER_63_1894 ();
 sg13g2_decap_4 FILLER_63_1901 ();
 sg13g2_fill_2 FILLER_63_1939 ();
 sg13g2_decap_4 FILLER_63_1967 ();
 sg13g2_fill_2 FILLER_63_1971 ();
 sg13g2_decap_8 FILLER_63_1981 ();
 sg13g2_decap_8 FILLER_63_1988 ();
 sg13g2_decap_8 FILLER_63_1995 ();
 sg13g2_fill_2 FILLER_63_2002 ();
 sg13g2_decap_4 FILLER_63_2062 ();
 sg13g2_fill_1 FILLER_63_2066 ();
 sg13g2_decap_8 FILLER_63_2124 ();
 sg13g2_fill_2 FILLER_63_2131 ();
 sg13g2_fill_1 FILLER_63_2133 ();
 sg13g2_decap_8 FILLER_63_2160 ();
 sg13g2_decap_4 FILLER_63_2167 ();
 sg13g2_fill_2 FILLER_63_2171 ();
 sg13g2_decap_8 FILLER_63_2199 ();
 sg13g2_decap_8 FILLER_63_2206 ();
 sg13g2_decap_8 FILLER_63_2213 ();
 sg13g2_decap_8 FILLER_63_2220 ();
 sg13g2_decap_8 FILLER_63_2227 ();
 sg13g2_decap_8 FILLER_63_2234 ();
 sg13g2_decap_8 FILLER_63_2241 ();
 sg13g2_decap_8 FILLER_63_2248 ();
 sg13g2_decap_8 FILLER_63_2255 ();
 sg13g2_decap_8 FILLER_63_2262 ();
 sg13g2_decap_8 FILLER_63_2269 ();
 sg13g2_decap_8 FILLER_63_2276 ();
 sg13g2_decap_8 FILLER_63_2283 ();
 sg13g2_decap_8 FILLER_63_2290 ();
 sg13g2_decap_8 FILLER_63_2297 ();
 sg13g2_decap_8 FILLER_63_2304 ();
 sg13g2_decap_8 FILLER_63_2311 ();
 sg13g2_decap_8 FILLER_63_2318 ();
 sg13g2_decap_8 FILLER_63_2325 ();
 sg13g2_decap_8 FILLER_63_2332 ();
 sg13g2_decap_8 FILLER_63_2339 ();
 sg13g2_decap_8 FILLER_63_2346 ();
 sg13g2_decap_8 FILLER_63_2353 ();
 sg13g2_decap_8 FILLER_63_2360 ();
 sg13g2_decap_8 FILLER_63_2367 ();
 sg13g2_decap_8 FILLER_63_2374 ();
 sg13g2_decap_8 FILLER_63_2381 ();
 sg13g2_decap_8 FILLER_63_2388 ();
 sg13g2_decap_8 FILLER_63_2395 ();
 sg13g2_decap_8 FILLER_63_2402 ();
 sg13g2_decap_8 FILLER_63_2409 ();
 sg13g2_decap_8 FILLER_63_2416 ();
 sg13g2_decap_8 FILLER_63_2423 ();
 sg13g2_decap_8 FILLER_63_2430 ();
 sg13g2_decap_8 FILLER_63_2437 ();
 sg13g2_decap_8 FILLER_63_2444 ();
 sg13g2_decap_8 FILLER_63_2451 ();
 sg13g2_decap_8 FILLER_63_2458 ();
 sg13g2_decap_8 FILLER_63_2465 ();
 sg13g2_decap_8 FILLER_63_2472 ();
 sg13g2_decap_8 FILLER_63_2479 ();
 sg13g2_decap_8 FILLER_63_2486 ();
 sg13g2_decap_8 FILLER_63_2493 ();
 sg13g2_decap_8 FILLER_63_2500 ();
 sg13g2_decap_8 FILLER_63_2507 ();
 sg13g2_decap_8 FILLER_63_2514 ();
 sg13g2_decap_8 FILLER_63_2521 ();
 sg13g2_decap_8 FILLER_63_2528 ();
 sg13g2_decap_8 FILLER_63_2535 ();
 sg13g2_decap_8 FILLER_63_2542 ();
 sg13g2_decap_8 FILLER_63_2549 ();
 sg13g2_decap_8 FILLER_63_2556 ();
 sg13g2_decap_8 FILLER_63_2563 ();
 sg13g2_decap_8 FILLER_63_2570 ();
 sg13g2_decap_8 FILLER_63_2577 ();
 sg13g2_decap_8 FILLER_63_2584 ();
 sg13g2_decap_8 FILLER_63_2591 ();
 sg13g2_decap_8 FILLER_63_2598 ();
 sg13g2_decap_8 FILLER_63_2605 ();
 sg13g2_decap_8 FILLER_63_2612 ();
 sg13g2_decap_8 FILLER_63_2619 ();
 sg13g2_decap_8 FILLER_63_2652 ();
 sg13g2_decap_8 FILLER_63_2659 ();
 sg13g2_decap_8 FILLER_63_2666 ();
 sg13g2_decap_8 FILLER_63_2673 ();
 sg13g2_decap_8 FILLER_63_2680 ();
 sg13g2_decap_4 FILLER_63_2687 ();
 sg13g2_decap_8 FILLER_63_2725 ();
 sg13g2_decap_8 FILLER_63_2732 ();
 sg13g2_decap_8 FILLER_63_2739 ();
 sg13g2_decap_8 FILLER_63_2746 ();
 sg13g2_decap_8 FILLER_63_2753 ();
 sg13g2_decap_8 FILLER_63_2760 ();
 sg13g2_decap_8 FILLER_63_2767 ();
 sg13g2_decap_8 FILLER_63_2774 ();
 sg13g2_decap_8 FILLER_63_2781 ();
 sg13g2_decap_8 FILLER_63_2788 ();
 sg13g2_decap_4 FILLER_63_2795 ();
 sg13g2_decap_8 FILLER_63_2825 ();
 sg13g2_decap_8 FILLER_63_2832 ();
 sg13g2_decap_4 FILLER_63_2839 ();
 sg13g2_fill_2 FILLER_63_2843 ();
 sg13g2_decap_8 FILLER_63_2871 ();
 sg13g2_decap_8 FILLER_63_2878 ();
 sg13g2_decap_8 FILLER_63_2885 ();
 sg13g2_decap_8 FILLER_63_2892 ();
 sg13g2_decap_8 FILLER_63_2899 ();
 sg13g2_decap_8 FILLER_63_2906 ();
 sg13g2_decap_8 FILLER_63_2913 ();
 sg13g2_decap_8 FILLER_63_2920 ();
 sg13g2_decap_8 FILLER_63_2927 ();
 sg13g2_decap_8 FILLER_63_2934 ();
 sg13g2_decap_8 FILLER_63_2941 ();
 sg13g2_decap_8 FILLER_63_2948 ();
 sg13g2_decap_8 FILLER_63_2955 ();
 sg13g2_decap_8 FILLER_63_2962 ();
 sg13g2_decap_8 FILLER_63_2969 ();
 sg13g2_decap_8 FILLER_63_2976 ();
 sg13g2_decap_8 FILLER_63_2983 ();
 sg13g2_decap_8 FILLER_63_2990 ();
 sg13g2_decap_8 FILLER_63_2997 ();
 sg13g2_decap_8 FILLER_63_3004 ();
 sg13g2_decap_8 FILLER_63_3011 ();
 sg13g2_decap_8 FILLER_63_3018 ();
 sg13g2_decap_8 FILLER_63_3025 ();
 sg13g2_decap_8 FILLER_63_3032 ();
 sg13g2_decap_8 FILLER_63_3039 ();
 sg13g2_decap_8 FILLER_63_3046 ();
 sg13g2_decap_8 FILLER_63_3053 ();
 sg13g2_decap_8 FILLER_63_3060 ();
 sg13g2_decap_8 FILLER_63_3067 ();
 sg13g2_decap_8 FILLER_63_3074 ();
 sg13g2_decap_8 FILLER_63_3081 ();
 sg13g2_decap_8 FILLER_63_3088 ();
 sg13g2_decap_8 FILLER_63_3095 ();
 sg13g2_decap_8 FILLER_63_3102 ();
 sg13g2_decap_8 FILLER_63_3109 ();
 sg13g2_decap_8 FILLER_63_3116 ();
 sg13g2_decap_8 FILLER_63_3123 ();
 sg13g2_decap_8 FILLER_63_3130 ();
 sg13g2_decap_8 FILLER_63_3137 ();
 sg13g2_decap_8 FILLER_63_3144 ();
 sg13g2_decap_8 FILLER_63_3151 ();
 sg13g2_decap_8 FILLER_63_3158 ();
 sg13g2_decap_8 FILLER_63_3165 ();
 sg13g2_decap_8 FILLER_63_3172 ();
 sg13g2_decap_8 FILLER_63_3179 ();
 sg13g2_decap_8 FILLER_63_3186 ();
 sg13g2_decap_8 FILLER_63_3193 ();
 sg13g2_decap_8 FILLER_63_3200 ();
 sg13g2_decap_8 FILLER_63_3207 ();
 sg13g2_decap_8 FILLER_63_3214 ();
 sg13g2_decap_8 FILLER_63_3221 ();
 sg13g2_decap_8 FILLER_63_3228 ();
 sg13g2_decap_8 FILLER_63_3235 ();
 sg13g2_decap_8 FILLER_63_3242 ();
 sg13g2_decap_8 FILLER_63_3249 ();
 sg13g2_decap_8 FILLER_63_3256 ();
 sg13g2_decap_8 FILLER_63_3263 ();
 sg13g2_decap_8 FILLER_63_3270 ();
 sg13g2_decap_8 FILLER_63_3277 ();
 sg13g2_decap_8 FILLER_63_3284 ();
 sg13g2_decap_8 FILLER_63_3291 ();
 sg13g2_decap_8 FILLER_63_3298 ();
 sg13g2_decap_8 FILLER_63_3305 ();
 sg13g2_decap_8 FILLER_63_3312 ();
 sg13g2_decap_8 FILLER_63_3319 ();
 sg13g2_decap_8 FILLER_63_3326 ();
 sg13g2_decap_8 FILLER_63_3333 ();
 sg13g2_decap_8 FILLER_63_3340 ();
 sg13g2_decap_8 FILLER_63_3347 ();
 sg13g2_decap_8 FILLER_63_3354 ();
 sg13g2_decap_8 FILLER_63_3361 ();
 sg13g2_decap_8 FILLER_63_3368 ();
 sg13g2_decap_8 FILLER_63_3375 ();
 sg13g2_decap_8 FILLER_63_3382 ();
 sg13g2_decap_8 FILLER_63_3389 ();
 sg13g2_decap_8 FILLER_63_3396 ();
 sg13g2_decap_8 FILLER_63_3403 ();
 sg13g2_decap_8 FILLER_63_3410 ();
 sg13g2_decap_8 FILLER_63_3417 ();
 sg13g2_decap_8 FILLER_63_3424 ();
 sg13g2_decap_8 FILLER_63_3431 ();
 sg13g2_decap_8 FILLER_63_3438 ();
 sg13g2_decap_8 FILLER_63_3445 ();
 sg13g2_decap_8 FILLER_63_3452 ();
 sg13g2_decap_8 FILLER_63_3459 ();
 sg13g2_decap_8 FILLER_63_3466 ();
 sg13g2_decap_8 FILLER_63_3473 ();
 sg13g2_decap_8 FILLER_63_3480 ();
 sg13g2_decap_8 FILLER_63_3487 ();
 sg13g2_decap_8 FILLER_63_3494 ();
 sg13g2_decap_8 FILLER_63_3501 ();
 sg13g2_decap_8 FILLER_63_3508 ();
 sg13g2_decap_8 FILLER_63_3515 ();
 sg13g2_decap_8 FILLER_63_3522 ();
 sg13g2_decap_8 FILLER_63_3529 ();
 sg13g2_decap_8 FILLER_63_3536 ();
 sg13g2_decap_8 FILLER_63_3543 ();
 sg13g2_decap_8 FILLER_63_3550 ();
 sg13g2_decap_8 FILLER_63_3557 ();
 sg13g2_decap_8 FILLER_63_3564 ();
 sg13g2_decap_8 FILLER_63_3571 ();
 sg13g2_fill_2 FILLER_63_3578 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_168 ();
 sg13g2_decap_8 FILLER_64_175 ();
 sg13g2_decap_8 FILLER_64_182 ();
 sg13g2_decap_8 FILLER_64_189 ();
 sg13g2_decap_8 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_decap_8 FILLER_64_217 ();
 sg13g2_decap_8 FILLER_64_224 ();
 sg13g2_decap_8 FILLER_64_231 ();
 sg13g2_decap_8 FILLER_64_238 ();
 sg13g2_decap_8 FILLER_64_245 ();
 sg13g2_decap_8 FILLER_64_252 ();
 sg13g2_decap_8 FILLER_64_259 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_273 ();
 sg13g2_decap_8 FILLER_64_280 ();
 sg13g2_decap_8 FILLER_64_287 ();
 sg13g2_decap_8 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_308 ();
 sg13g2_decap_8 FILLER_64_315 ();
 sg13g2_decap_8 FILLER_64_322 ();
 sg13g2_decap_8 FILLER_64_329 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_decap_8 FILLER_64_343 ();
 sg13g2_decap_8 FILLER_64_350 ();
 sg13g2_decap_8 FILLER_64_357 ();
 sg13g2_decap_8 FILLER_64_364 ();
 sg13g2_decap_8 FILLER_64_371 ();
 sg13g2_decap_8 FILLER_64_378 ();
 sg13g2_decap_8 FILLER_64_385 ();
 sg13g2_decap_8 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_399 ();
 sg13g2_decap_8 FILLER_64_406 ();
 sg13g2_decap_8 FILLER_64_413 ();
 sg13g2_decap_8 FILLER_64_420 ();
 sg13g2_decap_8 FILLER_64_466 ();
 sg13g2_decap_8 FILLER_64_473 ();
 sg13g2_decap_8 FILLER_64_480 ();
 sg13g2_fill_1 FILLER_64_487 ();
 sg13g2_decap_8 FILLER_64_519 ();
 sg13g2_decap_8 FILLER_64_526 ();
 sg13g2_fill_2 FILLER_64_533 ();
 sg13g2_decap_8 FILLER_64_584 ();
 sg13g2_decap_4 FILLER_64_591 ();
 sg13g2_fill_2 FILLER_64_595 ();
 sg13g2_decap_8 FILLER_64_662 ();
 sg13g2_decap_8 FILLER_64_669 ();
 sg13g2_decap_8 FILLER_64_676 ();
 sg13g2_decap_8 FILLER_64_683 ();
 sg13g2_decap_8 FILLER_64_690 ();
 sg13g2_decap_8 FILLER_64_701 ();
 sg13g2_decap_8 FILLER_64_708 ();
 sg13g2_decap_8 FILLER_64_715 ();
 sg13g2_decap_8 FILLER_64_722 ();
 sg13g2_decap_4 FILLER_64_729 ();
 sg13g2_fill_2 FILLER_64_733 ();
 sg13g2_decap_8 FILLER_64_740 ();
 sg13g2_fill_1 FILLER_64_747 ();
 sg13g2_fill_2 FILLER_64_774 ();
 sg13g2_fill_1 FILLER_64_776 ();
 sg13g2_fill_2 FILLER_64_781 ();
 sg13g2_decap_8 FILLER_64_821 ();
 sg13g2_fill_1 FILLER_64_928 ();
 sg13g2_fill_1 FILLER_64_981 ();
 sg13g2_decap_8 FILLER_64_995 ();
 sg13g2_fill_1 FILLER_64_1002 ();
 sg13g2_fill_2 FILLER_64_1014 ();
 sg13g2_decap_8 FILLER_64_1020 ();
 sg13g2_fill_2 FILLER_64_1027 ();
 sg13g2_fill_1 FILLER_64_1029 ();
 sg13g2_decap_8 FILLER_64_1056 ();
 sg13g2_decap_4 FILLER_64_1063 ();
 sg13g2_fill_2 FILLER_64_1067 ();
 sg13g2_fill_2 FILLER_64_1072 ();
 sg13g2_fill_2 FILLER_64_1085 ();
 sg13g2_decap_4 FILLER_64_1165 ();
 sg13g2_decap_8 FILLER_64_1270 ();
 sg13g2_decap_8 FILLER_64_1277 ();
 sg13g2_decap_8 FILLER_64_1284 ();
 sg13g2_decap_4 FILLER_64_1291 ();
 sg13g2_fill_2 FILLER_64_1295 ();
 sg13g2_fill_2 FILLER_64_1307 ();
 sg13g2_decap_8 FILLER_64_1333 ();
 sg13g2_decap_4 FILLER_64_1340 ();
 sg13g2_decap_8 FILLER_64_1378 ();
 sg13g2_fill_1 FILLER_64_1385 ();
 sg13g2_decap_8 FILLER_64_1418 ();
 sg13g2_decap_8 FILLER_64_1425 ();
 sg13g2_fill_1 FILLER_64_1432 ();
 sg13g2_decap_8 FILLER_64_1473 ();
 sg13g2_fill_2 FILLER_64_1480 ();
 sg13g2_fill_1 FILLER_64_1519 ();
 sg13g2_fill_2 FILLER_64_1526 ();
 sg13g2_fill_1 FILLER_64_1528 ();
 sg13g2_decap_8 FILLER_64_1543 ();
 sg13g2_decap_4 FILLER_64_1550 ();
 sg13g2_fill_1 FILLER_64_1554 ();
 sg13g2_fill_2 FILLER_64_1561 ();
 sg13g2_decap_8 FILLER_64_1595 ();
 sg13g2_decap_8 FILLER_64_1602 ();
 sg13g2_decap_8 FILLER_64_1609 ();
 sg13g2_decap_4 FILLER_64_1616 ();
 sg13g2_fill_1 FILLER_64_1620 ();
 sg13g2_decap_8 FILLER_64_1647 ();
 sg13g2_decap_8 FILLER_64_1654 ();
 sg13g2_decap_8 FILLER_64_1661 ();
 sg13g2_decap_8 FILLER_64_1668 ();
 sg13g2_fill_2 FILLER_64_1675 ();
 sg13g2_fill_1 FILLER_64_1677 ();
 sg13g2_fill_2 FILLER_64_1683 ();
 sg13g2_fill_1 FILLER_64_1685 ();
 sg13g2_decap_8 FILLER_64_1733 ();
 sg13g2_decap_8 FILLER_64_1740 ();
 sg13g2_decap_8 FILLER_64_1747 ();
 sg13g2_decap_8 FILLER_64_1754 ();
 sg13g2_decap_4 FILLER_64_1761 ();
 sg13g2_fill_2 FILLER_64_1765 ();
 sg13g2_decap_4 FILLER_64_1775 ();
 sg13g2_decap_8 FILLER_64_1785 ();
 sg13g2_decap_4 FILLER_64_1792 ();
 sg13g2_fill_2 FILLER_64_1796 ();
 sg13g2_decap_8 FILLER_64_1816 ();
 sg13g2_decap_8 FILLER_64_1823 ();
 sg13g2_decap_8 FILLER_64_1890 ();
 sg13g2_decap_4 FILLER_64_1897 ();
 sg13g2_fill_1 FILLER_64_1901 ();
 sg13g2_decap_8 FILLER_64_1980 ();
 sg13g2_decap_8 FILLER_64_1987 ();
 sg13g2_decap_4 FILLER_64_1994 ();
 sg13g2_fill_1 FILLER_64_1998 ();
 sg13g2_fill_1 FILLER_64_2017 ();
 sg13g2_decap_8 FILLER_64_2048 ();
 sg13g2_decap_8 FILLER_64_2055 ();
 sg13g2_decap_8 FILLER_64_2062 ();
 sg13g2_fill_2 FILLER_64_2069 ();
 sg13g2_fill_2 FILLER_64_2081 ();
 sg13g2_decap_8 FILLER_64_2116 ();
 sg13g2_decap_8 FILLER_64_2123 ();
 sg13g2_decap_8 FILLER_64_2130 ();
 sg13g2_decap_8 FILLER_64_2137 ();
 sg13g2_decap_8 FILLER_64_2144 ();
 sg13g2_decap_4 FILLER_64_2151 ();
 sg13g2_fill_1 FILLER_64_2155 ();
 sg13g2_fill_1 FILLER_64_2167 ();
 sg13g2_decap_8 FILLER_64_2200 ();
 sg13g2_decap_8 FILLER_64_2207 ();
 sg13g2_decap_8 FILLER_64_2214 ();
 sg13g2_decap_8 FILLER_64_2221 ();
 sg13g2_decap_8 FILLER_64_2228 ();
 sg13g2_decap_8 FILLER_64_2235 ();
 sg13g2_decap_8 FILLER_64_2242 ();
 sg13g2_decap_8 FILLER_64_2249 ();
 sg13g2_decap_8 FILLER_64_2256 ();
 sg13g2_decap_8 FILLER_64_2263 ();
 sg13g2_decap_8 FILLER_64_2270 ();
 sg13g2_decap_8 FILLER_64_2277 ();
 sg13g2_decap_8 FILLER_64_2284 ();
 sg13g2_decap_8 FILLER_64_2291 ();
 sg13g2_decap_8 FILLER_64_2298 ();
 sg13g2_decap_8 FILLER_64_2305 ();
 sg13g2_decap_8 FILLER_64_2312 ();
 sg13g2_decap_8 FILLER_64_2319 ();
 sg13g2_decap_8 FILLER_64_2326 ();
 sg13g2_decap_8 FILLER_64_2333 ();
 sg13g2_decap_8 FILLER_64_2340 ();
 sg13g2_decap_8 FILLER_64_2347 ();
 sg13g2_decap_8 FILLER_64_2354 ();
 sg13g2_decap_8 FILLER_64_2361 ();
 sg13g2_decap_8 FILLER_64_2368 ();
 sg13g2_decap_8 FILLER_64_2375 ();
 sg13g2_decap_8 FILLER_64_2382 ();
 sg13g2_decap_8 FILLER_64_2389 ();
 sg13g2_decap_8 FILLER_64_2396 ();
 sg13g2_decap_8 FILLER_64_2403 ();
 sg13g2_decap_8 FILLER_64_2410 ();
 sg13g2_decap_8 FILLER_64_2417 ();
 sg13g2_decap_8 FILLER_64_2424 ();
 sg13g2_decap_8 FILLER_64_2431 ();
 sg13g2_decap_8 FILLER_64_2438 ();
 sg13g2_decap_8 FILLER_64_2445 ();
 sg13g2_decap_8 FILLER_64_2452 ();
 sg13g2_decap_8 FILLER_64_2459 ();
 sg13g2_decap_8 FILLER_64_2466 ();
 sg13g2_decap_8 FILLER_64_2473 ();
 sg13g2_decap_8 FILLER_64_2480 ();
 sg13g2_decap_8 FILLER_64_2487 ();
 sg13g2_decap_8 FILLER_64_2494 ();
 sg13g2_decap_8 FILLER_64_2501 ();
 sg13g2_decap_8 FILLER_64_2508 ();
 sg13g2_decap_8 FILLER_64_2515 ();
 sg13g2_decap_8 FILLER_64_2522 ();
 sg13g2_decap_8 FILLER_64_2529 ();
 sg13g2_decap_8 FILLER_64_2536 ();
 sg13g2_decap_8 FILLER_64_2543 ();
 sg13g2_decap_8 FILLER_64_2550 ();
 sg13g2_decap_8 FILLER_64_2557 ();
 sg13g2_decap_8 FILLER_64_2564 ();
 sg13g2_decap_8 FILLER_64_2571 ();
 sg13g2_decap_8 FILLER_64_2578 ();
 sg13g2_decap_8 FILLER_64_2585 ();
 sg13g2_decap_8 FILLER_64_2592 ();
 sg13g2_decap_8 FILLER_64_2599 ();
 sg13g2_decap_8 FILLER_64_2606 ();
 sg13g2_decap_8 FILLER_64_2613 ();
 sg13g2_decap_8 FILLER_64_2620 ();
 sg13g2_fill_2 FILLER_64_2627 ();
 sg13g2_fill_1 FILLER_64_2629 ();
 sg13g2_decap_8 FILLER_64_2656 ();
 sg13g2_decap_8 FILLER_64_2663 ();
 sg13g2_decap_8 FILLER_64_2670 ();
 sg13g2_decap_8 FILLER_64_2677 ();
 sg13g2_decap_8 FILLER_64_2684 ();
 sg13g2_decap_8 FILLER_64_2691 ();
 sg13g2_decap_8 FILLER_64_2698 ();
 sg13g2_decap_4 FILLER_64_2705 ();
 sg13g2_fill_1 FILLER_64_2709 ();
 sg13g2_decap_8 FILLER_64_2715 ();
 sg13g2_decap_8 FILLER_64_2722 ();
 sg13g2_decap_8 FILLER_64_2729 ();
 sg13g2_decap_8 FILLER_64_2736 ();
 sg13g2_decap_8 FILLER_64_2743 ();
 sg13g2_decap_8 FILLER_64_2750 ();
 sg13g2_decap_8 FILLER_64_2757 ();
 sg13g2_decap_8 FILLER_64_2764 ();
 sg13g2_decap_8 FILLER_64_2771 ();
 sg13g2_decap_8 FILLER_64_2778 ();
 sg13g2_decap_8 FILLER_64_2785 ();
 sg13g2_decap_8 FILLER_64_2792 ();
 sg13g2_decap_8 FILLER_64_2799 ();
 sg13g2_fill_2 FILLER_64_2806 ();
 sg13g2_fill_1 FILLER_64_2808 ();
 sg13g2_decap_8 FILLER_64_2835 ();
 sg13g2_decap_4 FILLER_64_2842 ();
 sg13g2_fill_2 FILLER_64_2846 ();
 sg13g2_decap_8 FILLER_64_2874 ();
 sg13g2_decap_8 FILLER_64_2881 ();
 sg13g2_decap_8 FILLER_64_2888 ();
 sg13g2_decap_8 FILLER_64_2895 ();
 sg13g2_decap_8 FILLER_64_2902 ();
 sg13g2_decap_8 FILLER_64_2909 ();
 sg13g2_decap_8 FILLER_64_2916 ();
 sg13g2_decap_8 FILLER_64_2923 ();
 sg13g2_decap_8 FILLER_64_2930 ();
 sg13g2_decap_8 FILLER_64_2937 ();
 sg13g2_decap_8 FILLER_64_2944 ();
 sg13g2_decap_8 FILLER_64_2951 ();
 sg13g2_decap_8 FILLER_64_2958 ();
 sg13g2_decap_8 FILLER_64_2965 ();
 sg13g2_decap_8 FILLER_64_2972 ();
 sg13g2_decap_8 FILLER_64_2979 ();
 sg13g2_decap_8 FILLER_64_2986 ();
 sg13g2_decap_8 FILLER_64_2993 ();
 sg13g2_decap_8 FILLER_64_3000 ();
 sg13g2_decap_8 FILLER_64_3007 ();
 sg13g2_decap_8 FILLER_64_3014 ();
 sg13g2_decap_8 FILLER_64_3021 ();
 sg13g2_decap_8 FILLER_64_3028 ();
 sg13g2_decap_8 FILLER_64_3035 ();
 sg13g2_decap_8 FILLER_64_3042 ();
 sg13g2_decap_8 FILLER_64_3049 ();
 sg13g2_decap_8 FILLER_64_3056 ();
 sg13g2_decap_8 FILLER_64_3063 ();
 sg13g2_decap_8 FILLER_64_3070 ();
 sg13g2_decap_8 FILLER_64_3077 ();
 sg13g2_decap_8 FILLER_64_3084 ();
 sg13g2_decap_8 FILLER_64_3091 ();
 sg13g2_decap_8 FILLER_64_3098 ();
 sg13g2_decap_8 FILLER_64_3105 ();
 sg13g2_decap_8 FILLER_64_3112 ();
 sg13g2_decap_8 FILLER_64_3119 ();
 sg13g2_decap_8 FILLER_64_3126 ();
 sg13g2_decap_8 FILLER_64_3133 ();
 sg13g2_decap_8 FILLER_64_3140 ();
 sg13g2_decap_8 FILLER_64_3147 ();
 sg13g2_decap_8 FILLER_64_3154 ();
 sg13g2_decap_8 FILLER_64_3161 ();
 sg13g2_decap_8 FILLER_64_3168 ();
 sg13g2_decap_8 FILLER_64_3175 ();
 sg13g2_decap_8 FILLER_64_3182 ();
 sg13g2_decap_8 FILLER_64_3189 ();
 sg13g2_decap_8 FILLER_64_3196 ();
 sg13g2_decap_8 FILLER_64_3203 ();
 sg13g2_decap_8 FILLER_64_3210 ();
 sg13g2_decap_8 FILLER_64_3217 ();
 sg13g2_decap_8 FILLER_64_3224 ();
 sg13g2_decap_8 FILLER_64_3231 ();
 sg13g2_decap_8 FILLER_64_3238 ();
 sg13g2_decap_8 FILLER_64_3245 ();
 sg13g2_decap_8 FILLER_64_3252 ();
 sg13g2_decap_8 FILLER_64_3259 ();
 sg13g2_decap_8 FILLER_64_3266 ();
 sg13g2_decap_8 FILLER_64_3273 ();
 sg13g2_decap_8 FILLER_64_3280 ();
 sg13g2_decap_8 FILLER_64_3287 ();
 sg13g2_decap_8 FILLER_64_3294 ();
 sg13g2_decap_8 FILLER_64_3301 ();
 sg13g2_decap_8 FILLER_64_3308 ();
 sg13g2_decap_8 FILLER_64_3315 ();
 sg13g2_decap_8 FILLER_64_3322 ();
 sg13g2_decap_8 FILLER_64_3329 ();
 sg13g2_decap_8 FILLER_64_3336 ();
 sg13g2_decap_8 FILLER_64_3343 ();
 sg13g2_decap_8 FILLER_64_3350 ();
 sg13g2_decap_8 FILLER_64_3357 ();
 sg13g2_decap_8 FILLER_64_3364 ();
 sg13g2_decap_8 FILLER_64_3371 ();
 sg13g2_decap_8 FILLER_64_3378 ();
 sg13g2_decap_8 FILLER_64_3385 ();
 sg13g2_decap_8 FILLER_64_3392 ();
 sg13g2_decap_8 FILLER_64_3399 ();
 sg13g2_decap_8 FILLER_64_3406 ();
 sg13g2_decap_8 FILLER_64_3413 ();
 sg13g2_decap_8 FILLER_64_3420 ();
 sg13g2_decap_8 FILLER_64_3427 ();
 sg13g2_decap_8 FILLER_64_3434 ();
 sg13g2_decap_8 FILLER_64_3441 ();
 sg13g2_decap_8 FILLER_64_3448 ();
 sg13g2_decap_8 FILLER_64_3455 ();
 sg13g2_decap_8 FILLER_64_3462 ();
 sg13g2_decap_8 FILLER_64_3469 ();
 sg13g2_decap_8 FILLER_64_3476 ();
 sg13g2_decap_8 FILLER_64_3483 ();
 sg13g2_decap_8 FILLER_64_3490 ();
 sg13g2_decap_8 FILLER_64_3497 ();
 sg13g2_decap_8 FILLER_64_3504 ();
 sg13g2_decap_8 FILLER_64_3511 ();
 sg13g2_decap_8 FILLER_64_3518 ();
 sg13g2_decap_8 FILLER_64_3525 ();
 sg13g2_decap_8 FILLER_64_3532 ();
 sg13g2_decap_8 FILLER_64_3539 ();
 sg13g2_decap_8 FILLER_64_3546 ();
 sg13g2_decap_8 FILLER_64_3553 ();
 sg13g2_decap_8 FILLER_64_3560 ();
 sg13g2_decap_8 FILLER_64_3567 ();
 sg13g2_decap_4 FILLER_64_3574 ();
 sg13g2_fill_2 FILLER_64_3578 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_189 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_203 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_245 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_decap_8 FILLER_65_259 ();
 sg13g2_decap_8 FILLER_65_266 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_8 FILLER_65_280 ();
 sg13g2_decap_8 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_294 ();
 sg13g2_decap_8 FILLER_65_301 ();
 sg13g2_decap_8 FILLER_65_308 ();
 sg13g2_decap_8 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_decap_8 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_decap_8 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_65_406 ();
 sg13g2_decap_8 FILLER_65_413 ();
 sg13g2_decap_8 FILLER_65_420 ();
 sg13g2_decap_8 FILLER_65_427 ();
 sg13g2_fill_2 FILLER_65_434 ();
 sg13g2_decap_8 FILLER_65_484 ();
 sg13g2_decap_4 FILLER_65_491 ();
 sg13g2_fill_1 FILLER_65_495 ();
 sg13g2_decap_8 FILLER_65_512 ();
 sg13g2_decap_4 FILLER_65_519 ();
 sg13g2_fill_1 FILLER_65_528 ();
 sg13g2_decap_8 FILLER_65_533 ();
 sg13g2_decap_8 FILLER_65_540 ();
 sg13g2_fill_2 FILLER_65_547 ();
 sg13g2_fill_1 FILLER_65_549 ();
 sg13g2_decap_8 FILLER_65_576 ();
 sg13g2_decap_8 FILLER_65_583 ();
 sg13g2_fill_1 FILLER_65_590 ();
 sg13g2_fill_1 FILLER_65_632 ();
 sg13g2_decap_8 FILLER_65_642 ();
 sg13g2_decap_8 FILLER_65_649 ();
 sg13g2_decap_8 FILLER_65_656 ();
 sg13g2_decap_4 FILLER_65_663 ();
 sg13g2_fill_2 FILLER_65_667 ();
 sg13g2_decap_8 FILLER_65_698 ();
 sg13g2_decap_8 FILLER_65_705 ();
 sg13g2_fill_1 FILLER_65_712 ();
 sg13g2_decap_4 FILLER_65_717 ();
 sg13g2_fill_2 FILLER_65_729 ();
 sg13g2_fill_1 FILLER_65_731 ();
 sg13g2_fill_2 FILLER_65_758 ();
 sg13g2_fill_1 FILLER_65_760 ();
 sg13g2_decap_4 FILLER_65_799 ();
 sg13g2_fill_1 FILLER_65_803 ();
 sg13g2_decap_4 FILLER_65_856 ();
 sg13g2_fill_2 FILLER_65_893 ();
 sg13g2_decap_4 FILLER_65_961 ();
 sg13g2_fill_1 FILLER_65_965 ();
 sg13g2_fill_2 FILLER_65_973 ();
 sg13g2_fill_1 FILLER_65_990 ();
 sg13g2_fill_2 FILLER_65_1004 ();
 sg13g2_decap_8 FILLER_65_1032 ();
 sg13g2_decap_8 FILLER_65_1039 ();
 sg13g2_decap_8 FILLER_65_1046 ();
 sg13g2_decap_8 FILLER_65_1053 ();
 sg13g2_fill_2 FILLER_65_1060 ();
 sg13g2_fill_1 FILLER_65_1062 ();
 sg13g2_fill_2 FILLER_65_1099 ();
 sg13g2_fill_1 FILLER_65_1101 ();
 sg13g2_decap_4 FILLER_65_1141 ();
 sg13g2_fill_2 FILLER_65_1145 ();
 sg13g2_fill_2 FILLER_65_1173 ();
 sg13g2_fill_2 FILLER_65_1201 ();
 sg13g2_fill_1 FILLER_65_1203 ();
 sg13g2_decap_8 FILLER_65_1209 ();
 sg13g2_decap_4 FILLER_65_1216 ();
 sg13g2_fill_2 FILLER_65_1220 ();
 sg13g2_decap_8 FILLER_65_1259 ();
 sg13g2_fill_1 FILLER_65_1266 ();
 sg13g2_decap_8 FILLER_65_1310 ();
 sg13g2_decap_8 FILLER_65_1317 ();
 sg13g2_fill_2 FILLER_65_1324 ();
 sg13g2_fill_1 FILLER_65_1326 ();
 sg13g2_decap_8 FILLER_65_1379 ();
 sg13g2_decap_8 FILLER_65_1386 ();
 sg13g2_decap_8 FILLER_65_1393 ();
 sg13g2_decap_8 FILLER_65_1400 ();
 sg13g2_decap_8 FILLER_65_1407 ();
 sg13g2_decap_8 FILLER_65_1414 ();
 sg13g2_decap_8 FILLER_65_1421 ();
 sg13g2_fill_1 FILLER_65_1428 ();
 sg13g2_decap_8 FILLER_65_1467 ();
 sg13g2_fill_1 FILLER_65_1474 ();
 sg13g2_decap_4 FILLER_65_1526 ();
 sg13g2_fill_1 FILLER_65_1530 ();
 sg13g2_decap_8 FILLER_65_1539 ();
 sg13g2_fill_2 FILLER_65_1546 ();
 sg13g2_decap_8 FILLER_65_1600 ();
 sg13g2_decap_8 FILLER_65_1607 ();
 sg13g2_fill_1 FILLER_65_1614 ();
 sg13g2_decap_4 FILLER_65_1735 ();
 sg13g2_fill_1 FILLER_65_1771 ();
 sg13g2_decap_8 FILLER_65_1798 ();
 sg13g2_decap_8 FILLER_65_1805 ();
 sg13g2_decap_8 FILLER_65_1812 ();
 sg13g2_decap_8 FILLER_65_1819 ();
 sg13g2_fill_2 FILLER_65_1891 ();
 sg13g2_fill_1 FILLER_65_1893 ();
 sg13g2_decap_8 FILLER_65_1985 ();
 sg13g2_fill_1 FILLER_65_1992 ();
 sg13g2_decap_4 FILLER_65_2025 ();
 sg13g2_decap_8 FILLER_65_2037 ();
 sg13g2_decap_8 FILLER_65_2044 ();
 sg13g2_decap_8 FILLER_65_2051 ();
 sg13g2_decap_4 FILLER_65_2058 ();
 sg13g2_decap_8 FILLER_65_2067 ();
 sg13g2_decap_8 FILLER_65_2074 ();
 sg13g2_fill_2 FILLER_65_2081 ();
 sg13g2_decap_8 FILLER_65_2109 ();
 sg13g2_decap_8 FILLER_65_2116 ();
 sg13g2_decap_8 FILLER_65_2123 ();
 sg13g2_decap_8 FILLER_65_2130 ();
 sg13g2_decap_8 FILLER_65_2137 ();
 sg13g2_fill_1 FILLER_65_2144 ();
 sg13g2_fill_2 FILLER_65_2166 ();
 sg13g2_fill_1 FILLER_65_2168 ();
 sg13g2_decap_8 FILLER_65_2221 ();
 sg13g2_decap_8 FILLER_65_2228 ();
 sg13g2_decap_8 FILLER_65_2235 ();
 sg13g2_decap_8 FILLER_65_2242 ();
 sg13g2_decap_8 FILLER_65_2249 ();
 sg13g2_decap_8 FILLER_65_2256 ();
 sg13g2_decap_8 FILLER_65_2263 ();
 sg13g2_decap_8 FILLER_65_2270 ();
 sg13g2_decap_8 FILLER_65_2277 ();
 sg13g2_decap_8 FILLER_65_2284 ();
 sg13g2_decap_8 FILLER_65_2291 ();
 sg13g2_decap_8 FILLER_65_2298 ();
 sg13g2_decap_8 FILLER_65_2305 ();
 sg13g2_decap_8 FILLER_65_2312 ();
 sg13g2_decap_8 FILLER_65_2319 ();
 sg13g2_decap_8 FILLER_65_2326 ();
 sg13g2_decap_8 FILLER_65_2333 ();
 sg13g2_decap_8 FILLER_65_2340 ();
 sg13g2_decap_8 FILLER_65_2347 ();
 sg13g2_decap_8 FILLER_65_2354 ();
 sg13g2_decap_8 FILLER_65_2361 ();
 sg13g2_decap_8 FILLER_65_2368 ();
 sg13g2_decap_8 FILLER_65_2375 ();
 sg13g2_decap_8 FILLER_65_2382 ();
 sg13g2_decap_8 FILLER_65_2389 ();
 sg13g2_decap_8 FILLER_65_2396 ();
 sg13g2_decap_8 FILLER_65_2403 ();
 sg13g2_decap_8 FILLER_65_2410 ();
 sg13g2_decap_8 FILLER_65_2417 ();
 sg13g2_decap_8 FILLER_65_2424 ();
 sg13g2_decap_8 FILLER_65_2431 ();
 sg13g2_decap_8 FILLER_65_2438 ();
 sg13g2_decap_8 FILLER_65_2445 ();
 sg13g2_decap_8 FILLER_65_2452 ();
 sg13g2_decap_8 FILLER_65_2459 ();
 sg13g2_decap_8 FILLER_65_2466 ();
 sg13g2_decap_8 FILLER_65_2473 ();
 sg13g2_decap_8 FILLER_65_2480 ();
 sg13g2_decap_8 FILLER_65_2487 ();
 sg13g2_decap_8 FILLER_65_2494 ();
 sg13g2_decap_8 FILLER_65_2501 ();
 sg13g2_decap_8 FILLER_65_2508 ();
 sg13g2_decap_8 FILLER_65_2515 ();
 sg13g2_decap_8 FILLER_65_2522 ();
 sg13g2_decap_8 FILLER_65_2529 ();
 sg13g2_decap_8 FILLER_65_2536 ();
 sg13g2_decap_8 FILLER_65_2543 ();
 sg13g2_decap_8 FILLER_65_2550 ();
 sg13g2_decap_8 FILLER_65_2557 ();
 sg13g2_decap_8 FILLER_65_2564 ();
 sg13g2_decap_8 FILLER_65_2571 ();
 sg13g2_decap_8 FILLER_65_2578 ();
 sg13g2_decap_8 FILLER_65_2585 ();
 sg13g2_decap_8 FILLER_65_2592 ();
 sg13g2_decap_8 FILLER_65_2599 ();
 sg13g2_decap_8 FILLER_65_2606 ();
 sg13g2_decap_8 FILLER_65_2613 ();
 sg13g2_decap_8 FILLER_65_2620 ();
 sg13g2_decap_8 FILLER_65_2627 ();
 sg13g2_decap_8 FILLER_65_2634 ();
 sg13g2_decap_8 FILLER_65_2641 ();
 sg13g2_decap_8 FILLER_65_2648 ();
 sg13g2_decap_8 FILLER_65_2655 ();
 sg13g2_decap_8 FILLER_65_2662 ();
 sg13g2_decap_8 FILLER_65_2669 ();
 sg13g2_decap_8 FILLER_65_2676 ();
 sg13g2_decap_8 FILLER_65_2683 ();
 sg13g2_decap_8 FILLER_65_2690 ();
 sg13g2_decap_8 FILLER_65_2697 ();
 sg13g2_decap_8 FILLER_65_2704 ();
 sg13g2_decap_8 FILLER_65_2711 ();
 sg13g2_decap_8 FILLER_65_2718 ();
 sg13g2_decap_8 FILLER_65_2725 ();
 sg13g2_decap_8 FILLER_65_2732 ();
 sg13g2_decap_8 FILLER_65_2739 ();
 sg13g2_decap_8 FILLER_65_2746 ();
 sg13g2_decap_8 FILLER_65_2753 ();
 sg13g2_decap_8 FILLER_65_2760 ();
 sg13g2_decap_8 FILLER_65_2767 ();
 sg13g2_decap_8 FILLER_65_2774 ();
 sg13g2_decap_8 FILLER_65_2781 ();
 sg13g2_decap_8 FILLER_65_2788 ();
 sg13g2_decap_8 FILLER_65_2795 ();
 sg13g2_decap_8 FILLER_65_2802 ();
 sg13g2_decap_8 FILLER_65_2809 ();
 sg13g2_decap_8 FILLER_65_2816 ();
 sg13g2_decap_8 FILLER_65_2823 ();
 sg13g2_decap_8 FILLER_65_2830 ();
 sg13g2_decap_8 FILLER_65_2837 ();
 sg13g2_decap_8 FILLER_65_2844 ();
 sg13g2_decap_8 FILLER_65_2851 ();
 sg13g2_decap_8 FILLER_65_2858 ();
 sg13g2_decap_8 FILLER_65_2865 ();
 sg13g2_decap_8 FILLER_65_2872 ();
 sg13g2_decap_8 FILLER_65_2879 ();
 sg13g2_decap_8 FILLER_65_2886 ();
 sg13g2_decap_8 FILLER_65_2893 ();
 sg13g2_decap_8 FILLER_65_2900 ();
 sg13g2_decap_8 FILLER_65_2907 ();
 sg13g2_decap_8 FILLER_65_2914 ();
 sg13g2_decap_8 FILLER_65_2921 ();
 sg13g2_decap_8 FILLER_65_2928 ();
 sg13g2_decap_8 FILLER_65_2935 ();
 sg13g2_decap_8 FILLER_65_2942 ();
 sg13g2_decap_8 FILLER_65_2949 ();
 sg13g2_decap_8 FILLER_65_2956 ();
 sg13g2_decap_8 FILLER_65_2963 ();
 sg13g2_decap_8 FILLER_65_2970 ();
 sg13g2_decap_8 FILLER_65_2977 ();
 sg13g2_decap_8 FILLER_65_2984 ();
 sg13g2_decap_8 FILLER_65_2991 ();
 sg13g2_decap_8 FILLER_65_2998 ();
 sg13g2_decap_8 FILLER_65_3005 ();
 sg13g2_decap_8 FILLER_65_3012 ();
 sg13g2_decap_8 FILLER_65_3019 ();
 sg13g2_decap_8 FILLER_65_3026 ();
 sg13g2_decap_8 FILLER_65_3033 ();
 sg13g2_decap_8 FILLER_65_3040 ();
 sg13g2_decap_8 FILLER_65_3047 ();
 sg13g2_decap_8 FILLER_65_3054 ();
 sg13g2_decap_8 FILLER_65_3061 ();
 sg13g2_decap_8 FILLER_65_3068 ();
 sg13g2_decap_8 FILLER_65_3075 ();
 sg13g2_decap_8 FILLER_65_3082 ();
 sg13g2_decap_8 FILLER_65_3089 ();
 sg13g2_decap_8 FILLER_65_3096 ();
 sg13g2_decap_8 FILLER_65_3103 ();
 sg13g2_decap_8 FILLER_65_3110 ();
 sg13g2_decap_8 FILLER_65_3117 ();
 sg13g2_decap_8 FILLER_65_3124 ();
 sg13g2_decap_8 FILLER_65_3131 ();
 sg13g2_decap_8 FILLER_65_3138 ();
 sg13g2_decap_8 FILLER_65_3145 ();
 sg13g2_decap_8 FILLER_65_3152 ();
 sg13g2_decap_8 FILLER_65_3159 ();
 sg13g2_decap_8 FILLER_65_3166 ();
 sg13g2_decap_8 FILLER_65_3173 ();
 sg13g2_decap_8 FILLER_65_3180 ();
 sg13g2_decap_8 FILLER_65_3187 ();
 sg13g2_decap_8 FILLER_65_3194 ();
 sg13g2_decap_8 FILLER_65_3201 ();
 sg13g2_decap_8 FILLER_65_3208 ();
 sg13g2_decap_8 FILLER_65_3215 ();
 sg13g2_decap_8 FILLER_65_3222 ();
 sg13g2_decap_8 FILLER_65_3229 ();
 sg13g2_decap_8 FILLER_65_3236 ();
 sg13g2_decap_8 FILLER_65_3243 ();
 sg13g2_decap_8 FILLER_65_3250 ();
 sg13g2_decap_8 FILLER_65_3257 ();
 sg13g2_decap_8 FILLER_65_3264 ();
 sg13g2_decap_8 FILLER_65_3271 ();
 sg13g2_decap_8 FILLER_65_3278 ();
 sg13g2_decap_8 FILLER_65_3285 ();
 sg13g2_decap_8 FILLER_65_3292 ();
 sg13g2_decap_8 FILLER_65_3299 ();
 sg13g2_decap_8 FILLER_65_3306 ();
 sg13g2_decap_8 FILLER_65_3313 ();
 sg13g2_decap_8 FILLER_65_3320 ();
 sg13g2_decap_8 FILLER_65_3327 ();
 sg13g2_decap_8 FILLER_65_3334 ();
 sg13g2_decap_8 FILLER_65_3341 ();
 sg13g2_decap_8 FILLER_65_3348 ();
 sg13g2_decap_8 FILLER_65_3355 ();
 sg13g2_decap_8 FILLER_65_3362 ();
 sg13g2_decap_8 FILLER_65_3369 ();
 sg13g2_decap_8 FILLER_65_3376 ();
 sg13g2_decap_8 FILLER_65_3383 ();
 sg13g2_decap_8 FILLER_65_3390 ();
 sg13g2_decap_8 FILLER_65_3397 ();
 sg13g2_decap_8 FILLER_65_3404 ();
 sg13g2_decap_8 FILLER_65_3411 ();
 sg13g2_decap_8 FILLER_65_3418 ();
 sg13g2_decap_8 FILLER_65_3425 ();
 sg13g2_decap_8 FILLER_65_3432 ();
 sg13g2_decap_8 FILLER_65_3439 ();
 sg13g2_decap_8 FILLER_65_3446 ();
 sg13g2_decap_8 FILLER_65_3453 ();
 sg13g2_decap_8 FILLER_65_3460 ();
 sg13g2_decap_8 FILLER_65_3467 ();
 sg13g2_decap_8 FILLER_65_3474 ();
 sg13g2_decap_8 FILLER_65_3481 ();
 sg13g2_decap_8 FILLER_65_3488 ();
 sg13g2_decap_8 FILLER_65_3495 ();
 sg13g2_decap_8 FILLER_65_3502 ();
 sg13g2_decap_8 FILLER_65_3509 ();
 sg13g2_decap_8 FILLER_65_3516 ();
 sg13g2_decap_8 FILLER_65_3523 ();
 sg13g2_decap_8 FILLER_65_3530 ();
 sg13g2_decap_8 FILLER_65_3537 ();
 sg13g2_decap_8 FILLER_65_3544 ();
 sg13g2_decap_8 FILLER_65_3551 ();
 sg13g2_decap_8 FILLER_65_3558 ();
 sg13g2_decap_8 FILLER_65_3565 ();
 sg13g2_decap_8 FILLER_65_3572 ();
 sg13g2_fill_1 FILLER_65_3579 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_189 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_231 ();
 sg13g2_decap_8 FILLER_66_238 ();
 sg13g2_decap_8 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_252 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_decap_8 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_8 FILLER_66_280 ();
 sg13g2_decap_8 FILLER_66_287 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_decap_8 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_308 ();
 sg13g2_decap_8 FILLER_66_315 ();
 sg13g2_decap_8 FILLER_66_322 ();
 sg13g2_decap_8 FILLER_66_329 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_decap_8 FILLER_66_343 ();
 sg13g2_decap_8 FILLER_66_350 ();
 sg13g2_decap_8 FILLER_66_357 ();
 sg13g2_decap_8 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_decap_8 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_decap_8 FILLER_66_406 ();
 sg13g2_decap_8 FILLER_66_413 ();
 sg13g2_decap_8 FILLER_66_420 ();
 sg13g2_decap_4 FILLER_66_427 ();
 sg13g2_fill_2 FILLER_66_431 ();
 sg13g2_decap_4 FILLER_66_480 ();
 sg13g2_fill_2 FILLER_66_484 ();
 sg13g2_decap_8 FILLER_66_576 ();
 sg13g2_decap_8 FILLER_66_583 ();
 sg13g2_decap_4 FILLER_66_590 ();
 sg13g2_fill_2 FILLER_66_594 ();
 sg13g2_fill_2 FILLER_66_621 ();
 sg13g2_fill_1 FILLER_66_623 ();
 sg13g2_decap_8 FILLER_66_650 ();
 sg13g2_decap_8 FILLER_66_657 ();
 sg13g2_fill_1 FILLER_66_664 ();
 sg13g2_fill_1 FILLER_66_767 ();
 sg13g2_fill_2 FILLER_66_776 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_4 FILLER_66_807 ();
 sg13g2_fill_1 FILLER_66_811 ();
 sg13g2_decap_8 FILLER_66_832 ();
 sg13g2_fill_2 FILLER_66_839 ();
 sg13g2_fill_1 FILLER_66_845 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_decap_8 FILLER_66_857 ();
 sg13g2_fill_2 FILLER_66_864 ();
 sg13g2_fill_1 FILLER_66_869 ();
 sg13g2_decap_8 FILLER_66_926 ();
 sg13g2_fill_2 FILLER_66_933 ();
 sg13g2_fill_2 FILLER_66_991 ();
 sg13g2_fill_1 FILLER_66_993 ();
 sg13g2_decap_8 FILLER_66_1007 ();
 sg13g2_decap_8 FILLER_66_1044 ();
 sg13g2_decap_8 FILLER_66_1051 ();
 sg13g2_fill_1 FILLER_66_1058 ();
 sg13g2_decap_8 FILLER_66_1090 ();
 sg13g2_decap_8 FILLER_66_1097 ();
 sg13g2_decap_8 FILLER_66_1104 ();
 sg13g2_fill_2 FILLER_66_1111 ();
 sg13g2_fill_1 FILLER_66_1113 ();
 sg13g2_decap_4 FILLER_66_1140 ();
 sg13g2_decap_8 FILLER_66_1170 ();
 sg13g2_decap_8 FILLER_66_1177 ();
 sg13g2_decap_4 FILLER_66_1184 ();
 sg13g2_decap_8 FILLER_66_1193 ();
 sg13g2_decap_8 FILLER_66_1200 ();
 sg13g2_decap_4 FILLER_66_1207 ();
 sg13g2_fill_1 FILLER_66_1211 ();
 sg13g2_decap_8 FILLER_66_1218 ();
 sg13g2_fill_2 FILLER_66_1225 ();
 sg13g2_fill_2 FILLER_66_1276 ();
 sg13g2_decap_8 FILLER_66_1318 ();
 sg13g2_decap_8 FILLER_66_1325 ();
 sg13g2_decap_8 FILLER_66_1332 ();
 sg13g2_fill_1 FILLER_66_1339 ();
 sg13g2_decap_8 FILLER_66_1372 ();
 sg13g2_decap_4 FILLER_66_1379 ();
 sg13g2_decap_8 FILLER_66_1391 ();
 sg13g2_decap_8 FILLER_66_1398 ();
 sg13g2_decap_8 FILLER_66_1405 ();
 sg13g2_decap_8 FILLER_66_1412 ();
 sg13g2_decap_8 FILLER_66_1419 ();
 sg13g2_decap_4 FILLER_66_1426 ();
 sg13g2_decap_8 FILLER_66_1461 ();
 sg13g2_decap_8 FILLER_66_1468 ();
 sg13g2_decap_4 FILLER_66_1475 ();
 sg13g2_fill_2 FILLER_66_1479 ();
 sg13g2_decap_8 FILLER_66_1525 ();
 sg13g2_decap_8 FILLER_66_1532 ();
 sg13g2_decap_8 FILLER_66_1539 ();
 sg13g2_decap_8 FILLER_66_1546 ();
 sg13g2_fill_1 FILLER_66_1553 ();
 sg13g2_fill_1 FILLER_66_1559 ();
 sg13g2_decap_8 FILLER_66_1592 ();
 sg13g2_decap_8 FILLER_66_1599 ();
 sg13g2_decap_8 FILLER_66_1606 ();
 sg13g2_decap_4 FILLER_66_1613 ();
 sg13g2_fill_2 FILLER_66_1617 ();
 sg13g2_fill_2 FILLER_66_1648 ();
 sg13g2_decap_8 FILLER_66_1733 ();
 sg13g2_fill_2 FILLER_66_1740 ();
 sg13g2_decap_8 FILLER_66_1805 ();
 sg13g2_decap_8 FILLER_66_1812 ();
 sg13g2_fill_2 FILLER_66_1819 ();
 sg13g2_decap_4 FILLER_66_1899 ();
 sg13g2_decap_8 FILLER_66_1961 ();
 sg13g2_decap_8 FILLER_66_1968 ();
 sg13g2_decap_4 FILLER_66_1975 ();
 sg13g2_decap_4 FILLER_66_2013 ();
 sg13g2_fill_1 FILLER_66_2017 ();
 sg13g2_decap_8 FILLER_66_2049 ();
 sg13g2_fill_2 FILLER_66_2056 ();
 sg13g2_fill_1 FILLER_66_2058 ();
 sg13g2_fill_2 FILLER_66_2111 ();
 sg13g2_fill_1 FILLER_66_2121 ();
 sg13g2_decap_4 FILLER_66_2136 ();
 sg13g2_decap_8 FILLER_66_2145 ();
 sg13g2_fill_1 FILLER_66_2152 ();
 sg13g2_decap_8 FILLER_66_2213 ();
 sg13g2_decap_8 FILLER_66_2220 ();
 sg13g2_decap_8 FILLER_66_2227 ();
 sg13g2_decap_8 FILLER_66_2234 ();
 sg13g2_decap_8 FILLER_66_2241 ();
 sg13g2_decap_8 FILLER_66_2248 ();
 sg13g2_decap_8 FILLER_66_2255 ();
 sg13g2_decap_8 FILLER_66_2262 ();
 sg13g2_decap_8 FILLER_66_2269 ();
 sg13g2_decap_8 FILLER_66_2276 ();
 sg13g2_decap_8 FILLER_66_2283 ();
 sg13g2_decap_8 FILLER_66_2290 ();
 sg13g2_decap_8 FILLER_66_2297 ();
 sg13g2_decap_8 FILLER_66_2304 ();
 sg13g2_decap_8 FILLER_66_2311 ();
 sg13g2_decap_8 FILLER_66_2318 ();
 sg13g2_decap_8 FILLER_66_2325 ();
 sg13g2_decap_8 FILLER_66_2332 ();
 sg13g2_decap_8 FILLER_66_2339 ();
 sg13g2_decap_8 FILLER_66_2346 ();
 sg13g2_decap_8 FILLER_66_2353 ();
 sg13g2_decap_8 FILLER_66_2360 ();
 sg13g2_decap_8 FILLER_66_2367 ();
 sg13g2_decap_8 FILLER_66_2374 ();
 sg13g2_decap_8 FILLER_66_2381 ();
 sg13g2_decap_8 FILLER_66_2388 ();
 sg13g2_decap_8 FILLER_66_2395 ();
 sg13g2_decap_8 FILLER_66_2402 ();
 sg13g2_decap_8 FILLER_66_2409 ();
 sg13g2_decap_8 FILLER_66_2416 ();
 sg13g2_decap_8 FILLER_66_2423 ();
 sg13g2_decap_8 FILLER_66_2430 ();
 sg13g2_decap_8 FILLER_66_2437 ();
 sg13g2_decap_8 FILLER_66_2444 ();
 sg13g2_decap_8 FILLER_66_2451 ();
 sg13g2_decap_8 FILLER_66_2458 ();
 sg13g2_decap_8 FILLER_66_2465 ();
 sg13g2_decap_8 FILLER_66_2472 ();
 sg13g2_decap_8 FILLER_66_2479 ();
 sg13g2_decap_8 FILLER_66_2486 ();
 sg13g2_decap_8 FILLER_66_2493 ();
 sg13g2_decap_8 FILLER_66_2500 ();
 sg13g2_decap_8 FILLER_66_2507 ();
 sg13g2_decap_8 FILLER_66_2514 ();
 sg13g2_decap_8 FILLER_66_2521 ();
 sg13g2_decap_8 FILLER_66_2528 ();
 sg13g2_decap_8 FILLER_66_2535 ();
 sg13g2_decap_8 FILLER_66_2542 ();
 sg13g2_decap_8 FILLER_66_2549 ();
 sg13g2_decap_8 FILLER_66_2556 ();
 sg13g2_decap_8 FILLER_66_2563 ();
 sg13g2_decap_8 FILLER_66_2570 ();
 sg13g2_decap_8 FILLER_66_2577 ();
 sg13g2_decap_8 FILLER_66_2584 ();
 sg13g2_decap_8 FILLER_66_2591 ();
 sg13g2_decap_8 FILLER_66_2598 ();
 sg13g2_decap_8 FILLER_66_2605 ();
 sg13g2_decap_8 FILLER_66_2612 ();
 sg13g2_decap_8 FILLER_66_2619 ();
 sg13g2_decap_8 FILLER_66_2626 ();
 sg13g2_decap_8 FILLER_66_2633 ();
 sg13g2_decap_8 FILLER_66_2640 ();
 sg13g2_decap_8 FILLER_66_2647 ();
 sg13g2_decap_8 FILLER_66_2654 ();
 sg13g2_decap_8 FILLER_66_2661 ();
 sg13g2_decap_8 FILLER_66_2668 ();
 sg13g2_decap_8 FILLER_66_2675 ();
 sg13g2_decap_8 FILLER_66_2682 ();
 sg13g2_decap_8 FILLER_66_2689 ();
 sg13g2_decap_8 FILLER_66_2696 ();
 sg13g2_decap_8 FILLER_66_2703 ();
 sg13g2_decap_8 FILLER_66_2710 ();
 sg13g2_decap_8 FILLER_66_2717 ();
 sg13g2_decap_8 FILLER_66_2724 ();
 sg13g2_decap_8 FILLER_66_2731 ();
 sg13g2_decap_8 FILLER_66_2738 ();
 sg13g2_decap_8 FILLER_66_2745 ();
 sg13g2_decap_8 FILLER_66_2752 ();
 sg13g2_decap_8 FILLER_66_2759 ();
 sg13g2_decap_8 FILLER_66_2766 ();
 sg13g2_decap_8 FILLER_66_2773 ();
 sg13g2_decap_8 FILLER_66_2780 ();
 sg13g2_decap_8 FILLER_66_2787 ();
 sg13g2_decap_8 FILLER_66_2794 ();
 sg13g2_decap_8 FILLER_66_2801 ();
 sg13g2_decap_8 FILLER_66_2808 ();
 sg13g2_decap_8 FILLER_66_2815 ();
 sg13g2_decap_8 FILLER_66_2822 ();
 sg13g2_decap_8 FILLER_66_2829 ();
 sg13g2_decap_8 FILLER_66_2836 ();
 sg13g2_decap_8 FILLER_66_2843 ();
 sg13g2_decap_8 FILLER_66_2850 ();
 sg13g2_decap_8 FILLER_66_2857 ();
 sg13g2_decap_8 FILLER_66_2864 ();
 sg13g2_decap_8 FILLER_66_2871 ();
 sg13g2_decap_8 FILLER_66_2878 ();
 sg13g2_decap_8 FILLER_66_2885 ();
 sg13g2_decap_8 FILLER_66_2892 ();
 sg13g2_decap_8 FILLER_66_2899 ();
 sg13g2_decap_8 FILLER_66_2906 ();
 sg13g2_decap_8 FILLER_66_2913 ();
 sg13g2_decap_8 FILLER_66_2920 ();
 sg13g2_decap_8 FILLER_66_2927 ();
 sg13g2_decap_8 FILLER_66_2934 ();
 sg13g2_decap_8 FILLER_66_2941 ();
 sg13g2_decap_8 FILLER_66_2948 ();
 sg13g2_decap_8 FILLER_66_2955 ();
 sg13g2_decap_8 FILLER_66_2962 ();
 sg13g2_decap_8 FILLER_66_2969 ();
 sg13g2_decap_8 FILLER_66_2976 ();
 sg13g2_decap_8 FILLER_66_2983 ();
 sg13g2_decap_8 FILLER_66_2990 ();
 sg13g2_decap_8 FILLER_66_2997 ();
 sg13g2_decap_8 FILLER_66_3004 ();
 sg13g2_decap_8 FILLER_66_3011 ();
 sg13g2_decap_8 FILLER_66_3018 ();
 sg13g2_decap_8 FILLER_66_3025 ();
 sg13g2_decap_8 FILLER_66_3032 ();
 sg13g2_decap_8 FILLER_66_3039 ();
 sg13g2_decap_8 FILLER_66_3046 ();
 sg13g2_decap_8 FILLER_66_3053 ();
 sg13g2_decap_8 FILLER_66_3060 ();
 sg13g2_decap_8 FILLER_66_3067 ();
 sg13g2_decap_8 FILLER_66_3074 ();
 sg13g2_decap_8 FILLER_66_3081 ();
 sg13g2_decap_8 FILLER_66_3088 ();
 sg13g2_decap_8 FILLER_66_3095 ();
 sg13g2_decap_8 FILLER_66_3102 ();
 sg13g2_decap_8 FILLER_66_3109 ();
 sg13g2_decap_8 FILLER_66_3116 ();
 sg13g2_decap_8 FILLER_66_3123 ();
 sg13g2_decap_8 FILLER_66_3130 ();
 sg13g2_decap_8 FILLER_66_3137 ();
 sg13g2_decap_8 FILLER_66_3144 ();
 sg13g2_decap_8 FILLER_66_3151 ();
 sg13g2_decap_8 FILLER_66_3158 ();
 sg13g2_decap_8 FILLER_66_3165 ();
 sg13g2_decap_8 FILLER_66_3172 ();
 sg13g2_decap_8 FILLER_66_3179 ();
 sg13g2_decap_8 FILLER_66_3186 ();
 sg13g2_decap_8 FILLER_66_3193 ();
 sg13g2_decap_8 FILLER_66_3200 ();
 sg13g2_decap_8 FILLER_66_3207 ();
 sg13g2_decap_8 FILLER_66_3214 ();
 sg13g2_decap_8 FILLER_66_3221 ();
 sg13g2_decap_8 FILLER_66_3228 ();
 sg13g2_decap_8 FILLER_66_3235 ();
 sg13g2_decap_8 FILLER_66_3242 ();
 sg13g2_decap_8 FILLER_66_3249 ();
 sg13g2_decap_8 FILLER_66_3256 ();
 sg13g2_decap_8 FILLER_66_3263 ();
 sg13g2_decap_8 FILLER_66_3270 ();
 sg13g2_decap_8 FILLER_66_3277 ();
 sg13g2_decap_8 FILLER_66_3284 ();
 sg13g2_decap_8 FILLER_66_3291 ();
 sg13g2_decap_8 FILLER_66_3298 ();
 sg13g2_decap_8 FILLER_66_3305 ();
 sg13g2_decap_8 FILLER_66_3312 ();
 sg13g2_decap_8 FILLER_66_3319 ();
 sg13g2_decap_8 FILLER_66_3326 ();
 sg13g2_decap_8 FILLER_66_3333 ();
 sg13g2_decap_8 FILLER_66_3340 ();
 sg13g2_decap_8 FILLER_66_3347 ();
 sg13g2_decap_8 FILLER_66_3354 ();
 sg13g2_decap_8 FILLER_66_3361 ();
 sg13g2_decap_8 FILLER_66_3368 ();
 sg13g2_decap_8 FILLER_66_3375 ();
 sg13g2_decap_8 FILLER_66_3382 ();
 sg13g2_decap_8 FILLER_66_3389 ();
 sg13g2_decap_8 FILLER_66_3396 ();
 sg13g2_decap_8 FILLER_66_3403 ();
 sg13g2_decap_8 FILLER_66_3410 ();
 sg13g2_decap_8 FILLER_66_3417 ();
 sg13g2_decap_8 FILLER_66_3424 ();
 sg13g2_decap_8 FILLER_66_3431 ();
 sg13g2_decap_8 FILLER_66_3438 ();
 sg13g2_decap_8 FILLER_66_3445 ();
 sg13g2_decap_8 FILLER_66_3452 ();
 sg13g2_decap_8 FILLER_66_3459 ();
 sg13g2_decap_8 FILLER_66_3466 ();
 sg13g2_decap_8 FILLER_66_3473 ();
 sg13g2_decap_8 FILLER_66_3480 ();
 sg13g2_decap_8 FILLER_66_3487 ();
 sg13g2_decap_8 FILLER_66_3494 ();
 sg13g2_decap_8 FILLER_66_3501 ();
 sg13g2_decap_8 FILLER_66_3508 ();
 sg13g2_decap_8 FILLER_66_3515 ();
 sg13g2_decap_8 FILLER_66_3522 ();
 sg13g2_decap_8 FILLER_66_3529 ();
 sg13g2_decap_8 FILLER_66_3536 ();
 sg13g2_decap_8 FILLER_66_3543 ();
 sg13g2_decap_8 FILLER_66_3550 ();
 sg13g2_decap_8 FILLER_66_3557 ();
 sg13g2_decap_8 FILLER_66_3564 ();
 sg13g2_decap_8 FILLER_66_3571 ();
 sg13g2_fill_2 FILLER_66_3578 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_266 ();
 sg13g2_decap_8 FILLER_67_273 ();
 sg13g2_decap_8 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_287 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_decap_8 FILLER_67_301 ();
 sg13g2_decap_8 FILLER_67_308 ();
 sg13g2_decap_8 FILLER_67_315 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_329 ();
 sg13g2_decap_8 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_67_350 ();
 sg13g2_decap_8 FILLER_67_357 ();
 sg13g2_decap_8 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_decap_8 FILLER_67_406 ();
 sg13g2_decap_8 FILLER_67_413 ();
 sg13g2_decap_8 FILLER_67_420 ();
 sg13g2_decap_8 FILLER_67_427 ();
 sg13g2_decap_8 FILLER_67_434 ();
 sg13g2_decap_4 FILLER_67_441 ();
 sg13g2_decap_4 FILLER_67_487 ();
 sg13g2_fill_1 FILLER_67_491 ();
 sg13g2_fill_2 FILLER_67_507 ();
 sg13g2_decap_8 FILLER_67_577 ();
 sg13g2_decap_8 FILLER_67_584 ();
 sg13g2_decap_8 FILLER_67_591 ();
 sg13g2_decap_8 FILLER_67_598 ();
 sg13g2_fill_2 FILLER_67_605 ();
 sg13g2_fill_2 FILLER_67_624 ();
 sg13g2_decap_4 FILLER_67_629 ();
 sg13g2_fill_1 FILLER_67_693 ();
 sg13g2_decap_8 FILLER_67_702 ();
 sg13g2_decap_8 FILLER_67_709 ();
 sg13g2_decap_8 FILLER_67_746 ();
 sg13g2_fill_1 FILLER_67_753 ();
 sg13g2_decap_4 FILLER_67_758 ();
 sg13g2_fill_1 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_832 ();
 sg13g2_decap_8 FILLER_67_839 ();
 sg13g2_decap_8 FILLER_67_846 ();
 sg13g2_fill_1 FILLER_67_858 ();
 sg13g2_fill_1 FILLER_67_864 ();
 sg13g2_decap_8 FILLER_67_873 ();
 sg13g2_decap_8 FILLER_67_880 ();
 sg13g2_decap_4 FILLER_67_891 ();
 sg13g2_fill_2 FILLER_67_895 ();
 sg13g2_decap_8 FILLER_67_901 ();
 sg13g2_decap_4 FILLER_67_908 ();
 sg13g2_fill_1 FILLER_67_912 ();
 sg13g2_decap_8 FILLER_67_921 ();
 sg13g2_decap_8 FILLER_67_928 ();
 sg13g2_decap_8 FILLER_67_935 ();
 sg13g2_decap_8 FILLER_67_942 ();
 sg13g2_decap_4 FILLER_67_949 ();
 sg13g2_fill_1 FILLER_67_953 ();
 sg13g2_decap_8 FILLER_67_958 ();
 sg13g2_decap_8 FILLER_67_965 ();
 sg13g2_decap_4 FILLER_67_972 ();
 sg13g2_fill_2 FILLER_67_980 ();
 sg13g2_fill_1 FILLER_67_982 ();
 sg13g2_fill_1 FILLER_67_988 ();
 sg13g2_fill_1 FILLER_67_994 ();
 sg13g2_fill_1 FILLER_67_1005 ();
 sg13g2_decap_4 FILLER_67_1014 ();
 sg13g2_fill_1 FILLER_67_1018 ();
 sg13g2_fill_1 FILLER_67_1024 ();
 sg13g2_decap_8 FILLER_67_1091 ();
 sg13g2_decap_4 FILLER_67_1098 ();
 sg13g2_fill_1 FILLER_67_1102 ();
 sg13g2_decap_8 FILLER_67_1129 ();
 sg13g2_decap_8 FILLER_67_1136 ();
 sg13g2_fill_2 FILLER_67_1143 ();
 sg13g2_decap_8 FILLER_67_1171 ();
 sg13g2_decap_8 FILLER_67_1178 ();
 sg13g2_decap_8 FILLER_67_1185 ();
 sg13g2_decap_4 FILLER_67_1192 ();
 sg13g2_fill_1 FILLER_67_1196 ();
 sg13g2_decap_4 FILLER_67_1223 ();
 sg13g2_decap_8 FILLER_67_1259 ();
 sg13g2_decap_8 FILLER_67_1266 ();
 sg13g2_decap_4 FILLER_67_1273 ();
 sg13g2_fill_1 FILLER_67_1277 ();
 sg13g2_decap_8 FILLER_67_1317 ();
 sg13g2_decap_8 FILLER_67_1324 ();
 sg13g2_decap_4 FILLER_67_1331 ();
 sg13g2_fill_1 FILLER_67_1335 ();
 sg13g2_decap_8 FILLER_67_1362 ();
 sg13g2_decap_4 FILLER_67_1369 ();
 sg13g2_fill_1 FILLER_67_1373 ();
 sg13g2_fill_2 FILLER_67_1379 ();
 sg13g2_fill_1 FILLER_67_1381 ();
 sg13g2_decap_8 FILLER_67_1408 ();
 sg13g2_decap_8 FILLER_67_1415 ();
 sg13g2_fill_2 FILLER_67_1422 ();
 sg13g2_fill_1 FILLER_67_1424 ();
 sg13g2_decap_8 FILLER_67_1456 ();
 sg13g2_decap_8 FILLER_67_1463 ();
 sg13g2_decap_8 FILLER_67_1470 ();
 sg13g2_decap_8 FILLER_67_1477 ();
 sg13g2_fill_2 FILLER_67_1484 ();
 sg13g2_fill_1 FILLER_67_1486 ();
 sg13g2_fill_2 FILLER_67_1517 ();
 sg13g2_fill_1 FILLER_67_1519 ();
 sg13g2_decap_8 FILLER_67_1598 ();
 sg13g2_decap_8 FILLER_67_1605 ();
 sg13g2_decap_8 FILLER_67_1612 ();
 sg13g2_decap_4 FILLER_67_1619 ();
 sg13g2_decap_8 FILLER_67_1649 ();
 sg13g2_decap_8 FILLER_67_1656 ();
 sg13g2_decap_8 FILLER_67_1663 ();
 sg13g2_fill_1 FILLER_67_1670 ();
 sg13g2_fill_2 FILLER_67_1697 ();
 sg13g2_fill_1 FILLER_67_1699 ();
 sg13g2_decap_8 FILLER_67_1726 ();
 sg13g2_decap_4 FILLER_67_1733 ();
 sg13g2_fill_2 FILLER_67_1737 ();
 sg13g2_decap_8 FILLER_67_1806 ();
 sg13g2_decap_8 FILLER_67_1813 ();
 sg13g2_decap_8 FILLER_67_1820 ();
 sg13g2_fill_2 FILLER_67_1827 ();
 sg13g2_decap_8 FILLER_67_1881 ();
 sg13g2_decap_8 FILLER_67_1888 ();
 sg13g2_decap_8 FILLER_67_1895 ();
 sg13g2_decap_4 FILLER_67_1902 ();
 sg13g2_fill_2 FILLER_67_1906 ();
 sg13g2_fill_2 FILLER_67_1934 ();
 sg13g2_fill_1 FILLER_67_1936 ();
 sg13g2_decap_8 FILLER_67_1950 ();
 sg13g2_decap_8 FILLER_67_1957 ();
 sg13g2_decap_4 FILLER_67_1964 ();
 sg13g2_fill_1 FILLER_67_1968 ();
 sg13g2_decap_4 FILLER_67_2073 ();
 sg13g2_fill_2 FILLER_67_2077 ();
 sg13g2_decap_4 FILLER_67_2110 ();
 sg13g2_decap_8 FILLER_67_2147 ();
 sg13g2_decap_8 FILLER_67_2154 ();
 sg13g2_fill_1 FILLER_67_2161 ();
 sg13g2_decap_8 FILLER_67_2214 ();
 sg13g2_decap_8 FILLER_67_2221 ();
 sg13g2_decap_8 FILLER_67_2228 ();
 sg13g2_decap_8 FILLER_67_2235 ();
 sg13g2_decap_8 FILLER_67_2242 ();
 sg13g2_decap_8 FILLER_67_2249 ();
 sg13g2_decap_8 FILLER_67_2256 ();
 sg13g2_decap_8 FILLER_67_2263 ();
 sg13g2_decap_8 FILLER_67_2270 ();
 sg13g2_decap_8 FILLER_67_2277 ();
 sg13g2_decap_8 FILLER_67_2284 ();
 sg13g2_decap_8 FILLER_67_2291 ();
 sg13g2_decap_8 FILLER_67_2298 ();
 sg13g2_decap_8 FILLER_67_2305 ();
 sg13g2_decap_8 FILLER_67_2312 ();
 sg13g2_decap_8 FILLER_67_2319 ();
 sg13g2_decap_8 FILLER_67_2326 ();
 sg13g2_decap_8 FILLER_67_2333 ();
 sg13g2_decap_8 FILLER_67_2340 ();
 sg13g2_decap_8 FILLER_67_2347 ();
 sg13g2_decap_8 FILLER_67_2354 ();
 sg13g2_decap_8 FILLER_67_2361 ();
 sg13g2_decap_8 FILLER_67_2368 ();
 sg13g2_decap_8 FILLER_67_2375 ();
 sg13g2_decap_8 FILLER_67_2382 ();
 sg13g2_decap_8 FILLER_67_2389 ();
 sg13g2_decap_8 FILLER_67_2396 ();
 sg13g2_decap_8 FILLER_67_2403 ();
 sg13g2_decap_8 FILLER_67_2410 ();
 sg13g2_decap_8 FILLER_67_2417 ();
 sg13g2_decap_8 FILLER_67_2424 ();
 sg13g2_decap_8 FILLER_67_2431 ();
 sg13g2_decap_8 FILLER_67_2438 ();
 sg13g2_decap_8 FILLER_67_2445 ();
 sg13g2_decap_8 FILLER_67_2452 ();
 sg13g2_decap_8 FILLER_67_2459 ();
 sg13g2_decap_8 FILLER_67_2466 ();
 sg13g2_decap_8 FILLER_67_2473 ();
 sg13g2_decap_8 FILLER_67_2480 ();
 sg13g2_decap_8 FILLER_67_2487 ();
 sg13g2_decap_8 FILLER_67_2494 ();
 sg13g2_decap_8 FILLER_67_2501 ();
 sg13g2_decap_8 FILLER_67_2508 ();
 sg13g2_decap_8 FILLER_67_2515 ();
 sg13g2_decap_8 FILLER_67_2522 ();
 sg13g2_decap_8 FILLER_67_2529 ();
 sg13g2_decap_8 FILLER_67_2536 ();
 sg13g2_decap_8 FILLER_67_2543 ();
 sg13g2_decap_8 FILLER_67_2550 ();
 sg13g2_decap_8 FILLER_67_2557 ();
 sg13g2_decap_8 FILLER_67_2564 ();
 sg13g2_decap_8 FILLER_67_2571 ();
 sg13g2_decap_8 FILLER_67_2578 ();
 sg13g2_decap_8 FILLER_67_2585 ();
 sg13g2_decap_8 FILLER_67_2592 ();
 sg13g2_decap_8 FILLER_67_2599 ();
 sg13g2_decap_8 FILLER_67_2606 ();
 sg13g2_decap_8 FILLER_67_2613 ();
 sg13g2_decap_8 FILLER_67_2620 ();
 sg13g2_decap_8 FILLER_67_2627 ();
 sg13g2_decap_8 FILLER_67_2634 ();
 sg13g2_decap_8 FILLER_67_2641 ();
 sg13g2_decap_8 FILLER_67_2648 ();
 sg13g2_decap_8 FILLER_67_2655 ();
 sg13g2_decap_8 FILLER_67_2662 ();
 sg13g2_decap_8 FILLER_67_2669 ();
 sg13g2_decap_8 FILLER_67_2676 ();
 sg13g2_decap_8 FILLER_67_2683 ();
 sg13g2_decap_8 FILLER_67_2690 ();
 sg13g2_decap_8 FILLER_67_2697 ();
 sg13g2_decap_8 FILLER_67_2704 ();
 sg13g2_decap_8 FILLER_67_2711 ();
 sg13g2_decap_8 FILLER_67_2718 ();
 sg13g2_decap_8 FILLER_67_2725 ();
 sg13g2_decap_8 FILLER_67_2732 ();
 sg13g2_decap_8 FILLER_67_2739 ();
 sg13g2_decap_8 FILLER_67_2746 ();
 sg13g2_decap_8 FILLER_67_2753 ();
 sg13g2_decap_8 FILLER_67_2760 ();
 sg13g2_decap_8 FILLER_67_2767 ();
 sg13g2_decap_8 FILLER_67_2774 ();
 sg13g2_decap_8 FILLER_67_2781 ();
 sg13g2_decap_8 FILLER_67_2788 ();
 sg13g2_decap_8 FILLER_67_2795 ();
 sg13g2_decap_8 FILLER_67_2802 ();
 sg13g2_decap_8 FILLER_67_2809 ();
 sg13g2_decap_8 FILLER_67_2816 ();
 sg13g2_decap_8 FILLER_67_2823 ();
 sg13g2_decap_8 FILLER_67_2830 ();
 sg13g2_decap_8 FILLER_67_2837 ();
 sg13g2_decap_8 FILLER_67_2844 ();
 sg13g2_decap_8 FILLER_67_2851 ();
 sg13g2_decap_8 FILLER_67_2858 ();
 sg13g2_decap_8 FILLER_67_2865 ();
 sg13g2_decap_8 FILLER_67_2872 ();
 sg13g2_decap_8 FILLER_67_2879 ();
 sg13g2_decap_8 FILLER_67_2886 ();
 sg13g2_decap_8 FILLER_67_2893 ();
 sg13g2_decap_8 FILLER_67_2900 ();
 sg13g2_decap_8 FILLER_67_2907 ();
 sg13g2_decap_8 FILLER_67_2914 ();
 sg13g2_decap_8 FILLER_67_2921 ();
 sg13g2_decap_8 FILLER_67_2928 ();
 sg13g2_decap_8 FILLER_67_2935 ();
 sg13g2_decap_8 FILLER_67_2942 ();
 sg13g2_decap_8 FILLER_67_2949 ();
 sg13g2_decap_8 FILLER_67_2956 ();
 sg13g2_decap_8 FILLER_67_2963 ();
 sg13g2_decap_8 FILLER_67_2970 ();
 sg13g2_decap_8 FILLER_67_2977 ();
 sg13g2_decap_8 FILLER_67_2984 ();
 sg13g2_decap_8 FILLER_67_2991 ();
 sg13g2_decap_8 FILLER_67_2998 ();
 sg13g2_decap_8 FILLER_67_3005 ();
 sg13g2_decap_8 FILLER_67_3012 ();
 sg13g2_decap_8 FILLER_67_3019 ();
 sg13g2_decap_8 FILLER_67_3026 ();
 sg13g2_decap_8 FILLER_67_3033 ();
 sg13g2_decap_8 FILLER_67_3040 ();
 sg13g2_decap_8 FILLER_67_3047 ();
 sg13g2_decap_8 FILLER_67_3054 ();
 sg13g2_decap_8 FILLER_67_3061 ();
 sg13g2_decap_8 FILLER_67_3068 ();
 sg13g2_decap_8 FILLER_67_3075 ();
 sg13g2_decap_8 FILLER_67_3082 ();
 sg13g2_decap_8 FILLER_67_3089 ();
 sg13g2_decap_8 FILLER_67_3096 ();
 sg13g2_decap_8 FILLER_67_3103 ();
 sg13g2_decap_8 FILLER_67_3110 ();
 sg13g2_decap_8 FILLER_67_3117 ();
 sg13g2_decap_8 FILLER_67_3124 ();
 sg13g2_decap_8 FILLER_67_3131 ();
 sg13g2_decap_8 FILLER_67_3138 ();
 sg13g2_decap_8 FILLER_67_3145 ();
 sg13g2_decap_8 FILLER_67_3152 ();
 sg13g2_decap_8 FILLER_67_3159 ();
 sg13g2_decap_8 FILLER_67_3166 ();
 sg13g2_decap_8 FILLER_67_3173 ();
 sg13g2_decap_8 FILLER_67_3180 ();
 sg13g2_decap_8 FILLER_67_3187 ();
 sg13g2_decap_8 FILLER_67_3194 ();
 sg13g2_decap_8 FILLER_67_3201 ();
 sg13g2_decap_8 FILLER_67_3208 ();
 sg13g2_decap_8 FILLER_67_3215 ();
 sg13g2_decap_8 FILLER_67_3222 ();
 sg13g2_decap_8 FILLER_67_3229 ();
 sg13g2_decap_8 FILLER_67_3236 ();
 sg13g2_decap_8 FILLER_67_3243 ();
 sg13g2_decap_8 FILLER_67_3250 ();
 sg13g2_decap_8 FILLER_67_3257 ();
 sg13g2_decap_8 FILLER_67_3264 ();
 sg13g2_decap_8 FILLER_67_3271 ();
 sg13g2_decap_8 FILLER_67_3278 ();
 sg13g2_decap_8 FILLER_67_3285 ();
 sg13g2_decap_8 FILLER_67_3292 ();
 sg13g2_decap_8 FILLER_67_3299 ();
 sg13g2_decap_8 FILLER_67_3306 ();
 sg13g2_decap_8 FILLER_67_3313 ();
 sg13g2_decap_8 FILLER_67_3320 ();
 sg13g2_decap_8 FILLER_67_3327 ();
 sg13g2_decap_8 FILLER_67_3334 ();
 sg13g2_decap_8 FILLER_67_3341 ();
 sg13g2_decap_8 FILLER_67_3348 ();
 sg13g2_decap_8 FILLER_67_3355 ();
 sg13g2_decap_8 FILLER_67_3362 ();
 sg13g2_decap_8 FILLER_67_3369 ();
 sg13g2_decap_8 FILLER_67_3376 ();
 sg13g2_decap_8 FILLER_67_3383 ();
 sg13g2_decap_8 FILLER_67_3390 ();
 sg13g2_decap_8 FILLER_67_3397 ();
 sg13g2_decap_8 FILLER_67_3404 ();
 sg13g2_decap_8 FILLER_67_3411 ();
 sg13g2_decap_8 FILLER_67_3418 ();
 sg13g2_decap_8 FILLER_67_3425 ();
 sg13g2_decap_8 FILLER_67_3432 ();
 sg13g2_decap_8 FILLER_67_3439 ();
 sg13g2_decap_8 FILLER_67_3446 ();
 sg13g2_decap_8 FILLER_67_3453 ();
 sg13g2_decap_8 FILLER_67_3460 ();
 sg13g2_decap_8 FILLER_67_3467 ();
 sg13g2_decap_8 FILLER_67_3474 ();
 sg13g2_decap_8 FILLER_67_3481 ();
 sg13g2_decap_8 FILLER_67_3488 ();
 sg13g2_decap_8 FILLER_67_3495 ();
 sg13g2_decap_8 FILLER_67_3502 ();
 sg13g2_decap_8 FILLER_67_3509 ();
 sg13g2_decap_8 FILLER_67_3516 ();
 sg13g2_decap_8 FILLER_67_3523 ();
 sg13g2_decap_8 FILLER_67_3530 ();
 sg13g2_decap_8 FILLER_67_3537 ();
 sg13g2_decap_8 FILLER_67_3544 ();
 sg13g2_decap_8 FILLER_67_3551 ();
 sg13g2_decap_8 FILLER_67_3558 ();
 sg13g2_decap_8 FILLER_67_3565 ();
 sg13g2_decap_8 FILLER_67_3572 ();
 sg13g2_fill_1 FILLER_67_3579 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_196 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_decap_8 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_231 ();
 sg13g2_decap_8 FILLER_68_238 ();
 sg13g2_decap_8 FILLER_68_245 ();
 sg13g2_decap_8 FILLER_68_252 ();
 sg13g2_decap_8 FILLER_68_259 ();
 sg13g2_decap_8 FILLER_68_266 ();
 sg13g2_decap_8 FILLER_68_273 ();
 sg13g2_decap_8 FILLER_68_280 ();
 sg13g2_decap_8 FILLER_68_287 ();
 sg13g2_decap_8 FILLER_68_294 ();
 sg13g2_decap_8 FILLER_68_301 ();
 sg13g2_decap_8 FILLER_68_308 ();
 sg13g2_decap_8 FILLER_68_315 ();
 sg13g2_decap_8 FILLER_68_322 ();
 sg13g2_decap_8 FILLER_68_329 ();
 sg13g2_decap_8 FILLER_68_336 ();
 sg13g2_decap_8 FILLER_68_343 ();
 sg13g2_decap_8 FILLER_68_350 ();
 sg13g2_decap_8 FILLER_68_357 ();
 sg13g2_decap_8 FILLER_68_364 ();
 sg13g2_decap_8 FILLER_68_371 ();
 sg13g2_decap_8 FILLER_68_378 ();
 sg13g2_decap_8 FILLER_68_385 ();
 sg13g2_decap_8 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_decap_8 FILLER_68_406 ();
 sg13g2_decap_8 FILLER_68_413 ();
 sg13g2_decap_8 FILLER_68_420 ();
 sg13g2_decap_8 FILLER_68_427 ();
 sg13g2_decap_8 FILLER_68_434 ();
 sg13g2_decap_8 FILLER_68_441 ();
 sg13g2_fill_2 FILLER_68_453 ();
 sg13g2_decap_8 FILLER_68_481 ();
 sg13g2_decap_8 FILLER_68_488 ();
 sg13g2_decap_8 FILLER_68_495 ();
 sg13g2_fill_2 FILLER_68_510 ();
 sg13g2_fill_1 FILLER_68_512 ();
 sg13g2_fill_2 FILLER_68_521 ();
 sg13g2_fill_1 FILLER_68_523 ();
 sg13g2_decap_8 FILLER_68_540 ();
 sg13g2_fill_2 FILLER_68_547 ();
 sg13g2_decap_8 FILLER_68_575 ();
 sg13g2_decap_8 FILLER_68_582 ();
 sg13g2_fill_2 FILLER_68_589 ();
 sg13g2_fill_1 FILLER_68_591 ();
 sg13g2_fill_2 FILLER_68_618 ();
 sg13g2_decap_4 FILLER_68_636 ();
 sg13g2_decap_8 FILLER_68_671 ();
 sg13g2_decap_8 FILLER_68_678 ();
 sg13g2_fill_2 FILLER_68_685 ();
 sg13g2_decap_8 FILLER_68_713 ();
 sg13g2_decap_8 FILLER_68_720 ();
 sg13g2_fill_1 FILLER_68_727 ();
 sg13g2_decap_8 FILLER_68_736 ();
 sg13g2_fill_1 FILLER_68_743 ();
 sg13g2_decap_4 FILLER_68_770 ();
 sg13g2_fill_2 FILLER_68_774 ();
 sg13g2_decap_4 FILLER_68_780 ();
 sg13g2_fill_1 FILLER_68_875 ();
 sg13g2_decap_4 FILLER_68_881 ();
 sg13g2_fill_2 FILLER_68_885 ();
 sg13g2_decap_8 FILLER_68_895 ();
 sg13g2_decap_8 FILLER_68_902 ();
 sg13g2_decap_4 FILLER_68_909 ();
 sg13g2_fill_2 FILLER_68_913 ();
 sg13g2_fill_2 FILLER_68_941 ();
 sg13g2_fill_2 FILLER_68_995 ();
 sg13g2_fill_1 FILLER_68_997 ();
 sg13g2_fill_2 FILLER_68_1008 ();
 sg13g2_fill_1 FILLER_68_1010 ();
 sg13g2_fill_1 FILLER_68_1015 ();
 sg13g2_decap_8 FILLER_68_1034 ();
 sg13g2_decap_8 FILLER_68_1041 ();
 sg13g2_decap_8 FILLER_68_1048 ();
 sg13g2_decap_4 FILLER_68_1099 ();
 sg13g2_fill_2 FILLER_68_1103 ();
 sg13g2_fill_2 FILLER_68_1108 ();
 sg13g2_fill_1 FILLER_68_1110 ();
 sg13g2_decap_8 FILLER_68_1137 ();
 sg13g2_decap_8 FILLER_68_1144 ();
 sg13g2_decap_8 FILLER_68_1151 ();
 sg13g2_decap_8 FILLER_68_1158 ();
 sg13g2_decap_8 FILLER_68_1165 ();
 sg13g2_decap_8 FILLER_68_1172 ();
 sg13g2_decap_8 FILLER_68_1179 ();
 sg13g2_decap_4 FILLER_68_1186 ();
 sg13g2_fill_2 FILLER_68_1190 ();
 sg13g2_decap_8 FILLER_68_1247 ();
 sg13g2_fill_1 FILLER_68_1254 ();
 sg13g2_decap_8 FILLER_68_1265 ();
 sg13g2_decap_8 FILLER_68_1272 ();
 sg13g2_decap_8 FILLER_68_1305 ();
 sg13g2_decap_8 FILLER_68_1312 ();
 sg13g2_decap_8 FILLER_68_1319 ();
 sg13g2_decap_4 FILLER_68_1326 ();
 sg13g2_fill_1 FILLER_68_1330 ();
 sg13g2_fill_1 FILLER_68_1357 ();
 sg13g2_decap_8 FILLER_68_1410 ();
 sg13g2_decap_8 FILLER_68_1417 ();
 sg13g2_decap_8 FILLER_68_1424 ();
 sg13g2_decap_8 FILLER_68_1486 ();
 sg13g2_decap_4 FILLER_68_1493 ();
 sg13g2_fill_1 FILLER_68_1497 ();
 sg13g2_fill_1 FILLER_68_1524 ();
 sg13g2_decap_8 FILLER_68_1551 ();
 sg13g2_decap_8 FILLER_68_1558 ();
 sg13g2_decap_4 FILLER_68_1565 ();
 sg13g2_decap_8 FILLER_68_1595 ();
 sg13g2_decap_4 FILLER_68_1602 ();
 sg13g2_fill_2 FILLER_68_1606 ();
 sg13g2_decap_8 FILLER_68_1619 ();
 sg13g2_decap_4 FILLER_68_1626 ();
 sg13g2_fill_1 FILLER_68_1630 ();
 sg13g2_decap_8 FILLER_68_1657 ();
 sg13g2_decap_8 FILLER_68_1664 ();
 sg13g2_decap_8 FILLER_68_1671 ();
 sg13g2_decap_4 FILLER_68_1678 ();
 sg13g2_decap_8 FILLER_68_1716 ();
 sg13g2_decap_8 FILLER_68_1723 ();
 sg13g2_decap_8 FILLER_68_1730 ();
 sg13g2_decap_8 FILLER_68_1737 ();
 sg13g2_decap_8 FILLER_68_1744 ();
 sg13g2_decap_4 FILLER_68_1751 ();
 sg13g2_fill_1 FILLER_68_1755 ();
 sg13g2_decap_4 FILLER_68_1761 ();
 sg13g2_fill_1 FILLER_68_1765 ();
 sg13g2_decap_8 FILLER_68_1797 ();
 sg13g2_decap_8 FILLER_68_1804 ();
 sg13g2_decap_8 FILLER_68_1811 ();
 sg13g2_decap_8 FILLER_68_1818 ();
 sg13g2_decap_8 FILLER_68_1825 ();
 sg13g2_decap_8 FILLER_68_1832 ();
 sg13g2_fill_2 FILLER_68_1839 ();
 sg13g2_fill_1 FILLER_68_1841 ();
 sg13g2_fill_1 FILLER_68_1868 ();
 sg13g2_fill_2 FILLER_68_1879 ();
 sg13g2_decap_8 FILLER_68_1886 ();
 sg13g2_decap_8 FILLER_68_1893 ();
 sg13g2_decap_8 FILLER_68_1900 ();
 sg13g2_fill_2 FILLER_68_1907 ();
 sg13g2_fill_1 FILLER_68_1909 ();
 sg13g2_fill_2 FILLER_68_1916 ();
 sg13g2_fill_1 FILLER_68_1922 ();
 sg13g2_decap_8 FILLER_68_1928 ();
 sg13g2_decap_4 FILLER_68_1935 ();
 sg13g2_fill_2 FILLER_68_1939 ();
 sg13g2_fill_1 FILLER_68_1948 ();
 sg13g2_decap_8 FILLER_68_1960 ();
 sg13g2_decap_8 FILLER_68_1967 ();
 sg13g2_decap_8 FILLER_68_1974 ();
 sg13g2_decap_4 FILLER_68_1981 ();
 sg13g2_fill_1 FILLER_68_1985 ();
 sg13g2_decap_4 FILLER_68_2025 ();
 sg13g2_decap_8 FILLER_68_2055 ();
 sg13g2_fill_1 FILLER_68_2062 ();
 sg13g2_fill_1 FILLER_68_2150 ();
 sg13g2_decap_8 FILLER_68_2156 ();
 sg13g2_decap_8 FILLER_68_2163 ();
 sg13g2_fill_1 FILLER_68_2170 ();
 sg13g2_decap_8 FILLER_68_2205 ();
 sg13g2_decap_8 FILLER_68_2212 ();
 sg13g2_decap_8 FILLER_68_2219 ();
 sg13g2_decap_8 FILLER_68_2226 ();
 sg13g2_decap_8 FILLER_68_2233 ();
 sg13g2_decap_8 FILLER_68_2240 ();
 sg13g2_decap_8 FILLER_68_2247 ();
 sg13g2_decap_8 FILLER_68_2254 ();
 sg13g2_decap_8 FILLER_68_2261 ();
 sg13g2_decap_8 FILLER_68_2268 ();
 sg13g2_decap_8 FILLER_68_2275 ();
 sg13g2_decap_8 FILLER_68_2282 ();
 sg13g2_decap_8 FILLER_68_2289 ();
 sg13g2_decap_8 FILLER_68_2296 ();
 sg13g2_decap_8 FILLER_68_2303 ();
 sg13g2_decap_8 FILLER_68_2310 ();
 sg13g2_decap_8 FILLER_68_2317 ();
 sg13g2_decap_8 FILLER_68_2324 ();
 sg13g2_decap_8 FILLER_68_2331 ();
 sg13g2_decap_8 FILLER_68_2338 ();
 sg13g2_decap_8 FILLER_68_2345 ();
 sg13g2_decap_8 FILLER_68_2352 ();
 sg13g2_decap_8 FILLER_68_2359 ();
 sg13g2_decap_8 FILLER_68_2366 ();
 sg13g2_decap_8 FILLER_68_2373 ();
 sg13g2_decap_8 FILLER_68_2380 ();
 sg13g2_decap_8 FILLER_68_2387 ();
 sg13g2_decap_8 FILLER_68_2394 ();
 sg13g2_decap_8 FILLER_68_2401 ();
 sg13g2_decap_8 FILLER_68_2408 ();
 sg13g2_decap_8 FILLER_68_2415 ();
 sg13g2_decap_8 FILLER_68_2422 ();
 sg13g2_decap_8 FILLER_68_2429 ();
 sg13g2_decap_8 FILLER_68_2436 ();
 sg13g2_decap_8 FILLER_68_2443 ();
 sg13g2_decap_8 FILLER_68_2450 ();
 sg13g2_decap_8 FILLER_68_2457 ();
 sg13g2_decap_8 FILLER_68_2464 ();
 sg13g2_decap_8 FILLER_68_2471 ();
 sg13g2_decap_8 FILLER_68_2478 ();
 sg13g2_decap_8 FILLER_68_2485 ();
 sg13g2_decap_8 FILLER_68_2492 ();
 sg13g2_decap_8 FILLER_68_2499 ();
 sg13g2_decap_8 FILLER_68_2506 ();
 sg13g2_decap_8 FILLER_68_2513 ();
 sg13g2_decap_8 FILLER_68_2520 ();
 sg13g2_decap_8 FILLER_68_2527 ();
 sg13g2_decap_8 FILLER_68_2534 ();
 sg13g2_decap_8 FILLER_68_2541 ();
 sg13g2_decap_8 FILLER_68_2548 ();
 sg13g2_decap_8 FILLER_68_2555 ();
 sg13g2_decap_8 FILLER_68_2562 ();
 sg13g2_decap_8 FILLER_68_2569 ();
 sg13g2_decap_8 FILLER_68_2576 ();
 sg13g2_decap_8 FILLER_68_2583 ();
 sg13g2_decap_8 FILLER_68_2590 ();
 sg13g2_decap_8 FILLER_68_2597 ();
 sg13g2_decap_8 FILLER_68_2604 ();
 sg13g2_decap_8 FILLER_68_2611 ();
 sg13g2_decap_8 FILLER_68_2618 ();
 sg13g2_decap_8 FILLER_68_2625 ();
 sg13g2_decap_8 FILLER_68_2632 ();
 sg13g2_decap_8 FILLER_68_2639 ();
 sg13g2_decap_8 FILLER_68_2646 ();
 sg13g2_decap_8 FILLER_68_2653 ();
 sg13g2_decap_8 FILLER_68_2660 ();
 sg13g2_decap_8 FILLER_68_2667 ();
 sg13g2_decap_8 FILLER_68_2674 ();
 sg13g2_decap_8 FILLER_68_2681 ();
 sg13g2_decap_8 FILLER_68_2688 ();
 sg13g2_decap_8 FILLER_68_2695 ();
 sg13g2_decap_8 FILLER_68_2702 ();
 sg13g2_decap_8 FILLER_68_2709 ();
 sg13g2_decap_8 FILLER_68_2716 ();
 sg13g2_decap_8 FILLER_68_2723 ();
 sg13g2_decap_8 FILLER_68_2730 ();
 sg13g2_decap_8 FILLER_68_2737 ();
 sg13g2_decap_8 FILLER_68_2744 ();
 sg13g2_decap_8 FILLER_68_2751 ();
 sg13g2_decap_8 FILLER_68_2758 ();
 sg13g2_decap_8 FILLER_68_2765 ();
 sg13g2_decap_8 FILLER_68_2772 ();
 sg13g2_decap_8 FILLER_68_2779 ();
 sg13g2_decap_8 FILLER_68_2786 ();
 sg13g2_decap_8 FILLER_68_2793 ();
 sg13g2_decap_8 FILLER_68_2800 ();
 sg13g2_decap_8 FILLER_68_2807 ();
 sg13g2_decap_8 FILLER_68_2814 ();
 sg13g2_decap_8 FILLER_68_2821 ();
 sg13g2_decap_8 FILLER_68_2828 ();
 sg13g2_decap_8 FILLER_68_2835 ();
 sg13g2_decap_8 FILLER_68_2842 ();
 sg13g2_decap_8 FILLER_68_2849 ();
 sg13g2_decap_8 FILLER_68_2856 ();
 sg13g2_decap_8 FILLER_68_2863 ();
 sg13g2_decap_8 FILLER_68_2870 ();
 sg13g2_decap_8 FILLER_68_2877 ();
 sg13g2_decap_8 FILLER_68_2884 ();
 sg13g2_decap_8 FILLER_68_2891 ();
 sg13g2_decap_8 FILLER_68_2898 ();
 sg13g2_decap_8 FILLER_68_2905 ();
 sg13g2_decap_8 FILLER_68_2912 ();
 sg13g2_decap_8 FILLER_68_2919 ();
 sg13g2_decap_8 FILLER_68_2926 ();
 sg13g2_decap_8 FILLER_68_2933 ();
 sg13g2_decap_8 FILLER_68_2940 ();
 sg13g2_decap_8 FILLER_68_2947 ();
 sg13g2_decap_8 FILLER_68_2954 ();
 sg13g2_decap_8 FILLER_68_2961 ();
 sg13g2_decap_8 FILLER_68_2968 ();
 sg13g2_decap_8 FILLER_68_2975 ();
 sg13g2_decap_8 FILLER_68_2982 ();
 sg13g2_decap_8 FILLER_68_2989 ();
 sg13g2_decap_8 FILLER_68_2996 ();
 sg13g2_decap_8 FILLER_68_3003 ();
 sg13g2_decap_8 FILLER_68_3010 ();
 sg13g2_decap_8 FILLER_68_3017 ();
 sg13g2_decap_8 FILLER_68_3024 ();
 sg13g2_decap_8 FILLER_68_3031 ();
 sg13g2_decap_8 FILLER_68_3038 ();
 sg13g2_decap_8 FILLER_68_3045 ();
 sg13g2_decap_8 FILLER_68_3052 ();
 sg13g2_decap_8 FILLER_68_3059 ();
 sg13g2_decap_8 FILLER_68_3066 ();
 sg13g2_decap_8 FILLER_68_3073 ();
 sg13g2_decap_8 FILLER_68_3080 ();
 sg13g2_decap_8 FILLER_68_3087 ();
 sg13g2_decap_8 FILLER_68_3094 ();
 sg13g2_decap_8 FILLER_68_3101 ();
 sg13g2_decap_8 FILLER_68_3108 ();
 sg13g2_decap_8 FILLER_68_3115 ();
 sg13g2_decap_8 FILLER_68_3122 ();
 sg13g2_decap_8 FILLER_68_3129 ();
 sg13g2_decap_8 FILLER_68_3136 ();
 sg13g2_decap_8 FILLER_68_3143 ();
 sg13g2_decap_8 FILLER_68_3150 ();
 sg13g2_decap_8 FILLER_68_3157 ();
 sg13g2_decap_8 FILLER_68_3164 ();
 sg13g2_decap_8 FILLER_68_3171 ();
 sg13g2_decap_8 FILLER_68_3178 ();
 sg13g2_decap_8 FILLER_68_3185 ();
 sg13g2_decap_8 FILLER_68_3192 ();
 sg13g2_decap_8 FILLER_68_3199 ();
 sg13g2_decap_8 FILLER_68_3206 ();
 sg13g2_decap_8 FILLER_68_3213 ();
 sg13g2_decap_8 FILLER_68_3220 ();
 sg13g2_decap_8 FILLER_68_3227 ();
 sg13g2_decap_8 FILLER_68_3234 ();
 sg13g2_decap_8 FILLER_68_3241 ();
 sg13g2_decap_8 FILLER_68_3248 ();
 sg13g2_decap_8 FILLER_68_3255 ();
 sg13g2_decap_8 FILLER_68_3262 ();
 sg13g2_decap_8 FILLER_68_3269 ();
 sg13g2_decap_8 FILLER_68_3276 ();
 sg13g2_decap_8 FILLER_68_3283 ();
 sg13g2_decap_8 FILLER_68_3290 ();
 sg13g2_decap_8 FILLER_68_3297 ();
 sg13g2_decap_8 FILLER_68_3304 ();
 sg13g2_decap_8 FILLER_68_3311 ();
 sg13g2_decap_8 FILLER_68_3318 ();
 sg13g2_decap_8 FILLER_68_3325 ();
 sg13g2_decap_8 FILLER_68_3332 ();
 sg13g2_decap_8 FILLER_68_3339 ();
 sg13g2_decap_8 FILLER_68_3346 ();
 sg13g2_decap_8 FILLER_68_3353 ();
 sg13g2_decap_8 FILLER_68_3360 ();
 sg13g2_decap_8 FILLER_68_3367 ();
 sg13g2_decap_8 FILLER_68_3374 ();
 sg13g2_decap_8 FILLER_68_3381 ();
 sg13g2_decap_8 FILLER_68_3388 ();
 sg13g2_decap_8 FILLER_68_3395 ();
 sg13g2_decap_8 FILLER_68_3402 ();
 sg13g2_decap_8 FILLER_68_3409 ();
 sg13g2_decap_8 FILLER_68_3416 ();
 sg13g2_decap_8 FILLER_68_3423 ();
 sg13g2_decap_8 FILLER_68_3430 ();
 sg13g2_decap_8 FILLER_68_3437 ();
 sg13g2_decap_8 FILLER_68_3444 ();
 sg13g2_decap_8 FILLER_68_3451 ();
 sg13g2_decap_8 FILLER_68_3458 ();
 sg13g2_decap_8 FILLER_68_3465 ();
 sg13g2_decap_8 FILLER_68_3472 ();
 sg13g2_decap_8 FILLER_68_3479 ();
 sg13g2_decap_8 FILLER_68_3486 ();
 sg13g2_decap_8 FILLER_68_3493 ();
 sg13g2_decap_8 FILLER_68_3500 ();
 sg13g2_decap_8 FILLER_68_3507 ();
 sg13g2_decap_8 FILLER_68_3514 ();
 sg13g2_decap_8 FILLER_68_3521 ();
 sg13g2_decap_8 FILLER_68_3528 ();
 sg13g2_decap_8 FILLER_68_3535 ();
 sg13g2_decap_8 FILLER_68_3542 ();
 sg13g2_decap_8 FILLER_68_3549 ();
 sg13g2_decap_8 FILLER_68_3556 ();
 sg13g2_decap_8 FILLER_68_3563 ();
 sg13g2_decap_8 FILLER_68_3570 ();
 sg13g2_fill_2 FILLER_68_3577 ();
 sg13g2_fill_1 FILLER_68_3579 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_168 ();
 sg13g2_decap_8 FILLER_69_175 ();
 sg13g2_decap_8 FILLER_69_182 ();
 sg13g2_decap_8 FILLER_69_189 ();
 sg13g2_decap_8 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_203 ();
 sg13g2_decap_8 FILLER_69_210 ();
 sg13g2_decap_8 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_224 ();
 sg13g2_decap_8 FILLER_69_231 ();
 sg13g2_decap_8 FILLER_69_238 ();
 sg13g2_decap_8 FILLER_69_245 ();
 sg13g2_decap_8 FILLER_69_252 ();
 sg13g2_decap_8 FILLER_69_259 ();
 sg13g2_decap_8 FILLER_69_266 ();
 sg13g2_decap_8 FILLER_69_273 ();
 sg13g2_decap_8 FILLER_69_280 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_8 FILLER_69_294 ();
 sg13g2_decap_8 FILLER_69_301 ();
 sg13g2_decap_8 FILLER_69_308 ();
 sg13g2_decap_8 FILLER_69_315 ();
 sg13g2_decap_8 FILLER_69_322 ();
 sg13g2_decap_8 FILLER_69_329 ();
 sg13g2_decap_8 FILLER_69_336 ();
 sg13g2_decap_8 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_350 ();
 sg13g2_decap_8 FILLER_69_357 ();
 sg13g2_decap_8 FILLER_69_364 ();
 sg13g2_decap_8 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_378 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_decap_8 FILLER_69_406 ();
 sg13g2_decap_8 FILLER_69_413 ();
 sg13g2_decap_8 FILLER_69_420 ();
 sg13g2_decap_8 FILLER_69_427 ();
 sg13g2_decap_8 FILLER_69_434 ();
 sg13g2_decap_8 FILLER_69_441 ();
 sg13g2_decap_8 FILLER_69_448 ();
 sg13g2_fill_2 FILLER_69_455 ();
 sg13g2_fill_1 FILLER_69_457 ();
 sg13g2_decap_8 FILLER_69_463 ();
 sg13g2_decap_8 FILLER_69_470 ();
 sg13g2_decap_8 FILLER_69_477 ();
 sg13g2_decap_8 FILLER_69_484 ();
 sg13g2_decap_8 FILLER_69_491 ();
 sg13g2_decap_8 FILLER_69_498 ();
 sg13g2_decap_8 FILLER_69_505 ();
 sg13g2_decap_4 FILLER_69_512 ();
 sg13g2_fill_1 FILLER_69_516 ();
 sg13g2_fill_2 FILLER_69_530 ();
 sg13g2_fill_1 FILLER_69_532 ();
 sg13g2_decap_8 FILLER_69_559 ();
 sg13g2_decap_8 FILLER_69_566 ();
 sg13g2_decap_8 FILLER_69_573 ();
 sg13g2_decap_4 FILLER_69_580 ();
 sg13g2_fill_2 FILLER_69_584 ();
 sg13g2_fill_2 FILLER_69_594 ();
 sg13g2_decap_8 FILLER_69_630 ();
 sg13g2_decap_8 FILLER_69_672 ();
 sg13g2_decap_8 FILLER_69_679 ();
 sg13g2_fill_1 FILLER_69_686 ();
 sg13g2_fill_1 FILLER_69_718 ();
 sg13g2_fill_2 FILLER_69_745 ();
 sg13g2_decap_8 FILLER_69_755 ();
 sg13g2_decap_8 FILLER_69_762 ();
 sg13g2_decap_8 FILLER_69_769 ();
 sg13g2_decap_8 FILLER_69_776 ();
 sg13g2_decap_4 FILLER_69_796 ();
 sg13g2_fill_2 FILLER_69_800 ();
 sg13g2_decap_8 FILLER_69_805 ();
 sg13g2_decap_8 FILLER_69_812 ();
 sg13g2_decap_4 FILLER_69_819 ();
 sg13g2_decap_8 FILLER_69_828 ();
 sg13g2_fill_1 FILLER_69_867 ();
 sg13g2_fill_2 FILLER_69_891 ();
 sg13g2_fill_1 FILLER_69_893 ();
 sg13g2_fill_1 FILLER_69_902 ();
 sg13g2_decap_4 FILLER_69_911 ();
 sg13g2_fill_1 FILLER_69_915 ();
 sg13g2_fill_2 FILLER_69_924 ();
 sg13g2_fill_1 FILLER_69_926 ();
 sg13g2_decap_8 FILLER_69_953 ();
 sg13g2_decap_4 FILLER_69_964 ();
 sg13g2_fill_1 FILLER_69_968 ();
 sg13g2_fill_2 FILLER_69_977 ();
 sg13g2_fill_1 FILLER_69_979 ();
 sg13g2_decap_8 FILLER_69_984 ();
 sg13g2_fill_2 FILLER_69_991 ();
 sg13g2_decap_4 FILLER_69_998 ();
 sg13g2_fill_2 FILLER_69_1002 ();
 sg13g2_fill_2 FILLER_69_1045 ();
 sg13g2_fill_1 FILLER_69_1047 ();
 sg13g2_decap_4 FILLER_69_1092 ();
 sg13g2_decap_8 FILLER_69_1122 ();
 sg13g2_decap_8 FILLER_69_1129 ();
 sg13g2_decap_8 FILLER_69_1136 ();
 sg13g2_decap_4 FILLER_69_1143 ();
 sg13g2_fill_2 FILLER_69_1147 ();
 sg13g2_fill_1 FILLER_69_1182 ();
 sg13g2_decap_8 FILLER_69_1235 ();
 sg13g2_decap_4 FILLER_69_1242 ();
 sg13g2_fill_2 FILLER_69_1246 ();
 sg13g2_fill_2 FILLER_69_1274 ();
 sg13g2_fill_2 FILLER_69_1375 ();
 sg13g2_decap_8 FILLER_69_1429 ();
 sg13g2_fill_1 FILLER_69_1436 ();
 sg13g2_decap_8 FILLER_69_1463 ();
 sg13g2_decap_8 FILLER_69_1522 ();
 sg13g2_decap_8 FILLER_69_1529 ();
 sg13g2_decap_8 FILLER_69_1536 ();
 sg13g2_decap_8 FILLER_69_1543 ();
 sg13g2_decap_8 FILLER_69_1550 ();
 sg13g2_decap_8 FILLER_69_1588 ();
 sg13g2_fill_2 FILLER_69_1595 ();
 sg13g2_decap_4 FILLER_69_1641 ();
 sg13g2_decap_8 FILLER_69_1671 ();
 sg13g2_decap_4 FILLER_69_1678 ();
 sg13g2_decap_8 FILLER_69_1700 ();
 sg13g2_decap_8 FILLER_69_1707 ();
 sg13g2_decap_8 FILLER_69_1714 ();
 sg13g2_fill_1 FILLER_69_1721 ();
 sg13g2_fill_2 FILLER_69_1727 ();
 sg13g2_decap_8 FILLER_69_1742 ();
 sg13g2_decap_8 FILLER_69_1804 ();
 sg13g2_decap_8 FILLER_69_1811 ();
 sg13g2_decap_8 FILLER_69_1818 ();
 sg13g2_decap_8 FILLER_69_1825 ();
 sg13g2_decap_8 FILLER_69_1832 ();
 sg13g2_decap_8 FILLER_69_1839 ();
 sg13g2_decap_8 FILLER_69_1846 ();
 sg13g2_decap_8 FILLER_69_1853 ();
 sg13g2_fill_2 FILLER_69_1860 ();
 sg13g2_fill_1 FILLER_69_1862 ();
 sg13g2_fill_1 FILLER_69_1897 ();
 sg13g2_fill_2 FILLER_69_1958 ();
 sg13g2_decap_8 FILLER_69_1968 ();
 sg13g2_decap_8 FILLER_69_1975 ();
 sg13g2_decap_8 FILLER_69_1982 ();
 sg13g2_decap_8 FILLER_69_1989 ();
 sg13g2_fill_2 FILLER_69_2004 ();
 sg13g2_decap_8 FILLER_69_2032 ();
 sg13g2_decap_4 FILLER_69_2039 ();
 sg13g2_decap_8 FILLER_69_2048 ();
 sg13g2_decap_8 FILLER_69_2055 ();
 sg13g2_decap_8 FILLER_69_2062 ();
 sg13g2_decap_8 FILLER_69_2069 ();
 sg13g2_fill_2 FILLER_69_2076 ();
 sg13g2_fill_2 FILLER_69_2104 ();
 sg13g2_fill_1 FILLER_69_2106 ();
 sg13g2_decap_4 FILLER_69_2112 ();
 sg13g2_decap_4 FILLER_69_2155 ();
 sg13g2_decap_8 FILLER_69_2190 ();
 sg13g2_decap_8 FILLER_69_2197 ();
 sg13g2_decap_8 FILLER_69_2204 ();
 sg13g2_decap_8 FILLER_69_2211 ();
 sg13g2_decap_8 FILLER_69_2218 ();
 sg13g2_decap_8 FILLER_69_2225 ();
 sg13g2_decap_8 FILLER_69_2232 ();
 sg13g2_decap_8 FILLER_69_2239 ();
 sg13g2_decap_8 FILLER_69_2246 ();
 sg13g2_decap_8 FILLER_69_2253 ();
 sg13g2_decap_8 FILLER_69_2260 ();
 sg13g2_decap_8 FILLER_69_2267 ();
 sg13g2_decap_8 FILLER_69_2274 ();
 sg13g2_decap_8 FILLER_69_2281 ();
 sg13g2_decap_8 FILLER_69_2288 ();
 sg13g2_decap_8 FILLER_69_2295 ();
 sg13g2_decap_8 FILLER_69_2302 ();
 sg13g2_decap_8 FILLER_69_2309 ();
 sg13g2_decap_8 FILLER_69_2316 ();
 sg13g2_decap_8 FILLER_69_2323 ();
 sg13g2_decap_8 FILLER_69_2330 ();
 sg13g2_decap_8 FILLER_69_2337 ();
 sg13g2_decap_8 FILLER_69_2344 ();
 sg13g2_decap_8 FILLER_69_2351 ();
 sg13g2_decap_8 FILLER_69_2358 ();
 sg13g2_decap_8 FILLER_69_2365 ();
 sg13g2_decap_8 FILLER_69_2372 ();
 sg13g2_decap_8 FILLER_69_2379 ();
 sg13g2_decap_8 FILLER_69_2386 ();
 sg13g2_decap_8 FILLER_69_2393 ();
 sg13g2_decap_8 FILLER_69_2400 ();
 sg13g2_decap_8 FILLER_69_2407 ();
 sg13g2_decap_8 FILLER_69_2414 ();
 sg13g2_decap_8 FILLER_69_2421 ();
 sg13g2_decap_8 FILLER_69_2428 ();
 sg13g2_decap_8 FILLER_69_2435 ();
 sg13g2_decap_8 FILLER_69_2442 ();
 sg13g2_decap_8 FILLER_69_2449 ();
 sg13g2_decap_8 FILLER_69_2456 ();
 sg13g2_decap_8 FILLER_69_2463 ();
 sg13g2_decap_8 FILLER_69_2470 ();
 sg13g2_decap_8 FILLER_69_2477 ();
 sg13g2_decap_8 FILLER_69_2484 ();
 sg13g2_decap_8 FILLER_69_2491 ();
 sg13g2_decap_8 FILLER_69_2498 ();
 sg13g2_decap_8 FILLER_69_2505 ();
 sg13g2_decap_8 FILLER_69_2512 ();
 sg13g2_decap_8 FILLER_69_2519 ();
 sg13g2_decap_8 FILLER_69_2526 ();
 sg13g2_decap_8 FILLER_69_2533 ();
 sg13g2_decap_8 FILLER_69_2540 ();
 sg13g2_decap_8 FILLER_69_2547 ();
 sg13g2_decap_8 FILLER_69_2554 ();
 sg13g2_decap_8 FILLER_69_2561 ();
 sg13g2_decap_8 FILLER_69_2568 ();
 sg13g2_decap_8 FILLER_69_2575 ();
 sg13g2_decap_8 FILLER_69_2582 ();
 sg13g2_decap_8 FILLER_69_2589 ();
 sg13g2_decap_8 FILLER_69_2596 ();
 sg13g2_decap_8 FILLER_69_2603 ();
 sg13g2_decap_8 FILLER_69_2610 ();
 sg13g2_decap_8 FILLER_69_2617 ();
 sg13g2_decap_8 FILLER_69_2624 ();
 sg13g2_decap_8 FILLER_69_2631 ();
 sg13g2_decap_8 FILLER_69_2638 ();
 sg13g2_decap_8 FILLER_69_2645 ();
 sg13g2_decap_8 FILLER_69_2652 ();
 sg13g2_decap_8 FILLER_69_2659 ();
 sg13g2_decap_8 FILLER_69_2666 ();
 sg13g2_decap_8 FILLER_69_2673 ();
 sg13g2_decap_8 FILLER_69_2680 ();
 sg13g2_decap_8 FILLER_69_2687 ();
 sg13g2_decap_8 FILLER_69_2694 ();
 sg13g2_decap_8 FILLER_69_2701 ();
 sg13g2_decap_8 FILLER_69_2708 ();
 sg13g2_decap_8 FILLER_69_2715 ();
 sg13g2_decap_8 FILLER_69_2722 ();
 sg13g2_decap_8 FILLER_69_2729 ();
 sg13g2_decap_8 FILLER_69_2736 ();
 sg13g2_decap_8 FILLER_69_2743 ();
 sg13g2_decap_8 FILLER_69_2750 ();
 sg13g2_decap_8 FILLER_69_2757 ();
 sg13g2_decap_8 FILLER_69_2764 ();
 sg13g2_decap_8 FILLER_69_2771 ();
 sg13g2_decap_8 FILLER_69_2778 ();
 sg13g2_decap_8 FILLER_69_2785 ();
 sg13g2_decap_8 FILLER_69_2792 ();
 sg13g2_decap_8 FILLER_69_2799 ();
 sg13g2_decap_8 FILLER_69_2806 ();
 sg13g2_decap_8 FILLER_69_2813 ();
 sg13g2_decap_8 FILLER_69_2820 ();
 sg13g2_decap_8 FILLER_69_2827 ();
 sg13g2_decap_8 FILLER_69_2834 ();
 sg13g2_decap_8 FILLER_69_2841 ();
 sg13g2_decap_8 FILLER_69_2848 ();
 sg13g2_decap_8 FILLER_69_2855 ();
 sg13g2_decap_8 FILLER_69_2862 ();
 sg13g2_decap_8 FILLER_69_2869 ();
 sg13g2_decap_8 FILLER_69_2876 ();
 sg13g2_decap_8 FILLER_69_2883 ();
 sg13g2_decap_8 FILLER_69_2890 ();
 sg13g2_decap_8 FILLER_69_2897 ();
 sg13g2_decap_8 FILLER_69_2904 ();
 sg13g2_decap_8 FILLER_69_2911 ();
 sg13g2_decap_8 FILLER_69_2918 ();
 sg13g2_decap_8 FILLER_69_2925 ();
 sg13g2_decap_8 FILLER_69_2932 ();
 sg13g2_decap_8 FILLER_69_2939 ();
 sg13g2_decap_8 FILLER_69_2946 ();
 sg13g2_decap_8 FILLER_69_2953 ();
 sg13g2_decap_8 FILLER_69_2960 ();
 sg13g2_decap_8 FILLER_69_2967 ();
 sg13g2_decap_8 FILLER_69_2974 ();
 sg13g2_decap_8 FILLER_69_2981 ();
 sg13g2_decap_8 FILLER_69_2988 ();
 sg13g2_decap_8 FILLER_69_2995 ();
 sg13g2_decap_8 FILLER_69_3002 ();
 sg13g2_decap_8 FILLER_69_3009 ();
 sg13g2_decap_8 FILLER_69_3016 ();
 sg13g2_decap_8 FILLER_69_3023 ();
 sg13g2_decap_8 FILLER_69_3030 ();
 sg13g2_decap_8 FILLER_69_3037 ();
 sg13g2_decap_8 FILLER_69_3044 ();
 sg13g2_decap_8 FILLER_69_3051 ();
 sg13g2_decap_8 FILLER_69_3058 ();
 sg13g2_decap_8 FILLER_69_3065 ();
 sg13g2_decap_8 FILLER_69_3072 ();
 sg13g2_decap_8 FILLER_69_3079 ();
 sg13g2_decap_8 FILLER_69_3086 ();
 sg13g2_decap_8 FILLER_69_3093 ();
 sg13g2_decap_8 FILLER_69_3100 ();
 sg13g2_decap_8 FILLER_69_3107 ();
 sg13g2_decap_8 FILLER_69_3114 ();
 sg13g2_decap_8 FILLER_69_3121 ();
 sg13g2_decap_8 FILLER_69_3128 ();
 sg13g2_decap_8 FILLER_69_3135 ();
 sg13g2_decap_8 FILLER_69_3142 ();
 sg13g2_decap_8 FILLER_69_3149 ();
 sg13g2_decap_8 FILLER_69_3156 ();
 sg13g2_decap_8 FILLER_69_3163 ();
 sg13g2_decap_8 FILLER_69_3170 ();
 sg13g2_decap_8 FILLER_69_3177 ();
 sg13g2_decap_8 FILLER_69_3184 ();
 sg13g2_decap_8 FILLER_69_3191 ();
 sg13g2_decap_8 FILLER_69_3198 ();
 sg13g2_decap_8 FILLER_69_3205 ();
 sg13g2_decap_8 FILLER_69_3212 ();
 sg13g2_decap_8 FILLER_69_3219 ();
 sg13g2_decap_8 FILLER_69_3226 ();
 sg13g2_decap_8 FILLER_69_3233 ();
 sg13g2_decap_8 FILLER_69_3240 ();
 sg13g2_decap_8 FILLER_69_3247 ();
 sg13g2_decap_8 FILLER_69_3254 ();
 sg13g2_decap_8 FILLER_69_3261 ();
 sg13g2_decap_8 FILLER_69_3268 ();
 sg13g2_decap_8 FILLER_69_3275 ();
 sg13g2_decap_8 FILLER_69_3282 ();
 sg13g2_decap_8 FILLER_69_3289 ();
 sg13g2_decap_8 FILLER_69_3296 ();
 sg13g2_decap_8 FILLER_69_3303 ();
 sg13g2_decap_8 FILLER_69_3310 ();
 sg13g2_decap_8 FILLER_69_3317 ();
 sg13g2_decap_8 FILLER_69_3324 ();
 sg13g2_decap_8 FILLER_69_3331 ();
 sg13g2_decap_8 FILLER_69_3338 ();
 sg13g2_decap_8 FILLER_69_3345 ();
 sg13g2_decap_8 FILLER_69_3352 ();
 sg13g2_decap_8 FILLER_69_3359 ();
 sg13g2_decap_8 FILLER_69_3366 ();
 sg13g2_decap_8 FILLER_69_3373 ();
 sg13g2_decap_8 FILLER_69_3380 ();
 sg13g2_decap_8 FILLER_69_3387 ();
 sg13g2_decap_8 FILLER_69_3394 ();
 sg13g2_decap_8 FILLER_69_3401 ();
 sg13g2_decap_8 FILLER_69_3408 ();
 sg13g2_decap_8 FILLER_69_3415 ();
 sg13g2_decap_8 FILLER_69_3422 ();
 sg13g2_decap_8 FILLER_69_3429 ();
 sg13g2_decap_8 FILLER_69_3436 ();
 sg13g2_decap_8 FILLER_69_3443 ();
 sg13g2_decap_8 FILLER_69_3450 ();
 sg13g2_decap_8 FILLER_69_3457 ();
 sg13g2_decap_8 FILLER_69_3464 ();
 sg13g2_decap_8 FILLER_69_3471 ();
 sg13g2_decap_8 FILLER_69_3478 ();
 sg13g2_decap_8 FILLER_69_3485 ();
 sg13g2_decap_8 FILLER_69_3492 ();
 sg13g2_decap_8 FILLER_69_3499 ();
 sg13g2_decap_8 FILLER_69_3506 ();
 sg13g2_decap_8 FILLER_69_3513 ();
 sg13g2_decap_8 FILLER_69_3520 ();
 sg13g2_decap_8 FILLER_69_3527 ();
 sg13g2_decap_8 FILLER_69_3534 ();
 sg13g2_decap_8 FILLER_69_3541 ();
 sg13g2_decap_8 FILLER_69_3548 ();
 sg13g2_decap_8 FILLER_69_3555 ();
 sg13g2_decap_8 FILLER_69_3562 ();
 sg13g2_decap_8 FILLER_69_3569 ();
 sg13g2_decap_4 FILLER_69_3576 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_8 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_196 ();
 sg13g2_decap_8 FILLER_70_203 ();
 sg13g2_decap_8 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_217 ();
 sg13g2_decap_8 FILLER_70_224 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_decap_8 FILLER_70_252 ();
 sg13g2_decap_8 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_266 ();
 sg13g2_decap_8 FILLER_70_273 ();
 sg13g2_decap_8 FILLER_70_280 ();
 sg13g2_decap_8 FILLER_70_287 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_decap_8 FILLER_70_301 ();
 sg13g2_decap_8 FILLER_70_308 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_322 ();
 sg13g2_decap_8 FILLER_70_329 ();
 sg13g2_decap_8 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_8 FILLER_70_371 ();
 sg13g2_decap_8 FILLER_70_378 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_392 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_decap_8 FILLER_70_406 ();
 sg13g2_decap_8 FILLER_70_413 ();
 sg13g2_decap_8 FILLER_70_420 ();
 sg13g2_decap_8 FILLER_70_427 ();
 sg13g2_decap_8 FILLER_70_434 ();
 sg13g2_decap_8 FILLER_70_441 ();
 sg13g2_decap_8 FILLER_70_448 ();
 sg13g2_decap_8 FILLER_70_455 ();
 sg13g2_decap_8 FILLER_70_462 ();
 sg13g2_decap_8 FILLER_70_469 ();
 sg13g2_decap_8 FILLER_70_476 ();
 sg13g2_decap_8 FILLER_70_483 ();
 sg13g2_decap_8 FILLER_70_490 ();
 sg13g2_decap_8 FILLER_70_497 ();
 sg13g2_decap_8 FILLER_70_504 ();
 sg13g2_decap_8 FILLER_70_511 ();
 sg13g2_decap_8 FILLER_70_518 ();
 sg13g2_decap_8 FILLER_70_525 ();
 sg13g2_decap_8 FILLER_70_532 ();
 sg13g2_decap_8 FILLER_70_539 ();
 sg13g2_decap_8 FILLER_70_546 ();
 sg13g2_decap_8 FILLER_70_553 ();
 sg13g2_decap_8 FILLER_70_560 ();
 sg13g2_decap_8 FILLER_70_567 ();
 sg13g2_fill_2 FILLER_70_605 ();
 sg13g2_decap_8 FILLER_70_633 ();
 sg13g2_decap_8 FILLER_70_679 ();
 sg13g2_fill_2 FILLER_70_686 ();
 sg13g2_fill_1 FILLER_70_688 ();
 sg13g2_fill_2 FILLER_70_731 ();
 sg13g2_decap_8 FILLER_70_759 ();
 sg13g2_decap_4 FILLER_70_766 ();
 sg13g2_decap_8 FILLER_70_822 ();
 sg13g2_decap_8 FILLER_70_829 ();
 sg13g2_decap_8 FILLER_70_836 ();
 sg13g2_fill_1 FILLER_70_843 ();
 sg13g2_fill_1 FILLER_70_855 ();
 sg13g2_fill_2 FILLER_70_882 ();
 sg13g2_fill_1 FILLER_70_915 ();
 sg13g2_decap_4 FILLER_70_933 ();
 sg13g2_fill_1 FILLER_70_937 ();
 sg13g2_decap_8 FILLER_70_942 ();
 sg13g2_decap_4 FILLER_70_949 ();
 sg13g2_fill_1 FILLER_70_1026 ();
 sg13g2_fill_2 FILLER_70_1053 ();
 sg13g2_decap_8 FILLER_70_1116 ();
 sg13g2_decap_8 FILLER_70_1123 ();
 sg13g2_decap_8 FILLER_70_1130 ();
 sg13g2_fill_1 FILLER_70_1137 ();
 sg13g2_fill_1 FILLER_70_1168 ();
 sg13g2_fill_1 FILLER_70_1208 ();
 sg13g2_decap_8 FILLER_70_1235 ();
 sg13g2_decap_8 FILLER_70_1242 ();
 sg13g2_decap_8 FILLER_70_1249 ();
 sg13g2_decap_8 FILLER_70_1256 ();
 sg13g2_decap_8 FILLER_70_1263 ();
 sg13g2_fill_2 FILLER_70_1270 ();
 sg13g2_fill_1 FILLER_70_1280 ();
 sg13g2_fill_2 FILLER_70_1307 ();
 sg13g2_fill_1 FILLER_70_1309 ();
 sg13g2_decap_8 FILLER_70_1315 ();
 sg13g2_decap_8 FILLER_70_1322 ();
 sg13g2_decap_8 FILLER_70_1368 ();
 sg13g2_decap_8 FILLER_70_1375 ();
 sg13g2_decap_8 FILLER_70_1382 ();
 sg13g2_decap_8 FILLER_70_1389 ();
 sg13g2_decap_8 FILLER_70_1401 ();
 sg13g2_decap_4 FILLER_70_1408 ();
 sg13g2_fill_2 FILLER_70_1412 ();
 sg13g2_decap_8 FILLER_70_1418 ();
 sg13g2_decap_8 FILLER_70_1425 ();
 sg13g2_decap_4 FILLER_70_1432 ();
 sg13g2_fill_1 FILLER_70_1436 ();
 sg13g2_decap_8 FILLER_70_1463 ();
 sg13g2_decap_8 FILLER_70_1470 ();
 sg13g2_decap_8 FILLER_70_1477 ();
 sg13g2_fill_1 FILLER_70_1484 ();
 sg13g2_decap_8 FILLER_70_1511 ();
 sg13g2_decap_4 FILLER_70_1518 ();
 sg13g2_decap_8 FILLER_70_1582 ();
 sg13g2_decap_8 FILLER_70_1634 ();
 sg13g2_fill_1 FILLER_70_1641 ();
 sg13g2_decap_8 FILLER_70_1658 ();
 sg13g2_fill_2 FILLER_70_1665 ();
 sg13g2_fill_1 FILLER_70_1667 ();
 sg13g2_fill_2 FILLER_70_1700 ();
 sg13g2_fill_1 FILLER_70_1702 ();
 sg13g2_fill_2 FILLER_70_1755 ();
 sg13g2_decap_4 FILLER_70_1783 ();
 sg13g2_fill_2 FILLER_70_1816 ();
 sg13g2_decap_8 FILLER_70_1852 ();
 sg13g2_fill_1 FILLER_70_1859 ();
 sg13g2_fill_2 FILLER_70_1938 ();
 sg13g2_fill_1 FILLER_70_1940 ();
 sg13g2_decap_4 FILLER_70_1951 ();
 sg13g2_decap_8 FILLER_70_1966 ();
 sg13g2_decap_8 FILLER_70_1973 ();
 sg13g2_decap_8 FILLER_70_1980 ();
 sg13g2_decap_4 FILLER_70_1987 ();
 sg13g2_fill_2 FILLER_70_1991 ();
 sg13g2_fill_2 FILLER_70_2031 ();
 sg13g2_decap_8 FILLER_70_2041 ();
 sg13g2_fill_1 FILLER_70_2048 ();
 sg13g2_decap_8 FILLER_70_2065 ();
 sg13g2_fill_1 FILLER_70_2072 ();
 sg13g2_fill_1 FILLER_70_2092 ();
 sg13g2_decap_8 FILLER_70_2119 ();
 sg13g2_fill_2 FILLER_70_2126 ();
 sg13g2_fill_1 FILLER_70_2128 ();
 sg13g2_decap_8 FILLER_70_2207 ();
 sg13g2_decap_8 FILLER_70_2214 ();
 sg13g2_decap_8 FILLER_70_2221 ();
 sg13g2_decap_8 FILLER_70_2228 ();
 sg13g2_decap_8 FILLER_70_2235 ();
 sg13g2_decap_8 FILLER_70_2242 ();
 sg13g2_decap_8 FILLER_70_2249 ();
 sg13g2_decap_8 FILLER_70_2256 ();
 sg13g2_decap_8 FILLER_70_2263 ();
 sg13g2_decap_8 FILLER_70_2270 ();
 sg13g2_decap_8 FILLER_70_2277 ();
 sg13g2_decap_8 FILLER_70_2284 ();
 sg13g2_decap_8 FILLER_70_2291 ();
 sg13g2_decap_8 FILLER_70_2298 ();
 sg13g2_decap_8 FILLER_70_2305 ();
 sg13g2_decap_8 FILLER_70_2312 ();
 sg13g2_decap_8 FILLER_70_2319 ();
 sg13g2_decap_8 FILLER_70_2326 ();
 sg13g2_decap_8 FILLER_70_2333 ();
 sg13g2_decap_8 FILLER_70_2340 ();
 sg13g2_decap_8 FILLER_70_2347 ();
 sg13g2_decap_8 FILLER_70_2354 ();
 sg13g2_decap_8 FILLER_70_2361 ();
 sg13g2_decap_8 FILLER_70_2368 ();
 sg13g2_decap_8 FILLER_70_2375 ();
 sg13g2_decap_8 FILLER_70_2382 ();
 sg13g2_decap_8 FILLER_70_2389 ();
 sg13g2_decap_8 FILLER_70_2396 ();
 sg13g2_decap_8 FILLER_70_2403 ();
 sg13g2_decap_8 FILLER_70_2410 ();
 sg13g2_decap_8 FILLER_70_2417 ();
 sg13g2_decap_8 FILLER_70_2424 ();
 sg13g2_decap_8 FILLER_70_2431 ();
 sg13g2_decap_8 FILLER_70_2438 ();
 sg13g2_decap_8 FILLER_70_2445 ();
 sg13g2_decap_8 FILLER_70_2452 ();
 sg13g2_decap_8 FILLER_70_2459 ();
 sg13g2_decap_8 FILLER_70_2466 ();
 sg13g2_decap_8 FILLER_70_2473 ();
 sg13g2_decap_8 FILLER_70_2480 ();
 sg13g2_decap_8 FILLER_70_2487 ();
 sg13g2_decap_8 FILLER_70_2494 ();
 sg13g2_decap_8 FILLER_70_2501 ();
 sg13g2_decap_8 FILLER_70_2508 ();
 sg13g2_decap_8 FILLER_70_2515 ();
 sg13g2_decap_8 FILLER_70_2522 ();
 sg13g2_decap_8 FILLER_70_2529 ();
 sg13g2_decap_8 FILLER_70_2536 ();
 sg13g2_decap_8 FILLER_70_2543 ();
 sg13g2_decap_8 FILLER_70_2550 ();
 sg13g2_decap_8 FILLER_70_2557 ();
 sg13g2_decap_8 FILLER_70_2564 ();
 sg13g2_decap_8 FILLER_70_2571 ();
 sg13g2_decap_8 FILLER_70_2578 ();
 sg13g2_decap_8 FILLER_70_2585 ();
 sg13g2_decap_8 FILLER_70_2592 ();
 sg13g2_decap_8 FILLER_70_2599 ();
 sg13g2_decap_8 FILLER_70_2606 ();
 sg13g2_decap_8 FILLER_70_2613 ();
 sg13g2_decap_8 FILLER_70_2620 ();
 sg13g2_decap_8 FILLER_70_2627 ();
 sg13g2_decap_8 FILLER_70_2634 ();
 sg13g2_decap_8 FILLER_70_2641 ();
 sg13g2_decap_8 FILLER_70_2648 ();
 sg13g2_decap_8 FILLER_70_2655 ();
 sg13g2_decap_8 FILLER_70_2662 ();
 sg13g2_decap_8 FILLER_70_2669 ();
 sg13g2_decap_8 FILLER_70_2676 ();
 sg13g2_decap_8 FILLER_70_2683 ();
 sg13g2_decap_8 FILLER_70_2690 ();
 sg13g2_decap_8 FILLER_70_2697 ();
 sg13g2_decap_8 FILLER_70_2704 ();
 sg13g2_decap_8 FILLER_70_2711 ();
 sg13g2_decap_8 FILLER_70_2718 ();
 sg13g2_decap_8 FILLER_70_2725 ();
 sg13g2_decap_8 FILLER_70_2732 ();
 sg13g2_decap_8 FILLER_70_2739 ();
 sg13g2_decap_8 FILLER_70_2746 ();
 sg13g2_decap_8 FILLER_70_2753 ();
 sg13g2_decap_8 FILLER_70_2760 ();
 sg13g2_decap_8 FILLER_70_2767 ();
 sg13g2_decap_8 FILLER_70_2774 ();
 sg13g2_decap_8 FILLER_70_2781 ();
 sg13g2_decap_8 FILLER_70_2788 ();
 sg13g2_decap_8 FILLER_70_2795 ();
 sg13g2_decap_8 FILLER_70_2802 ();
 sg13g2_decap_8 FILLER_70_2809 ();
 sg13g2_decap_8 FILLER_70_2816 ();
 sg13g2_decap_8 FILLER_70_2823 ();
 sg13g2_decap_8 FILLER_70_2830 ();
 sg13g2_decap_8 FILLER_70_2837 ();
 sg13g2_decap_8 FILLER_70_2844 ();
 sg13g2_decap_8 FILLER_70_2851 ();
 sg13g2_decap_8 FILLER_70_2858 ();
 sg13g2_decap_8 FILLER_70_2865 ();
 sg13g2_decap_8 FILLER_70_2872 ();
 sg13g2_decap_8 FILLER_70_2879 ();
 sg13g2_decap_8 FILLER_70_2886 ();
 sg13g2_decap_8 FILLER_70_2893 ();
 sg13g2_decap_8 FILLER_70_2900 ();
 sg13g2_decap_8 FILLER_70_2907 ();
 sg13g2_decap_8 FILLER_70_2914 ();
 sg13g2_decap_8 FILLER_70_2921 ();
 sg13g2_decap_8 FILLER_70_2928 ();
 sg13g2_decap_8 FILLER_70_2935 ();
 sg13g2_decap_8 FILLER_70_2942 ();
 sg13g2_decap_8 FILLER_70_2949 ();
 sg13g2_decap_8 FILLER_70_2956 ();
 sg13g2_decap_8 FILLER_70_2963 ();
 sg13g2_decap_8 FILLER_70_2970 ();
 sg13g2_decap_8 FILLER_70_2977 ();
 sg13g2_decap_8 FILLER_70_2984 ();
 sg13g2_decap_8 FILLER_70_2991 ();
 sg13g2_decap_8 FILLER_70_2998 ();
 sg13g2_decap_8 FILLER_70_3005 ();
 sg13g2_decap_8 FILLER_70_3012 ();
 sg13g2_decap_8 FILLER_70_3019 ();
 sg13g2_decap_8 FILLER_70_3026 ();
 sg13g2_decap_8 FILLER_70_3033 ();
 sg13g2_decap_8 FILLER_70_3040 ();
 sg13g2_decap_8 FILLER_70_3047 ();
 sg13g2_decap_8 FILLER_70_3054 ();
 sg13g2_decap_8 FILLER_70_3061 ();
 sg13g2_decap_8 FILLER_70_3068 ();
 sg13g2_decap_8 FILLER_70_3075 ();
 sg13g2_decap_8 FILLER_70_3082 ();
 sg13g2_decap_8 FILLER_70_3089 ();
 sg13g2_decap_8 FILLER_70_3096 ();
 sg13g2_decap_8 FILLER_70_3103 ();
 sg13g2_decap_8 FILLER_70_3110 ();
 sg13g2_decap_8 FILLER_70_3117 ();
 sg13g2_decap_8 FILLER_70_3124 ();
 sg13g2_decap_8 FILLER_70_3131 ();
 sg13g2_decap_8 FILLER_70_3138 ();
 sg13g2_decap_8 FILLER_70_3145 ();
 sg13g2_decap_8 FILLER_70_3152 ();
 sg13g2_decap_8 FILLER_70_3159 ();
 sg13g2_decap_8 FILLER_70_3166 ();
 sg13g2_decap_8 FILLER_70_3173 ();
 sg13g2_decap_8 FILLER_70_3180 ();
 sg13g2_decap_8 FILLER_70_3187 ();
 sg13g2_decap_8 FILLER_70_3194 ();
 sg13g2_decap_8 FILLER_70_3201 ();
 sg13g2_decap_8 FILLER_70_3208 ();
 sg13g2_decap_8 FILLER_70_3215 ();
 sg13g2_decap_8 FILLER_70_3222 ();
 sg13g2_decap_8 FILLER_70_3229 ();
 sg13g2_decap_8 FILLER_70_3236 ();
 sg13g2_decap_8 FILLER_70_3243 ();
 sg13g2_decap_8 FILLER_70_3250 ();
 sg13g2_decap_8 FILLER_70_3257 ();
 sg13g2_decap_8 FILLER_70_3264 ();
 sg13g2_decap_8 FILLER_70_3271 ();
 sg13g2_decap_8 FILLER_70_3278 ();
 sg13g2_decap_8 FILLER_70_3285 ();
 sg13g2_decap_8 FILLER_70_3292 ();
 sg13g2_decap_8 FILLER_70_3299 ();
 sg13g2_decap_8 FILLER_70_3306 ();
 sg13g2_decap_8 FILLER_70_3313 ();
 sg13g2_decap_8 FILLER_70_3320 ();
 sg13g2_decap_8 FILLER_70_3327 ();
 sg13g2_decap_8 FILLER_70_3334 ();
 sg13g2_decap_8 FILLER_70_3341 ();
 sg13g2_decap_8 FILLER_70_3348 ();
 sg13g2_decap_8 FILLER_70_3355 ();
 sg13g2_decap_8 FILLER_70_3362 ();
 sg13g2_decap_8 FILLER_70_3369 ();
 sg13g2_decap_8 FILLER_70_3376 ();
 sg13g2_decap_8 FILLER_70_3383 ();
 sg13g2_decap_8 FILLER_70_3390 ();
 sg13g2_decap_8 FILLER_70_3397 ();
 sg13g2_decap_8 FILLER_70_3404 ();
 sg13g2_decap_8 FILLER_70_3411 ();
 sg13g2_decap_8 FILLER_70_3418 ();
 sg13g2_decap_8 FILLER_70_3425 ();
 sg13g2_decap_8 FILLER_70_3432 ();
 sg13g2_decap_8 FILLER_70_3439 ();
 sg13g2_decap_8 FILLER_70_3446 ();
 sg13g2_decap_8 FILLER_70_3453 ();
 sg13g2_decap_8 FILLER_70_3460 ();
 sg13g2_decap_8 FILLER_70_3467 ();
 sg13g2_decap_8 FILLER_70_3474 ();
 sg13g2_decap_8 FILLER_70_3481 ();
 sg13g2_decap_8 FILLER_70_3488 ();
 sg13g2_decap_8 FILLER_70_3495 ();
 sg13g2_decap_8 FILLER_70_3502 ();
 sg13g2_decap_8 FILLER_70_3509 ();
 sg13g2_decap_8 FILLER_70_3516 ();
 sg13g2_decap_8 FILLER_70_3523 ();
 sg13g2_decap_8 FILLER_70_3530 ();
 sg13g2_decap_8 FILLER_70_3537 ();
 sg13g2_decap_8 FILLER_70_3544 ();
 sg13g2_decap_8 FILLER_70_3551 ();
 sg13g2_decap_8 FILLER_70_3558 ();
 sg13g2_decap_8 FILLER_70_3565 ();
 sg13g2_decap_8 FILLER_70_3572 ();
 sg13g2_fill_1 FILLER_70_3579 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_203 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_245 ();
 sg13g2_decap_8 FILLER_71_252 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_decap_8 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_273 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_decap_8 FILLER_71_315 ();
 sg13g2_decap_8 FILLER_71_322 ();
 sg13g2_decap_8 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_decap_8 FILLER_71_350 ();
 sg13g2_decap_8 FILLER_71_357 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_399 ();
 sg13g2_decap_8 FILLER_71_406 ();
 sg13g2_decap_8 FILLER_71_413 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_decap_8 FILLER_71_427 ();
 sg13g2_decap_8 FILLER_71_434 ();
 sg13g2_decap_8 FILLER_71_441 ();
 sg13g2_decap_8 FILLER_71_448 ();
 sg13g2_decap_8 FILLER_71_455 ();
 sg13g2_decap_8 FILLER_71_462 ();
 sg13g2_decap_8 FILLER_71_469 ();
 sg13g2_decap_8 FILLER_71_476 ();
 sg13g2_decap_8 FILLER_71_483 ();
 sg13g2_decap_8 FILLER_71_490 ();
 sg13g2_decap_8 FILLER_71_497 ();
 sg13g2_decap_8 FILLER_71_504 ();
 sg13g2_decap_8 FILLER_71_511 ();
 sg13g2_decap_8 FILLER_71_518 ();
 sg13g2_decap_8 FILLER_71_525 ();
 sg13g2_decap_8 FILLER_71_532 ();
 sg13g2_decap_8 FILLER_71_539 ();
 sg13g2_decap_8 FILLER_71_546 ();
 sg13g2_decap_8 FILLER_71_553 ();
 sg13g2_decap_8 FILLER_71_560 ();
 sg13g2_decap_8 FILLER_71_567 ();
 sg13g2_decap_4 FILLER_71_574 ();
 sg13g2_decap_8 FILLER_71_617 ();
 sg13g2_decap_8 FILLER_71_624 ();
 sg13g2_decap_8 FILLER_71_631 ();
 sg13g2_decap_8 FILLER_71_638 ();
 sg13g2_fill_1 FILLER_71_645 ();
 sg13g2_fill_2 FILLER_71_659 ();
 sg13g2_fill_1 FILLER_71_661 ();
 sg13g2_decap_8 FILLER_71_674 ();
 sg13g2_decap_8 FILLER_71_681 ();
 sg13g2_decap_4 FILLER_71_688 ();
 sg13g2_fill_1 FILLER_71_692 ();
 sg13g2_fill_1 FILLER_71_719 ();
 sg13g2_decap_8 FILLER_71_751 ();
 sg13g2_decap_8 FILLER_71_758 ();
 sg13g2_fill_1 FILLER_71_765 ();
 sg13g2_fill_1 FILLER_71_774 ();
 sg13g2_decap_4 FILLER_71_831 ();
 sg13g2_fill_1 FILLER_71_835 ();
 sg13g2_fill_2 FILLER_71_893 ();
 sg13g2_fill_1 FILLER_71_900 ();
 sg13g2_fill_1 FILLER_71_932 ();
 sg13g2_decap_8 FILLER_71_989 ();
 sg13g2_decap_8 FILLER_71_996 ();
 sg13g2_decap_8 FILLER_71_1031 ();
 sg13g2_decap_4 FILLER_71_1038 ();
 sg13g2_fill_2 FILLER_71_1042 ();
 sg13g2_decap_4 FILLER_71_1090 ();
 sg13g2_fill_1 FILLER_71_1094 ();
 sg13g2_decap_8 FILLER_71_1099 ();
 sg13g2_fill_2 FILLER_71_1106 ();
 sg13g2_decap_4 FILLER_71_1121 ();
 sg13g2_fill_2 FILLER_71_1125 ();
 sg13g2_decap_4 FILLER_71_1160 ();
 sg13g2_fill_2 FILLER_71_1164 ();
 sg13g2_fill_2 FILLER_71_1174 ();
 sg13g2_fill_1 FILLER_71_1176 ();
 sg13g2_decap_8 FILLER_71_1198 ();
 sg13g2_decap_8 FILLER_71_1205 ();
 sg13g2_decap_8 FILLER_71_1212 ();
 sg13g2_fill_1 FILLER_71_1219 ();
 sg13g2_fill_1 FILLER_71_1224 ();
 sg13g2_decap_8 FILLER_71_1251 ();
 sg13g2_fill_1 FILLER_71_1261 ();
 sg13g2_fill_2 FILLER_71_1291 ();
 sg13g2_decap_4 FILLER_71_1301 ();
 sg13g2_decap_8 FILLER_71_1331 ();
 sg13g2_decap_8 FILLER_71_1411 ();
 sg13g2_decap_4 FILLER_71_1418 ();
 sg13g2_fill_2 FILLER_71_1422 ();
 sg13g2_fill_1 FILLER_71_1505 ();
 sg13g2_fill_1 FILLER_71_1532 ();
 sg13g2_decap_8 FILLER_71_1551 ();
 sg13g2_fill_1 FILLER_71_1558 ();
 sg13g2_fill_2 FILLER_71_1585 ();
 sg13g2_fill_1 FILLER_71_1587 ();
 sg13g2_decap_8 FILLER_71_1626 ();
 sg13g2_decap_8 FILLER_71_1633 ();
 sg13g2_decap_8 FILLER_71_1640 ();
 sg13g2_decap_4 FILLER_71_1647 ();
 sg13g2_decap_4 FILLER_71_1717 ();
 sg13g2_decap_4 FILLER_71_1725 ();
 sg13g2_fill_2 FILLER_71_1755 ();
 sg13g2_decap_8 FILLER_71_1801 ();
 sg13g2_decap_4 FILLER_71_1808 ();
 sg13g2_fill_2 FILLER_71_1812 ();
 sg13g2_fill_2 FILLER_71_1852 ();
 sg13g2_fill_1 FILLER_71_1906 ();
 sg13g2_decap_4 FILLER_71_1955 ();
 sg13g2_fill_2 FILLER_71_1980 ();
 sg13g2_fill_1 FILLER_71_1982 ();
 sg13g2_fill_2 FILLER_71_2009 ();
 sg13g2_fill_1 FILLER_71_2011 ();
 sg13g2_decap_8 FILLER_71_2052 ();
 sg13g2_decap_8 FILLER_71_2059 ();
 sg13g2_decap_4 FILLER_71_2066 ();
 sg13g2_decap_8 FILLER_71_2137 ();
 sg13g2_decap_8 FILLER_71_2184 ();
 sg13g2_decap_8 FILLER_71_2191 ();
 sg13g2_decap_8 FILLER_71_2198 ();
 sg13g2_decap_8 FILLER_71_2205 ();
 sg13g2_decap_8 FILLER_71_2212 ();
 sg13g2_decap_8 FILLER_71_2219 ();
 sg13g2_decap_8 FILLER_71_2226 ();
 sg13g2_decap_8 FILLER_71_2233 ();
 sg13g2_decap_8 FILLER_71_2240 ();
 sg13g2_decap_8 FILLER_71_2247 ();
 sg13g2_decap_8 FILLER_71_2254 ();
 sg13g2_decap_8 FILLER_71_2261 ();
 sg13g2_decap_8 FILLER_71_2268 ();
 sg13g2_decap_8 FILLER_71_2275 ();
 sg13g2_decap_8 FILLER_71_2282 ();
 sg13g2_decap_8 FILLER_71_2289 ();
 sg13g2_decap_8 FILLER_71_2296 ();
 sg13g2_decap_8 FILLER_71_2303 ();
 sg13g2_decap_8 FILLER_71_2310 ();
 sg13g2_decap_8 FILLER_71_2317 ();
 sg13g2_decap_8 FILLER_71_2324 ();
 sg13g2_decap_8 FILLER_71_2331 ();
 sg13g2_decap_8 FILLER_71_2338 ();
 sg13g2_decap_8 FILLER_71_2345 ();
 sg13g2_decap_8 FILLER_71_2352 ();
 sg13g2_decap_8 FILLER_71_2359 ();
 sg13g2_decap_8 FILLER_71_2366 ();
 sg13g2_decap_8 FILLER_71_2373 ();
 sg13g2_decap_8 FILLER_71_2380 ();
 sg13g2_decap_8 FILLER_71_2387 ();
 sg13g2_decap_8 FILLER_71_2394 ();
 sg13g2_decap_8 FILLER_71_2401 ();
 sg13g2_decap_8 FILLER_71_2408 ();
 sg13g2_decap_8 FILLER_71_2415 ();
 sg13g2_decap_8 FILLER_71_2422 ();
 sg13g2_decap_8 FILLER_71_2429 ();
 sg13g2_decap_8 FILLER_71_2436 ();
 sg13g2_decap_8 FILLER_71_2443 ();
 sg13g2_decap_8 FILLER_71_2450 ();
 sg13g2_decap_8 FILLER_71_2457 ();
 sg13g2_decap_8 FILLER_71_2464 ();
 sg13g2_decap_8 FILLER_71_2471 ();
 sg13g2_decap_8 FILLER_71_2478 ();
 sg13g2_decap_8 FILLER_71_2485 ();
 sg13g2_decap_8 FILLER_71_2492 ();
 sg13g2_decap_8 FILLER_71_2499 ();
 sg13g2_decap_8 FILLER_71_2506 ();
 sg13g2_decap_8 FILLER_71_2513 ();
 sg13g2_decap_8 FILLER_71_2520 ();
 sg13g2_decap_8 FILLER_71_2527 ();
 sg13g2_decap_8 FILLER_71_2534 ();
 sg13g2_decap_8 FILLER_71_2541 ();
 sg13g2_decap_8 FILLER_71_2548 ();
 sg13g2_decap_8 FILLER_71_2555 ();
 sg13g2_decap_8 FILLER_71_2562 ();
 sg13g2_decap_8 FILLER_71_2569 ();
 sg13g2_decap_8 FILLER_71_2576 ();
 sg13g2_decap_8 FILLER_71_2583 ();
 sg13g2_decap_8 FILLER_71_2590 ();
 sg13g2_decap_8 FILLER_71_2597 ();
 sg13g2_decap_8 FILLER_71_2604 ();
 sg13g2_decap_8 FILLER_71_2611 ();
 sg13g2_decap_8 FILLER_71_2618 ();
 sg13g2_decap_8 FILLER_71_2625 ();
 sg13g2_decap_8 FILLER_71_2632 ();
 sg13g2_decap_8 FILLER_71_2639 ();
 sg13g2_decap_8 FILLER_71_2646 ();
 sg13g2_decap_8 FILLER_71_2653 ();
 sg13g2_decap_8 FILLER_71_2660 ();
 sg13g2_decap_8 FILLER_71_2667 ();
 sg13g2_decap_8 FILLER_71_2674 ();
 sg13g2_decap_8 FILLER_71_2681 ();
 sg13g2_decap_8 FILLER_71_2688 ();
 sg13g2_decap_8 FILLER_71_2695 ();
 sg13g2_decap_8 FILLER_71_2702 ();
 sg13g2_decap_8 FILLER_71_2709 ();
 sg13g2_decap_8 FILLER_71_2716 ();
 sg13g2_decap_8 FILLER_71_2723 ();
 sg13g2_decap_8 FILLER_71_2730 ();
 sg13g2_decap_8 FILLER_71_2737 ();
 sg13g2_decap_8 FILLER_71_2744 ();
 sg13g2_decap_8 FILLER_71_2751 ();
 sg13g2_decap_8 FILLER_71_2758 ();
 sg13g2_decap_8 FILLER_71_2765 ();
 sg13g2_decap_8 FILLER_71_2772 ();
 sg13g2_decap_8 FILLER_71_2779 ();
 sg13g2_decap_8 FILLER_71_2786 ();
 sg13g2_decap_8 FILLER_71_2793 ();
 sg13g2_decap_8 FILLER_71_2800 ();
 sg13g2_decap_8 FILLER_71_2807 ();
 sg13g2_decap_8 FILLER_71_2814 ();
 sg13g2_decap_8 FILLER_71_2821 ();
 sg13g2_decap_8 FILLER_71_2828 ();
 sg13g2_decap_8 FILLER_71_2835 ();
 sg13g2_decap_8 FILLER_71_2842 ();
 sg13g2_decap_8 FILLER_71_2849 ();
 sg13g2_decap_8 FILLER_71_2856 ();
 sg13g2_decap_8 FILLER_71_2863 ();
 sg13g2_decap_8 FILLER_71_2870 ();
 sg13g2_decap_8 FILLER_71_2877 ();
 sg13g2_decap_8 FILLER_71_2884 ();
 sg13g2_decap_8 FILLER_71_2891 ();
 sg13g2_decap_8 FILLER_71_2898 ();
 sg13g2_decap_8 FILLER_71_2905 ();
 sg13g2_decap_8 FILLER_71_2912 ();
 sg13g2_decap_8 FILLER_71_2919 ();
 sg13g2_decap_8 FILLER_71_2926 ();
 sg13g2_decap_8 FILLER_71_2933 ();
 sg13g2_decap_8 FILLER_71_2940 ();
 sg13g2_decap_8 FILLER_71_2947 ();
 sg13g2_decap_8 FILLER_71_2954 ();
 sg13g2_decap_8 FILLER_71_2961 ();
 sg13g2_decap_8 FILLER_71_2968 ();
 sg13g2_decap_8 FILLER_71_2975 ();
 sg13g2_decap_8 FILLER_71_2982 ();
 sg13g2_decap_8 FILLER_71_2989 ();
 sg13g2_decap_8 FILLER_71_2996 ();
 sg13g2_decap_8 FILLER_71_3003 ();
 sg13g2_decap_8 FILLER_71_3010 ();
 sg13g2_decap_8 FILLER_71_3017 ();
 sg13g2_decap_8 FILLER_71_3024 ();
 sg13g2_decap_8 FILLER_71_3031 ();
 sg13g2_decap_8 FILLER_71_3038 ();
 sg13g2_decap_8 FILLER_71_3045 ();
 sg13g2_decap_8 FILLER_71_3052 ();
 sg13g2_decap_8 FILLER_71_3059 ();
 sg13g2_decap_8 FILLER_71_3066 ();
 sg13g2_decap_8 FILLER_71_3073 ();
 sg13g2_decap_8 FILLER_71_3080 ();
 sg13g2_decap_8 FILLER_71_3087 ();
 sg13g2_decap_8 FILLER_71_3094 ();
 sg13g2_decap_8 FILLER_71_3101 ();
 sg13g2_decap_8 FILLER_71_3108 ();
 sg13g2_decap_8 FILLER_71_3115 ();
 sg13g2_decap_8 FILLER_71_3122 ();
 sg13g2_decap_8 FILLER_71_3129 ();
 sg13g2_decap_8 FILLER_71_3136 ();
 sg13g2_decap_8 FILLER_71_3143 ();
 sg13g2_decap_8 FILLER_71_3150 ();
 sg13g2_decap_8 FILLER_71_3157 ();
 sg13g2_decap_8 FILLER_71_3164 ();
 sg13g2_decap_8 FILLER_71_3171 ();
 sg13g2_decap_8 FILLER_71_3178 ();
 sg13g2_decap_8 FILLER_71_3185 ();
 sg13g2_decap_8 FILLER_71_3192 ();
 sg13g2_decap_8 FILLER_71_3199 ();
 sg13g2_decap_8 FILLER_71_3206 ();
 sg13g2_decap_8 FILLER_71_3213 ();
 sg13g2_decap_8 FILLER_71_3220 ();
 sg13g2_decap_8 FILLER_71_3227 ();
 sg13g2_decap_8 FILLER_71_3234 ();
 sg13g2_decap_8 FILLER_71_3241 ();
 sg13g2_decap_8 FILLER_71_3248 ();
 sg13g2_decap_8 FILLER_71_3255 ();
 sg13g2_decap_8 FILLER_71_3262 ();
 sg13g2_decap_8 FILLER_71_3269 ();
 sg13g2_decap_8 FILLER_71_3276 ();
 sg13g2_decap_8 FILLER_71_3283 ();
 sg13g2_decap_8 FILLER_71_3290 ();
 sg13g2_decap_8 FILLER_71_3297 ();
 sg13g2_decap_8 FILLER_71_3304 ();
 sg13g2_decap_8 FILLER_71_3311 ();
 sg13g2_decap_8 FILLER_71_3318 ();
 sg13g2_decap_8 FILLER_71_3325 ();
 sg13g2_decap_8 FILLER_71_3332 ();
 sg13g2_decap_8 FILLER_71_3339 ();
 sg13g2_decap_8 FILLER_71_3346 ();
 sg13g2_decap_8 FILLER_71_3353 ();
 sg13g2_decap_8 FILLER_71_3360 ();
 sg13g2_decap_8 FILLER_71_3367 ();
 sg13g2_decap_8 FILLER_71_3374 ();
 sg13g2_decap_8 FILLER_71_3381 ();
 sg13g2_decap_8 FILLER_71_3388 ();
 sg13g2_decap_8 FILLER_71_3395 ();
 sg13g2_decap_8 FILLER_71_3402 ();
 sg13g2_decap_8 FILLER_71_3409 ();
 sg13g2_decap_8 FILLER_71_3416 ();
 sg13g2_decap_8 FILLER_71_3423 ();
 sg13g2_decap_8 FILLER_71_3430 ();
 sg13g2_decap_8 FILLER_71_3437 ();
 sg13g2_decap_8 FILLER_71_3444 ();
 sg13g2_decap_8 FILLER_71_3451 ();
 sg13g2_decap_8 FILLER_71_3458 ();
 sg13g2_decap_8 FILLER_71_3465 ();
 sg13g2_decap_8 FILLER_71_3472 ();
 sg13g2_decap_8 FILLER_71_3479 ();
 sg13g2_decap_8 FILLER_71_3486 ();
 sg13g2_decap_8 FILLER_71_3493 ();
 sg13g2_decap_8 FILLER_71_3500 ();
 sg13g2_decap_8 FILLER_71_3507 ();
 sg13g2_decap_8 FILLER_71_3514 ();
 sg13g2_decap_8 FILLER_71_3521 ();
 sg13g2_decap_8 FILLER_71_3528 ();
 sg13g2_decap_8 FILLER_71_3535 ();
 sg13g2_decap_8 FILLER_71_3542 ();
 sg13g2_decap_8 FILLER_71_3549 ();
 sg13g2_decap_8 FILLER_71_3556 ();
 sg13g2_decap_8 FILLER_71_3563 ();
 sg13g2_decap_8 FILLER_71_3570 ();
 sg13g2_fill_2 FILLER_71_3577 ();
 sg13g2_fill_1 FILLER_71_3579 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_252 ();
 sg13g2_decap_8 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_280 ();
 sg13g2_decap_8 FILLER_72_287 ();
 sg13g2_decap_8 FILLER_72_294 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_8 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_343 ();
 sg13g2_decap_8 FILLER_72_350 ();
 sg13g2_decap_8 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_decap_8 FILLER_72_406 ();
 sg13g2_decap_8 FILLER_72_413 ();
 sg13g2_decap_8 FILLER_72_420 ();
 sg13g2_decap_8 FILLER_72_427 ();
 sg13g2_decap_8 FILLER_72_434 ();
 sg13g2_decap_8 FILLER_72_441 ();
 sg13g2_decap_8 FILLER_72_448 ();
 sg13g2_decap_8 FILLER_72_455 ();
 sg13g2_decap_8 FILLER_72_462 ();
 sg13g2_decap_8 FILLER_72_469 ();
 sg13g2_decap_8 FILLER_72_476 ();
 sg13g2_decap_8 FILLER_72_483 ();
 sg13g2_decap_8 FILLER_72_490 ();
 sg13g2_decap_8 FILLER_72_497 ();
 sg13g2_decap_8 FILLER_72_504 ();
 sg13g2_decap_8 FILLER_72_511 ();
 sg13g2_decap_8 FILLER_72_518 ();
 sg13g2_decap_8 FILLER_72_525 ();
 sg13g2_decap_8 FILLER_72_532 ();
 sg13g2_decap_8 FILLER_72_539 ();
 sg13g2_decap_8 FILLER_72_546 ();
 sg13g2_decap_8 FILLER_72_553 ();
 sg13g2_decap_8 FILLER_72_560 ();
 sg13g2_decap_8 FILLER_72_567 ();
 sg13g2_fill_2 FILLER_72_574 ();
 sg13g2_fill_1 FILLER_72_576 ();
 sg13g2_decap_8 FILLER_72_619 ();
 sg13g2_decap_8 FILLER_72_626 ();
 sg13g2_decap_4 FILLER_72_633 ();
 sg13g2_fill_1 FILLER_72_637 ();
 sg13g2_decap_8 FILLER_72_669 ();
 sg13g2_decap_8 FILLER_72_676 ();
 sg13g2_fill_1 FILLER_72_721 ();
 sg13g2_fill_1 FILLER_72_727 ();
 sg13g2_decap_8 FILLER_72_736 ();
 sg13g2_decap_8 FILLER_72_743 ();
 sg13g2_decap_4 FILLER_72_750 ();
 sg13g2_fill_2 FILLER_72_754 ();
 sg13g2_decap_8 FILLER_72_821 ();
 sg13g2_decap_8 FILLER_72_828 ();
 sg13g2_decap_8 FILLER_72_835 ();
 sg13g2_decap_8 FILLER_72_842 ();
 sg13g2_fill_2 FILLER_72_849 ();
 sg13g2_fill_1 FILLER_72_851 ();
 sg13g2_decap_4 FILLER_72_860 ();
 sg13g2_fill_2 FILLER_72_864 ();
 sg13g2_fill_2 FILLER_72_870 ();
 sg13g2_fill_1 FILLER_72_872 ();
 sg13g2_decap_8 FILLER_72_877 ();
 sg13g2_decap_8 FILLER_72_884 ();
 sg13g2_decap_8 FILLER_72_891 ();
 sg13g2_fill_2 FILLER_72_898 ();
 sg13g2_fill_2 FILLER_72_907 ();
 sg13g2_fill_1 FILLER_72_909 ();
 sg13g2_decap_4 FILLER_72_945 ();
 sg13g2_decap_8 FILLER_72_1031 ();
 sg13g2_decap_8 FILLER_72_1042 ();
 sg13g2_fill_2 FILLER_72_1115 ();
 sg13g2_decap_8 FILLER_72_1125 ();
 sg13g2_fill_2 FILLER_72_1132 ();
 sg13g2_decap_4 FILLER_72_1160 ();
 sg13g2_decap_4 FILLER_72_1194 ();
 sg13g2_fill_2 FILLER_72_1198 ();
 sg13g2_decap_4 FILLER_72_1205 ();
 sg13g2_fill_1 FILLER_72_1217 ();
 sg13g2_decap_8 FILLER_72_1223 ();
 sg13g2_fill_1 FILLER_72_1230 ();
 sg13g2_fill_2 FILLER_72_1314 ();
 sg13g2_fill_2 FILLER_72_1346 ();
 sg13g2_fill_1 FILLER_72_1348 ();
 sg13g2_fill_2 FILLER_72_1352 ();
 sg13g2_fill_1 FILLER_72_1354 ();
 sg13g2_fill_1 FILLER_72_1407 ();
 sg13g2_fill_1 FILLER_72_1421 ();
 sg13g2_fill_2 FILLER_72_1482 ();
 sg13g2_fill_2 FILLER_72_1523 ();
 sg13g2_decap_8 FILLER_72_1577 ();
 sg13g2_decap_4 FILLER_72_1584 ();
 sg13g2_decap_4 FILLER_72_1614 ();
 sg13g2_decap_8 FILLER_72_1623 ();
 sg13g2_fill_1 FILLER_72_1643 ();
 sg13g2_fill_2 FILLER_72_1649 ();
 sg13g2_decap_8 FILLER_72_1677 ();
 sg13g2_fill_1 FILLER_72_1684 ();
 sg13g2_decap_8 FILLER_72_1715 ();
 sg13g2_decap_4 FILLER_72_1722 ();
 sg13g2_fill_2 FILLER_72_1726 ();
 sg13g2_decap_8 FILLER_72_1733 ();
 sg13g2_decap_8 FILLER_72_1740 ();
 sg13g2_fill_2 FILLER_72_1747 ();
 sg13g2_decap_8 FILLER_72_1841 ();
 sg13g2_decap_8 FILLER_72_1848 ();
 sg13g2_decap_8 FILLER_72_1855 ();
 sg13g2_fill_1 FILLER_72_1862 ();
 sg13g2_decap_8 FILLER_72_1889 ();
 sg13g2_fill_1 FILLER_72_1896 ();
 sg13g2_fill_1 FILLER_72_1923 ();
 sg13g2_fill_2 FILLER_72_1950 ();
 sg13g2_fill_2 FILLER_72_2012 ();
 sg13g2_fill_2 FILLER_72_2073 ();
 sg13g2_fill_1 FILLER_72_2075 ();
 sg13g2_decap_8 FILLER_72_2135 ();
 sg13g2_decap_8 FILLER_72_2142 ();
 sg13g2_decap_8 FILLER_72_2149 ();
 sg13g2_decap_8 FILLER_72_2156 ();
 sg13g2_decap_8 FILLER_72_2163 ();
 sg13g2_decap_8 FILLER_72_2170 ();
 sg13g2_decap_8 FILLER_72_2177 ();
 sg13g2_decap_8 FILLER_72_2184 ();
 sg13g2_decap_8 FILLER_72_2191 ();
 sg13g2_decap_8 FILLER_72_2198 ();
 sg13g2_decap_8 FILLER_72_2205 ();
 sg13g2_decap_8 FILLER_72_2212 ();
 sg13g2_decap_8 FILLER_72_2219 ();
 sg13g2_decap_8 FILLER_72_2226 ();
 sg13g2_decap_8 FILLER_72_2233 ();
 sg13g2_decap_8 FILLER_72_2240 ();
 sg13g2_decap_8 FILLER_72_2247 ();
 sg13g2_decap_8 FILLER_72_2254 ();
 sg13g2_decap_8 FILLER_72_2261 ();
 sg13g2_decap_8 FILLER_72_2268 ();
 sg13g2_decap_8 FILLER_72_2275 ();
 sg13g2_decap_8 FILLER_72_2282 ();
 sg13g2_decap_8 FILLER_72_2289 ();
 sg13g2_decap_8 FILLER_72_2296 ();
 sg13g2_decap_8 FILLER_72_2303 ();
 sg13g2_decap_8 FILLER_72_2310 ();
 sg13g2_decap_8 FILLER_72_2317 ();
 sg13g2_decap_8 FILLER_72_2324 ();
 sg13g2_decap_8 FILLER_72_2331 ();
 sg13g2_decap_8 FILLER_72_2338 ();
 sg13g2_decap_8 FILLER_72_2345 ();
 sg13g2_decap_8 FILLER_72_2352 ();
 sg13g2_decap_8 FILLER_72_2359 ();
 sg13g2_decap_8 FILLER_72_2366 ();
 sg13g2_decap_8 FILLER_72_2373 ();
 sg13g2_decap_8 FILLER_72_2380 ();
 sg13g2_decap_8 FILLER_72_2387 ();
 sg13g2_decap_8 FILLER_72_2394 ();
 sg13g2_decap_8 FILLER_72_2401 ();
 sg13g2_decap_8 FILLER_72_2408 ();
 sg13g2_decap_8 FILLER_72_2415 ();
 sg13g2_decap_8 FILLER_72_2422 ();
 sg13g2_decap_8 FILLER_72_2429 ();
 sg13g2_decap_8 FILLER_72_2436 ();
 sg13g2_decap_8 FILLER_72_2443 ();
 sg13g2_decap_8 FILLER_72_2450 ();
 sg13g2_decap_8 FILLER_72_2457 ();
 sg13g2_decap_8 FILLER_72_2464 ();
 sg13g2_decap_8 FILLER_72_2471 ();
 sg13g2_decap_8 FILLER_72_2478 ();
 sg13g2_decap_8 FILLER_72_2485 ();
 sg13g2_decap_8 FILLER_72_2492 ();
 sg13g2_decap_8 FILLER_72_2499 ();
 sg13g2_decap_8 FILLER_72_2506 ();
 sg13g2_decap_8 FILLER_72_2513 ();
 sg13g2_decap_8 FILLER_72_2520 ();
 sg13g2_decap_8 FILLER_72_2527 ();
 sg13g2_decap_8 FILLER_72_2534 ();
 sg13g2_decap_8 FILLER_72_2541 ();
 sg13g2_decap_8 FILLER_72_2548 ();
 sg13g2_decap_8 FILLER_72_2555 ();
 sg13g2_decap_8 FILLER_72_2562 ();
 sg13g2_decap_8 FILLER_72_2569 ();
 sg13g2_decap_8 FILLER_72_2576 ();
 sg13g2_decap_8 FILLER_72_2583 ();
 sg13g2_decap_8 FILLER_72_2590 ();
 sg13g2_decap_8 FILLER_72_2597 ();
 sg13g2_decap_8 FILLER_72_2604 ();
 sg13g2_decap_8 FILLER_72_2611 ();
 sg13g2_decap_8 FILLER_72_2618 ();
 sg13g2_decap_8 FILLER_72_2625 ();
 sg13g2_decap_8 FILLER_72_2632 ();
 sg13g2_decap_8 FILLER_72_2639 ();
 sg13g2_decap_8 FILLER_72_2646 ();
 sg13g2_decap_8 FILLER_72_2653 ();
 sg13g2_decap_8 FILLER_72_2660 ();
 sg13g2_decap_8 FILLER_72_2667 ();
 sg13g2_decap_8 FILLER_72_2674 ();
 sg13g2_decap_8 FILLER_72_2681 ();
 sg13g2_decap_8 FILLER_72_2688 ();
 sg13g2_decap_8 FILLER_72_2695 ();
 sg13g2_decap_8 FILLER_72_2702 ();
 sg13g2_decap_8 FILLER_72_2709 ();
 sg13g2_decap_8 FILLER_72_2716 ();
 sg13g2_decap_8 FILLER_72_2723 ();
 sg13g2_decap_8 FILLER_72_2730 ();
 sg13g2_decap_8 FILLER_72_2737 ();
 sg13g2_decap_8 FILLER_72_2744 ();
 sg13g2_decap_8 FILLER_72_2751 ();
 sg13g2_decap_8 FILLER_72_2758 ();
 sg13g2_decap_8 FILLER_72_2765 ();
 sg13g2_decap_8 FILLER_72_2772 ();
 sg13g2_decap_8 FILLER_72_2779 ();
 sg13g2_decap_8 FILLER_72_2786 ();
 sg13g2_decap_8 FILLER_72_2793 ();
 sg13g2_decap_8 FILLER_72_2800 ();
 sg13g2_decap_8 FILLER_72_2807 ();
 sg13g2_decap_8 FILLER_72_2814 ();
 sg13g2_decap_8 FILLER_72_2821 ();
 sg13g2_decap_8 FILLER_72_2828 ();
 sg13g2_decap_8 FILLER_72_2835 ();
 sg13g2_decap_8 FILLER_72_2842 ();
 sg13g2_decap_8 FILLER_72_2849 ();
 sg13g2_decap_8 FILLER_72_2856 ();
 sg13g2_decap_8 FILLER_72_2863 ();
 sg13g2_decap_8 FILLER_72_2870 ();
 sg13g2_decap_8 FILLER_72_2877 ();
 sg13g2_decap_8 FILLER_72_2884 ();
 sg13g2_decap_8 FILLER_72_2891 ();
 sg13g2_decap_8 FILLER_72_2898 ();
 sg13g2_decap_8 FILLER_72_2905 ();
 sg13g2_decap_8 FILLER_72_2912 ();
 sg13g2_decap_8 FILLER_72_2919 ();
 sg13g2_decap_8 FILLER_72_2926 ();
 sg13g2_decap_8 FILLER_72_2933 ();
 sg13g2_decap_8 FILLER_72_2940 ();
 sg13g2_decap_8 FILLER_72_2947 ();
 sg13g2_decap_8 FILLER_72_2954 ();
 sg13g2_decap_8 FILLER_72_2961 ();
 sg13g2_decap_8 FILLER_72_2968 ();
 sg13g2_decap_8 FILLER_72_2975 ();
 sg13g2_decap_8 FILLER_72_2982 ();
 sg13g2_decap_8 FILLER_72_2989 ();
 sg13g2_decap_8 FILLER_72_2996 ();
 sg13g2_decap_8 FILLER_72_3003 ();
 sg13g2_decap_8 FILLER_72_3010 ();
 sg13g2_decap_8 FILLER_72_3017 ();
 sg13g2_decap_8 FILLER_72_3024 ();
 sg13g2_decap_8 FILLER_72_3031 ();
 sg13g2_decap_8 FILLER_72_3038 ();
 sg13g2_decap_8 FILLER_72_3045 ();
 sg13g2_decap_8 FILLER_72_3052 ();
 sg13g2_decap_8 FILLER_72_3059 ();
 sg13g2_decap_8 FILLER_72_3066 ();
 sg13g2_decap_8 FILLER_72_3073 ();
 sg13g2_decap_8 FILLER_72_3080 ();
 sg13g2_decap_8 FILLER_72_3087 ();
 sg13g2_decap_8 FILLER_72_3094 ();
 sg13g2_decap_8 FILLER_72_3101 ();
 sg13g2_decap_8 FILLER_72_3108 ();
 sg13g2_decap_8 FILLER_72_3115 ();
 sg13g2_decap_8 FILLER_72_3122 ();
 sg13g2_decap_8 FILLER_72_3129 ();
 sg13g2_decap_8 FILLER_72_3136 ();
 sg13g2_decap_8 FILLER_72_3143 ();
 sg13g2_decap_8 FILLER_72_3150 ();
 sg13g2_decap_8 FILLER_72_3157 ();
 sg13g2_decap_8 FILLER_72_3164 ();
 sg13g2_decap_8 FILLER_72_3171 ();
 sg13g2_decap_8 FILLER_72_3178 ();
 sg13g2_decap_8 FILLER_72_3185 ();
 sg13g2_decap_8 FILLER_72_3192 ();
 sg13g2_decap_8 FILLER_72_3199 ();
 sg13g2_decap_8 FILLER_72_3206 ();
 sg13g2_decap_8 FILLER_72_3213 ();
 sg13g2_decap_8 FILLER_72_3220 ();
 sg13g2_decap_8 FILLER_72_3227 ();
 sg13g2_decap_8 FILLER_72_3234 ();
 sg13g2_decap_8 FILLER_72_3241 ();
 sg13g2_decap_8 FILLER_72_3248 ();
 sg13g2_decap_8 FILLER_72_3255 ();
 sg13g2_decap_8 FILLER_72_3262 ();
 sg13g2_decap_8 FILLER_72_3269 ();
 sg13g2_decap_8 FILLER_72_3276 ();
 sg13g2_decap_8 FILLER_72_3283 ();
 sg13g2_decap_8 FILLER_72_3290 ();
 sg13g2_decap_8 FILLER_72_3297 ();
 sg13g2_decap_8 FILLER_72_3304 ();
 sg13g2_decap_8 FILLER_72_3311 ();
 sg13g2_decap_8 FILLER_72_3318 ();
 sg13g2_decap_8 FILLER_72_3325 ();
 sg13g2_decap_8 FILLER_72_3332 ();
 sg13g2_decap_8 FILLER_72_3339 ();
 sg13g2_decap_8 FILLER_72_3346 ();
 sg13g2_decap_8 FILLER_72_3353 ();
 sg13g2_decap_8 FILLER_72_3360 ();
 sg13g2_decap_8 FILLER_72_3367 ();
 sg13g2_decap_8 FILLER_72_3374 ();
 sg13g2_decap_8 FILLER_72_3381 ();
 sg13g2_decap_8 FILLER_72_3388 ();
 sg13g2_decap_8 FILLER_72_3395 ();
 sg13g2_decap_8 FILLER_72_3402 ();
 sg13g2_decap_8 FILLER_72_3409 ();
 sg13g2_decap_8 FILLER_72_3416 ();
 sg13g2_decap_8 FILLER_72_3423 ();
 sg13g2_decap_8 FILLER_72_3430 ();
 sg13g2_decap_8 FILLER_72_3437 ();
 sg13g2_decap_8 FILLER_72_3444 ();
 sg13g2_decap_8 FILLER_72_3451 ();
 sg13g2_decap_8 FILLER_72_3458 ();
 sg13g2_decap_8 FILLER_72_3465 ();
 sg13g2_decap_8 FILLER_72_3472 ();
 sg13g2_decap_8 FILLER_72_3479 ();
 sg13g2_decap_8 FILLER_72_3486 ();
 sg13g2_decap_8 FILLER_72_3493 ();
 sg13g2_decap_8 FILLER_72_3500 ();
 sg13g2_decap_8 FILLER_72_3507 ();
 sg13g2_decap_8 FILLER_72_3514 ();
 sg13g2_decap_8 FILLER_72_3521 ();
 sg13g2_decap_8 FILLER_72_3528 ();
 sg13g2_decap_8 FILLER_72_3535 ();
 sg13g2_decap_8 FILLER_72_3542 ();
 sg13g2_decap_8 FILLER_72_3549 ();
 sg13g2_decap_8 FILLER_72_3556 ();
 sg13g2_decap_8 FILLER_72_3563 ();
 sg13g2_decap_8 FILLER_72_3570 ();
 sg13g2_fill_2 FILLER_72_3577 ();
 sg13g2_fill_1 FILLER_72_3579 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_8 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_decap_8 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_245 ();
 sg13g2_decap_8 FILLER_73_252 ();
 sg13g2_decap_8 FILLER_73_259 ();
 sg13g2_decap_8 FILLER_73_266 ();
 sg13g2_decap_8 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_decap_8 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_322 ();
 sg13g2_decap_8 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_73_336 ();
 sg13g2_decap_8 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_350 ();
 sg13g2_decap_8 FILLER_73_357 ();
 sg13g2_decap_8 FILLER_73_364 ();
 sg13g2_decap_8 FILLER_73_371 ();
 sg13g2_decap_8 FILLER_73_378 ();
 sg13g2_decap_8 FILLER_73_385 ();
 sg13g2_decap_8 FILLER_73_392 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_decap_8 FILLER_73_427 ();
 sg13g2_decap_8 FILLER_73_434 ();
 sg13g2_decap_8 FILLER_73_441 ();
 sg13g2_decap_8 FILLER_73_448 ();
 sg13g2_decap_8 FILLER_73_455 ();
 sg13g2_decap_8 FILLER_73_462 ();
 sg13g2_decap_8 FILLER_73_469 ();
 sg13g2_decap_8 FILLER_73_476 ();
 sg13g2_decap_8 FILLER_73_483 ();
 sg13g2_decap_8 FILLER_73_490 ();
 sg13g2_decap_8 FILLER_73_497 ();
 sg13g2_decap_8 FILLER_73_504 ();
 sg13g2_decap_8 FILLER_73_511 ();
 sg13g2_decap_8 FILLER_73_518 ();
 sg13g2_decap_8 FILLER_73_525 ();
 sg13g2_decap_8 FILLER_73_532 ();
 sg13g2_decap_8 FILLER_73_539 ();
 sg13g2_decap_8 FILLER_73_546 ();
 sg13g2_decap_8 FILLER_73_553 ();
 sg13g2_decap_8 FILLER_73_560 ();
 sg13g2_decap_8 FILLER_73_567 ();
 sg13g2_decap_4 FILLER_73_574 ();
 sg13g2_decap_8 FILLER_73_616 ();
 sg13g2_fill_1 FILLER_73_623 ();
 sg13g2_decap_8 FILLER_73_674 ();
 sg13g2_decap_8 FILLER_73_681 ();
 sg13g2_decap_8 FILLER_73_700 ();
 sg13g2_decap_8 FILLER_73_711 ();
 sg13g2_decap_8 FILLER_73_718 ();
 sg13g2_decap_8 FILLER_73_725 ();
 sg13g2_fill_2 FILLER_73_732 ();
 sg13g2_fill_1 FILLER_73_734 ();
 sg13g2_fill_1 FILLER_73_761 ();
 sg13g2_fill_2 FILLER_73_769 ();
 sg13g2_decap_8 FILLER_73_787 ();
 sg13g2_fill_2 FILLER_73_794 ();
 sg13g2_fill_1 FILLER_73_796 ();
 sg13g2_decap_8 FILLER_73_820 ();
 sg13g2_fill_2 FILLER_73_827 ();
 sg13g2_fill_1 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_847 ();
 sg13g2_decap_8 FILLER_73_854 ();
 sg13g2_fill_2 FILLER_73_861 ();
 sg13g2_fill_1 FILLER_73_863 ();
 sg13g2_decap_4 FILLER_73_869 ();
 sg13g2_fill_2 FILLER_73_873 ();
 sg13g2_fill_2 FILLER_73_901 ();
 sg13g2_fill_2 FILLER_73_910 ();
 sg13g2_fill_2 FILLER_73_917 ();
 sg13g2_fill_1 FILLER_73_924 ();
 sg13g2_decap_8 FILLER_73_959 ();
 sg13g2_fill_2 FILLER_73_966 ();
 sg13g2_fill_1 FILLER_73_968 ();
 sg13g2_decap_8 FILLER_73_973 ();
 sg13g2_fill_2 FILLER_73_980 ();
 sg13g2_decap_8 FILLER_73_986 ();
 sg13g2_decap_8 FILLER_73_993 ();
 sg13g2_decap_4 FILLER_73_1000 ();
 sg13g2_fill_2 FILLER_73_1004 ();
 sg13g2_fill_2 FILLER_73_1010 ();
 sg13g2_fill_2 FILLER_73_1017 ();
 sg13g2_decap_8 FILLER_73_1045 ();
 sg13g2_decap_8 FILLER_73_1052 ();
 sg13g2_fill_2 FILLER_73_1059 ();
 sg13g2_decap_4 FILLER_73_1066 ();
 sg13g2_decap_8 FILLER_73_1110 ();
 sg13g2_decap_8 FILLER_73_1117 ();
 sg13g2_decap_8 FILLER_73_1124 ();
 sg13g2_decap_8 FILLER_73_1131 ();
 sg13g2_decap_8 FILLER_73_1138 ();
 sg13g2_decap_8 FILLER_73_1149 ();
 sg13g2_decap_8 FILLER_73_1156 ();
 sg13g2_fill_1 FILLER_73_1163 ();
 sg13g2_decap_4 FILLER_73_1246 ();
 sg13g2_fill_1 FILLER_73_1250 ();
 sg13g2_decap_8 FILLER_73_1289 ();
 sg13g2_fill_2 FILLER_73_1296 ();
 sg13g2_fill_1 FILLER_73_1302 ();
 sg13g2_fill_2 FILLER_73_1337 ();
 sg13g2_decap_8 FILLER_73_1360 ();
 sg13g2_fill_2 FILLER_73_1367 ();
 sg13g2_fill_2 FILLER_73_1373 ();
 sg13g2_fill_2 FILLER_73_1379 ();
 sg13g2_fill_2 FILLER_73_1444 ();
 sg13g2_decap_8 FILLER_73_1475 ();
 sg13g2_decap_8 FILLER_73_1482 ();
 sg13g2_fill_1 FILLER_73_1529 ();
 sg13g2_decap_8 FILLER_73_1590 ();
 sg13g2_fill_2 FILLER_73_1597 ();
 sg13g2_decap_4 FILLER_73_1603 ();
 sg13g2_fill_1 FILLER_73_1607 ();
 sg13g2_fill_1 FILLER_73_1634 ();
 sg13g2_fill_2 FILLER_73_1686 ();
 sg13g2_fill_1 FILLER_73_1700 ();
 sg13g2_decap_8 FILLER_73_1779 ();
 sg13g2_decap_8 FILLER_73_1786 ();
 sg13g2_decap_8 FILLER_73_1793 ();
 sg13g2_fill_1 FILLER_73_1832 ();
 sg13g2_decap_8 FILLER_73_1837 ();
 sg13g2_decap_8 FILLER_73_1844 ();
 sg13g2_decap_8 FILLER_73_1851 ();
 sg13g2_decap_8 FILLER_73_1858 ();
 sg13g2_decap_8 FILLER_73_1865 ();
 sg13g2_decap_8 FILLER_73_1872 ();
 sg13g2_decap_8 FILLER_73_1879 ();
 sg13g2_decap_8 FILLER_73_1886 ();
 sg13g2_decap_8 FILLER_73_1893 ();
 sg13g2_decap_4 FILLER_73_1900 ();
 sg13g2_decap_4 FILLER_73_1909 ();
 sg13g2_decap_8 FILLER_73_1996 ();
 sg13g2_decap_8 FILLER_73_2003 ();
 sg13g2_decap_8 FILLER_73_2010 ();
 sg13g2_fill_1 FILLER_73_2017 ();
 sg13g2_decap_8 FILLER_73_2055 ();
 sg13g2_decap_8 FILLER_73_2062 ();
 sg13g2_fill_2 FILLER_73_2069 ();
 sg13g2_fill_1 FILLER_73_2071 ();
 sg13g2_decap_8 FILLER_73_2130 ();
 sg13g2_decap_8 FILLER_73_2137 ();
 sg13g2_decap_8 FILLER_73_2144 ();
 sg13g2_decap_8 FILLER_73_2151 ();
 sg13g2_decap_8 FILLER_73_2158 ();
 sg13g2_decap_8 FILLER_73_2165 ();
 sg13g2_decap_8 FILLER_73_2172 ();
 sg13g2_decap_8 FILLER_73_2179 ();
 sg13g2_decap_8 FILLER_73_2186 ();
 sg13g2_decap_8 FILLER_73_2193 ();
 sg13g2_decap_8 FILLER_73_2200 ();
 sg13g2_decap_8 FILLER_73_2207 ();
 sg13g2_decap_8 FILLER_73_2214 ();
 sg13g2_decap_8 FILLER_73_2221 ();
 sg13g2_decap_8 FILLER_73_2228 ();
 sg13g2_decap_8 FILLER_73_2235 ();
 sg13g2_decap_8 FILLER_73_2242 ();
 sg13g2_decap_8 FILLER_73_2249 ();
 sg13g2_decap_8 FILLER_73_2256 ();
 sg13g2_decap_8 FILLER_73_2263 ();
 sg13g2_decap_8 FILLER_73_2270 ();
 sg13g2_decap_8 FILLER_73_2277 ();
 sg13g2_decap_8 FILLER_73_2284 ();
 sg13g2_decap_8 FILLER_73_2291 ();
 sg13g2_decap_8 FILLER_73_2298 ();
 sg13g2_decap_8 FILLER_73_2305 ();
 sg13g2_decap_8 FILLER_73_2312 ();
 sg13g2_decap_8 FILLER_73_2319 ();
 sg13g2_decap_8 FILLER_73_2326 ();
 sg13g2_decap_8 FILLER_73_2333 ();
 sg13g2_decap_8 FILLER_73_2340 ();
 sg13g2_decap_8 FILLER_73_2347 ();
 sg13g2_decap_8 FILLER_73_2354 ();
 sg13g2_decap_8 FILLER_73_2361 ();
 sg13g2_decap_8 FILLER_73_2368 ();
 sg13g2_decap_8 FILLER_73_2375 ();
 sg13g2_decap_8 FILLER_73_2382 ();
 sg13g2_decap_8 FILLER_73_2389 ();
 sg13g2_decap_8 FILLER_73_2396 ();
 sg13g2_decap_8 FILLER_73_2403 ();
 sg13g2_decap_8 FILLER_73_2410 ();
 sg13g2_decap_8 FILLER_73_2417 ();
 sg13g2_decap_8 FILLER_73_2424 ();
 sg13g2_decap_8 FILLER_73_2431 ();
 sg13g2_decap_8 FILLER_73_2438 ();
 sg13g2_decap_8 FILLER_73_2445 ();
 sg13g2_decap_8 FILLER_73_2452 ();
 sg13g2_decap_8 FILLER_73_2459 ();
 sg13g2_decap_8 FILLER_73_2466 ();
 sg13g2_decap_8 FILLER_73_2473 ();
 sg13g2_decap_8 FILLER_73_2480 ();
 sg13g2_decap_8 FILLER_73_2487 ();
 sg13g2_decap_8 FILLER_73_2494 ();
 sg13g2_decap_8 FILLER_73_2501 ();
 sg13g2_decap_8 FILLER_73_2508 ();
 sg13g2_decap_8 FILLER_73_2515 ();
 sg13g2_decap_8 FILLER_73_2522 ();
 sg13g2_decap_8 FILLER_73_2529 ();
 sg13g2_decap_8 FILLER_73_2536 ();
 sg13g2_decap_8 FILLER_73_2543 ();
 sg13g2_decap_8 FILLER_73_2550 ();
 sg13g2_decap_8 FILLER_73_2557 ();
 sg13g2_decap_8 FILLER_73_2564 ();
 sg13g2_decap_8 FILLER_73_2571 ();
 sg13g2_decap_8 FILLER_73_2578 ();
 sg13g2_decap_8 FILLER_73_2585 ();
 sg13g2_decap_8 FILLER_73_2592 ();
 sg13g2_decap_8 FILLER_73_2599 ();
 sg13g2_decap_8 FILLER_73_2606 ();
 sg13g2_decap_8 FILLER_73_2613 ();
 sg13g2_decap_8 FILLER_73_2620 ();
 sg13g2_decap_8 FILLER_73_2627 ();
 sg13g2_decap_8 FILLER_73_2634 ();
 sg13g2_decap_8 FILLER_73_2641 ();
 sg13g2_decap_8 FILLER_73_2648 ();
 sg13g2_decap_8 FILLER_73_2655 ();
 sg13g2_decap_8 FILLER_73_2662 ();
 sg13g2_decap_8 FILLER_73_2669 ();
 sg13g2_decap_8 FILLER_73_2676 ();
 sg13g2_decap_8 FILLER_73_2683 ();
 sg13g2_decap_8 FILLER_73_2690 ();
 sg13g2_decap_8 FILLER_73_2697 ();
 sg13g2_decap_8 FILLER_73_2704 ();
 sg13g2_decap_8 FILLER_73_2711 ();
 sg13g2_decap_8 FILLER_73_2718 ();
 sg13g2_decap_8 FILLER_73_2725 ();
 sg13g2_decap_8 FILLER_73_2732 ();
 sg13g2_decap_8 FILLER_73_2739 ();
 sg13g2_decap_8 FILLER_73_2746 ();
 sg13g2_decap_8 FILLER_73_2753 ();
 sg13g2_decap_8 FILLER_73_2760 ();
 sg13g2_decap_8 FILLER_73_2767 ();
 sg13g2_decap_8 FILLER_73_2774 ();
 sg13g2_decap_8 FILLER_73_2781 ();
 sg13g2_decap_8 FILLER_73_2788 ();
 sg13g2_decap_8 FILLER_73_2795 ();
 sg13g2_decap_8 FILLER_73_2802 ();
 sg13g2_decap_8 FILLER_73_2809 ();
 sg13g2_decap_8 FILLER_73_2816 ();
 sg13g2_decap_8 FILLER_73_2823 ();
 sg13g2_decap_8 FILLER_73_2830 ();
 sg13g2_decap_8 FILLER_73_2837 ();
 sg13g2_decap_8 FILLER_73_2844 ();
 sg13g2_decap_8 FILLER_73_2851 ();
 sg13g2_decap_8 FILLER_73_2858 ();
 sg13g2_decap_8 FILLER_73_2865 ();
 sg13g2_decap_8 FILLER_73_2872 ();
 sg13g2_decap_8 FILLER_73_2879 ();
 sg13g2_decap_8 FILLER_73_2886 ();
 sg13g2_decap_8 FILLER_73_2893 ();
 sg13g2_decap_8 FILLER_73_2900 ();
 sg13g2_decap_8 FILLER_73_2907 ();
 sg13g2_decap_8 FILLER_73_2914 ();
 sg13g2_decap_8 FILLER_73_2921 ();
 sg13g2_decap_8 FILLER_73_2928 ();
 sg13g2_decap_8 FILLER_73_2935 ();
 sg13g2_decap_8 FILLER_73_2942 ();
 sg13g2_decap_8 FILLER_73_2949 ();
 sg13g2_decap_8 FILLER_73_2956 ();
 sg13g2_decap_8 FILLER_73_2963 ();
 sg13g2_decap_8 FILLER_73_2970 ();
 sg13g2_decap_8 FILLER_73_2977 ();
 sg13g2_decap_8 FILLER_73_2984 ();
 sg13g2_decap_8 FILLER_73_2991 ();
 sg13g2_decap_8 FILLER_73_2998 ();
 sg13g2_decap_8 FILLER_73_3005 ();
 sg13g2_decap_8 FILLER_73_3012 ();
 sg13g2_decap_8 FILLER_73_3019 ();
 sg13g2_decap_8 FILLER_73_3026 ();
 sg13g2_decap_8 FILLER_73_3033 ();
 sg13g2_decap_8 FILLER_73_3040 ();
 sg13g2_decap_8 FILLER_73_3047 ();
 sg13g2_decap_8 FILLER_73_3054 ();
 sg13g2_decap_8 FILLER_73_3061 ();
 sg13g2_decap_8 FILLER_73_3068 ();
 sg13g2_decap_8 FILLER_73_3075 ();
 sg13g2_decap_8 FILLER_73_3082 ();
 sg13g2_decap_8 FILLER_73_3089 ();
 sg13g2_decap_8 FILLER_73_3096 ();
 sg13g2_decap_8 FILLER_73_3103 ();
 sg13g2_decap_8 FILLER_73_3110 ();
 sg13g2_decap_8 FILLER_73_3117 ();
 sg13g2_decap_8 FILLER_73_3124 ();
 sg13g2_decap_8 FILLER_73_3131 ();
 sg13g2_decap_8 FILLER_73_3138 ();
 sg13g2_decap_8 FILLER_73_3145 ();
 sg13g2_decap_8 FILLER_73_3152 ();
 sg13g2_decap_8 FILLER_73_3159 ();
 sg13g2_decap_8 FILLER_73_3166 ();
 sg13g2_decap_8 FILLER_73_3173 ();
 sg13g2_decap_8 FILLER_73_3180 ();
 sg13g2_decap_8 FILLER_73_3187 ();
 sg13g2_decap_8 FILLER_73_3194 ();
 sg13g2_decap_8 FILLER_73_3201 ();
 sg13g2_decap_8 FILLER_73_3208 ();
 sg13g2_decap_8 FILLER_73_3215 ();
 sg13g2_decap_8 FILLER_73_3222 ();
 sg13g2_decap_8 FILLER_73_3229 ();
 sg13g2_decap_8 FILLER_73_3236 ();
 sg13g2_decap_8 FILLER_73_3243 ();
 sg13g2_decap_8 FILLER_73_3250 ();
 sg13g2_decap_8 FILLER_73_3257 ();
 sg13g2_decap_8 FILLER_73_3264 ();
 sg13g2_decap_8 FILLER_73_3271 ();
 sg13g2_decap_8 FILLER_73_3278 ();
 sg13g2_decap_8 FILLER_73_3285 ();
 sg13g2_decap_8 FILLER_73_3292 ();
 sg13g2_decap_8 FILLER_73_3299 ();
 sg13g2_decap_8 FILLER_73_3306 ();
 sg13g2_decap_8 FILLER_73_3313 ();
 sg13g2_decap_8 FILLER_73_3320 ();
 sg13g2_decap_8 FILLER_73_3327 ();
 sg13g2_decap_8 FILLER_73_3334 ();
 sg13g2_decap_8 FILLER_73_3341 ();
 sg13g2_decap_8 FILLER_73_3348 ();
 sg13g2_decap_8 FILLER_73_3355 ();
 sg13g2_decap_8 FILLER_73_3362 ();
 sg13g2_decap_8 FILLER_73_3369 ();
 sg13g2_decap_8 FILLER_73_3376 ();
 sg13g2_decap_8 FILLER_73_3383 ();
 sg13g2_decap_8 FILLER_73_3390 ();
 sg13g2_decap_8 FILLER_73_3397 ();
 sg13g2_decap_8 FILLER_73_3404 ();
 sg13g2_decap_8 FILLER_73_3411 ();
 sg13g2_decap_8 FILLER_73_3418 ();
 sg13g2_decap_8 FILLER_73_3425 ();
 sg13g2_decap_8 FILLER_73_3432 ();
 sg13g2_decap_8 FILLER_73_3439 ();
 sg13g2_decap_8 FILLER_73_3446 ();
 sg13g2_decap_8 FILLER_73_3453 ();
 sg13g2_decap_8 FILLER_73_3460 ();
 sg13g2_decap_8 FILLER_73_3467 ();
 sg13g2_decap_8 FILLER_73_3474 ();
 sg13g2_decap_8 FILLER_73_3481 ();
 sg13g2_decap_8 FILLER_73_3488 ();
 sg13g2_decap_8 FILLER_73_3495 ();
 sg13g2_decap_8 FILLER_73_3502 ();
 sg13g2_decap_8 FILLER_73_3509 ();
 sg13g2_decap_8 FILLER_73_3516 ();
 sg13g2_decap_8 FILLER_73_3523 ();
 sg13g2_decap_8 FILLER_73_3530 ();
 sg13g2_decap_8 FILLER_73_3537 ();
 sg13g2_decap_8 FILLER_73_3544 ();
 sg13g2_decap_8 FILLER_73_3551 ();
 sg13g2_decap_8 FILLER_73_3558 ();
 sg13g2_decap_8 FILLER_73_3565 ();
 sg13g2_decap_8 FILLER_73_3572 ();
 sg13g2_fill_1 FILLER_73_3579 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_8 FILLER_74_252 ();
 sg13g2_decap_8 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_266 ();
 sg13g2_decap_8 FILLER_74_273 ();
 sg13g2_decap_8 FILLER_74_280 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_decap_8 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_decap_8 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_322 ();
 sg13g2_decap_8 FILLER_74_329 ();
 sg13g2_decap_8 FILLER_74_336 ();
 sg13g2_decap_8 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_decap_8 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_decap_8 FILLER_74_406 ();
 sg13g2_decap_8 FILLER_74_413 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_decap_8 FILLER_74_427 ();
 sg13g2_decap_8 FILLER_74_434 ();
 sg13g2_decap_8 FILLER_74_441 ();
 sg13g2_decap_8 FILLER_74_448 ();
 sg13g2_decap_8 FILLER_74_455 ();
 sg13g2_decap_8 FILLER_74_462 ();
 sg13g2_decap_8 FILLER_74_469 ();
 sg13g2_decap_8 FILLER_74_476 ();
 sg13g2_decap_8 FILLER_74_483 ();
 sg13g2_decap_8 FILLER_74_490 ();
 sg13g2_decap_8 FILLER_74_497 ();
 sg13g2_decap_8 FILLER_74_504 ();
 sg13g2_decap_8 FILLER_74_511 ();
 sg13g2_decap_8 FILLER_74_518 ();
 sg13g2_decap_8 FILLER_74_525 ();
 sg13g2_decap_8 FILLER_74_532 ();
 sg13g2_decap_8 FILLER_74_539 ();
 sg13g2_decap_8 FILLER_74_546 ();
 sg13g2_decap_8 FILLER_74_553 ();
 sg13g2_decap_8 FILLER_74_560 ();
 sg13g2_decap_8 FILLER_74_567 ();
 sg13g2_fill_2 FILLER_74_611 ();
 sg13g2_fill_1 FILLER_74_613 ();
 sg13g2_decap_8 FILLER_74_647 ();
 sg13g2_fill_1 FILLER_74_654 ();
 sg13g2_fill_1 FILLER_74_676 ();
 sg13g2_fill_2 FILLER_74_708 ();
 sg13g2_fill_1 FILLER_74_710 ();
 sg13g2_decap_8 FILLER_74_719 ();
 sg13g2_decap_8 FILLER_74_726 ();
 sg13g2_decap_4 FILLER_74_733 ();
 sg13g2_fill_1 FILLER_74_737 ();
 sg13g2_decap_8 FILLER_74_764 ();
 sg13g2_fill_2 FILLER_74_771 ();
 sg13g2_fill_1 FILLER_74_773 ();
 sg13g2_decap_8 FILLER_74_783 ();
 sg13g2_fill_2 FILLER_74_790 ();
 sg13g2_fill_1 FILLER_74_792 ();
 sg13g2_decap_8 FILLER_74_806 ();
 sg13g2_decap_4 FILLER_74_813 ();
 sg13g2_fill_2 FILLER_74_817 ();
 sg13g2_fill_2 FILLER_74_857 ();
 sg13g2_fill_1 FILLER_74_859 ();
 sg13g2_fill_2 FILLER_74_901 ();
 sg13g2_decap_4 FILLER_74_945 ();
 sg13g2_fill_1 FILLER_74_949 ();
 sg13g2_fill_2 FILLER_74_976 ();
 sg13g2_fill_2 FILLER_74_1004 ();
 sg13g2_fill_1 FILLER_74_1006 ();
 sg13g2_decap_8 FILLER_74_1020 ();
 sg13g2_fill_1 FILLER_74_1027 ();
 sg13g2_decap_8 FILLER_74_1059 ();
 sg13g2_decap_8 FILLER_74_1066 ();
 sg13g2_decap_4 FILLER_74_1073 ();
 sg13g2_decap_8 FILLER_74_1113 ();
 sg13g2_decap_8 FILLER_74_1120 ();
 sg13g2_fill_1 FILLER_74_1127 ();
 sg13g2_fill_2 FILLER_74_1195 ();
 sg13g2_fill_1 FILLER_74_1205 ();
 sg13g2_decap_8 FILLER_74_1210 ();
 sg13g2_fill_2 FILLER_74_1222 ();
 sg13g2_decap_4 FILLER_74_1238 ();
 sg13g2_fill_2 FILLER_74_1242 ();
 sg13g2_decap_4 FILLER_74_1252 ();
 sg13g2_decap_8 FILLER_74_1259 ();
 sg13g2_fill_2 FILLER_74_1266 ();
 sg13g2_decap_8 FILLER_74_1276 ();
 sg13g2_decap_4 FILLER_74_1283 ();
 sg13g2_fill_1 FILLER_74_1287 ();
 sg13g2_fill_2 FILLER_74_1343 ();
 sg13g2_fill_1 FILLER_74_1349 ();
 sg13g2_decap_4 FILLER_74_1384 ();
 sg13g2_fill_1 FILLER_74_1388 ();
 sg13g2_fill_1 FILLER_74_1400 ();
 sg13g2_decap_8 FILLER_74_1432 ();
 sg13g2_fill_2 FILLER_74_1439 ();
 sg13g2_decap_8 FILLER_74_1451 ();
 sg13g2_decap_8 FILLER_74_1458 ();
 sg13g2_fill_1 FILLER_74_1465 ();
 sg13g2_decap_4 FILLER_74_1492 ();
 sg13g2_fill_2 FILLER_74_1496 ();
 sg13g2_decap_8 FILLER_74_1553 ();
 sg13g2_decap_4 FILLER_74_1560 ();
 sg13g2_decap_8 FILLER_74_1567 ();
 sg13g2_decap_8 FILLER_74_1574 ();
 sg13g2_decap_8 FILLER_74_1581 ();
 sg13g2_decap_8 FILLER_74_1588 ();
 sg13g2_decap_8 FILLER_74_1595 ();
 sg13g2_decap_8 FILLER_74_1602 ();
 sg13g2_decap_4 FILLER_74_1609 ();
 sg13g2_fill_1 FILLER_74_1613 ();
 sg13g2_fill_2 FILLER_74_1739 ();
 sg13g2_decap_8 FILLER_74_1753 ();
 sg13g2_fill_2 FILLER_74_1760 ();
 sg13g2_fill_1 FILLER_74_1762 ();
 sg13g2_decap_8 FILLER_74_1767 ();
 sg13g2_fill_2 FILLER_74_1774 ();
 sg13g2_decap_8 FILLER_74_1780 ();
 sg13g2_fill_2 FILLER_74_1787 ();
 sg13g2_fill_1 FILLER_74_1789 ();
 sg13g2_decap_4 FILLER_74_1793 ();
 sg13g2_fill_2 FILLER_74_1797 ();
 sg13g2_decap_4 FILLER_74_1809 ();
 sg13g2_decap_8 FILLER_74_1826 ();
 sg13g2_decap_8 FILLER_74_1833 ();
 sg13g2_decap_8 FILLER_74_1840 ();
 sg13g2_decap_8 FILLER_74_1847 ();
 sg13g2_decap_8 FILLER_74_1854 ();
 sg13g2_decap_8 FILLER_74_1861 ();
 sg13g2_decap_8 FILLER_74_1868 ();
 sg13g2_decap_8 FILLER_74_1875 ();
 sg13g2_decap_8 FILLER_74_1882 ();
 sg13g2_decap_8 FILLER_74_1889 ();
 sg13g2_decap_8 FILLER_74_1896 ();
 sg13g2_decap_8 FILLER_74_1903 ();
 sg13g2_decap_8 FILLER_74_1910 ();
 sg13g2_decap_8 FILLER_74_1917 ();
 sg13g2_decap_4 FILLER_74_1929 ();
 sg13g2_decap_8 FILLER_74_1985 ();
 sg13g2_decap_8 FILLER_74_1992 ();
 sg13g2_decap_8 FILLER_74_1999 ();
 sg13g2_fill_2 FILLER_74_2006 ();
 sg13g2_decap_8 FILLER_74_2047 ();
 sg13g2_decap_8 FILLER_74_2054 ();
 sg13g2_decap_8 FILLER_74_2061 ();
 sg13g2_decap_8 FILLER_74_2068 ();
 sg13g2_decap_8 FILLER_74_2075 ();
 sg13g2_fill_2 FILLER_74_2082 ();
 sg13g2_fill_1 FILLER_74_2084 ();
 sg13g2_decap_8 FILLER_74_2137 ();
 sg13g2_decap_8 FILLER_74_2144 ();
 sg13g2_decap_8 FILLER_74_2151 ();
 sg13g2_decap_8 FILLER_74_2158 ();
 sg13g2_decap_8 FILLER_74_2165 ();
 sg13g2_decap_8 FILLER_74_2172 ();
 sg13g2_decap_8 FILLER_74_2179 ();
 sg13g2_decap_8 FILLER_74_2186 ();
 sg13g2_decap_8 FILLER_74_2193 ();
 sg13g2_decap_8 FILLER_74_2200 ();
 sg13g2_decap_8 FILLER_74_2207 ();
 sg13g2_decap_8 FILLER_74_2214 ();
 sg13g2_decap_8 FILLER_74_2221 ();
 sg13g2_decap_8 FILLER_74_2228 ();
 sg13g2_decap_8 FILLER_74_2235 ();
 sg13g2_decap_8 FILLER_74_2242 ();
 sg13g2_decap_8 FILLER_74_2249 ();
 sg13g2_decap_8 FILLER_74_2256 ();
 sg13g2_decap_8 FILLER_74_2263 ();
 sg13g2_decap_8 FILLER_74_2270 ();
 sg13g2_decap_8 FILLER_74_2277 ();
 sg13g2_decap_8 FILLER_74_2284 ();
 sg13g2_decap_8 FILLER_74_2291 ();
 sg13g2_decap_8 FILLER_74_2298 ();
 sg13g2_decap_8 FILLER_74_2305 ();
 sg13g2_decap_8 FILLER_74_2312 ();
 sg13g2_decap_8 FILLER_74_2319 ();
 sg13g2_decap_8 FILLER_74_2326 ();
 sg13g2_decap_8 FILLER_74_2333 ();
 sg13g2_decap_8 FILLER_74_2340 ();
 sg13g2_decap_8 FILLER_74_2347 ();
 sg13g2_decap_8 FILLER_74_2354 ();
 sg13g2_decap_8 FILLER_74_2361 ();
 sg13g2_decap_8 FILLER_74_2368 ();
 sg13g2_decap_8 FILLER_74_2375 ();
 sg13g2_decap_8 FILLER_74_2382 ();
 sg13g2_decap_8 FILLER_74_2389 ();
 sg13g2_decap_8 FILLER_74_2396 ();
 sg13g2_decap_8 FILLER_74_2403 ();
 sg13g2_decap_8 FILLER_74_2410 ();
 sg13g2_decap_8 FILLER_74_2417 ();
 sg13g2_decap_8 FILLER_74_2424 ();
 sg13g2_decap_8 FILLER_74_2431 ();
 sg13g2_decap_8 FILLER_74_2438 ();
 sg13g2_decap_8 FILLER_74_2445 ();
 sg13g2_decap_8 FILLER_74_2452 ();
 sg13g2_decap_8 FILLER_74_2459 ();
 sg13g2_decap_8 FILLER_74_2466 ();
 sg13g2_decap_8 FILLER_74_2473 ();
 sg13g2_decap_8 FILLER_74_2480 ();
 sg13g2_decap_8 FILLER_74_2487 ();
 sg13g2_decap_8 FILLER_74_2494 ();
 sg13g2_decap_8 FILLER_74_2501 ();
 sg13g2_decap_8 FILLER_74_2508 ();
 sg13g2_decap_8 FILLER_74_2515 ();
 sg13g2_decap_8 FILLER_74_2522 ();
 sg13g2_decap_8 FILLER_74_2529 ();
 sg13g2_decap_8 FILLER_74_2536 ();
 sg13g2_decap_8 FILLER_74_2543 ();
 sg13g2_decap_8 FILLER_74_2550 ();
 sg13g2_decap_8 FILLER_74_2557 ();
 sg13g2_decap_8 FILLER_74_2564 ();
 sg13g2_decap_8 FILLER_74_2571 ();
 sg13g2_decap_8 FILLER_74_2578 ();
 sg13g2_decap_8 FILLER_74_2585 ();
 sg13g2_decap_8 FILLER_74_2592 ();
 sg13g2_decap_8 FILLER_74_2599 ();
 sg13g2_decap_8 FILLER_74_2606 ();
 sg13g2_decap_8 FILLER_74_2613 ();
 sg13g2_decap_8 FILLER_74_2620 ();
 sg13g2_decap_8 FILLER_74_2627 ();
 sg13g2_decap_8 FILLER_74_2634 ();
 sg13g2_decap_8 FILLER_74_2641 ();
 sg13g2_decap_8 FILLER_74_2648 ();
 sg13g2_decap_8 FILLER_74_2655 ();
 sg13g2_decap_8 FILLER_74_2662 ();
 sg13g2_decap_8 FILLER_74_2669 ();
 sg13g2_decap_8 FILLER_74_2676 ();
 sg13g2_decap_8 FILLER_74_2683 ();
 sg13g2_decap_8 FILLER_74_2690 ();
 sg13g2_decap_8 FILLER_74_2697 ();
 sg13g2_decap_8 FILLER_74_2704 ();
 sg13g2_decap_8 FILLER_74_2711 ();
 sg13g2_decap_8 FILLER_74_2718 ();
 sg13g2_decap_8 FILLER_74_2725 ();
 sg13g2_decap_8 FILLER_74_2732 ();
 sg13g2_decap_8 FILLER_74_2739 ();
 sg13g2_decap_8 FILLER_74_2746 ();
 sg13g2_decap_8 FILLER_74_2753 ();
 sg13g2_decap_8 FILLER_74_2760 ();
 sg13g2_decap_8 FILLER_74_2767 ();
 sg13g2_decap_8 FILLER_74_2774 ();
 sg13g2_decap_8 FILLER_74_2781 ();
 sg13g2_decap_8 FILLER_74_2788 ();
 sg13g2_decap_8 FILLER_74_2795 ();
 sg13g2_decap_8 FILLER_74_2802 ();
 sg13g2_decap_8 FILLER_74_2809 ();
 sg13g2_decap_8 FILLER_74_2816 ();
 sg13g2_decap_8 FILLER_74_2823 ();
 sg13g2_decap_8 FILLER_74_2830 ();
 sg13g2_decap_8 FILLER_74_2837 ();
 sg13g2_decap_8 FILLER_74_2844 ();
 sg13g2_decap_8 FILLER_74_2851 ();
 sg13g2_decap_8 FILLER_74_2858 ();
 sg13g2_decap_8 FILLER_74_2865 ();
 sg13g2_decap_8 FILLER_74_2872 ();
 sg13g2_decap_8 FILLER_74_2879 ();
 sg13g2_decap_8 FILLER_74_2886 ();
 sg13g2_decap_8 FILLER_74_2893 ();
 sg13g2_decap_8 FILLER_74_2900 ();
 sg13g2_decap_8 FILLER_74_2907 ();
 sg13g2_decap_8 FILLER_74_2914 ();
 sg13g2_decap_8 FILLER_74_2921 ();
 sg13g2_decap_8 FILLER_74_2928 ();
 sg13g2_decap_8 FILLER_74_2935 ();
 sg13g2_decap_8 FILLER_74_2942 ();
 sg13g2_decap_8 FILLER_74_2949 ();
 sg13g2_decap_8 FILLER_74_2956 ();
 sg13g2_decap_8 FILLER_74_2963 ();
 sg13g2_decap_8 FILLER_74_2970 ();
 sg13g2_decap_8 FILLER_74_2977 ();
 sg13g2_decap_8 FILLER_74_2984 ();
 sg13g2_decap_8 FILLER_74_2991 ();
 sg13g2_decap_8 FILLER_74_2998 ();
 sg13g2_decap_8 FILLER_74_3005 ();
 sg13g2_decap_8 FILLER_74_3012 ();
 sg13g2_decap_8 FILLER_74_3019 ();
 sg13g2_decap_8 FILLER_74_3026 ();
 sg13g2_decap_8 FILLER_74_3033 ();
 sg13g2_decap_8 FILLER_74_3040 ();
 sg13g2_decap_8 FILLER_74_3047 ();
 sg13g2_decap_8 FILLER_74_3054 ();
 sg13g2_decap_8 FILLER_74_3061 ();
 sg13g2_decap_8 FILLER_74_3068 ();
 sg13g2_decap_8 FILLER_74_3075 ();
 sg13g2_decap_8 FILLER_74_3082 ();
 sg13g2_decap_8 FILLER_74_3089 ();
 sg13g2_decap_8 FILLER_74_3096 ();
 sg13g2_decap_8 FILLER_74_3103 ();
 sg13g2_decap_8 FILLER_74_3110 ();
 sg13g2_decap_8 FILLER_74_3117 ();
 sg13g2_decap_8 FILLER_74_3124 ();
 sg13g2_decap_8 FILLER_74_3131 ();
 sg13g2_decap_8 FILLER_74_3138 ();
 sg13g2_decap_8 FILLER_74_3145 ();
 sg13g2_decap_8 FILLER_74_3152 ();
 sg13g2_decap_8 FILLER_74_3159 ();
 sg13g2_decap_8 FILLER_74_3166 ();
 sg13g2_decap_8 FILLER_74_3173 ();
 sg13g2_decap_8 FILLER_74_3180 ();
 sg13g2_decap_8 FILLER_74_3187 ();
 sg13g2_decap_8 FILLER_74_3194 ();
 sg13g2_decap_8 FILLER_74_3201 ();
 sg13g2_decap_8 FILLER_74_3208 ();
 sg13g2_decap_8 FILLER_74_3215 ();
 sg13g2_decap_8 FILLER_74_3222 ();
 sg13g2_decap_8 FILLER_74_3229 ();
 sg13g2_decap_8 FILLER_74_3236 ();
 sg13g2_decap_8 FILLER_74_3243 ();
 sg13g2_decap_8 FILLER_74_3250 ();
 sg13g2_decap_8 FILLER_74_3257 ();
 sg13g2_decap_8 FILLER_74_3264 ();
 sg13g2_decap_8 FILLER_74_3271 ();
 sg13g2_decap_8 FILLER_74_3278 ();
 sg13g2_decap_8 FILLER_74_3285 ();
 sg13g2_decap_8 FILLER_74_3292 ();
 sg13g2_decap_8 FILLER_74_3299 ();
 sg13g2_decap_8 FILLER_74_3306 ();
 sg13g2_decap_8 FILLER_74_3313 ();
 sg13g2_decap_8 FILLER_74_3320 ();
 sg13g2_decap_8 FILLER_74_3327 ();
 sg13g2_decap_8 FILLER_74_3334 ();
 sg13g2_decap_8 FILLER_74_3341 ();
 sg13g2_decap_8 FILLER_74_3348 ();
 sg13g2_decap_8 FILLER_74_3355 ();
 sg13g2_decap_8 FILLER_74_3362 ();
 sg13g2_decap_8 FILLER_74_3369 ();
 sg13g2_decap_8 FILLER_74_3376 ();
 sg13g2_decap_8 FILLER_74_3383 ();
 sg13g2_decap_8 FILLER_74_3390 ();
 sg13g2_decap_8 FILLER_74_3397 ();
 sg13g2_decap_8 FILLER_74_3404 ();
 sg13g2_decap_8 FILLER_74_3411 ();
 sg13g2_decap_8 FILLER_74_3418 ();
 sg13g2_decap_8 FILLER_74_3425 ();
 sg13g2_decap_8 FILLER_74_3432 ();
 sg13g2_decap_8 FILLER_74_3439 ();
 sg13g2_decap_8 FILLER_74_3446 ();
 sg13g2_decap_8 FILLER_74_3453 ();
 sg13g2_decap_8 FILLER_74_3460 ();
 sg13g2_decap_8 FILLER_74_3467 ();
 sg13g2_decap_8 FILLER_74_3474 ();
 sg13g2_decap_8 FILLER_74_3481 ();
 sg13g2_decap_8 FILLER_74_3488 ();
 sg13g2_decap_8 FILLER_74_3495 ();
 sg13g2_decap_8 FILLER_74_3502 ();
 sg13g2_decap_8 FILLER_74_3509 ();
 sg13g2_decap_8 FILLER_74_3516 ();
 sg13g2_decap_8 FILLER_74_3523 ();
 sg13g2_decap_8 FILLER_74_3530 ();
 sg13g2_decap_8 FILLER_74_3537 ();
 sg13g2_decap_8 FILLER_74_3544 ();
 sg13g2_decap_8 FILLER_74_3551 ();
 sg13g2_decap_8 FILLER_74_3558 ();
 sg13g2_decap_8 FILLER_74_3565 ();
 sg13g2_decap_8 FILLER_74_3572 ();
 sg13g2_fill_1 FILLER_74_3579 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_329 ();
 sg13g2_decap_8 FILLER_75_336 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_350 ();
 sg13g2_decap_8 FILLER_75_357 ();
 sg13g2_decap_8 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_378 ();
 sg13g2_decap_8 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_decap_8 FILLER_75_406 ();
 sg13g2_decap_8 FILLER_75_413 ();
 sg13g2_decap_8 FILLER_75_420 ();
 sg13g2_decap_8 FILLER_75_427 ();
 sg13g2_decap_8 FILLER_75_434 ();
 sg13g2_decap_8 FILLER_75_441 ();
 sg13g2_decap_8 FILLER_75_448 ();
 sg13g2_decap_8 FILLER_75_455 ();
 sg13g2_decap_8 FILLER_75_462 ();
 sg13g2_decap_8 FILLER_75_469 ();
 sg13g2_decap_8 FILLER_75_476 ();
 sg13g2_decap_8 FILLER_75_483 ();
 sg13g2_decap_8 FILLER_75_490 ();
 sg13g2_decap_8 FILLER_75_497 ();
 sg13g2_decap_8 FILLER_75_504 ();
 sg13g2_decap_8 FILLER_75_511 ();
 sg13g2_decap_8 FILLER_75_518 ();
 sg13g2_decap_8 FILLER_75_525 ();
 sg13g2_decap_8 FILLER_75_532 ();
 sg13g2_decap_8 FILLER_75_539 ();
 sg13g2_decap_8 FILLER_75_546 ();
 sg13g2_decap_8 FILLER_75_553 ();
 sg13g2_decap_8 FILLER_75_560 ();
 sg13g2_decap_8 FILLER_75_567 ();
 sg13g2_decap_4 FILLER_75_574 ();
 sg13g2_fill_2 FILLER_75_578 ();
 sg13g2_fill_2 FILLER_75_635 ();
 sg13g2_decap_4 FILLER_75_671 ();
 sg13g2_fill_1 FILLER_75_685 ();
 sg13g2_fill_2 FILLER_75_694 ();
 sg13g2_decap_4 FILLER_75_734 ();
 sg13g2_fill_2 FILLER_75_743 ();
 sg13g2_fill_1 FILLER_75_745 ();
 sg13g2_fill_2 FILLER_75_750 ();
 sg13g2_decap_8 FILLER_75_757 ();
 sg13g2_decap_8 FILLER_75_764 ();
 sg13g2_decap_8 FILLER_75_771 ();
 sg13g2_decap_8 FILLER_75_809 ();
 sg13g2_decap_8 FILLER_75_816 ();
 sg13g2_decap_4 FILLER_75_823 ();
 sg13g2_fill_1 FILLER_75_827 ();
 sg13g2_decap_8 FILLER_75_854 ();
 sg13g2_decap_8 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_fill_1 FILLER_75_875 ();
 sg13g2_decap_8 FILLER_75_888 ();
 sg13g2_decap_8 FILLER_75_895 ();
 sg13g2_decap_8 FILLER_75_902 ();
 sg13g2_decap_4 FILLER_75_909 ();
 sg13g2_fill_2 FILLER_75_913 ();
 sg13g2_fill_1 FILLER_75_919 ();
 sg13g2_decap_8 FILLER_75_933 ();
 sg13g2_decap_8 FILLER_75_940 ();
 sg13g2_decap_8 FILLER_75_947 ();
 sg13g2_fill_2 FILLER_75_954 ();
 sg13g2_fill_1 FILLER_75_956 ();
 sg13g2_fill_1 FILLER_75_983 ();
 sg13g2_decap_8 FILLER_75_994 ();
 sg13g2_decap_4 FILLER_75_1001 ();
 sg13g2_fill_2 FILLER_75_1005 ();
 sg13g2_fill_2 FILLER_75_1015 ();
 sg13g2_fill_1 FILLER_75_1017 ();
 sg13g2_fill_1 FILLER_75_1039 ();
 sg13g2_decap_8 FILLER_75_1066 ();
 sg13g2_decap_8 FILLER_75_1073 ();
 sg13g2_fill_2 FILLER_75_1106 ();
 sg13g2_decap_4 FILLER_75_1121 ();
 sg13g2_decap_4 FILLER_75_1164 ();
 sg13g2_fill_2 FILLER_75_1173 ();
 sg13g2_fill_2 FILLER_75_1183 ();
 sg13g2_decap_8 FILLER_75_1215 ();
 sg13g2_fill_1 FILLER_75_1222 ();
 sg13g2_fill_2 FILLER_75_1249 ();
 sg13g2_decap_8 FILLER_75_1266 ();
 sg13g2_fill_2 FILLER_75_1273 ();
 sg13g2_fill_1 FILLER_75_1275 ();
 sg13g2_decap_4 FILLER_75_1302 ();
 sg13g2_fill_1 FILLER_75_1311 ();
 sg13g2_decap_4 FILLER_75_1321 ();
 sg13g2_fill_1 FILLER_75_1325 ();
 sg13g2_decap_8 FILLER_75_1360 ();
 sg13g2_fill_2 FILLER_75_1367 ();
 sg13g2_decap_8 FILLER_75_1373 ();
 sg13g2_decap_4 FILLER_75_1380 ();
 sg13g2_fill_2 FILLER_75_1384 ();
 sg13g2_fill_1 FILLER_75_1391 ();
 sg13g2_fill_2 FILLER_75_1395 ();
 sg13g2_fill_2 FILLER_75_1406 ();
 sg13g2_fill_1 FILLER_75_1408 ();
 sg13g2_decap_8 FILLER_75_1417 ();
 sg13g2_decap_8 FILLER_75_1424 ();
 sg13g2_decap_8 FILLER_75_1435 ();
 sg13g2_decap_8 FILLER_75_1442 ();
 sg13g2_fill_2 FILLER_75_1449 ();
 sg13g2_fill_2 FILLER_75_1464 ();
 sg13g2_fill_1 FILLER_75_1466 ();
 sg13g2_decap_8 FILLER_75_1493 ();
 sg13g2_decap_4 FILLER_75_1500 ();
 sg13g2_decap_8 FILLER_75_1545 ();
 sg13g2_decap_8 FILLER_75_1552 ();
 sg13g2_decap_8 FILLER_75_1559 ();
 sg13g2_decap_8 FILLER_75_1566 ();
 sg13g2_decap_8 FILLER_75_1573 ();
 sg13g2_decap_8 FILLER_75_1580 ();
 sg13g2_decap_8 FILLER_75_1587 ();
 sg13g2_decap_8 FILLER_75_1594 ();
 sg13g2_decap_8 FILLER_75_1601 ();
 sg13g2_decap_8 FILLER_75_1608 ();
 sg13g2_decap_4 FILLER_75_1615 ();
 sg13g2_fill_2 FILLER_75_1626 ();
 sg13g2_fill_1 FILLER_75_1628 ();
 sg13g2_decap_8 FILLER_75_1633 ();
 sg13g2_decap_8 FILLER_75_1640 ();
 sg13g2_fill_2 FILLER_75_1647 ();
 sg13g2_fill_1 FILLER_75_1649 ();
 sg13g2_fill_2 FILLER_75_1654 ();
 sg13g2_decap_8 FILLER_75_1682 ();
 sg13g2_fill_2 FILLER_75_1693 ();
 sg13g2_decap_4 FILLER_75_1700 ();
 sg13g2_fill_2 FILLER_75_1704 ();
 sg13g2_decap_8 FILLER_75_1744 ();
 sg13g2_decap_8 FILLER_75_1751 ();
 sg13g2_decap_4 FILLER_75_1758 ();
 sg13g2_fill_1 FILLER_75_1762 ();
 sg13g2_decap_8 FILLER_75_1820 ();
 sg13g2_decap_8 FILLER_75_1827 ();
 sg13g2_decap_8 FILLER_75_1834 ();
 sg13g2_decap_8 FILLER_75_1841 ();
 sg13g2_decap_8 FILLER_75_1848 ();
 sg13g2_decap_8 FILLER_75_1855 ();
 sg13g2_decap_8 FILLER_75_1862 ();
 sg13g2_decap_8 FILLER_75_1869 ();
 sg13g2_decap_8 FILLER_75_1876 ();
 sg13g2_decap_8 FILLER_75_1883 ();
 sg13g2_decap_8 FILLER_75_1890 ();
 sg13g2_decap_8 FILLER_75_1897 ();
 sg13g2_decap_8 FILLER_75_1904 ();
 sg13g2_decap_8 FILLER_75_1911 ();
 sg13g2_decap_8 FILLER_75_1918 ();
 sg13g2_decap_4 FILLER_75_1925 ();
 sg13g2_fill_1 FILLER_75_1929 ();
 sg13g2_fill_1 FILLER_75_1956 ();
 sg13g2_decap_8 FILLER_75_1983 ();
 sg13g2_decap_8 FILLER_75_1990 ();
 sg13g2_decap_8 FILLER_75_1997 ();
 sg13g2_decap_8 FILLER_75_2004 ();
 sg13g2_fill_1 FILLER_75_2011 ();
 sg13g2_decap_8 FILLER_75_2064 ();
 sg13g2_decap_8 FILLER_75_2071 ();
 sg13g2_decap_8 FILLER_75_2078 ();
 sg13g2_decap_8 FILLER_75_2085 ();
 sg13g2_fill_1 FILLER_75_2092 ();
 sg13g2_decap_8 FILLER_75_2119 ();
 sg13g2_decap_8 FILLER_75_2126 ();
 sg13g2_decap_8 FILLER_75_2133 ();
 sg13g2_decap_8 FILLER_75_2140 ();
 sg13g2_decap_8 FILLER_75_2147 ();
 sg13g2_decap_8 FILLER_75_2154 ();
 sg13g2_decap_8 FILLER_75_2161 ();
 sg13g2_decap_8 FILLER_75_2168 ();
 sg13g2_decap_8 FILLER_75_2175 ();
 sg13g2_decap_8 FILLER_75_2182 ();
 sg13g2_decap_8 FILLER_75_2189 ();
 sg13g2_decap_8 FILLER_75_2196 ();
 sg13g2_decap_8 FILLER_75_2203 ();
 sg13g2_decap_8 FILLER_75_2210 ();
 sg13g2_decap_8 FILLER_75_2217 ();
 sg13g2_decap_8 FILLER_75_2224 ();
 sg13g2_decap_8 FILLER_75_2231 ();
 sg13g2_decap_8 FILLER_75_2238 ();
 sg13g2_decap_8 FILLER_75_2245 ();
 sg13g2_decap_8 FILLER_75_2252 ();
 sg13g2_decap_8 FILLER_75_2259 ();
 sg13g2_decap_8 FILLER_75_2266 ();
 sg13g2_decap_8 FILLER_75_2273 ();
 sg13g2_decap_8 FILLER_75_2280 ();
 sg13g2_decap_8 FILLER_75_2287 ();
 sg13g2_decap_8 FILLER_75_2294 ();
 sg13g2_decap_8 FILLER_75_2301 ();
 sg13g2_decap_8 FILLER_75_2308 ();
 sg13g2_decap_8 FILLER_75_2315 ();
 sg13g2_decap_8 FILLER_75_2322 ();
 sg13g2_decap_8 FILLER_75_2329 ();
 sg13g2_decap_8 FILLER_75_2336 ();
 sg13g2_decap_8 FILLER_75_2343 ();
 sg13g2_decap_8 FILLER_75_2350 ();
 sg13g2_decap_8 FILLER_75_2357 ();
 sg13g2_decap_8 FILLER_75_2364 ();
 sg13g2_decap_8 FILLER_75_2371 ();
 sg13g2_decap_8 FILLER_75_2378 ();
 sg13g2_decap_8 FILLER_75_2385 ();
 sg13g2_decap_8 FILLER_75_2392 ();
 sg13g2_decap_8 FILLER_75_2399 ();
 sg13g2_decap_8 FILLER_75_2406 ();
 sg13g2_decap_8 FILLER_75_2413 ();
 sg13g2_decap_8 FILLER_75_2420 ();
 sg13g2_decap_8 FILLER_75_2427 ();
 sg13g2_decap_8 FILLER_75_2434 ();
 sg13g2_decap_8 FILLER_75_2441 ();
 sg13g2_decap_8 FILLER_75_2448 ();
 sg13g2_decap_8 FILLER_75_2455 ();
 sg13g2_decap_8 FILLER_75_2462 ();
 sg13g2_decap_8 FILLER_75_2469 ();
 sg13g2_decap_8 FILLER_75_2476 ();
 sg13g2_decap_8 FILLER_75_2483 ();
 sg13g2_decap_8 FILLER_75_2490 ();
 sg13g2_decap_8 FILLER_75_2497 ();
 sg13g2_decap_8 FILLER_75_2504 ();
 sg13g2_decap_8 FILLER_75_2511 ();
 sg13g2_decap_8 FILLER_75_2518 ();
 sg13g2_decap_8 FILLER_75_2525 ();
 sg13g2_decap_8 FILLER_75_2532 ();
 sg13g2_decap_8 FILLER_75_2539 ();
 sg13g2_decap_8 FILLER_75_2546 ();
 sg13g2_decap_8 FILLER_75_2553 ();
 sg13g2_decap_8 FILLER_75_2560 ();
 sg13g2_decap_8 FILLER_75_2567 ();
 sg13g2_decap_8 FILLER_75_2574 ();
 sg13g2_decap_8 FILLER_75_2581 ();
 sg13g2_decap_8 FILLER_75_2588 ();
 sg13g2_decap_8 FILLER_75_2595 ();
 sg13g2_decap_8 FILLER_75_2602 ();
 sg13g2_decap_8 FILLER_75_2609 ();
 sg13g2_decap_8 FILLER_75_2616 ();
 sg13g2_decap_8 FILLER_75_2623 ();
 sg13g2_decap_8 FILLER_75_2630 ();
 sg13g2_decap_8 FILLER_75_2637 ();
 sg13g2_decap_8 FILLER_75_2644 ();
 sg13g2_decap_8 FILLER_75_2651 ();
 sg13g2_decap_8 FILLER_75_2658 ();
 sg13g2_decap_8 FILLER_75_2665 ();
 sg13g2_decap_8 FILLER_75_2672 ();
 sg13g2_decap_8 FILLER_75_2679 ();
 sg13g2_decap_8 FILLER_75_2686 ();
 sg13g2_decap_8 FILLER_75_2693 ();
 sg13g2_decap_8 FILLER_75_2700 ();
 sg13g2_decap_8 FILLER_75_2707 ();
 sg13g2_decap_8 FILLER_75_2714 ();
 sg13g2_decap_8 FILLER_75_2721 ();
 sg13g2_decap_8 FILLER_75_2728 ();
 sg13g2_decap_8 FILLER_75_2735 ();
 sg13g2_decap_8 FILLER_75_2742 ();
 sg13g2_decap_8 FILLER_75_2749 ();
 sg13g2_decap_8 FILLER_75_2756 ();
 sg13g2_decap_8 FILLER_75_2763 ();
 sg13g2_decap_8 FILLER_75_2770 ();
 sg13g2_decap_8 FILLER_75_2777 ();
 sg13g2_decap_8 FILLER_75_2784 ();
 sg13g2_decap_8 FILLER_75_2791 ();
 sg13g2_decap_8 FILLER_75_2798 ();
 sg13g2_decap_8 FILLER_75_2805 ();
 sg13g2_decap_8 FILLER_75_2812 ();
 sg13g2_decap_8 FILLER_75_2819 ();
 sg13g2_decap_8 FILLER_75_2826 ();
 sg13g2_decap_8 FILLER_75_2833 ();
 sg13g2_decap_8 FILLER_75_2840 ();
 sg13g2_decap_8 FILLER_75_2847 ();
 sg13g2_decap_8 FILLER_75_2854 ();
 sg13g2_decap_8 FILLER_75_2861 ();
 sg13g2_decap_8 FILLER_75_2868 ();
 sg13g2_decap_8 FILLER_75_2875 ();
 sg13g2_decap_8 FILLER_75_2882 ();
 sg13g2_decap_8 FILLER_75_2889 ();
 sg13g2_decap_8 FILLER_75_2896 ();
 sg13g2_decap_8 FILLER_75_2903 ();
 sg13g2_decap_8 FILLER_75_2910 ();
 sg13g2_decap_8 FILLER_75_2917 ();
 sg13g2_decap_8 FILLER_75_2924 ();
 sg13g2_decap_8 FILLER_75_2931 ();
 sg13g2_decap_8 FILLER_75_2938 ();
 sg13g2_decap_8 FILLER_75_2945 ();
 sg13g2_decap_8 FILLER_75_2952 ();
 sg13g2_decap_8 FILLER_75_2959 ();
 sg13g2_decap_8 FILLER_75_2966 ();
 sg13g2_decap_8 FILLER_75_2973 ();
 sg13g2_decap_8 FILLER_75_2980 ();
 sg13g2_decap_8 FILLER_75_2987 ();
 sg13g2_decap_8 FILLER_75_2994 ();
 sg13g2_decap_8 FILLER_75_3001 ();
 sg13g2_decap_8 FILLER_75_3008 ();
 sg13g2_decap_8 FILLER_75_3015 ();
 sg13g2_decap_8 FILLER_75_3022 ();
 sg13g2_decap_8 FILLER_75_3029 ();
 sg13g2_decap_8 FILLER_75_3036 ();
 sg13g2_decap_8 FILLER_75_3043 ();
 sg13g2_decap_8 FILLER_75_3050 ();
 sg13g2_decap_8 FILLER_75_3057 ();
 sg13g2_decap_8 FILLER_75_3064 ();
 sg13g2_decap_8 FILLER_75_3071 ();
 sg13g2_decap_8 FILLER_75_3078 ();
 sg13g2_decap_8 FILLER_75_3085 ();
 sg13g2_decap_8 FILLER_75_3092 ();
 sg13g2_decap_8 FILLER_75_3099 ();
 sg13g2_decap_8 FILLER_75_3106 ();
 sg13g2_decap_8 FILLER_75_3113 ();
 sg13g2_decap_8 FILLER_75_3120 ();
 sg13g2_decap_8 FILLER_75_3127 ();
 sg13g2_decap_8 FILLER_75_3134 ();
 sg13g2_decap_8 FILLER_75_3141 ();
 sg13g2_decap_8 FILLER_75_3148 ();
 sg13g2_decap_8 FILLER_75_3155 ();
 sg13g2_decap_8 FILLER_75_3162 ();
 sg13g2_decap_8 FILLER_75_3169 ();
 sg13g2_decap_8 FILLER_75_3176 ();
 sg13g2_decap_8 FILLER_75_3183 ();
 sg13g2_decap_8 FILLER_75_3190 ();
 sg13g2_decap_8 FILLER_75_3197 ();
 sg13g2_decap_8 FILLER_75_3204 ();
 sg13g2_decap_8 FILLER_75_3211 ();
 sg13g2_decap_8 FILLER_75_3218 ();
 sg13g2_decap_8 FILLER_75_3225 ();
 sg13g2_decap_8 FILLER_75_3232 ();
 sg13g2_decap_8 FILLER_75_3239 ();
 sg13g2_decap_8 FILLER_75_3246 ();
 sg13g2_decap_8 FILLER_75_3253 ();
 sg13g2_decap_8 FILLER_75_3260 ();
 sg13g2_decap_8 FILLER_75_3267 ();
 sg13g2_decap_8 FILLER_75_3274 ();
 sg13g2_decap_8 FILLER_75_3281 ();
 sg13g2_decap_8 FILLER_75_3288 ();
 sg13g2_decap_8 FILLER_75_3295 ();
 sg13g2_decap_8 FILLER_75_3302 ();
 sg13g2_decap_8 FILLER_75_3309 ();
 sg13g2_decap_8 FILLER_75_3316 ();
 sg13g2_decap_8 FILLER_75_3323 ();
 sg13g2_decap_8 FILLER_75_3330 ();
 sg13g2_decap_8 FILLER_75_3337 ();
 sg13g2_decap_8 FILLER_75_3344 ();
 sg13g2_decap_8 FILLER_75_3351 ();
 sg13g2_decap_8 FILLER_75_3358 ();
 sg13g2_decap_8 FILLER_75_3365 ();
 sg13g2_decap_8 FILLER_75_3372 ();
 sg13g2_decap_8 FILLER_75_3379 ();
 sg13g2_decap_8 FILLER_75_3386 ();
 sg13g2_decap_8 FILLER_75_3393 ();
 sg13g2_decap_8 FILLER_75_3400 ();
 sg13g2_decap_8 FILLER_75_3407 ();
 sg13g2_decap_8 FILLER_75_3414 ();
 sg13g2_decap_8 FILLER_75_3421 ();
 sg13g2_decap_8 FILLER_75_3428 ();
 sg13g2_decap_8 FILLER_75_3435 ();
 sg13g2_decap_8 FILLER_75_3442 ();
 sg13g2_decap_8 FILLER_75_3449 ();
 sg13g2_decap_8 FILLER_75_3456 ();
 sg13g2_decap_8 FILLER_75_3463 ();
 sg13g2_decap_8 FILLER_75_3470 ();
 sg13g2_decap_8 FILLER_75_3477 ();
 sg13g2_decap_8 FILLER_75_3484 ();
 sg13g2_decap_8 FILLER_75_3491 ();
 sg13g2_decap_8 FILLER_75_3498 ();
 sg13g2_decap_8 FILLER_75_3505 ();
 sg13g2_decap_8 FILLER_75_3512 ();
 sg13g2_decap_8 FILLER_75_3519 ();
 sg13g2_decap_8 FILLER_75_3526 ();
 sg13g2_decap_8 FILLER_75_3533 ();
 sg13g2_decap_8 FILLER_75_3540 ();
 sg13g2_decap_8 FILLER_75_3547 ();
 sg13g2_decap_8 FILLER_75_3554 ();
 sg13g2_decap_8 FILLER_75_3561 ();
 sg13g2_decap_8 FILLER_75_3568 ();
 sg13g2_decap_4 FILLER_75_3575 ();
 sg13g2_fill_1 FILLER_75_3579 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_413 ();
 sg13g2_decap_8 FILLER_76_420 ();
 sg13g2_decap_8 FILLER_76_427 ();
 sg13g2_decap_8 FILLER_76_434 ();
 sg13g2_decap_8 FILLER_76_441 ();
 sg13g2_decap_8 FILLER_76_448 ();
 sg13g2_decap_8 FILLER_76_455 ();
 sg13g2_decap_8 FILLER_76_462 ();
 sg13g2_decap_8 FILLER_76_469 ();
 sg13g2_decap_8 FILLER_76_476 ();
 sg13g2_decap_8 FILLER_76_483 ();
 sg13g2_decap_8 FILLER_76_490 ();
 sg13g2_decap_8 FILLER_76_497 ();
 sg13g2_decap_8 FILLER_76_504 ();
 sg13g2_decap_8 FILLER_76_511 ();
 sg13g2_decap_8 FILLER_76_518 ();
 sg13g2_decap_8 FILLER_76_525 ();
 sg13g2_decap_8 FILLER_76_532 ();
 sg13g2_decap_8 FILLER_76_539 ();
 sg13g2_decap_8 FILLER_76_546 ();
 sg13g2_decap_8 FILLER_76_553 ();
 sg13g2_decap_8 FILLER_76_560 ();
 sg13g2_decap_8 FILLER_76_567 ();
 sg13g2_decap_8 FILLER_76_574 ();
 sg13g2_decap_8 FILLER_76_581 ();
 sg13g2_fill_1 FILLER_76_588 ();
 sg13g2_decap_8 FILLER_76_613 ();
 sg13g2_decap_8 FILLER_76_620 ();
 sg13g2_decap_8 FILLER_76_627 ();
 sg13g2_decap_8 FILLER_76_634 ();
 sg13g2_decap_8 FILLER_76_641 ();
 sg13g2_decap_8 FILLER_76_648 ();
 sg13g2_fill_2 FILLER_76_655 ();
 sg13g2_fill_2 FILLER_76_701 ();
 sg13g2_fill_2 FILLER_76_716 ();
 sg13g2_decap_8 FILLER_76_770 ();
 sg13g2_decap_8 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_784 ();
 sg13g2_fill_1 FILLER_76_791 ();
 sg13g2_decap_4 FILLER_76_864 ();
 sg13g2_fill_1 FILLER_76_868 ();
 sg13g2_fill_2 FILLER_76_882 ();
 sg13g2_decap_8 FILLER_76_892 ();
 sg13g2_decap_8 FILLER_76_899 ();
 sg13g2_fill_2 FILLER_76_906 ();
 sg13g2_fill_1 FILLER_76_908 ();
 sg13g2_decap_8 FILLER_76_935 ();
 sg13g2_decap_8 FILLER_76_942 ();
 sg13g2_decap_8 FILLER_76_949 ();
 sg13g2_decap_4 FILLER_76_956 ();
 sg13g2_fill_2 FILLER_76_976 ();
 sg13g2_fill_1 FILLER_76_978 ();
 sg13g2_decap_8 FILLER_76_1000 ();
 sg13g2_decap_8 FILLER_76_1007 ();
 sg13g2_decap_4 FILLER_76_1014 ();
 sg13g2_fill_1 FILLER_76_1018 ();
 sg13g2_fill_1 FILLER_76_1034 ();
 sg13g2_decap_8 FILLER_76_1069 ();
 sg13g2_decap_8 FILLER_76_1076 ();
 sg13g2_fill_1 FILLER_76_1083 ();
 sg13g2_fill_2 FILLER_76_1122 ();
 sg13g2_fill_1 FILLER_76_1124 ();
 sg13g2_decap_8 FILLER_76_1175 ();
 sg13g2_decap_4 FILLER_76_1182 ();
 sg13g2_fill_2 FILLER_76_1186 ();
 sg13g2_decap_8 FILLER_76_1214 ();
 sg13g2_decap_8 FILLER_76_1221 ();
 sg13g2_decap_4 FILLER_76_1228 ();
 sg13g2_fill_1 FILLER_76_1232 ();
 sg13g2_decap_8 FILLER_76_1275 ();
 sg13g2_decap_4 FILLER_76_1282 ();
 sg13g2_fill_1 FILLER_76_1286 ();
 sg13g2_decap_8 FILLER_76_1296 ();
 sg13g2_fill_2 FILLER_76_1303 ();
 sg13g2_fill_1 FILLER_76_1305 ();
 sg13g2_decap_8 FILLER_76_1309 ();
 sg13g2_decap_8 FILLER_76_1316 ();
 sg13g2_decap_8 FILLER_76_1323 ();
 sg13g2_decap_8 FILLER_76_1330 ();
 sg13g2_decap_8 FILLER_76_1340 ();
 sg13g2_decap_8 FILLER_76_1347 ();
 sg13g2_decap_8 FILLER_76_1354 ();
 sg13g2_decap_8 FILLER_76_1361 ();
 sg13g2_decap_8 FILLER_76_1368 ();
 sg13g2_fill_1 FILLER_76_1375 ();
 sg13g2_decap_4 FILLER_76_1381 ();
 sg13g2_fill_2 FILLER_76_1393 ();
 sg13g2_fill_1 FILLER_76_1403 ();
 sg13g2_decap_4 FILLER_76_1412 ();
 sg13g2_fill_1 FILLER_76_1416 ();
 sg13g2_decap_8 FILLER_76_1462 ();
 sg13g2_fill_2 FILLER_76_1469 ();
 sg13g2_fill_1 FILLER_76_1471 ();
 sg13g2_fill_1 FILLER_76_1476 ();
 sg13g2_decap_8 FILLER_76_1485 ();
 sg13g2_decap_8 FILLER_76_1492 ();
 sg13g2_decap_8 FILLER_76_1499 ();
 sg13g2_decap_4 FILLER_76_1506 ();
 sg13g2_decap_8 FILLER_76_1539 ();
 sg13g2_decap_8 FILLER_76_1546 ();
 sg13g2_decap_8 FILLER_76_1553 ();
 sg13g2_decap_8 FILLER_76_1560 ();
 sg13g2_decap_8 FILLER_76_1567 ();
 sg13g2_decap_8 FILLER_76_1574 ();
 sg13g2_decap_8 FILLER_76_1581 ();
 sg13g2_decap_8 FILLER_76_1588 ();
 sg13g2_decap_8 FILLER_76_1595 ();
 sg13g2_decap_8 FILLER_76_1602 ();
 sg13g2_decap_8 FILLER_76_1609 ();
 sg13g2_decap_8 FILLER_76_1616 ();
 sg13g2_decap_8 FILLER_76_1623 ();
 sg13g2_decap_8 FILLER_76_1630 ();
 sg13g2_decap_8 FILLER_76_1637 ();
 sg13g2_decap_8 FILLER_76_1644 ();
 sg13g2_decap_4 FILLER_76_1651 ();
 sg13g2_fill_2 FILLER_76_1655 ();
 sg13g2_decap_4 FILLER_76_1660 ();
 sg13g2_fill_2 FILLER_76_1664 ();
 sg13g2_decap_8 FILLER_76_1670 ();
 sg13g2_decap_8 FILLER_76_1677 ();
 sg13g2_decap_8 FILLER_76_1684 ();
 sg13g2_decap_8 FILLER_76_1691 ();
 sg13g2_decap_8 FILLER_76_1698 ();
 sg13g2_decap_4 FILLER_76_1705 ();
 sg13g2_fill_2 FILLER_76_1709 ();
 sg13g2_decap_8 FILLER_76_1715 ();
 sg13g2_fill_2 FILLER_76_1722 ();
 sg13g2_decap_8 FILLER_76_1728 ();
 sg13g2_decap_8 FILLER_76_1735 ();
 sg13g2_decap_8 FILLER_76_1742 ();
 sg13g2_decap_8 FILLER_76_1749 ();
 sg13g2_decap_8 FILLER_76_1756 ();
 sg13g2_decap_8 FILLER_76_1763 ();
 sg13g2_decap_8 FILLER_76_1770 ();
 sg13g2_decap_8 FILLER_76_1777 ();
 sg13g2_decap_8 FILLER_76_1784 ();
 sg13g2_decap_8 FILLER_76_1791 ();
 sg13g2_fill_2 FILLER_76_1798 ();
 sg13g2_decap_8 FILLER_76_1804 ();
 sg13g2_decap_8 FILLER_76_1811 ();
 sg13g2_decap_8 FILLER_76_1818 ();
 sg13g2_decap_8 FILLER_76_1825 ();
 sg13g2_decap_8 FILLER_76_1832 ();
 sg13g2_decap_8 FILLER_76_1839 ();
 sg13g2_decap_8 FILLER_76_1846 ();
 sg13g2_decap_8 FILLER_76_1853 ();
 sg13g2_decap_8 FILLER_76_1860 ();
 sg13g2_decap_8 FILLER_76_1867 ();
 sg13g2_decap_8 FILLER_76_1874 ();
 sg13g2_decap_8 FILLER_76_1881 ();
 sg13g2_decap_8 FILLER_76_1888 ();
 sg13g2_decap_8 FILLER_76_1895 ();
 sg13g2_decap_8 FILLER_76_1902 ();
 sg13g2_decap_8 FILLER_76_1909 ();
 sg13g2_decap_8 FILLER_76_1916 ();
 sg13g2_decap_8 FILLER_76_1923 ();
 sg13g2_decap_8 FILLER_76_1930 ();
 sg13g2_decap_8 FILLER_76_1937 ();
 sg13g2_decap_4 FILLER_76_1944 ();
 sg13g2_fill_1 FILLER_76_1948 ();
 sg13g2_decap_8 FILLER_76_1975 ();
 sg13g2_decap_8 FILLER_76_1982 ();
 sg13g2_decap_8 FILLER_76_1989 ();
 sg13g2_decap_8 FILLER_76_1996 ();
 sg13g2_decap_8 FILLER_76_2003 ();
 sg13g2_decap_4 FILLER_76_2010 ();
 sg13g2_decap_8 FILLER_76_2066 ();
 sg13g2_decap_8 FILLER_76_2073 ();
 sg13g2_decap_8 FILLER_76_2080 ();
 sg13g2_decap_8 FILLER_76_2087 ();
 sg13g2_decap_8 FILLER_76_2094 ();
 sg13g2_decap_8 FILLER_76_2101 ();
 sg13g2_decap_8 FILLER_76_2108 ();
 sg13g2_decap_8 FILLER_76_2115 ();
 sg13g2_decap_8 FILLER_76_2122 ();
 sg13g2_decap_8 FILLER_76_2129 ();
 sg13g2_decap_8 FILLER_76_2136 ();
 sg13g2_decap_8 FILLER_76_2143 ();
 sg13g2_decap_8 FILLER_76_2150 ();
 sg13g2_decap_8 FILLER_76_2157 ();
 sg13g2_decap_8 FILLER_76_2164 ();
 sg13g2_decap_8 FILLER_76_2171 ();
 sg13g2_decap_8 FILLER_76_2178 ();
 sg13g2_decap_8 FILLER_76_2185 ();
 sg13g2_decap_8 FILLER_76_2192 ();
 sg13g2_decap_8 FILLER_76_2199 ();
 sg13g2_decap_8 FILLER_76_2206 ();
 sg13g2_decap_8 FILLER_76_2213 ();
 sg13g2_decap_8 FILLER_76_2220 ();
 sg13g2_decap_8 FILLER_76_2227 ();
 sg13g2_decap_8 FILLER_76_2234 ();
 sg13g2_decap_8 FILLER_76_2241 ();
 sg13g2_decap_8 FILLER_76_2248 ();
 sg13g2_decap_8 FILLER_76_2255 ();
 sg13g2_decap_8 FILLER_76_2262 ();
 sg13g2_decap_8 FILLER_76_2269 ();
 sg13g2_decap_8 FILLER_76_2276 ();
 sg13g2_decap_8 FILLER_76_2283 ();
 sg13g2_decap_8 FILLER_76_2290 ();
 sg13g2_decap_8 FILLER_76_2297 ();
 sg13g2_decap_8 FILLER_76_2304 ();
 sg13g2_decap_8 FILLER_76_2311 ();
 sg13g2_decap_8 FILLER_76_2318 ();
 sg13g2_decap_8 FILLER_76_2325 ();
 sg13g2_decap_8 FILLER_76_2332 ();
 sg13g2_decap_8 FILLER_76_2339 ();
 sg13g2_decap_8 FILLER_76_2346 ();
 sg13g2_decap_8 FILLER_76_2353 ();
 sg13g2_decap_8 FILLER_76_2360 ();
 sg13g2_decap_8 FILLER_76_2367 ();
 sg13g2_decap_8 FILLER_76_2374 ();
 sg13g2_decap_8 FILLER_76_2381 ();
 sg13g2_decap_8 FILLER_76_2388 ();
 sg13g2_decap_8 FILLER_76_2395 ();
 sg13g2_decap_8 FILLER_76_2402 ();
 sg13g2_decap_8 FILLER_76_2409 ();
 sg13g2_decap_8 FILLER_76_2416 ();
 sg13g2_decap_8 FILLER_76_2423 ();
 sg13g2_decap_8 FILLER_76_2430 ();
 sg13g2_decap_8 FILLER_76_2437 ();
 sg13g2_decap_8 FILLER_76_2444 ();
 sg13g2_decap_8 FILLER_76_2451 ();
 sg13g2_decap_8 FILLER_76_2458 ();
 sg13g2_decap_8 FILLER_76_2465 ();
 sg13g2_decap_8 FILLER_76_2472 ();
 sg13g2_decap_8 FILLER_76_2479 ();
 sg13g2_decap_8 FILLER_76_2486 ();
 sg13g2_decap_8 FILLER_76_2493 ();
 sg13g2_decap_8 FILLER_76_2500 ();
 sg13g2_decap_8 FILLER_76_2507 ();
 sg13g2_decap_8 FILLER_76_2514 ();
 sg13g2_decap_8 FILLER_76_2521 ();
 sg13g2_decap_8 FILLER_76_2528 ();
 sg13g2_decap_8 FILLER_76_2535 ();
 sg13g2_decap_8 FILLER_76_2542 ();
 sg13g2_decap_8 FILLER_76_2549 ();
 sg13g2_decap_8 FILLER_76_2556 ();
 sg13g2_decap_8 FILLER_76_2563 ();
 sg13g2_decap_8 FILLER_76_2570 ();
 sg13g2_decap_8 FILLER_76_2577 ();
 sg13g2_decap_8 FILLER_76_2584 ();
 sg13g2_decap_8 FILLER_76_2591 ();
 sg13g2_decap_8 FILLER_76_2598 ();
 sg13g2_decap_8 FILLER_76_2605 ();
 sg13g2_decap_8 FILLER_76_2612 ();
 sg13g2_decap_8 FILLER_76_2619 ();
 sg13g2_decap_8 FILLER_76_2626 ();
 sg13g2_decap_8 FILLER_76_2633 ();
 sg13g2_decap_8 FILLER_76_2640 ();
 sg13g2_decap_8 FILLER_76_2647 ();
 sg13g2_decap_8 FILLER_76_2654 ();
 sg13g2_decap_8 FILLER_76_2661 ();
 sg13g2_decap_8 FILLER_76_2668 ();
 sg13g2_decap_8 FILLER_76_2675 ();
 sg13g2_decap_8 FILLER_76_2682 ();
 sg13g2_decap_8 FILLER_76_2689 ();
 sg13g2_decap_8 FILLER_76_2696 ();
 sg13g2_decap_8 FILLER_76_2703 ();
 sg13g2_decap_8 FILLER_76_2710 ();
 sg13g2_decap_8 FILLER_76_2717 ();
 sg13g2_decap_8 FILLER_76_2724 ();
 sg13g2_decap_8 FILLER_76_2731 ();
 sg13g2_decap_8 FILLER_76_2738 ();
 sg13g2_decap_8 FILLER_76_2745 ();
 sg13g2_decap_8 FILLER_76_2752 ();
 sg13g2_decap_8 FILLER_76_2759 ();
 sg13g2_decap_8 FILLER_76_2766 ();
 sg13g2_decap_8 FILLER_76_2773 ();
 sg13g2_decap_8 FILLER_76_2780 ();
 sg13g2_decap_8 FILLER_76_2787 ();
 sg13g2_decap_8 FILLER_76_2794 ();
 sg13g2_decap_8 FILLER_76_2801 ();
 sg13g2_decap_8 FILLER_76_2808 ();
 sg13g2_decap_8 FILLER_76_2815 ();
 sg13g2_decap_8 FILLER_76_2822 ();
 sg13g2_decap_8 FILLER_76_2829 ();
 sg13g2_decap_8 FILLER_76_2836 ();
 sg13g2_decap_8 FILLER_76_2843 ();
 sg13g2_decap_8 FILLER_76_2850 ();
 sg13g2_decap_8 FILLER_76_2857 ();
 sg13g2_decap_8 FILLER_76_2864 ();
 sg13g2_decap_8 FILLER_76_2871 ();
 sg13g2_decap_8 FILLER_76_2878 ();
 sg13g2_decap_8 FILLER_76_2885 ();
 sg13g2_decap_8 FILLER_76_2892 ();
 sg13g2_decap_8 FILLER_76_2899 ();
 sg13g2_decap_8 FILLER_76_2906 ();
 sg13g2_decap_8 FILLER_76_2913 ();
 sg13g2_decap_8 FILLER_76_2920 ();
 sg13g2_decap_8 FILLER_76_2927 ();
 sg13g2_decap_8 FILLER_76_2934 ();
 sg13g2_decap_8 FILLER_76_2941 ();
 sg13g2_decap_8 FILLER_76_2948 ();
 sg13g2_decap_8 FILLER_76_2955 ();
 sg13g2_decap_8 FILLER_76_2962 ();
 sg13g2_decap_8 FILLER_76_2969 ();
 sg13g2_decap_8 FILLER_76_2976 ();
 sg13g2_decap_8 FILLER_76_2983 ();
 sg13g2_decap_8 FILLER_76_2990 ();
 sg13g2_decap_8 FILLER_76_2997 ();
 sg13g2_decap_8 FILLER_76_3004 ();
 sg13g2_decap_8 FILLER_76_3011 ();
 sg13g2_decap_8 FILLER_76_3018 ();
 sg13g2_decap_8 FILLER_76_3025 ();
 sg13g2_decap_8 FILLER_76_3032 ();
 sg13g2_decap_8 FILLER_76_3039 ();
 sg13g2_decap_8 FILLER_76_3046 ();
 sg13g2_decap_8 FILLER_76_3053 ();
 sg13g2_decap_8 FILLER_76_3060 ();
 sg13g2_decap_8 FILLER_76_3067 ();
 sg13g2_decap_8 FILLER_76_3074 ();
 sg13g2_decap_8 FILLER_76_3081 ();
 sg13g2_decap_8 FILLER_76_3088 ();
 sg13g2_decap_8 FILLER_76_3095 ();
 sg13g2_decap_8 FILLER_76_3102 ();
 sg13g2_decap_8 FILLER_76_3109 ();
 sg13g2_decap_8 FILLER_76_3116 ();
 sg13g2_decap_8 FILLER_76_3123 ();
 sg13g2_decap_8 FILLER_76_3130 ();
 sg13g2_decap_8 FILLER_76_3137 ();
 sg13g2_decap_8 FILLER_76_3144 ();
 sg13g2_decap_8 FILLER_76_3151 ();
 sg13g2_decap_8 FILLER_76_3158 ();
 sg13g2_decap_8 FILLER_76_3165 ();
 sg13g2_decap_8 FILLER_76_3172 ();
 sg13g2_decap_8 FILLER_76_3179 ();
 sg13g2_decap_8 FILLER_76_3186 ();
 sg13g2_decap_8 FILLER_76_3193 ();
 sg13g2_decap_8 FILLER_76_3200 ();
 sg13g2_decap_8 FILLER_76_3207 ();
 sg13g2_decap_8 FILLER_76_3214 ();
 sg13g2_decap_8 FILLER_76_3221 ();
 sg13g2_decap_8 FILLER_76_3228 ();
 sg13g2_decap_8 FILLER_76_3235 ();
 sg13g2_decap_8 FILLER_76_3242 ();
 sg13g2_decap_8 FILLER_76_3249 ();
 sg13g2_decap_8 FILLER_76_3256 ();
 sg13g2_decap_8 FILLER_76_3263 ();
 sg13g2_decap_8 FILLER_76_3270 ();
 sg13g2_decap_8 FILLER_76_3277 ();
 sg13g2_decap_8 FILLER_76_3284 ();
 sg13g2_decap_8 FILLER_76_3291 ();
 sg13g2_decap_8 FILLER_76_3298 ();
 sg13g2_decap_8 FILLER_76_3305 ();
 sg13g2_decap_8 FILLER_76_3312 ();
 sg13g2_decap_8 FILLER_76_3319 ();
 sg13g2_decap_8 FILLER_76_3326 ();
 sg13g2_decap_8 FILLER_76_3333 ();
 sg13g2_decap_8 FILLER_76_3340 ();
 sg13g2_decap_8 FILLER_76_3347 ();
 sg13g2_decap_8 FILLER_76_3354 ();
 sg13g2_decap_8 FILLER_76_3361 ();
 sg13g2_decap_8 FILLER_76_3368 ();
 sg13g2_decap_8 FILLER_76_3375 ();
 sg13g2_decap_8 FILLER_76_3382 ();
 sg13g2_decap_8 FILLER_76_3389 ();
 sg13g2_decap_8 FILLER_76_3396 ();
 sg13g2_decap_8 FILLER_76_3403 ();
 sg13g2_decap_8 FILLER_76_3410 ();
 sg13g2_decap_8 FILLER_76_3417 ();
 sg13g2_decap_8 FILLER_76_3424 ();
 sg13g2_decap_8 FILLER_76_3431 ();
 sg13g2_decap_8 FILLER_76_3438 ();
 sg13g2_decap_8 FILLER_76_3445 ();
 sg13g2_decap_8 FILLER_76_3452 ();
 sg13g2_decap_8 FILLER_76_3459 ();
 sg13g2_decap_8 FILLER_76_3466 ();
 sg13g2_decap_8 FILLER_76_3473 ();
 sg13g2_decap_8 FILLER_76_3480 ();
 sg13g2_decap_8 FILLER_76_3487 ();
 sg13g2_decap_8 FILLER_76_3494 ();
 sg13g2_decap_8 FILLER_76_3501 ();
 sg13g2_decap_8 FILLER_76_3508 ();
 sg13g2_decap_8 FILLER_76_3515 ();
 sg13g2_decap_8 FILLER_76_3522 ();
 sg13g2_decap_8 FILLER_76_3529 ();
 sg13g2_decap_8 FILLER_76_3536 ();
 sg13g2_decap_8 FILLER_76_3543 ();
 sg13g2_decap_8 FILLER_76_3550 ();
 sg13g2_decap_8 FILLER_76_3557 ();
 sg13g2_decap_8 FILLER_76_3564 ();
 sg13g2_decap_8 FILLER_76_3571 ();
 sg13g2_fill_2 FILLER_76_3578 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_448 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_8 FILLER_77_462 ();
 sg13g2_decap_8 FILLER_77_469 ();
 sg13g2_decap_8 FILLER_77_476 ();
 sg13g2_decap_8 FILLER_77_483 ();
 sg13g2_decap_8 FILLER_77_490 ();
 sg13g2_decap_8 FILLER_77_497 ();
 sg13g2_decap_8 FILLER_77_504 ();
 sg13g2_decap_8 FILLER_77_511 ();
 sg13g2_decap_8 FILLER_77_518 ();
 sg13g2_decap_8 FILLER_77_525 ();
 sg13g2_decap_8 FILLER_77_532 ();
 sg13g2_decap_8 FILLER_77_539 ();
 sg13g2_decap_8 FILLER_77_546 ();
 sg13g2_decap_8 FILLER_77_553 ();
 sg13g2_decap_8 FILLER_77_560 ();
 sg13g2_decap_8 FILLER_77_567 ();
 sg13g2_decap_8 FILLER_77_574 ();
 sg13g2_decap_8 FILLER_77_581 ();
 sg13g2_decap_4 FILLER_77_588 ();
 sg13g2_fill_1 FILLER_77_597 ();
 sg13g2_decap_8 FILLER_77_603 ();
 sg13g2_decap_8 FILLER_77_610 ();
 sg13g2_decap_8 FILLER_77_617 ();
 sg13g2_decap_8 FILLER_77_624 ();
 sg13g2_decap_8 FILLER_77_631 ();
 sg13g2_decap_8 FILLER_77_638 ();
 sg13g2_decap_8 FILLER_77_645 ();
 sg13g2_decap_8 FILLER_77_652 ();
 sg13g2_decap_4 FILLER_77_659 ();
 sg13g2_fill_1 FILLER_77_663 ();
 sg13g2_fill_2 FILLER_77_737 ();
 sg13g2_fill_1 FILLER_77_739 ();
 sg13g2_fill_2 FILLER_77_753 ();
 sg13g2_decap_4 FILLER_77_794 ();
 sg13g2_fill_1 FILLER_77_803 ();
 sg13g2_fill_1 FILLER_77_809 ();
 sg13g2_fill_2 FILLER_77_836 ();
 sg13g2_fill_1 FILLER_77_838 ();
 sg13g2_fill_2 FILLER_77_855 ();
 sg13g2_fill_1 FILLER_77_857 ();
 sg13g2_fill_2 FILLER_77_932 ();
 sg13g2_fill_1 FILLER_77_934 ();
 sg13g2_decap_8 FILLER_77_939 ();
 sg13g2_decap_4 FILLER_77_946 ();
 sg13g2_fill_2 FILLER_77_950 ();
 sg13g2_decap_8 FILLER_77_992 ();
 sg13g2_fill_2 FILLER_77_999 ();
 sg13g2_fill_1 FILLER_77_1016 ();
 sg13g2_decap_8 FILLER_77_1051 ();
 sg13g2_decap_8 FILLER_77_1058 ();
 sg13g2_decap_8 FILLER_77_1065 ();
 sg13g2_fill_2 FILLER_77_1072 ();
 sg13g2_fill_1 FILLER_77_1074 ();
 sg13g2_decap_8 FILLER_77_1101 ();
 sg13g2_decap_8 FILLER_77_1108 ();
 sg13g2_fill_1 FILLER_77_1115 ();
 sg13g2_fill_2 FILLER_77_1123 ();
 sg13g2_decap_8 FILLER_77_1181 ();
 sg13g2_fill_1 FILLER_77_1188 ();
 sg13g2_decap_8 FILLER_77_1215 ();
 sg13g2_decap_8 FILLER_77_1222 ();
 sg13g2_decap_4 FILLER_77_1229 ();
 sg13g2_fill_1 FILLER_77_1233 ();
 sg13g2_decap_4 FILLER_77_1238 ();
 sg13g2_fill_2 FILLER_77_1297 ();
 sg13g2_decap_4 FILLER_77_1323 ();
 sg13g2_fill_2 FILLER_77_1327 ();
 sg13g2_fill_2 FILLER_77_1359 ();
 sg13g2_fill_1 FILLER_77_1421 ();
 sg13g2_decap_8 FILLER_77_1487 ();
 sg13g2_decap_8 FILLER_77_1494 ();
 sg13g2_decap_8 FILLER_77_1501 ();
 sg13g2_decap_8 FILLER_77_1508 ();
 sg13g2_decap_8 FILLER_77_1515 ();
 sg13g2_decap_8 FILLER_77_1522 ();
 sg13g2_decap_8 FILLER_77_1529 ();
 sg13g2_decap_8 FILLER_77_1536 ();
 sg13g2_decap_8 FILLER_77_1543 ();
 sg13g2_decap_8 FILLER_77_1550 ();
 sg13g2_decap_8 FILLER_77_1557 ();
 sg13g2_decap_8 FILLER_77_1564 ();
 sg13g2_decap_8 FILLER_77_1571 ();
 sg13g2_decap_8 FILLER_77_1578 ();
 sg13g2_decap_8 FILLER_77_1585 ();
 sg13g2_decap_8 FILLER_77_1592 ();
 sg13g2_decap_8 FILLER_77_1599 ();
 sg13g2_decap_8 FILLER_77_1606 ();
 sg13g2_decap_8 FILLER_77_1613 ();
 sg13g2_decap_8 FILLER_77_1620 ();
 sg13g2_decap_8 FILLER_77_1627 ();
 sg13g2_decap_8 FILLER_77_1634 ();
 sg13g2_decap_8 FILLER_77_1641 ();
 sg13g2_decap_8 FILLER_77_1648 ();
 sg13g2_decap_8 FILLER_77_1655 ();
 sg13g2_decap_8 FILLER_77_1662 ();
 sg13g2_decap_8 FILLER_77_1669 ();
 sg13g2_decap_8 FILLER_77_1676 ();
 sg13g2_decap_8 FILLER_77_1683 ();
 sg13g2_decap_8 FILLER_77_1690 ();
 sg13g2_decap_8 FILLER_77_1697 ();
 sg13g2_decap_8 FILLER_77_1704 ();
 sg13g2_decap_8 FILLER_77_1711 ();
 sg13g2_decap_8 FILLER_77_1718 ();
 sg13g2_decap_8 FILLER_77_1725 ();
 sg13g2_decap_8 FILLER_77_1732 ();
 sg13g2_decap_8 FILLER_77_1739 ();
 sg13g2_decap_8 FILLER_77_1746 ();
 sg13g2_decap_8 FILLER_77_1753 ();
 sg13g2_decap_8 FILLER_77_1760 ();
 sg13g2_decap_8 FILLER_77_1767 ();
 sg13g2_decap_8 FILLER_77_1774 ();
 sg13g2_decap_8 FILLER_77_1781 ();
 sg13g2_decap_8 FILLER_77_1788 ();
 sg13g2_decap_8 FILLER_77_1795 ();
 sg13g2_decap_8 FILLER_77_1802 ();
 sg13g2_decap_8 FILLER_77_1809 ();
 sg13g2_decap_8 FILLER_77_1816 ();
 sg13g2_decap_8 FILLER_77_1823 ();
 sg13g2_decap_8 FILLER_77_1830 ();
 sg13g2_decap_8 FILLER_77_1837 ();
 sg13g2_decap_8 FILLER_77_1844 ();
 sg13g2_decap_8 FILLER_77_1851 ();
 sg13g2_decap_8 FILLER_77_1858 ();
 sg13g2_decap_8 FILLER_77_1865 ();
 sg13g2_decap_8 FILLER_77_1872 ();
 sg13g2_decap_8 FILLER_77_1879 ();
 sg13g2_decap_8 FILLER_77_1886 ();
 sg13g2_decap_8 FILLER_77_1893 ();
 sg13g2_decap_8 FILLER_77_1900 ();
 sg13g2_decap_8 FILLER_77_1907 ();
 sg13g2_decap_8 FILLER_77_1914 ();
 sg13g2_decap_8 FILLER_77_1921 ();
 sg13g2_decap_8 FILLER_77_1928 ();
 sg13g2_decap_8 FILLER_77_1935 ();
 sg13g2_decap_8 FILLER_77_1942 ();
 sg13g2_decap_8 FILLER_77_1949 ();
 sg13g2_decap_8 FILLER_77_1956 ();
 sg13g2_decap_8 FILLER_77_1963 ();
 sg13g2_decap_8 FILLER_77_1970 ();
 sg13g2_decap_8 FILLER_77_1977 ();
 sg13g2_decap_8 FILLER_77_1984 ();
 sg13g2_decap_8 FILLER_77_1991 ();
 sg13g2_decap_8 FILLER_77_1998 ();
 sg13g2_decap_8 FILLER_77_2005 ();
 sg13g2_decap_8 FILLER_77_2012 ();
 sg13g2_fill_1 FILLER_77_2019 ();
 sg13g2_decap_8 FILLER_77_2046 ();
 sg13g2_decap_8 FILLER_77_2053 ();
 sg13g2_decap_8 FILLER_77_2060 ();
 sg13g2_decap_8 FILLER_77_2067 ();
 sg13g2_decap_8 FILLER_77_2074 ();
 sg13g2_decap_8 FILLER_77_2081 ();
 sg13g2_decap_8 FILLER_77_2088 ();
 sg13g2_decap_8 FILLER_77_2095 ();
 sg13g2_decap_8 FILLER_77_2102 ();
 sg13g2_decap_8 FILLER_77_2109 ();
 sg13g2_decap_8 FILLER_77_2116 ();
 sg13g2_decap_8 FILLER_77_2123 ();
 sg13g2_decap_8 FILLER_77_2130 ();
 sg13g2_decap_8 FILLER_77_2137 ();
 sg13g2_decap_8 FILLER_77_2144 ();
 sg13g2_decap_8 FILLER_77_2151 ();
 sg13g2_decap_8 FILLER_77_2158 ();
 sg13g2_decap_8 FILLER_77_2165 ();
 sg13g2_decap_8 FILLER_77_2172 ();
 sg13g2_decap_8 FILLER_77_2179 ();
 sg13g2_decap_8 FILLER_77_2186 ();
 sg13g2_decap_8 FILLER_77_2193 ();
 sg13g2_decap_8 FILLER_77_2200 ();
 sg13g2_decap_8 FILLER_77_2207 ();
 sg13g2_decap_8 FILLER_77_2214 ();
 sg13g2_decap_8 FILLER_77_2221 ();
 sg13g2_decap_8 FILLER_77_2228 ();
 sg13g2_decap_8 FILLER_77_2235 ();
 sg13g2_decap_8 FILLER_77_2242 ();
 sg13g2_decap_8 FILLER_77_2249 ();
 sg13g2_decap_8 FILLER_77_2256 ();
 sg13g2_decap_8 FILLER_77_2263 ();
 sg13g2_decap_8 FILLER_77_2270 ();
 sg13g2_decap_8 FILLER_77_2277 ();
 sg13g2_decap_8 FILLER_77_2284 ();
 sg13g2_decap_8 FILLER_77_2291 ();
 sg13g2_decap_8 FILLER_77_2298 ();
 sg13g2_decap_8 FILLER_77_2305 ();
 sg13g2_decap_8 FILLER_77_2312 ();
 sg13g2_decap_8 FILLER_77_2319 ();
 sg13g2_decap_8 FILLER_77_2326 ();
 sg13g2_decap_8 FILLER_77_2333 ();
 sg13g2_decap_8 FILLER_77_2340 ();
 sg13g2_decap_8 FILLER_77_2347 ();
 sg13g2_decap_8 FILLER_77_2354 ();
 sg13g2_decap_8 FILLER_77_2361 ();
 sg13g2_decap_8 FILLER_77_2368 ();
 sg13g2_decap_8 FILLER_77_2375 ();
 sg13g2_decap_8 FILLER_77_2382 ();
 sg13g2_decap_8 FILLER_77_2389 ();
 sg13g2_decap_8 FILLER_77_2396 ();
 sg13g2_decap_8 FILLER_77_2403 ();
 sg13g2_decap_8 FILLER_77_2410 ();
 sg13g2_decap_8 FILLER_77_2417 ();
 sg13g2_decap_8 FILLER_77_2424 ();
 sg13g2_decap_8 FILLER_77_2431 ();
 sg13g2_decap_8 FILLER_77_2438 ();
 sg13g2_decap_8 FILLER_77_2445 ();
 sg13g2_decap_8 FILLER_77_2452 ();
 sg13g2_decap_8 FILLER_77_2459 ();
 sg13g2_decap_8 FILLER_77_2466 ();
 sg13g2_decap_8 FILLER_77_2473 ();
 sg13g2_decap_8 FILLER_77_2480 ();
 sg13g2_decap_8 FILLER_77_2487 ();
 sg13g2_decap_8 FILLER_77_2494 ();
 sg13g2_decap_8 FILLER_77_2501 ();
 sg13g2_decap_8 FILLER_77_2508 ();
 sg13g2_decap_8 FILLER_77_2515 ();
 sg13g2_decap_8 FILLER_77_2522 ();
 sg13g2_decap_8 FILLER_77_2529 ();
 sg13g2_decap_8 FILLER_77_2536 ();
 sg13g2_decap_8 FILLER_77_2543 ();
 sg13g2_decap_8 FILLER_77_2550 ();
 sg13g2_decap_8 FILLER_77_2557 ();
 sg13g2_decap_8 FILLER_77_2564 ();
 sg13g2_decap_8 FILLER_77_2571 ();
 sg13g2_decap_8 FILLER_77_2578 ();
 sg13g2_decap_8 FILLER_77_2585 ();
 sg13g2_decap_8 FILLER_77_2592 ();
 sg13g2_decap_8 FILLER_77_2599 ();
 sg13g2_decap_8 FILLER_77_2606 ();
 sg13g2_decap_8 FILLER_77_2613 ();
 sg13g2_decap_8 FILLER_77_2620 ();
 sg13g2_decap_8 FILLER_77_2627 ();
 sg13g2_decap_8 FILLER_77_2634 ();
 sg13g2_decap_8 FILLER_77_2641 ();
 sg13g2_decap_8 FILLER_77_2648 ();
 sg13g2_decap_8 FILLER_77_2655 ();
 sg13g2_decap_8 FILLER_77_2662 ();
 sg13g2_decap_8 FILLER_77_2669 ();
 sg13g2_decap_8 FILLER_77_2676 ();
 sg13g2_decap_8 FILLER_77_2683 ();
 sg13g2_decap_8 FILLER_77_2690 ();
 sg13g2_decap_8 FILLER_77_2697 ();
 sg13g2_decap_8 FILLER_77_2704 ();
 sg13g2_decap_8 FILLER_77_2711 ();
 sg13g2_decap_8 FILLER_77_2718 ();
 sg13g2_decap_8 FILLER_77_2725 ();
 sg13g2_decap_8 FILLER_77_2732 ();
 sg13g2_decap_8 FILLER_77_2739 ();
 sg13g2_decap_8 FILLER_77_2746 ();
 sg13g2_decap_8 FILLER_77_2753 ();
 sg13g2_decap_8 FILLER_77_2760 ();
 sg13g2_decap_8 FILLER_77_2767 ();
 sg13g2_decap_8 FILLER_77_2774 ();
 sg13g2_decap_8 FILLER_77_2781 ();
 sg13g2_decap_8 FILLER_77_2788 ();
 sg13g2_decap_8 FILLER_77_2795 ();
 sg13g2_decap_8 FILLER_77_2802 ();
 sg13g2_decap_8 FILLER_77_2809 ();
 sg13g2_decap_8 FILLER_77_2816 ();
 sg13g2_decap_8 FILLER_77_2823 ();
 sg13g2_decap_8 FILLER_77_2830 ();
 sg13g2_decap_8 FILLER_77_2837 ();
 sg13g2_decap_8 FILLER_77_2844 ();
 sg13g2_decap_8 FILLER_77_2851 ();
 sg13g2_decap_8 FILLER_77_2858 ();
 sg13g2_decap_8 FILLER_77_2865 ();
 sg13g2_decap_8 FILLER_77_2872 ();
 sg13g2_decap_8 FILLER_77_2879 ();
 sg13g2_decap_8 FILLER_77_2886 ();
 sg13g2_decap_8 FILLER_77_2893 ();
 sg13g2_decap_8 FILLER_77_2900 ();
 sg13g2_decap_8 FILLER_77_2907 ();
 sg13g2_decap_8 FILLER_77_2914 ();
 sg13g2_decap_8 FILLER_77_2921 ();
 sg13g2_decap_8 FILLER_77_2928 ();
 sg13g2_decap_8 FILLER_77_2935 ();
 sg13g2_decap_8 FILLER_77_2942 ();
 sg13g2_decap_8 FILLER_77_2949 ();
 sg13g2_decap_8 FILLER_77_2956 ();
 sg13g2_decap_8 FILLER_77_2963 ();
 sg13g2_decap_8 FILLER_77_2970 ();
 sg13g2_decap_8 FILLER_77_2977 ();
 sg13g2_decap_8 FILLER_77_2984 ();
 sg13g2_decap_8 FILLER_77_2991 ();
 sg13g2_decap_8 FILLER_77_2998 ();
 sg13g2_decap_8 FILLER_77_3005 ();
 sg13g2_decap_8 FILLER_77_3012 ();
 sg13g2_decap_8 FILLER_77_3019 ();
 sg13g2_decap_8 FILLER_77_3026 ();
 sg13g2_decap_8 FILLER_77_3033 ();
 sg13g2_decap_8 FILLER_77_3040 ();
 sg13g2_decap_8 FILLER_77_3047 ();
 sg13g2_decap_8 FILLER_77_3054 ();
 sg13g2_decap_8 FILLER_77_3061 ();
 sg13g2_decap_8 FILLER_77_3068 ();
 sg13g2_decap_8 FILLER_77_3075 ();
 sg13g2_decap_8 FILLER_77_3082 ();
 sg13g2_decap_8 FILLER_77_3089 ();
 sg13g2_decap_8 FILLER_77_3096 ();
 sg13g2_decap_8 FILLER_77_3103 ();
 sg13g2_decap_8 FILLER_77_3110 ();
 sg13g2_decap_8 FILLER_77_3117 ();
 sg13g2_decap_8 FILLER_77_3124 ();
 sg13g2_decap_8 FILLER_77_3131 ();
 sg13g2_decap_8 FILLER_77_3138 ();
 sg13g2_decap_8 FILLER_77_3145 ();
 sg13g2_decap_8 FILLER_77_3152 ();
 sg13g2_decap_8 FILLER_77_3159 ();
 sg13g2_decap_8 FILLER_77_3166 ();
 sg13g2_decap_8 FILLER_77_3173 ();
 sg13g2_decap_8 FILLER_77_3180 ();
 sg13g2_decap_8 FILLER_77_3187 ();
 sg13g2_decap_8 FILLER_77_3194 ();
 sg13g2_decap_8 FILLER_77_3201 ();
 sg13g2_decap_8 FILLER_77_3208 ();
 sg13g2_decap_8 FILLER_77_3215 ();
 sg13g2_decap_8 FILLER_77_3222 ();
 sg13g2_decap_8 FILLER_77_3229 ();
 sg13g2_decap_8 FILLER_77_3236 ();
 sg13g2_decap_8 FILLER_77_3243 ();
 sg13g2_decap_8 FILLER_77_3250 ();
 sg13g2_decap_8 FILLER_77_3257 ();
 sg13g2_decap_8 FILLER_77_3264 ();
 sg13g2_decap_8 FILLER_77_3271 ();
 sg13g2_decap_8 FILLER_77_3278 ();
 sg13g2_decap_8 FILLER_77_3285 ();
 sg13g2_decap_8 FILLER_77_3292 ();
 sg13g2_decap_8 FILLER_77_3299 ();
 sg13g2_decap_8 FILLER_77_3306 ();
 sg13g2_decap_8 FILLER_77_3313 ();
 sg13g2_decap_8 FILLER_77_3320 ();
 sg13g2_decap_8 FILLER_77_3327 ();
 sg13g2_decap_8 FILLER_77_3334 ();
 sg13g2_decap_8 FILLER_77_3341 ();
 sg13g2_decap_8 FILLER_77_3348 ();
 sg13g2_decap_8 FILLER_77_3355 ();
 sg13g2_decap_8 FILLER_77_3362 ();
 sg13g2_decap_8 FILLER_77_3369 ();
 sg13g2_decap_8 FILLER_77_3376 ();
 sg13g2_decap_8 FILLER_77_3383 ();
 sg13g2_decap_8 FILLER_77_3390 ();
 sg13g2_decap_8 FILLER_77_3397 ();
 sg13g2_decap_8 FILLER_77_3404 ();
 sg13g2_decap_8 FILLER_77_3411 ();
 sg13g2_decap_8 FILLER_77_3418 ();
 sg13g2_decap_8 FILLER_77_3425 ();
 sg13g2_decap_8 FILLER_77_3432 ();
 sg13g2_decap_8 FILLER_77_3439 ();
 sg13g2_decap_8 FILLER_77_3446 ();
 sg13g2_decap_8 FILLER_77_3453 ();
 sg13g2_decap_8 FILLER_77_3460 ();
 sg13g2_decap_8 FILLER_77_3467 ();
 sg13g2_decap_8 FILLER_77_3474 ();
 sg13g2_decap_8 FILLER_77_3481 ();
 sg13g2_decap_8 FILLER_77_3488 ();
 sg13g2_decap_8 FILLER_77_3495 ();
 sg13g2_decap_8 FILLER_77_3502 ();
 sg13g2_decap_8 FILLER_77_3509 ();
 sg13g2_decap_8 FILLER_77_3516 ();
 sg13g2_decap_8 FILLER_77_3523 ();
 sg13g2_decap_8 FILLER_77_3530 ();
 sg13g2_decap_8 FILLER_77_3537 ();
 sg13g2_decap_8 FILLER_77_3544 ();
 sg13g2_decap_8 FILLER_77_3551 ();
 sg13g2_decap_8 FILLER_77_3558 ();
 sg13g2_decap_8 FILLER_77_3565 ();
 sg13g2_decap_8 FILLER_77_3572 ();
 sg13g2_fill_1 FILLER_77_3579 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_decap_8 FILLER_78_448 ();
 sg13g2_decap_8 FILLER_78_455 ();
 sg13g2_decap_8 FILLER_78_462 ();
 sg13g2_decap_8 FILLER_78_469 ();
 sg13g2_decap_8 FILLER_78_476 ();
 sg13g2_decap_8 FILLER_78_483 ();
 sg13g2_decap_8 FILLER_78_490 ();
 sg13g2_decap_8 FILLER_78_497 ();
 sg13g2_decap_8 FILLER_78_504 ();
 sg13g2_decap_8 FILLER_78_511 ();
 sg13g2_decap_8 FILLER_78_518 ();
 sg13g2_decap_8 FILLER_78_525 ();
 sg13g2_decap_8 FILLER_78_532 ();
 sg13g2_decap_8 FILLER_78_539 ();
 sg13g2_decap_8 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_553 ();
 sg13g2_decap_8 FILLER_78_560 ();
 sg13g2_decap_8 FILLER_78_567 ();
 sg13g2_decap_8 FILLER_78_574 ();
 sg13g2_decap_8 FILLER_78_581 ();
 sg13g2_decap_8 FILLER_78_588 ();
 sg13g2_decap_8 FILLER_78_595 ();
 sg13g2_decap_8 FILLER_78_602 ();
 sg13g2_decap_8 FILLER_78_609 ();
 sg13g2_decap_8 FILLER_78_616 ();
 sg13g2_decap_8 FILLER_78_623 ();
 sg13g2_decap_8 FILLER_78_630 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_decap_8 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_651 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_fill_1 FILLER_78_672 ();
 sg13g2_fill_1 FILLER_78_770 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_fill_2 FILLER_78_833 ();
 sg13g2_decap_4 FILLER_78_842 ();
 sg13g2_fill_1 FILLER_78_942 ();
 sg13g2_decap_4 FILLER_78_985 ();
 sg13g2_decap_4 FILLER_78_1106 ();
 sg13g2_decap_8 FILLER_78_1172 ();
 sg13g2_decap_8 FILLER_78_1179 ();
 sg13g2_fill_2 FILLER_78_1186 ();
 sg13g2_fill_1 FILLER_78_1188 ();
 sg13g2_decap_8 FILLER_78_1215 ();
 sg13g2_decap_8 FILLER_78_1222 ();
 sg13g2_decap_8 FILLER_78_1229 ();
 sg13g2_fill_2 FILLER_78_1240 ();
 sg13g2_fill_1 FILLER_78_1242 ();
 sg13g2_fill_2 FILLER_78_1362 ();
 sg13g2_fill_1 FILLER_78_1364 ();
 sg13g2_fill_1 FILLER_78_1391 ();
 sg13g2_fill_2 FILLER_78_1429 ();
 sg13g2_decap_8 FILLER_78_1459 ();
 sg13g2_decap_8 FILLER_78_1466 ();
 sg13g2_decap_8 FILLER_78_1473 ();
 sg13g2_decap_8 FILLER_78_1480 ();
 sg13g2_decap_8 FILLER_78_1487 ();
 sg13g2_decap_8 FILLER_78_1494 ();
 sg13g2_decap_8 FILLER_78_1501 ();
 sg13g2_decap_8 FILLER_78_1508 ();
 sg13g2_decap_8 FILLER_78_1515 ();
 sg13g2_decap_8 FILLER_78_1522 ();
 sg13g2_decap_8 FILLER_78_1529 ();
 sg13g2_decap_8 FILLER_78_1536 ();
 sg13g2_decap_8 FILLER_78_1543 ();
 sg13g2_decap_8 FILLER_78_1550 ();
 sg13g2_decap_8 FILLER_78_1557 ();
 sg13g2_decap_8 FILLER_78_1564 ();
 sg13g2_decap_8 FILLER_78_1571 ();
 sg13g2_decap_8 FILLER_78_1578 ();
 sg13g2_decap_8 FILLER_78_1585 ();
 sg13g2_decap_8 FILLER_78_1592 ();
 sg13g2_decap_8 FILLER_78_1599 ();
 sg13g2_decap_8 FILLER_78_1606 ();
 sg13g2_decap_8 FILLER_78_1613 ();
 sg13g2_decap_8 FILLER_78_1620 ();
 sg13g2_decap_8 FILLER_78_1627 ();
 sg13g2_decap_8 FILLER_78_1634 ();
 sg13g2_decap_8 FILLER_78_1641 ();
 sg13g2_decap_8 FILLER_78_1648 ();
 sg13g2_decap_8 FILLER_78_1655 ();
 sg13g2_decap_8 FILLER_78_1662 ();
 sg13g2_decap_8 FILLER_78_1669 ();
 sg13g2_decap_8 FILLER_78_1676 ();
 sg13g2_decap_8 FILLER_78_1683 ();
 sg13g2_decap_8 FILLER_78_1690 ();
 sg13g2_decap_8 FILLER_78_1697 ();
 sg13g2_decap_8 FILLER_78_1704 ();
 sg13g2_decap_8 FILLER_78_1711 ();
 sg13g2_decap_8 FILLER_78_1718 ();
 sg13g2_decap_8 FILLER_78_1725 ();
 sg13g2_decap_8 FILLER_78_1732 ();
 sg13g2_decap_8 FILLER_78_1739 ();
 sg13g2_decap_8 FILLER_78_1746 ();
 sg13g2_decap_8 FILLER_78_1753 ();
 sg13g2_decap_8 FILLER_78_1760 ();
 sg13g2_decap_8 FILLER_78_1767 ();
 sg13g2_decap_8 FILLER_78_1774 ();
 sg13g2_decap_8 FILLER_78_1781 ();
 sg13g2_decap_8 FILLER_78_1788 ();
 sg13g2_decap_8 FILLER_78_1795 ();
 sg13g2_decap_8 FILLER_78_1802 ();
 sg13g2_decap_8 FILLER_78_1809 ();
 sg13g2_decap_8 FILLER_78_1816 ();
 sg13g2_decap_8 FILLER_78_1823 ();
 sg13g2_decap_8 FILLER_78_1830 ();
 sg13g2_decap_8 FILLER_78_1837 ();
 sg13g2_decap_8 FILLER_78_1844 ();
 sg13g2_decap_8 FILLER_78_1851 ();
 sg13g2_decap_8 FILLER_78_1858 ();
 sg13g2_decap_8 FILLER_78_1865 ();
 sg13g2_decap_8 FILLER_78_1872 ();
 sg13g2_decap_8 FILLER_78_1879 ();
 sg13g2_decap_8 FILLER_78_1886 ();
 sg13g2_decap_8 FILLER_78_1893 ();
 sg13g2_decap_8 FILLER_78_1900 ();
 sg13g2_decap_8 FILLER_78_1907 ();
 sg13g2_decap_8 FILLER_78_1914 ();
 sg13g2_decap_8 FILLER_78_1921 ();
 sg13g2_decap_8 FILLER_78_1928 ();
 sg13g2_decap_8 FILLER_78_1935 ();
 sg13g2_decap_8 FILLER_78_1942 ();
 sg13g2_decap_8 FILLER_78_1949 ();
 sg13g2_decap_8 FILLER_78_1956 ();
 sg13g2_decap_8 FILLER_78_1963 ();
 sg13g2_decap_8 FILLER_78_1970 ();
 sg13g2_decap_8 FILLER_78_1977 ();
 sg13g2_decap_8 FILLER_78_1984 ();
 sg13g2_decap_8 FILLER_78_1991 ();
 sg13g2_decap_8 FILLER_78_1998 ();
 sg13g2_decap_8 FILLER_78_2005 ();
 sg13g2_decap_8 FILLER_78_2012 ();
 sg13g2_decap_8 FILLER_78_2019 ();
 sg13g2_decap_8 FILLER_78_2026 ();
 sg13g2_decap_8 FILLER_78_2033 ();
 sg13g2_decap_8 FILLER_78_2040 ();
 sg13g2_decap_8 FILLER_78_2047 ();
 sg13g2_decap_8 FILLER_78_2054 ();
 sg13g2_decap_8 FILLER_78_2061 ();
 sg13g2_decap_8 FILLER_78_2068 ();
 sg13g2_decap_8 FILLER_78_2075 ();
 sg13g2_decap_8 FILLER_78_2082 ();
 sg13g2_decap_8 FILLER_78_2089 ();
 sg13g2_decap_8 FILLER_78_2096 ();
 sg13g2_decap_8 FILLER_78_2103 ();
 sg13g2_decap_8 FILLER_78_2110 ();
 sg13g2_decap_8 FILLER_78_2117 ();
 sg13g2_decap_8 FILLER_78_2124 ();
 sg13g2_decap_8 FILLER_78_2131 ();
 sg13g2_decap_8 FILLER_78_2138 ();
 sg13g2_decap_8 FILLER_78_2145 ();
 sg13g2_decap_8 FILLER_78_2152 ();
 sg13g2_decap_8 FILLER_78_2159 ();
 sg13g2_decap_8 FILLER_78_2166 ();
 sg13g2_decap_8 FILLER_78_2173 ();
 sg13g2_decap_8 FILLER_78_2180 ();
 sg13g2_decap_8 FILLER_78_2187 ();
 sg13g2_decap_8 FILLER_78_2194 ();
 sg13g2_decap_8 FILLER_78_2201 ();
 sg13g2_decap_8 FILLER_78_2208 ();
 sg13g2_decap_8 FILLER_78_2215 ();
 sg13g2_decap_8 FILLER_78_2222 ();
 sg13g2_decap_8 FILLER_78_2229 ();
 sg13g2_decap_8 FILLER_78_2236 ();
 sg13g2_decap_8 FILLER_78_2243 ();
 sg13g2_decap_8 FILLER_78_2250 ();
 sg13g2_decap_8 FILLER_78_2257 ();
 sg13g2_decap_8 FILLER_78_2264 ();
 sg13g2_decap_8 FILLER_78_2271 ();
 sg13g2_decap_8 FILLER_78_2278 ();
 sg13g2_decap_8 FILLER_78_2285 ();
 sg13g2_decap_8 FILLER_78_2292 ();
 sg13g2_decap_8 FILLER_78_2299 ();
 sg13g2_decap_8 FILLER_78_2306 ();
 sg13g2_decap_8 FILLER_78_2313 ();
 sg13g2_decap_8 FILLER_78_2320 ();
 sg13g2_decap_8 FILLER_78_2327 ();
 sg13g2_decap_8 FILLER_78_2334 ();
 sg13g2_decap_8 FILLER_78_2341 ();
 sg13g2_decap_8 FILLER_78_2348 ();
 sg13g2_decap_8 FILLER_78_2355 ();
 sg13g2_decap_8 FILLER_78_2362 ();
 sg13g2_decap_8 FILLER_78_2369 ();
 sg13g2_decap_8 FILLER_78_2376 ();
 sg13g2_decap_8 FILLER_78_2383 ();
 sg13g2_decap_8 FILLER_78_2390 ();
 sg13g2_decap_8 FILLER_78_2397 ();
 sg13g2_decap_8 FILLER_78_2404 ();
 sg13g2_decap_8 FILLER_78_2411 ();
 sg13g2_decap_8 FILLER_78_2418 ();
 sg13g2_decap_8 FILLER_78_2425 ();
 sg13g2_decap_8 FILLER_78_2432 ();
 sg13g2_decap_8 FILLER_78_2439 ();
 sg13g2_decap_8 FILLER_78_2446 ();
 sg13g2_decap_8 FILLER_78_2453 ();
 sg13g2_decap_8 FILLER_78_2460 ();
 sg13g2_decap_8 FILLER_78_2467 ();
 sg13g2_decap_8 FILLER_78_2474 ();
 sg13g2_decap_8 FILLER_78_2481 ();
 sg13g2_decap_8 FILLER_78_2488 ();
 sg13g2_decap_8 FILLER_78_2495 ();
 sg13g2_decap_8 FILLER_78_2502 ();
 sg13g2_decap_8 FILLER_78_2509 ();
 sg13g2_decap_8 FILLER_78_2516 ();
 sg13g2_decap_8 FILLER_78_2523 ();
 sg13g2_decap_8 FILLER_78_2530 ();
 sg13g2_decap_8 FILLER_78_2537 ();
 sg13g2_decap_8 FILLER_78_2544 ();
 sg13g2_decap_8 FILLER_78_2551 ();
 sg13g2_decap_8 FILLER_78_2558 ();
 sg13g2_decap_8 FILLER_78_2565 ();
 sg13g2_decap_8 FILLER_78_2572 ();
 sg13g2_decap_8 FILLER_78_2579 ();
 sg13g2_decap_8 FILLER_78_2586 ();
 sg13g2_decap_8 FILLER_78_2593 ();
 sg13g2_decap_8 FILLER_78_2600 ();
 sg13g2_decap_8 FILLER_78_2607 ();
 sg13g2_decap_8 FILLER_78_2614 ();
 sg13g2_decap_8 FILLER_78_2621 ();
 sg13g2_decap_8 FILLER_78_2628 ();
 sg13g2_decap_8 FILLER_78_2635 ();
 sg13g2_decap_8 FILLER_78_2642 ();
 sg13g2_decap_8 FILLER_78_2649 ();
 sg13g2_decap_8 FILLER_78_2656 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_decap_8 FILLER_78_2670 ();
 sg13g2_decap_8 FILLER_78_2677 ();
 sg13g2_decap_8 FILLER_78_2684 ();
 sg13g2_decap_8 FILLER_78_2691 ();
 sg13g2_decap_8 FILLER_78_2698 ();
 sg13g2_decap_8 FILLER_78_2705 ();
 sg13g2_decap_8 FILLER_78_2712 ();
 sg13g2_decap_8 FILLER_78_2719 ();
 sg13g2_decap_8 FILLER_78_2726 ();
 sg13g2_decap_8 FILLER_78_2733 ();
 sg13g2_decap_8 FILLER_78_2740 ();
 sg13g2_decap_8 FILLER_78_2747 ();
 sg13g2_decap_8 FILLER_78_2754 ();
 sg13g2_decap_8 FILLER_78_2761 ();
 sg13g2_decap_8 FILLER_78_2768 ();
 sg13g2_decap_8 FILLER_78_2775 ();
 sg13g2_decap_8 FILLER_78_2782 ();
 sg13g2_decap_8 FILLER_78_2789 ();
 sg13g2_decap_8 FILLER_78_2796 ();
 sg13g2_decap_8 FILLER_78_2803 ();
 sg13g2_decap_8 FILLER_78_2810 ();
 sg13g2_decap_8 FILLER_78_2817 ();
 sg13g2_decap_8 FILLER_78_2824 ();
 sg13g2_decap_8 FILLER_78_2831 ();
 sg13g2_decap_8 FILLER_78_2838 ();
 sg13g2_decap_8 FILLER_78_2845 ();
 sg13g2_decap_8 FILLER_78_2852 ();
 sg13g2_decap_8 FILLER_78_2859 ();
 sg13g2_decap_8 FILLER_78_2866 ();
 sg13g2_decap_8 FILLER_78_2873 ();
 sg13g2_decap_8 FILLER_78_2880 ();
 sg13g2_decap_8 FILLER_78_2887 ();
 sg13g2_decap_8 FILLER_78_2894 ();
 sg13g2_decap_8 FILLER_78_2901 ();
 sg13g2_decap_8 FILLER_78_2908 ();
 sg13g2_decap_8 FILLER_78_2915 ();
 sg13g2_decap_8 FILLER_78_2922 ();
 sg13g2_decap_8 FILLER_78_2929 ();
 sg13g2_decap_8 FILLER_78_2936 ();
 sg13g2_decap_8 FILLER_78_2943 ();
 sg13g2_decap_8 FILLER_78_2950 ();
 sg13g2_decap_8 FILLER_78_2957 ();
 sg13g2_decap_8 FILLER_78_2964 ();
 sg13g2_decap_8 FILLER_78_2971 ();
 sg13g2_decap_8 FILLER_78_2978 ();
 sg13g2_decap_8 FILLER_78_2985 ();
 sg13g2_decap_8 FILLER_78_2992 ();
 sg13g2_decap_8 FILLER_78_2999 ();
 sg13g2_decap_8 FILLER_78_3006 ();
 sg13g2_decap_8 FILLER_78_3013 ();
 sg13g2_decap_8 FILLER_78_3020 ();
 sg13g2_decap_8 FILLER_78_3027 ();
 sg13g2_decap_8 FILLER_78_3034 ();
 sg13g2_decap_8 FILLER_78_3041 ();
 sg13g2_decap_8 FILLER_78_3048 ();
 sg13g2_decap_8 FILLER_78_3055 ();
 sg13g2_decap_8 FILLER_78_3062 ();
 sg13g2_decap_8 FILLER_78_3069 ();
 sg13g2_decap_8 FILLER_78_3076 ();
 sg13g2_decap_8 FILLER_78_3083 ();
 sg13g2_decap_8 FILLER_78_3090 ();
 sg13g2_decap_8 FILLER_78_3097 ();
 sg13g2_decap_8 FILLER_78_3104 ();
 sg13g2_decap_8 FILLER_78_3111 ();
 sg13g2_decap_8 FILLER_78_3118 ();
 sg13g2_decap_8 FILLER_78_3125 ();
 sg13g2_decap_8 FILLER_78_3132 ();
 sg13g2_decap_8 FILLER_78_3139 ();
 sg13g2_decap_8 FILLER_78_3146 ();
 sg13g2_decap_8 FILLER_78_3153 ();
 sg13g2_decap_8 FILLER_78_3160 ();
 sg13g2_decap_8 FILLER_78_3167 ();
 sg13g2_decap_8 FILLER_78_3174 ();
 sg13g2_decap_8 FILLER_78_3181 ();
 sg13g2_decap_8 FILLER_78_3188 ();
 sg13g2_decap_8 FILLER_78_3195 ();
 sg13g2_decap_8 FILLER_78_3202 ();
 sg13g2_decap_8 FILLER_78_3209 ();
 sg13g2_decap_8 FILLER_78_3216 ();
 sg13g2_decap_8 FILLER_78_3223 ();
 sg13g2_decap_8 FILLER_78_3230 ();
 sg13g2_decap_8 FILLER_78_3237 ();
 sg13g2_decap_8 FILLER_78_3244 ();
 sg13g2_decap_8 FILLER_78_3251 ();
 sg13g2_decap_8 FILLER_78_3258 ();
 sg13g2_decap_8 FILLER_78_3265 ();
 sg13g2_decap_8 FILLER_78_3272 ();
 sg13g2_decap_8 FILLER_78_3279 ();
 sg13g2_decap_8 FILLER_78_3286 ();
 sg13g2_decap_8 FILLER_78_3293 ();
 sg13g2_decap_8 FILLER_78_3300 ();
 sg13g2_decap_8 FILLER_78_3307 ();
 sg13g2_decap_8 FILLER_78_3314 ();
 sg13g2_decap_8 FILLER_78_3321 ();
 sg13g2_decap_8 FILLER_78_3328 ();
 sg13g2_decap_8 FILLER_78_3335 ();
 sg13g2_decap_8 FILLER_78_3342 ();
 sg13g2_decap_8 FILLER_78_3349 ();
 sg13g2_decap_8 FILLER_78_3356 ();
 sg13g2_decap_8 FILLER_78_3363 ();
 sg13g2_decap_8 FILLER_78_3370 ();
 sg13g2_decap_8 FILLER_78_3377 ();
 sg13g2_decap_8 FILLER_78_3384 ();
 sg13g2_decap_8 FILLER_78_3391 ();
 sg13g2_decap_8 FILLER_78_3398 ();
 sg13g2_decap_8 FILLER_78_3405 ();
 sg13g2_decap_8 FILLER_78_3412 ();
 sg13g2_decap_8 FILLER_78_3419 ();
 sg13g2_decap_8 FILLER_78_3426 ();
 sg13g2_decap_8 FILLER_78_3433 ();
 sg13g2_decap_8 FILLER_78_3440 ();
 sg13g2_decap_8 FILLER_78_3447 ();
 sg13g2_decap_8 FILLER_78_3454 ();
 sg13g2_decap_8 FILLER_78_3461 ();
 sg13g2_decap_8 FILLER_78_3468 ();
 sg13g2_decap_8 FILLER_78_3475 ();
 sg13g2_decap_8 FILLER_78_3482 ();
 sg13g2_decap_8 FILLER_78_3489 ();
 sg13g2_decap_8 FILLER_78_3496 ();
 sg13g2_decap_8 FILLER_78_3503 ();
 sg13g2_decap_8 FILLER_78_3510 ();
 sg13g2_decap_8 FILLER_78_3517 ();
 sg13g2_decap_8 FILLER_78_3524 ();
 sg13g2_decap_8 FILLER_78_3531 ();
 sg13g2_decap_8 FILLER_78_3538 ();
 sg13g2_decap_8 FILLER_78_3545 ();
 sg13g2_decap_8 FILLER_78_3552 ();
 sg13g2_decap_8 FILLER_78_3559 ();
 sg13g2_decap_8 FILLER_78_3566 ();
 sg13g2_decap_8 FILLER_78_3573 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_354 ();
 sg13g2_decap_8 FILLER_79_361 ();
 sg13g2_decap_8 FILLER_79_368 ();
 sg13g2_decap_8 FILLER_79_375 ();
 sg13g2_decap_8 FILLER_79_382 ();
 sg13g2_decap_8 FILLER_79_389 ();
 sg13g2_decap_8 FILLER_79_396 ();
 sg13g2_decap_8 FILLER_79_403 ();
 sg13g2_decap_8 FILLER_79_410 ();
 sg13g2_decap_8 FILLER_79_417 ();
 sg13g2_decap_8 FILLER_79_424 ();
 sg13g2_decap_8 FILLER_79_431 ();
 sg13g2_decap_8 FILLER_79_438 ();
 sg13g2_decap_8 FILLER_79_445 ();
 sg13g2_decap_8 FILLER_79_452 ();
 sg13g2_decap_8 FILLER_79_459 ();
 sg13g2_decap_8 FILLER_79_466 ();
 sg13g2_decap_8 FILLER_79_473 ();
 sg13g2_decap_8 FILLER_79_480 ();
 sg13g2_decap_8 FILLER_79_487 ();
 sg13g2_decap_8 FILLER_79_494 ();
 sg13g2_decap_8 FILLER_79_501 ();
 sg13g2_decap_8 FILLER_79_508 ();
 sg13g2_decap_8 FILLER_79_515 ();
 sg13g2_decap_8 FILLER_79_522 ();
 sg13g2_decap_8 FILLER_79_529 ();
 sg13g2_decap_8 FILLER_79_536 ();
 sg13g2_decap_8 FILLER_79_543 ();
 sg13g2_decap_8 FILLER_79_550 ();
 sg13g2_decap_8 FILLER_79_557 ();
 sg13g2_decap_8 FILLER_79_564 ();
 sg13g2_decap_8 FILLER_79_571 ();
 sg13g2_decap_8 FILLER_79_578 ();
 sg13g2_decap_8 FILLER_79_585 ();
 sg13g2_decap_8 FILLER_79_592 ();
 sg13g2_decap_8 FILLER_79_599 ();
 sg13g2_decap_8 FILLER_79_606 ();
 sg13g2_decap_8 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_620 ();
 sg13g2_decap_8 FILLER_79_627 ();
 sg13g2_decap_8 FILLER_79_634 ();
 sg13g2_decap_8 FILLER_79_641 ();
 sg13g2_decap_8 FILLER_79_648 ();
 sg13g2_decap_8 FILLER_79_655 ();
 sg13g2_decap_8 FILLER_79_662 ();
 sg13g2_decap_8 FILLER_79_669 ();
 sg13g2_decap_4 FILLER_79_676 ();
 sg13g2_fill_1 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_712 ();
 sg13g2_fill_2 FILLER_79_719 ();
 sg13g2_decap_8 FILLER_79_765 ();
 sg13g2_decap_4 FILLER_79_772 ();
 sg13g2_fill_1 FILLER_79_776 ();
 sg13g2_decap_8 FILLER_79_842 ();
 sg13g2_fill_2 FILLER_79_849 ();
 sg13g2_fill_1 FILLER_79_851 ();
 sg13g2_decap_8 FILLER_79_907 ();
 sg13g2_decap_8 FILLER_79_914 ();
 sg13g2_decap_4 FILLER_79_921 ();
 sg13g2_fill_1 FILLER_79_925 ();
 sg13g2_decap_8 FILLER_79_983 ();
 sg13g2_decap_8 FILLER_79_990 ();
 sg13g2_fill_1 FILLER_79_1004 ();
 sg13g2_fill_1 FILLER_79_1021 ();
 sg13g2_decap_8 FILLER_79_1056 ();
 sg13g2_decap_8 FILLER_79_1063 ();
 sg13g2_fill_1 FILLER_79_1070 ();
 sg13g2_decap_8 FILLER_79_1105 ();
 sg13g2_decap_8 FILLER_79_1112 ();
 sg13g2_fill_2 FILLER_79_1119 ();
 sg13g2_fill_1 FILLER_79_1121 ();
 sg13g2_decap_8 FILLER_79_1163 ();
 sg13g2_decap_8 FILLER_79_1170 ();
 sg13g2_decap_8 FILLER_79_1177 ();
 sg13g2_decap_4 FILLER_79_1184 ();
 sg13g2_fill_1 FILLER_79_1188 ();
 sg13g2_decap_8 FILLER_79_1215 ();
 sg13g2_fill_1 FILLER_79_1222 ();
 sg13g2_decap_8 FILLER_79_1321 ();
 sg13g2_decap_4 FILLER_79_1328 ();
 sg13g2_decap_8 FILLER_79_1362 ();
 sg13g2_fill_2 FILLER_79_1369 ();
 sg13g2_fill_1 FILLER_79_1375 ();
 sg13g2_decap_8 FILLER_79_1458 ();
 sg13g2_decap_8 FILLER_79_1465 ();
 sg13g2_decap_8 FILLER_79_1472 ();
 sg13g2_decap_8 FILLER_79_1479 ();
 sg13g2_decap_8 FILLER_79_1486 ();
 sg13g2_decap_8 FILLER_79_1493 ();
 sg13g2_decap_8 FILLER_79_1500 ();
 sg13g2_decap_8 FILLER_79_1507 ();
 sg13g2_decap_8 FILLER_79_1514 ();
 sg13g2_decap_8 FILLER_79_1521 ();
 sg13g2_decap_8 FILLER_79_1528 ();
 sg13g2_decap_8 FILLER_79_1535 ();
 sg13g2_decap_8 FILLER_79_1542 ();
 sg13g2_decap_8 FILLER_79_1549 ();
 sg13g2_decap_8 FILLER_79_1556 ();
 sg13g2_decap_8 FILLER_79_1563 ();
 sg13g2_decap_8 FILLER_79_1570 ();
 sg13g2_decap_8 FILLER_79_1577 ();
 sg13g2_decap_8 FILLER_79_1584 ();
 sg13g2_decap_8 FILLER_79_1591 ();
 sg13g2_decap_8 FILLER_79_1598 ();
 sg13g2_decap_8 FILLER_79_1605 ();
 sg13g2_decap_8 FILLER_79_1612 ();
 sg13g2_decap_8 FILLER_79_1619 ();
 sg13g2_decap_8 FILLER_79_1626 ();
 sg13g2_decap_8 FILLER_79_1633 ();
 sg13g2_decap_8 FILLER_79_1640 ();
 sg13g2_decap_8 FILLER_79_1647 ();
 sg13g2_decap_8 FILLER_79_1654 ();
 sg13g2_decap_8 FILLER_79_1661 ();
 sg13g2_decap_8 FILLER_79_1668 ();
 sg13g2_decap_8 FILLER_79_1675 ();
 sg13g2_decap_8 FILLER_79_1682 ();
 sg13g2_decap_8 FILLER_79_1689 ();
 sg13g2_decap_8 FILLER_79_1696 ();
 sg13g2_decap_8 FILLER_79_1703 ();
 sg13g2_decap_8 FILLER_79_1710 ();
 sg13g2_decap_8 FILLER_79_1717 ();
 sg13g2_decap_8 FILLER_79_1724 ();
 sg13g2_decap_8 FILLER_79_1731 ();
 sg13g2_decap_8 FILLER_79_1738 ();
 sg13g2_decap_8 FILLER_79_1745 ();
 sg13g2_decap_8 FILLER_79_1752 ();
 sg13g2_decap_8 FILLER_79_1759 ();
 sg13g2_decap_8 FILLER_79_1766 ();
 sg13g2_decap_8 FILLER_79_1773 ();
 sg13g2_decap_8 FILLER_79_1780 ();
 sg13g2_decap_8 FILLER_79_1787 ();
 sg13g2_decap_8 FILLER_79_1794 ();
 sg13g2_decap_8 FILLER_79_1801 ();
 sg13g2_decap_8 FILLER_79_1808 ();
 sg13g2_decap_8 FILLER_79_1815 ();
 sg13g2_decap_8 FILLER_79_1822 ();
 sg13g2_decap_8 FILLER_79_1829 ();
 sg13g2_decap_8 FILLER_79_1836 ();
 sg13g2_decap_8 FILLER_79_1843 ();
 sg13g2_decap_8 FILLER_79_1850 ();
 sg13g2_decap_8 FILLER_79_1857 ();
 sg13g2_decap_8 FILLER_79_1864 ();
 sg13g2_decap_8 FILLER_79_1871 ();
 sg13g2_decap_8 FILLER_79_1878 ();
 sg13g2_decap_8 FILLER_79_1885 ();
 sg13g2_decap_8 FILLER_79_1892 ();
 sg13g2_decap_8 FILLER_79_1899 ();
 sg13g2_decap_8 FILLER_79_1906 ();
 sg13g2_decap_8 FILLER_79_1913 ();
 sg13g2_decap_8 FILLER_79_1920 ();
 sg13g2_decap_8 FILLER_79_1927 ();
 sg13g2_decap_8 FILLER_79_1934 ();
 sg13g2_decap_8 FILLER_79_1941 ();
 sg13g2_decap_8 FILLER_79_1948 ();
 sg13g2_decap_8 FILLER_79_1955 ();
 sg13g2_decap_8 FILLER_79_1962 ();
 sg13g2_decap_8 FILLER_79_1969 ();
 sg13g2_decap_8 FILLER_79_1976 ();
 sg13g2_decap_8 FILLER_79_1983 ();
 sg13g2_decap_8 FILLER_79_1990 ();
 sg13g2_decap_8 FILLER_79_1997 ();
 sg13g2_decap_8 FILLER_79_2004 ();
 sg13g2_decap_8 FILLER_79_2011 ();
 sg13g2_decap_8 FILLER_79_2018 ();
 sg13g2_decap_8 FILLER_79_2025 ();
 sg13g2_decap_8 FILLER_79_2032 ();
 sg13g2_decap_8 FILLER_79_2039 ();
 sg13g2_decap_8 FILLER_79_2046 ();
 sg13g2_decap_8 FILLER_79_2053 ();
 sg13g2_decap_8 FILLER_79_2060 ();
 sg13g2_decap_8 FILLER_79_2067 ();
 sg13g2_decap_8 FILLER_79_2074 ();
 sg13g2_decap_8 FILLER_79_2081 ();
 sg13g2_decap_8 FILLER_79_2088 ();
 sg13g2_decap_8 FILLER_79_2095 ();
 sg13g2_decap_8 FILLER_79_2102 ();
 sg13g2_decap_8 FILLER_79_2109 ();
 sg13g2_decap_8 FILLER_79_2116 ();
 sg13g2_decap_8 FILLER_79_2123 ();
 sg13g2_decap_8 FILLER_79_2130 ();
 sg13g2_decap_8 FILLER_79_2137 ();
 sg13g2_decap_8 FILLER_79_2144 ();
 sg13g2_decap_8 FILLER_79_2151 ();
 sg13g2_decap_8 FILLER_79_2158 ();
 sg13g2_decap_8 FILLER_79_2165 ();
 sg13g2_decap_8 FILLER_79_2172 ();
 sg13g2_decap_8 FILLER_79_2179 ();
 sg13g2_decap_8 FILLER_79_2186 ();
 sg13g2_decap_8 FILLER_79_2193 ();
 sg13g2_decap_8 FILLER_79_2200 ();
 sg13g2_decap_8 FILLER_79_2207 ();
 sg13g2_decap_8 FILLER_79_2214 ();
 sg13g2_decap_8 FILLER_79_2221 ();
 sg13g2_decap_8 FILLER_79_2228 ();
 sg13g2_decap_8 FILLER_79_2235 ();
 sg13g2_decap_8 FILLER_79_2242 ();
 sg13g2_decap_8 FILLER_79_2249 ();
 sg13g2_decap_8 FILLER_79_2256 ();
 sg13g2_decap_8 FILLER_79_2263 ();
 sg13g2_decap_8 FILLER_79_2270 ();
 sg13g2_decap_8 FILLER_79_2277 ();
 sg13g2_decap_8 FILLER_79_2284 ();
 sg13g2_decap_8 FILLER_79_2291 ();
 sg13g2_decap_8 FILLER_79_2298 ();
 sg13g2_decap_8 FILLER_79_2305 ();
 sg13g2_decap_8 FILLER_79_2312 ();
 sg13g2_decap_8 FILLER_79_2319 ();
 sg13g2_decap_8 FILLER_79_2326 ();
 sg13g2_decap_8 FILLER_79_2333 ();
 sg13g2_decap_8 FILLER_79_2340 ();
 sg13g2_decap_8 FILLER_79_2347 ();
 sg13g2_decap_8 FILLER_79_2354 ();
 sg13g2_decap_8 FILLER_79_2361 ();
 sg13g2_decap_8 FILLER_79_2368 ();
 sg13g2_decap_8 FILLER_79_2375 ();
 sg13g2_decap_8 FILLER_79_2382 ();
 sg13g2_decap_8 FILLER_79_2389 ();
 sg13g2_decap_8 FILLER_79_2396 ();
 sg13g2_decap_8 FILLER_79_2403 ();
 sg13g2_decap_8 FILLER_79_2410 ();
 sg13g2_decap_8 FILLER_79_2417 ();
 sg13g2_decap_8 FILLER_79_2424 ();
 sg13g2_decap_8 FILLER_79_2431 ();
 sg13g2_decap_8 FILLER_79_2438 ();
 sg13g2_decap_8 FILLER_79_2445 ();
 sg13g2_decap_8 FILLER_79_2452 ();
 sg13g2_decap_8 FILLER_79_2459 ();
 sg13g2_decap_8 FILLER_79_2466 ();
 sg13g2_decap_8 FILLER_79_2473 ();
 sg13g2_decap_8 FILLER_79_2480 ();
 sg13g2_decap_8 FILLER_79_2487 ();
 sg13g2_decap_8 FILLER_79_2494 ();
 sg13g2_decap_8 FILLER_79_2501 ();
 sg13g2_decap_8 FILLER_79_2508 ();
 sg13g2_decap_8 FILLER_79_2515 ();
 sg13g2_decap_8 FILLER_79_2522 ();
 sg13g2_decap_8 FILLER_79_2529 ();
 sg13g2_decap_8 FILLER_79_2536 ();
 sg13g2_decap_8 FILLER_79_2543 ();
 sg13g2_decap_8 FILLER_79_2550 ();
 sg13g2_decap_8 FILLER_79_2557 ();
 sg13g2_decap_8 FILLER_79_2564 ();
 sg13g2_decap_8 FILLER_79_2571 ();
 sg13g2_decap_8 FILLER_79_2578 ();
 sg13g2_decap_8 FILLER_79_2585 ();
 sg13g2_decap_8 FILLER_79_2592 ();
 sg13g2_decap_8 FILLER_79_2599 ();
 sg13g2_decap_8 FILLER_79_2606 ();
 sg13g2_decap_8 FILLER_79_2613 ();
 sg13g2_decap_8 FILLER_79_2620 ();
 sg13g2_decap_8 FILLER_79_2627 ();
 sg13g2_decap_8 FILLER_79_2634 ();
 sg13g2_decap_8 FILLER_79_2641 ();
 sg13g2_decap_8 FILLER_79_2648 ();
 sg13g2_decap_8 FILLER_79_2655 ();
 sg13g2_decap_8 FILLER_79_2662 ();
 sg13g2_decap_8 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_79_2676 ();
 sg13g2_decap_8 FILLER_79_2683 ();
 sg13g2_decap_8 FILLER_79_2690 ();
 sg13g2_decap_8 FILLER_79_2697 ();
 sg13g2_decap_8 FILLER_79_2704 ();
 sg13g2_decap_8 FILLER_79_2711 ();
 sg13g2_decap_8 FILLER_79_2718 ();
 sg13g2_decap_8 FILLER_79_2725 ();
 sg13g2_decap_8 FILLER_79_2732 ();
 sg13g2_decap_8 FILLER_79_2739 ();
 sg13g2_decap_8 FILLER_79_2746 ();
 sg13g2_decap_8 FILLER_79_2753 ();
 sg13g2_decap_8 FILLER_79_2760 ();
 sg13g2_decap_8 FILLER_79_2767 ();
 sg13g2_decap_8 FILLER_79_2774 ();
 sg13g2_decap_8 FILLER_79_2781 ();
 sg13g2_decap_8 FILLER_79_2788 ();
 sg13g2_decap_8 FILLER_79_2795 ();
 sg13g2_decap_8 FILLER_79_2802 ();
 sg13g2_decap_8 FILLER_79_2809 ();
 sg13g2_decap_8 FILLER_79_2816 ();
 sg13g2_decap_8 FILLER_79_2823 ();
 sg13g2_decap_8 FILLER_79_2830 ();
 sg13g2_decap_8 FILLER_79_2837 ();
 sg13g2_decap_8 FILLER_79_2844 ();
 sg13g2_decap_8 FILLER_79_2851 ();
 sg13g2_decap_8 FILLER_79_2858 ();
 sg13g2_decap_8 FILLER_79_2865 ();
 sg13g2_decap_8 FILLER_79_2872 ();
 sg13g2_decap_8 FILLER_79_2879 ();
 sg13g2_decap_8 FILLER_79_2886 ();
 sg13g2_decap_8 FILLER_79_2893 ();
 sg13g2_decap_8 FILLER_79_2900 ();
 sg13g2_decap_8 FILLER_79_2907 ();
 sg13g2_decap_8 FILLER_79_2914 ();
 sg13g2_decap_8 FILLER_79_2921 ();
 sg13g2_decap_8 FILLER_79_2928 ();
 sg13g2_decap_8 FILLER_79_2935 ();
 sg13g2_decap_8 FILLER_79_2942 ();
 sg13g2_decap_8 FILLER_79_2949 ();
 sg13g2_decap_8 FILLER_79_2956 ();
 sg13g2_decap_8 FILLER_79_2963 ();
 sg13g2_decap_8 FILLER_79_2970 ();
 sg13g2_decap_8 FILLER_79_2977 ();
 sg13g2_decap_8 FILLER_79_2984 ();
 sg13g2_decap_8 FILLER_79_2991 ();
 sg13g2_decap_8 FILLER_79_2998 ();
 sg13g2_decap_8 FILLER_79_3005 ();
 sg13g2_decap_8 FILLER_79_3012 ();
 sg13g2_decap_8 FILLER_79_3019 ();
 sg13g2_decap_8 FILLER_79_3026 ();
 sg13g2_decap_8 FILLER_79_3033 ();
 sg13g2_decap_8 FILLER_79_3040 ();
 sg13g2_decap_8 FILLER_79_3047 ();
 sg13g2_decap_8 FILLER_79_3054 ();
 sg13g2_decap_8 FILLER_79_3061 ();
 sg13g2_decap_8 FILLER_79_3068 ();
 sg13g2_decap_8 FILLER_79_3075 ();
 sg13g2_decap_8 FILLER_79_3082 ();
 sg13g2_decap_8 FILLER_79_3089 ();
 sg13g2_decap_8 FILLER_79_3096 ();
 sg13g2_decap_8 FILLER_79_3103 ();
 sg13g2_decap_8 FILLER_79_3110 ();
 sg13g2_decap_8 FILLER_79_3117 ();
 sg13g2_decap_8 FILLER_79_3124 ();
 sg13g2_decap_8 FILLER_79_3131 ();
 sg13g2_decap_8 FILLER_79_3138 ();
 sg13g2_decap_8 FILLER_79_3145 ();
 sg13g2_decap_8 FILLER_79_3152 ();
 sg13g2_decap_8 FILLER_79_3159 ();
 sg13g2_decap_8 FILLER_79_3166 ();
 sg13g2_decap_8 FILLER_79_3173 ();
 sg13g2_decap_8 FILLER_79_3180 ();
 sg13g2_decap_8 FILLER_79_3187 ();
 sg13g2_decap_8 FILLER_79_3194 ();
 sg13g2_decap_8 FILLER_79_3201 ();
 sg13g2_decap_8 FILLER_79_3208 ();
 sg13g2_decap_8 FILLER_79_3215 ();
 sg13g2_decap_8 FILLER_79_3222 ();
 sg13g2_decap_8 FILLER_79_3229 ();
 sg13g2_decap_8 FILLER_79_3236 ();
 sg13g2_decap_8 FILLER_79_3243 ();
 sg13g2_decap_8 FILLER_79_3250 ();
 sg13g2_decap_8 FILLER_79_3257 ();
 sg13g2_decap_8 FILLER_79_3264 ();
 sg13g2_decap_8 FILLER_79_3271 ();
 sg13g2_decap_8 FILLER_79_3278 ();
 sg13g2_decap_8 FILLER_79_3285 ();
 sg13g2_decap_8 FILLER_79_3292 ();
 sg13g2_decap_8 FILLER_79_3299 ();
 sg13g2_decap_8 FILLER_79_3306 ();
 sg13g2_decap_8 FILLER_79_3313 ();
 sg13g2_decap_8 FILLER_79_3320 ();
 sg13g2_decap_8 FILLER_79_3327 ();
 sg13g2_decap_8 FILLER_79_3334 ();
 sg13g2_decap_8 FILLER_79_3341 ();
 sg13g2_decap_8 FILLER_79_3348 ();
 sg13g2_decap_8 FILLER_79_3355 ();
 sg13g2_decap_8 FILLER_79_3362 ();
 sg13g2_decap_8 FILLER_79_3369 ();
 sg13g2_decap_8 FILLER_79_3376 ();
 sg13g2_decap_8 FILLER_79_3383 ();
 sg13g2_decap_8 FILLER_79_3390 ();
 sg13g2_decap_8 FILLER_79_3397 ();
 sg13g2_decap_8 FILLER_79_3404 ();
 sg13g2_decap_8 FILLER_79_3411 ();
 sg13g2_decap_8 FILLER_79_3418 ();
 sg13g2_decap_8 FILLER_79_3425 ();
 sg13g2_decap_8 FILLER_79_3432 ();
 sg13g2_decap_8 FILLER_79_3439 ();
 sg13g2_decap_8 FILLER_79_3446 ();
 sg13g2_decap_8 FILLER_79_3453 ();
 sg13g2_decap_8 FILLER_79_3460 ();
 sg13g2_decap_8 FILLER_79_3467 ();
 sg13g2_decap_8 FILLER_79_3474 ();
 sg13g2_decap_8 FILLER_79_3481 ();
 sg13g2_decap_8 FILLER_79_3488 ();
 sg13g2_decap_8 FILLER_79_3495 ();
 sg13g2_decap_8 FILLER_79_3502 ();
 sg13g2_decap_8 FILLER_79_3509 ();
 sg13g2_decap_8 FILLER_79_3516 ();
 sg13g2_decap_8 FILLER_79_3523 ();
 sg13g2_decap_8 FILLER_79_3530 ();
 sg13g2_decap_8 FILLER_79_3537 ();
 sg13g2_decap_8 FILLER_79_3544 ();
 sg13g2_decap_8 FILLER_79_3551 ();
 sg13g2_decap_8 FILLER_79_3558 ();
 sg13g2_decap_8 FILLER_79_3565 ();
 sg13g2_decap_8 FILLER_79_3572 ();
 sg13g2_fill_1 FILLER_79_3579 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_8 FILLER_80_164 ();
 sg13g2_decap_8 FILLER_80_171 ();
 sg13g2_decap_8 FILLER_80_178 ();
 sg13g2_decap_8 FILLER_80_185 ();
 sg13g2_decap_8 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_213 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_227 ();
 sg13g2_decap_8 FILLER_80_234 ();
 sg13g2_decap_8 FILLER_80_241 ();
 sg13g2_decap_8 FILLER_80_248 ();
 sg13g2_decap_8 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_fill_2 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_8 FILLER_80_306 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_fill_1 FILLER_80_327 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_decap_8 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_389 ();
 sg13g2_decap_8 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_403 ();
 sg13g2_decap_8 FILLER_80_410 ();
 sg13g2_decap_8 FILLER_80_417 ();
 sg13g2_decap_8 FILLER_80_424 ();
 sg13g2_decap_8 FILLER_80_431 ();
 sg13g2_decap_8 FILLER_80_438 ();
 sg13g2_decap_8 FILLER_80_445 ();
 sg13g2_decap_8 FILLER_80_452 ();
 sg13g2_decap_8 FILLER_80_459 ();
 sg13g2_decap_8 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_473 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_decap_8 FILLER_80_529 ();
 sg13g2_decap_8 FILLER_80_536 ();
 sg13g2_decap_8 FILLER_80_543 ();
 sg13g2_decap_8 FILLER_80_550 ();
 sg13g2_decap_8 FILLER_80_557 ();
 sg13g2_decap_8 FILLER_80_564 ();
 sg13g2_decap_8 FILLER_80_571 ();
 sg13g2_decap_8 FILLER_80_578 ();
 sg13g2_decap_8 FILLER_80_585 ();
 sg13g2_decap_8 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_599 ();
 sg13g2_decap_8 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_613 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_4 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_705 ();
 sg13g2_decap_8 FILLER_80_712 ();
 sg13g2_decap_8 FILLER_80_719 ();
 sg13g2_decap_4 FILLER_80_726 ();
 sg13g2_decap_8 FILLER_80_755 ();
 sg13g2_decap_8 FILLER_80_762 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_776 ();
 sg13g2_decap_4 FILLER_80_783 ();
 sg13g2_decap_8 FILLER_80_827 ();
 sg13g2_decap_8 FILLER_80_834 ();
 sg13g2_decap_8 FILLER_80_841 ();
 sg13g2_decap_8 FILLER_80_848 ();
 sg13g2_decap_8 FILLER_80_855 ();
 sg13g2_decap_8 FILLER_80_894 ();
 sg13g2_decap_8 FILLER_80_901 ();
 sg13g2_decap_8 FILLER_80_908 ();
 sg13g2_decap_8 FILLER_80_915 ();
 sg13g2_decap_8 FILLER_80_922 ();
 sg13g2_fill_2 FILLER_80_929 ();
 sg13g2_fill_1 FILLER_80_931 ();
 sg13g2_fill_2 FILLER_80_937 ();
 sg13g2_fill_1 FILLER_80_939 ();
 sg13g2_fill_2 FILLER_80_961 ();
 sg13g2_fill_1 FILLER_80_963 ();
 sg13g2_decap_8 FILLER_80_974 ();
 sg13g2_decap_8 FILLER_80_981 ();
 sg13g2_decap_8 FILLER_80_988 ();
 sg13g2_decap_8 FILLER_80_995 ();
 sg13g2_decap_8 FILLER_80_1002 ();
 sg13g2_fill_2 FILLER_80_1009 ();
 sg13g2_fill_1 FILLER_80_1011 ();
 sg13g2_fill_2 FILLER_80_1030 ();
 sg13g2_fill_1 FILLER_80_1032 ();
 sg13g2_decap_8 FILLER_80_1045 ();
 sg13g2_decap_8 FILLER_80_1052 ();
 sg13g2_decap_8 FILLER_80_1059 ();
 sg13g2_decap_8 FILLER_80_1066 ();
 sg13g2_fill_2 FILLER_80_1073 ();
 sg13g2_fill_1 FILLER_80_1075 ();
 sg13g2_decap_8 FILLER_80_1102 ();
 sg13g2_decap_8 FILLER_80_1109 ();
 sg13g2_decap_8 FILLER_80_1116 ();
 sg13g2_fill_2 FILLER_80_1123 ();
 sg13g2_fill_2 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1153 ();
 sg13g2_decap_8 FILLER_80_1160 ();
 sg13g2_decap_8 FILLER_80_1167 ();
 sg13g2_decap_8 FILLER_80_1174 ();
 sg13g2_decap_8 FILLER_80_1181 ();
 sg13g2_decap_8 FILLER_80_1188 ();
 sg13g2_decap_8 FILLER_80_1195 ();
 sg13g2_decap_8 FILLER_80_1202 ();
 sg13g2_decap_8 FILLER_80_1209 ();
 sg13g2_decap_8 FILLER_80_1216 ();
 sg13g2_decap_8 FILLER_80_1223 ();
 sg13g2_decap_8 FILLER_80_1230 ();
 sg13g2_decap_8 FILLER_80_1237 ();
 sg13g2_decap_8 FILLER_80_1244 ();
 sg13g2_fill_2 FILLER_80_1251 ();
 sg13g2_fill_2 FILLER_80_1257 ();
 sg13g2_fill_1 FILLER_80_1259 ();
 sg13g2_decap_4 FILLER_80_1264 ();
 sg13g2_fill_1 FILLER_80_1268 ();
 sg13g2_decap_4 FILLER_80_1281 ();
 sg13g2_decap_8 FILLER_80_1288 ();
 sg13g2_fill_1 FILLER_80_1299 ();
 sg13g2_decap_8 FILLER_80_1305 ();
 sg13g2_decap_8 FILLER_80_1312 ();
 sg13g2_decap_8 FILLER_80_1319 ();
 sg13g2_decap_8 FILLER_80_1326 ();
 sg13g2_fill_2 FILLER_80_1333 ();
 sg13g2_fill_1 FILLER_80_1335 ();
 sg13g2_decap_8 FILLER_80_1340 ();
 sg13g2_decap_8 FILLER_80_1351 ();
 sg13g2_decap_8 FILLER_80_1358 ();
 sg13g2_decap_8 FILLER_80_1365 ();
 sg13g2_decap_8 FILLER_80_1372 ();
 sg13g2_decap_8 FILLER_80_1379 ();
 sg13g2_decap_4 FILLER_80_1386 ();
 sg13g2_fill_1 FILLER_80_1390 ();
 sg13g2_decap_8 FILLER_80_1398 ();
 sg13g2_fill_1 FILLER_80_1405 ();
 sg13g2_fill_1 FILLER_80_1414 ();
 sg13g2_fill_2 FILLER_80_1420 ();
 sg13g2_decap_8 FILLER_80_1429 ();
 sg13g2_decap_8 FILLER_80_1436 ();
 sg13g2_decap_8 FILLER_80_1452 ();
 sg13g2_decap_8 FILLER_80_1459 ();
 sg13g2_decap_8 FILLER_80_1466 ();
 sg13g2_decap_8 FILLER_80_1473 ();
 sg13g2_decap_8 FILLER_80_1480 ();
 sg13g2_decap_8 FILLER_80_1487 ();
 sg13g2_decap_8 FILLER_80_1494 ();
 sg13g2_decap_8 FILLER_80_1501 ();
 sg13g2_decap_8 FILLER_80_1508 ();
 sg13g2_decap_8 FILLER_80_1515 ();
 sg13g2_decap_8 FILLER_80_1522 ();
 sg13g2_decap_8 FILLER_80_1529 ();
 sg13g2_decap_8 FILLER_80_1536 ();
 sg13g2_decap_8 FILLER_80_1543 ();
 sg13g2_decap_8 FILLER_80_1550 ();
 sg13g2_decap_8 FILLER_80_1557 ();
 sg13g2_decap_8 FILLER_80_1564 ();
 sg13g2_decap_8 FILLER_80_1571 ();
 sg13g2_decap_8 FILLER_80_1578 ();
 sg13g2_decap_8 FILLER_80_1585 ();
 sg13g2_decap_8 FILLER_80_1592 ();
 sg13g2_decap_8 FILLER_80_1599 ();
 sg13g2_decap_8 FILLER_80_1606 ();
 sg13g2_decap_8 FILLER_80_1613 ();
 sg13g2_decap_8 FILLER_80_1620 ();
 sg13g2_decap_8 FILLER_80_1627 ();
 sg13g2_decap_8 FILLER_80_1634 ();
 sg13g2_decap_8 FILLER_80_1641 ();
 sg13g2_decap_8 FILLER_80_1648 ();
 sg13g2_decap_8 FILLER_80_1655 ();
 sg13g2_decap_8 FILLER_80_1662 ();
 sg13g2_decap_8 FILLER_80_1669 ();
 sg13g2_decap_8 FILLER_80_1676 ();
 sg13g2_decap_8 FILLER_80_1683 ();
 sg13g2_decap_8 FILLER_80_1690 ();
 sg13g2_decap_8 FILLER_80_1697 ();
 sg13g2_decap_8 FILLER_80_1704 ();
 sg13g2_decap_8 FILLER_80_1711 ();
 sg13g2_decap_8 FILLER_80_1718 ();
 sg13g2_decap_8 FILLER_80_1725 ();
 sg13g2_decap_8 FILLER_80_1732 ();
 sg13g2_decap_8 FILLER_80_1739 ();
 sg13g2_decap_8 FILLER_80_1746 ();
 sg13g2_decap_8 FILLER_80_1753 ();
 sg13g2_decap_8 FILLER_80_1760 ();
 sg13g2_decap_8 FILLER_80_1767 ();
 sg13g2_decap_8 FILLER_80_1774 ();
 sg13g2_decap_8 FILLER_80_1781 ();
 sg13g2_decap_8 FILLER_80_1788 ();
 sg13g2_decap_8 FILLER_80_1795 ();
 sg13g2_decap_8 FILLER_80_1802 ();
 sg13g2_decap_8 FILLER_80_1809 ();
 sg13g2_decap_8 FILLER_80_1816 ();
 sg13g2_decap_8 FILLER_80_1823 ();
 sg13g2_decap_8 FILLER_80_1830 ();
 sg13g2_decap_8 FILLER_80_1837 ();
 sg13g2_decap_8 FILLER_80_1844 ();
 sg13g2_decap_8 FILLER_80_1851 ();
 sg13g2_decap_8 FILLER_80_1858 ();
 sg13g2_decap_8 FILLER_80_1865 ();
 sg13g2_decap_8 FILLER_80_1872 ();
 sg13g2_decap_8 FILLER_80_1879 ();
 sg13g2_decap_8 FILLER_80_1886 ();
 sg13g2_decap_8 FILLER_80_1893 ();
 sg13g2_decap_8 FILLER_80_1900 ();
 sg13g2_decap_8 FILLER_80_1907 ();
 sg13g2_decap_8 FILLER_80_1914 ();
 sg13g2_decap_8 FILLER_80_1921 ();
 sg13g2_decap_8 FILLER_80_1928 ();
 sg13g2_decap_8 FILLER_80_1935 ();
 sg13g2_decap_8 FILLER_80_1942 ();
 sg13g2_decap_8 FILLER_80_1949 ();
 sg13g2_decap_8 FILLER_80_1956 ();
 sg13g2_decap_8 FILLER_80_1963 ();
 sg13g2_decap_8 FILLER_80_1970 ();
 sg13g2_decap_8 FILLER_80_1977 ();
 sg13g2_decap_8 FILLER_80_1984 ();
 sg13g2_decap_8 FILLER_80_1991 ();
 sg13g2_decap_8 FILLER_80_1998 ();
 sg13g2_decap_8 FILLER_80_2005 ();
 sg13g2_decap_8 FILLER_80_2012 ();
 sg13g2_decap_8 FILLER_80_2019 ();
 sg13g2_decap_8 FILLER_80_2026 ();
 sg13g2_decap_8 FILLER_80_2033 ();
 sg13g2_decap_8 FILLER_80_2040 ();
 sg13g2_decap_8 FILLER_80_2047 ();
 sg13g2_decap_8 FILLER_80_2054 ();
 sg13g2_decap_8 FILLER_80_2061 ();
 sg13g2_decap_8 FILLER_80_2068 ();
 sg13g2_decap_8 FILLER_80_2075 ();
 sg13g2_decap_8 FILLER_80_2082 ();
 sg13g2_decap_8 FILLER_80_2089 ();
 sg13g2_decap_8 FILLER_80_2096 ();
 sg13g2_decap_8 FILLER_80_2103 ();
 sg13g2_decap_8 FILLER_80_2110 ();
 sg13g2_decap_8 FILLER_80_2117 ();
 sg13g2_decap_8 FILLER_80_2124 ();
 sg13g2_decap_8 FILLER_80_2131 ();
 sg13g2_decap_8 FILLER_80_2138 ();
 sg13g2_decap_8 FILLER_80_2145 ();
 sg13g2_decap_8 FILLER_80_2152 ();
 sg13g2_decap_8 FILLER_80_2159 ();
 sg13g2_decap_8 FILLER_80_2166 ();
 sg13g2_decap_8 FILLER_80_2173 ();
 sg13g2_decap_8 FILLER_80_2180 ();
 sg13g2_decap_8 FILLER_80_2187 ();
 sg13g2_decap_8 FILLER_80_2194 ();
 sg13g2_decap_8 FILLER_80_2201 ();
 sg13g2_decap_8 FILLER_80_2208 ();
 sg13g2_decap_8 FILLER_80_2215 ();
 sg13g2_decap_8 FILLER_80_2222 ();
 sg13g2_decap_8 FILLER_80_2229 ();
 sg13g2_decap_8 FILLER_80_2236 ();
 sg13g2_decap_8 FILLER_80_2243 ();
 sg13g2_decap_8 FILLER_80_2250 ();
 sg13g2_decap_8 FILLER_80_2257 ();
 sg13g2_decap_8 FILLER_80_2264 ();
 sg13g2_decap_8 FILLER_80_2271 ();
 sg13g2_decap_8 FILLER_80_2278 ();
 sg13g2_decap_8 FILLER_80_2285 ();
 sg13g2_decap_8 FILLER_80_2292 ();
 sg13g2_decap_8 FILLER_80_2299 ();
 sg13g2_decap_8 FILLER_80_2306 ();
 sg13g2_decap_8 FILLER_80_2313 ();
 sg13g2_decap_8 FILLER_80_2320 ();
 sg13g2_decap_8 FILLER_80_2327 ();
 sg13g2_decap_8 FILLER_80_2334 ();
 sg13g2_decap_8 FILLER_80_2341 ();
 sg13g2_decap_8 FILLER_80_2348 ();
 sg13g2_decap_8 FILLER_80_2355 ();
 sg13g2_decap_8 FILLER_80_2362 ();
 sg13g2_decap_8 FILLER_80_2369 ();
 sg13g2_decap_8 FILLER_80_2376 ();
 sg13g2_decap_8 FILLER_80_2383 ();
 sg13g2_decap_8 FILLER_80_2390 ();
 sg13g2_decap_8 FILLER_80_2397 ();
 sg13g2_decap_8 FILLER_80_2404 ();
 sg13g2_decap_8 FILLER_80_2411 ();
 sg13g2_decap_8 FILLER_80_2418 ();
 sg13g2_decap_8 FILLER_80_2425 ();
 sg13g2_decap_8 FILLER_80_2432 ();
 sg13g2_decap_8 FILLER_80_2439 ();
 sg13g2_decap_8 FILLER_80_2446 ();
 sg13g2_decap_8 FILLER_80_2453 ();
 sg13g2_decap_8 FILLER_80_2460 ();
 sg13g2_decap_8 FILLER_80_2467 ();
 sg13g2_decap_8 FILLER_80_2474 ();
 sg13g2_decap_8 FILLER_80_2481 ();
 sg13g2_decap_8 FILLER_80_2488 ();
 sg13g2_decap_8 FILLER_80_2495 ();
 sg13g2_decap_8 FILLER_80_2502 ();
 sg13g2_decap_8 FILLER_80_2509 ();
 sg13g2_decap_8 FILLER_80_2516 ();
 sg13g2_decap_8 FILLER_80_2523 ();
 sg13g2_decap_8 FILLER_80_2530 ();
 sg13g2_decap_8 FILLER_80_2537 ();
 sg13g2_decap_8 FILLER_80_2544 ();
 sg13g2_decap_8 FILLER_80_2551 ();
 sg13g2_decap_8 FILLER_80_2558 ();
 sg13g2_decap_8 FILLER_80_2565 ();
 sg13g2_decap_8 FILLER_80_2572 ();
 sg13g2_decap_8 FILLER_80_2579 ();
 sg13g2_decap_8 FILLER_80_2586 ();
 sg13g2_decap_8 FILLER_80_2593 ();
 sg13g2_decap_8 FILLER_80_2600 ();
 sg13g2_decap_8 FILLER_80_2607 ();
 sg13g2_decap_8 FILLER_80_2614 ();
 sg13g2_decap_8 FILLER_80_2621 ();
 sg13g2_decap_8 FILLER_80_2628 ();
 sg13g2_decap_8 FILLER_80_2635 ();
 sg13g2_decap_8 FILLER_80_2642 ();
 sg13g2_decap_8 FILLER_80_2649 ();
 sg13g2_decap_8 FILLER_80_2656 ();
 sg13g2_decap_8 FILLER_80_2663 ();
 sg13g2_decap_8 FILLER_80_2670 ();
 sg13g2_decap_8 FILLER_80_2677 ();
 sg13g2_decap_8 FILLER_80_2684 ();
 sg13g2_decap_8 FILLER_80_2691 ();
 sg13g2_decap_8 FILLER_80_2698 ();
 sg13g2_decap_8 FILLER_80_2705 ();
 sg13g2_decap_8 FILLER_80_2712 ();
 sg13g2_decap_8 FILLER_80_2719 ();
 sg13g2_decap_8 FILLER_80_2726 ();
 sg13g2_decap_8 FILLER_80_2733 ();
 sg13g2_decap_8 FILLER_80_2740 ();
 sg13g2_decap_8 FILLER_80_2747 ();
 sg13g2_decap_8 FILLER_80_2754 ();
 sg13g2_decap_8 FILLER_80_2761 ();
 sg13g2_decap_8 FILLER_80_2768 ();
 sg13g2_decap_8 FILLER_80_2775 ();
 sg13g2_decap_8 FILLER_80_2782 ();
 sg13g2_decap_8 FILLER_80_2789 ();
 sg13g2_decap_8 FILLER_80_2796 ();
 sg13g2_decap_8 FILLER_80_2803 ();
 sg13g2_decap_8 FILLER_80_2810 ();
 sg13g2_decap_8 FILLER_80_2817 ();
 sg13g2_decap_8 FILLER_80_2824 ();
 sg13g2_decap_8 FILLER_80_2831 ();
 sg13g2_decap_8 FILLER_80_2838 ();
 sg13g2_decap_8 FILLER_80_2845 ();
 sg13g2_decap_8 FILLER_80_2852 ();
 sg13g2_decap_8 FILLER_80_2859 ();
 sg13g2_decap_8 FILLER_80_2866 ();
 sg13g2_decap_8 FILLER_80_2873 ();
 sg13g2_decap_8 FILLER_80_2880 ();
 sg13g2_decap_8 FILLER_80_2887 ();
 sg13g2_decap_8 FILLER_80_2894 ();
 sg13g2_decap_8 FILLER_80_2901 ();
 sg13g2_decap_8 FILLER_80_2908 ();
 sg13g2_decap_8 FILLER_80_2915 ();
 sg13g2_decap_8 FILLER_80_2922 ();
 sg13g2_decap_8 FILLER_80_2929 ();
 sg13g2_decap_8 FILLER_80_2936 ();
 sg13g2_decap_8 FILLER_80_2943 ();
 sg13g2_decap_8 FILLER_80_2950 ();
 sg13g2_decap_8 FILLER_80_2957 ();
 sg13g2_decap_8 FILLER_80_2964 ();
 sg13g2_decap_8 FILLER_80_2971 ();
 sg13g2_decap_8 FILLER_80_2978 ();
 sg13g2_decap_8 FILLER_80_2985 ();
 sg13g2_decap_8 FILLER_80_2992 ();
 sg13g2_decap_8 FILLER_80_2999 ();
 sg13g2_decap_8 FILLER_80_3006 ();
 sg13g2_decap_8 FILLER_80_3013 ();
 sg13g2_decap_8 FILLER_80_3020 ();
 sg13g2_decap_8 FILLER_80_3027 ();
 sg13g2_decap_8 FILLER_80_3034 ();
 sg13g2_decap_8 FILLER_80_3041 ();
 sg13g2_decap_8 FILLER_80_3048 ();
 sg13g2_decap_8 FILLER_80_3055 ();
 sg13g2_decap_8 FILLER_80_3062 ();
 sg13g2_decap_8 FILLER_80_3069 ();
 sg13g2_decap_8 FILLER_80_3076 ();
 sg13g2_decap_8 FILLER_80_3083 ();
 sg13g2_decap_8 FILLER_80_3090 ();
 sg13g2_decap_8 FILLER_80_3097 ();
 sg13g2_decap_8 FILLER_80_3104 ();
 sg13g2_decap_8 FILLER_80_3111 ();
 sg13g2_decap_8 FILLER_80_3118 ();
 sg13g2_decap_8 FILLER_80_3125 ();
 sg13g2_decap_8 FILLER_80_3132 ();
 sg13g2_decap_8 FILLER_80_3139 ();
 sg13g2_decap_8 FILLER_80_3146 ();
 sg13g2_decap_8 FILLER_80_3153 ();
 sg13g2_decap_8 FILLER_80_3160 ();
 sg13g2_decap_8 FILLER_80_3167 ();
 sg13g2_decap_8 FILLER_80_3174 ();
 sg13g2_decap_8 FILLER_80_3181 ();
 sg13g2_decap_8 FILLER_80_3188 ();
 sg13g2_decap_8 FILLER_80_3195 ();
 sg13g2_decap_8 FILLER_80_3202 ();
 sg13g2_decap_8 FILLER_80_3209 ();
 sg13g2_decap_8 FILLER_80_3216 ();
 sg13g2_decap_8 FILLER_80_3223 ();
 sg13g2_decap_8 FILLER_80_3230 ();
 sg13g2_decap_8 FILLER_80_3237 ();
 sg13g2_decap_8 FILLER_80_3244 ();
 sg13g2_decap_8 FILLER_80_3251 ();
 sg13g2_decap_8 FILLER_80_3258 ();
 sg13g2_decap_8 FILLER_80_3265 ();
 sg13g2_decap_8 FILLER_80_3272 ();
 sg13g2_decap_8 FILLER_80_3279 ();
 sg13g2_decap_8 FILLER_80_3286 ();
 sg13g2_decap_8 FILLER_80_3293 ();
 sg13g2_decap_8 FILLER_80_3300 ();
 sg13g2_decap_8 FILLER_80_3307 ();
 sg13g2_decap_8 FILLER_80_3314 ();
 sg13g2_decap_8 FILLER_80_3321 ();
 sg13g2_decap_8 FILLER_80_3328 ();
 sg13g2_decap_8 FILLER_80_3335 ();
 sg13g2_decap_8 FILLER_80_3342 ();
 sg13g2_decap_8 FILLER_80_3349 ();
 sg13g2_decap_8 FILLER_80_3356 ();
 sg13g2_decap_8 FILLER_80_3363 ();
 sg13g2_decap_8 FILLER_80_3370 ();
 sg13g2_decap_8 FILLER_80_3377 ();
 sg13g2_decap_8 FILLER_80_3384 ();
 sg13g2_decap_8 FILLER_80_3391 ();
 sg13g2_decap_8 FILLER_80_3398 ();
 sg13g2_decap_8 FILLER_80_3405 ();
 sg13g2_decap_8 FILLER_80_3412 ();
 sg13g2_decap_8 FILLER_80_3419 ();
 sg13g2_decap_8 FILLER_80_3426 ();
 sg13g2_decap_8 FILLER_80_3433 ();
 sg13g2_decap_8 FILLER_80_3440 ();
 sg13g2_decap_8 FILLER_80_3447 ();
 sg13g2_decap_8 FILLER_80_3454 ();
 sg13g2_decap_8 FILLER_80_3461 ();
 sg13g2_decap_8 FILLER_80_3468 ();
 sg13g2_decap_8 FILLER_80_3475 ();
 sg13g2_decap_8 FILLER_80_3482 ();
 sg13g2_decap_8 FILLER_80_3489 ();
 sg13g2_decap_8 FILLER_80_3496 ();
 sg13g2_decap_8 FILLER_80_3503 ();
 sg13g2_decap_8 FILLER_80_3510 ();
 sg13g2_decap_8 FILLER_80_3517 ();
 sg13g2_decap_8 FILLER_80_3524 ();
 sg13g2_decap_8 FILLER_80_3531 ();
 sg13g2_decap_8 FILLER_80_3538 ();
 sg13g2_decap_8 FILLER_80_3545 ();
 sg13g2_decap_8 FILLER_80_3552 ();
 sg13g2_decap_8 FILLER_80_3559 ();
 sg13g2_decap_8 FILLER_80_3566 ();
 sg13g2_decap_8 FILLER_80_3573 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net940;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule

module tt_um_rejunity_vga_test01 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire \center_x[0] ;
 wire \center_x[1] ;
 wire \center_x[2] ;
 wire \center_x[3] ;
 wire \center_x[4] ;
 wire \center_x[5] ;
 wire \center_y[0] ;
 wire \envelopeA[0] ;
 wire \frame_counter[7] ;
 wire \frame_counter[8] ;
 wire \frame_counter[9] ;
 wire frame_counter_frac;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire noise;
 wire \noise_counter[0] ;
 wire \noise_counter[1] ;
 wire \noise_counter[2] ;
 wire note;
 wire note2;
 wire \note2_counter[0] ;
 wire \note2_counter[1] ;
 wire \note2_counter[2] ;
 wire \note2_counter[3] ;
 wire \note2_counter[4] ;
 wire \note2_counter[5] ;
 wire \note2_counter[6] ;
 wire \note2_counter[7] ;
 wire \note2_counter[8] ;
 wire \note2_freq[0] ;
 wire \note2_freq[1] ;
 wire \note2_freq[3] ;
 wire \note2_freq[4] ;
 wire \note2_freq[5] ;
 wire \note2_freq[6] ;
 wire \note2_freq[7] ;
 wire \note2_freq[8] ;
 wire \note_counter[0] ;
 wire \note_counter[1] ;
 wire \note_counter[2] ;
 wire \note_counter[3] ;
 wire \note_counter[4] ;
 wire \note_counter[5] ;
 wire \note_counter[6] ;
 wire \note_counter[7] ;
 wire \note_freq[0] ;
 wire \note_freq[1] ;
 wire \note_freq[2] ;
 wire \note_freq[4] ;
 wire \note_freq[5] ;
 wire \note_freq[6] ;
 wire \note_freq[7] ;
 wire \r1[0] ;
 wire \r1[10] ;
 wire \r1[11] ;
 wire \r1[12] ;
 wire \r1[13] ;
 wire \r1[14] ;
 wire \r1[15] ;
 wire \r1[16] ;
 wire \r1[17] ;
 wire \r1[1] ;
 wire \r1[2] ;
 wire \r1[3] ;
 wire \r1[4] ;
 wire \r1[5] ;
 wire \r1[6] ;
 wire \r1[7] ;
 wire \r1[8] ;
 wire \r1[9] ;
 wire \r2[0] ;
 wire \r2[10] ;
 wire \r2[11] ;
 wire \r2[12] ;
 wire \r2[13] ;
 wire \r2[14] ;
 wire \r2[15] ;
 wire \r2[16] ;
 wire \r2[17] ;
 wire \r2[18] ;
 wire \r2[1] ;
 wire \r2[2] ;
 wire \r2[3] ;
 wire \r2[4] ;
 wire \r2[5] ;
 wire \r2[6] ;
 wire \r2[7] ;
 wire \r2[8] ;
 wire \r2[9] ;
 wire \title_r[0] ;
 wire \title_r[10] ;
 wire \title_r[11] ;
 wire \title_r[12] ;
 wire \title_r[13] ;
 wire \title_r[1] ;
 wire \title_r[2] ;
 wire \title_r[3] ;
 wire \title_r[4] ;
 wire \title_r[5] ;
 wire \title_r[6] ;
 wire \title_r[7] ;
 wire \title_r[8] ;
 wire \title_r[9] ;
 wire \title_r_pixels_in_scanline[0] ;
 wire \title_r_pixels_in_scanline[1] ;
 wire \title_r_pixels_in_scanline[2] ;
 wire \title_r_pixels_in_scanline[3] ;
 wire \title_r_pixels_in_scanline[4] ;
 wire \title_r_pixels_in_scanline[5] ;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire clknet_0_clk;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net1;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;

 sg13g2_inv_1 _3843_ (.Y(_2356_),
    .A(\title_r[10] ));
 sg13g2_inv_1 _3844_ (.Y(_2367_),
    .A(\title_r[9] ));
 sg13g2_inv_1 _3845_ (.Y(_2377_),
    .A(net162));
 sg13g2_inv_2 _3846_ (.Y(_2388_),
    .A(net229));
 sg13g2_inv_4 _3847_ (.A(net854),
    .Y(_2397_));
 sg13g2_inv_4 _3848_ (.A(net863),
    .Y(_2407_));
 sg13g2_inv_2 _3849_ (.Y(_2416_),
    .A(net869));
 sg13g2_inv_2 _3850_ (.Y(_2427_),
    .A(net875));
 sg13g2_inv_4 _3851_ (.A(net878),
    .Y(_2437_));
 sg13g2_inv_2 _3852_ (.Y(_2445_),
    .A(net888));
 sg13g2_inv_1 _3853_ (.Y(_2456_),
    .A(\center_y[0] ));
 sg13g2_inv_1 _3854_ (.Y(_2465_),
    .A(note));
 sg13g2_inv_1 _3855_ (.Y(_2473_),
    .A(net219));
 sg13g2_inv_1 _3856_ (.Y(_2480_),
    .A(\note_counter[6] ));
 sg13g2_inv_1 _3857_ (.Y(_2490_),
    .A(\note_counter[4] ));
 sg13g2_inv_1 _3858_ (.Y(_2500_),
    .A(\note_counter[2] ));
 sg13g2_inv_1 _3859_ (.Y(_2507_),
    .A(note2));
 sg13g2_inv_1 _3860_ (.Y(_2514_),
    .A(net216));
 sg13g2_inv_1 _3861_ (.Y(_2522_),
    .A(\note2_counter[7] ));
 sg13g2_inv_1 _3862_ (.Y(_2529_),
    .A(\note2_counter[6] ));
 sg13g2_inv_1 _3863_ (.Y(_2536_),
    .A(\note2_counter[5] ));
 sg13g2_inv_1 _3864_ (.Y(_2543_),
    .A(\note2_counter[4] ));
 sg13g2_inv_1 _3865_ (.Y(_2550_),
    .A(net243));
 sg13g2_inv_2 _3866_ (.Y(_2557_),
    .A(net221));
 sg13g2_inv_2 _3867_ (.Y(_2568_),
    .A(net916));
 sg13g2_inv_2 _3868_ (.Y(_2579_),
    .A(net914));
 sg13g2_inv_2 _3869_ (.Y(_2590_),
    .A(net908));
 sg13g2_inv_2 _3870_ (.Y(_2601_),
    .A(net905));
 sg13g2_inv_1 _3871_ (.Y(_2611_),
    .A(net899));
 sg13g2_inv_2 _3872_ (.Y(_2622_),
    .A(\hvsync_gen.hpos[9] ));
 sg13g2_inv_2 _3873_ (.Y(_2633_),
    .A(net896));
 sg13g2_inv_1 _3874_ (.Y(_2644_),
    .A(net837));
 sg13g2_inv_1 _3875_ (.Y(_2654_),
    .A(net831));
 sg13g2_inv_1 _3876_ (.Y(_2664_),
    .A(net833));
 sg13g2_inv_1 _3877_ (.Y(_2675_),
    .A(net259));
 sg13g2_inv_2 _3878_ (.Y(_2685_),
    .A(net926));
 sg13g2_inv_4 _3879_ (.A(_0020_),
    .Y(_2695_));
 sg13g2_inv_1 _3880_ (.Y(_2705_),
    .A(\note2_freq[5] ));
 sg13g2_inv_1 _3881_ (.Y(_2716_),
    .A(\note2_freq[4] ));
 sg13g2_inv_1 _3882_ (.Y(_2726_),
    .A(\note2_freq[3] ));
 sg13g2_inv_1 _3883_ (.Y(_2737_),
    .A(\note_freq[4] ));
 sg13g2_inv_1 _3884_ (.Y(_2747_),
    .A(\note_freq[1] ));
 sg13g2_inv_1 _3885_ (.Y(_2757_),
    .A(\note_freq[2] ));
 sg13g2_inv_1 _3886_ (.Y(_2767_),
    .A(_0031_));
 sg13g2_inv_1 _3887_ (.Y(_2778_),
    .A(\r1[10] ));
 sg13g2_inv_1 _3888_ (.Y(_2789_),
    .A(_0038_));
 sg13g2_inv_1 _3889_ (.Y(_2799_),
    .A(_0037_));
 sg13g2_inv_1 _3890_ (.Y(_2810_),
    .A(_0039_));
 sg13g2_inv_1 _3891_ (.Y(_2820_),
    .A(_0040_));
 sg13g2_inv_1 _3892_ (.Y(_2831_),
    .A(_0041_));
 sg13g2_inv_1 _3893_ (.Y(_2841_),
    .A(\r1[1] ));
 sg13g2_inv_1 _3894_ (.Y(_2851_),
    .A(_0043_));
 sg13g2_inv_1 _3895_ (.Y(_2861_),
    .A(_0044_));
 sg13g2_inv_1 _3896_ (.Y(_2871_),
    .A(_0045_));
 sg13g2_inv_1 _3897_ (.Y(_2881_),
    .A(\r2[13] ));
 sg13g2_inv_1 _3898_ (.Y(_2892_),
    .A(_0047_));
 sg13g2_inv_1 _3899_ (.Y(_2902_),
    .A(\r2[11] ));
 sg13g2_inv_1 _3900_ (.Y(_2911_),
    .A(_0048_));
 sg13g2_inv_1 _3901_ (.Y(_2921_),
    .A(_0049_));
 sg13g2_inv_1 _3902_ (.Y(_2930_),
    .A(_0050_));
 sg13g2_inv_1 _3903_ (.Y(_2940_),
    .A(\r2[7] ));
 sg13g2_inv_1 _3904_ (.Y(_2949_),
    .A(_0052_));
 sg13g2_inv_1 _3905_ (.Y(_2959_),
    .A(_0054_));
 sg13g2_inv_2 _3906_ (.Y(_2969_),
    .A(net892));
 sg13g2_inv_1 _3907_ (.Y(_2979_),
    .A(\r1[16] ));
 sg13g2_inv_1 _3908_ (.Y(_2989_),
    .A(net248));
 sg13g2_inv_1 _3909_ (.Y(_2998_),
    .A(_0016_));
 sg13g2_inv_1 _3910_ (.Y(_3007_),
    .A(\title_r_pixels_in_scanline[0] ));
 sg13g2_inv_2 _3911_ (.Y(_3015_),
    .A(_0019_));
 sg13g2_inv_1 _3912_ (.Y(_3024_),
    .A(_0021_));
 sg13g2_nor2_2 _3913_ (.A(_2675_),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_3032_));
 sg13g2_nand2_1 _3914_ (.Y(_3040_),
    .A(net838),
    .B(_3032_));
 sg13g2_nand2_1 _3915_ (.Y(_3045_),
    .A(net832),
    .B(net827));
 sg13g2_nand4_1 _3916_ (.B(_2644_),
    .C(_2664_),
    .A(net835),
    .Y(_3046_),
    .D(net830));
 sg13g2_nor3_1 _3917_ (.A(_3040_),
    .B(net234),
    .C(_3046_),
    .Y(_0011_));
 sg13g2_nor2_1 _3918_ (.A(_2622_),
    .B(\hvsync_gen.hpos[8] ),
    .Y(_3047_));
 sg13g2_nand2_1 _3919_ (.Y(_3048_),
    .A(net897),
    .B(net900));
 sg13g2_nand4_1 _3920_ (.B(net903),
    .C(net898),
    .A(net907),
    .Y(_3049_),
    .D(net900));
 sg13g2_a21oi_1 _3921_ (.A1(_3047_),
    .A2(_3049_),
    .Y(_3050_),
    .B1(net213));
 sg13g2_nor2_1 _3922_ (.A(net898),
    .B(net896),
    .Y(_3051_));
 sg13g2_nor2_1 _3923_ (.A(_2622_),
    .B(_3051_),
    .Y(_3052_));
 sg13g2_o21ai_1 _3924_ (.B1(\hvsync_gen.hpos[9] ),
    .Y(_3053_),
    .A1(net897),
    .A2(\hvsync_gen.hpos[8] ));
 sg13g2_nor2_1 _3925_ (.A(_2622_),
    .B(_2633_),
    .Y(_3054_));
 sg13g2_nor4_1 _3926_ (.A(net907),
    .B(net903),
    .C(net900),
    .D(_3054_),
    .Y(_3055_));
 sg13g2_nor3_2 _3927_ (.A(net214),
    .B(_3053_),
    .C(_3055_),
    .Y(_0010_));
 sg13g2_nand4_1 _3928_ (.B(_2568_),
    .C(_2579_),
    .A(_2557_),
    .Y(_3056_),
    .D(_2601_));
 sg13g2_nor3_2 _3929_ (.A(net911),
    .B(net907),
    .C(_3056_),
    .Y(_3057_));
 sg13g2_nor2_2 _3930_ (.A(net897),
    .B(net901),
    .Y(_3058_));
 sg13g2_nor2_1 _3931_ (.A(\hvsync_gen.hpos[9] ),
    .B(net896),
    .Y(_3059_));
 sg13g2_and3_1 _3932_ (.X(_3060_),
    .A(_3057_),
    .B(_3058_),
    .C(_3059_));
 sg13g2_nand3_1 _3933_ (.B(_3058_),
    .C(_3059_),
    .A(_3057_),
    .Y(_3061_));
 sg13g2_nor4_2 _3934_ (.A(net831),
    .B(net833),
    .C(net830),
    .Y(_3062_),
    .D(net826));
 sg13g2_nor2_1 _3935_ (.A(net840),
    .B(net838),
    .Y(_3063_));
 sg13g2_nor4_1 _3936_ (.A(net840),
    .B(net838),
    .C(net835),
    .D(net837),
    .Y(_3064_));
 sg13g2_nor2_1 _3937_ (.A(\hvsync_gen.vpos[8] ),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_3065_));
 sg13g2_nand3_1 _3938_ (.B(_3064_),
    .C(_3065_),
    .A(_3062_),
    .Y(_3066_));
 sg13g2_nor2_1 _3939_ (.A(net767),
    .B(_3066_),
    .Y(_3067_));
 sg13g2_or2_2 _3940_ (.X(_3068_),
    .B(_3066_),
    .A(net767));
 sg13g2_nand4_1 _3941_ (.B(net879),
    .C(net885),
    .A(net849),
    .Y(_3069_),
    .D(net894));
 sg13g2_or3_1 _3942_ (.A(net818),
    .B(net817),
    .C(_3069_),
    .X(_3070_));
 sg13g2_nor2_1 _3943_ (.A(net861),
    .B(_3070_),
    .Y(_3071_));
 sg13g2_a21oi_1 _3944_ (.A1(net861),
    .A2(_3070_),
    .Y(_3072_),
    .B1(_3068_));
 sg13g2_nand2b_1 _3945_ (.Y(_3073_),
    .B(_3072_),
    .A_N(_3071_));
 sg13g2_o21ai_1 _3946_ (.B1(_3073_),
    .Y(_3074_),
    .A1(net861),
    .A2(net753));
 sg13g2_inv_1 _3947_ (.Y(_3075_),
    .A(_3074_));
 sg13g2_nand2_2 _3948_ (.Y(_0002_),
    .A(net926),
    .B(_3074_));
 sg13g2_nor2_1 _3949_ (.A(_0032_),
    .B(_3069_),
    .Y(_3076_));
 sg13g2_and2_1 _3950_ (.A(_0032_),
    .B(_3069_),
    .X(_3077_));
 sg13g2_nor3_1 _3951_ (.A(_3068_),
    .B(_3076_),
    .C(_3077_),
    .Y(_3078_));
 sg13g2_inv_1 _3952_ (.Y(_3079_),
    .A(_3078_));
 sg13g2_o21ai_1 _3953_ (.B1(_3079_),
    .Y(_3080_),
    .A1(_0032_),
    .A2(net753));
 sg13g2_inv_1 _3954_ (.Y(_3081_),
    .A(_3080_));
 sg13g2_xnor2_1 _3955_ (.Y(_3082_),
    .A(net262),
    .B(_3076_));
 sg13g2_nand2_1 _3956_ (.Y(_3083_),
    .A(net753),
    .B(_3082_));
 sg13g2_o21ai_1 _3957_ (.B1(_3083_),
    .Y(_3084_),
    .A1(_0031_),
    .A2(net753));
 sg13g2_and2_1 _3958_ (.A(net926),
    .B(_3084_),
    .X(_3085_));
 sg13g2_nor2_1 _3959_ (.A(_0002_),
    .B(_3080_),
    .Y(_3086_));
 sg13g2_a21oi_1 _3960_ (.A1(_3081_),
    .A2(_3085_),
    .Y(_0006_),
    .B1(_3086_));
 sg13g2_nor2_2 _3961_ (.A(net853),
    .B(_0002_),
    .Y(_3087_));
 sg13g2_nor3_1 _3962_ (.A(net853),
    .B(_0002_),
    .C(_3080_),
    .Y(_3088_));
 sg13g2_o21ai_1 _3963_ (.B1(_3081_),
    .Y(_0005_),
    .A1(_3085_),
    .A2(_3087_));
 sg13g2_xnor2_1 _3964_ (.Y(_3089_),
    .A(net853),
    .B(_3071_));
 sg13g2_nand2_1 _3965_ (.Y(_3090_),
    .A(net753),
    .B(_3089_));
 sg13g2_o21ai_1 _3966_ (.B1(_3090_),
    .Y(_3091_),
    .A1(net853),
    .A2(net753));
 sg13g2_nor3_1 _3967_ (.A(_0002_),
    .B(_3084_),
    .C(_3091_),
    .Y(_3092_));
 sg13g2_nor3_1 _3968_ (.A(net920),
    .B(_3081_),
    .C(_3092_),
    .Y(_3093_));
 sg13g2_a21oi_1 _3969_ (.A1(_3081_),
    .A2(_3092_),
    .Y(_0007_),
    .B1(_3093_));
 sg13g2_a21oi_1 _3970_ (.A1(net926),
    .A2(_3080_),
    .Y(_3094_),
    .B1(_3085_));
 sg13g2_or2_1 _3971_ (.X(_0009_),
    .B(_3094_),
    .A(_3088_));
 sg13g2_inv_1 _3972_ (.Y(_0008_),
    .A(_0009_));
 sg13g2_nor2_1 _3973_ (.A(_2397_),
    .B(_2407_),
    .Y(_3095_));
 sg13g2_nand2_2 _3974_ (.Y(_3096_),
    .A(net854),
    .B(net862));
 sg13g2_or3_2 _3975_ (.A(_3068_),
    .B(_3070_),
    .C(_3096_),
    .X(_3097_));
 sg13g2_nor2_1 _3976_ (.A(_0030_),
    .B(_3097_),
    .Y(_3098_));
 sg13g2_o21ai_1 _3977_ (.B1(net926),
    .Y(_3099_),
    .A1(_0030_),
    .A2(_3097_));
 sg13g2_a21oi_2 _3978_ (.B1(_3099_),
    .Y(_3100_),
    .A2(_3097_),
    .A1(_0030_));
 sg13g2_nand2_1 _3979_ (.Y(_0185_),
    .A(_3087_),
    .B(_3100_));
 sg13g2_nand3_1 _3980_ (.B(_3075_),
    .C(_3091_),
    .A(net926),
    .Y(_3101_));
 sg13g2_or2_1 _3981_ (.X(_0184_),
    .B(_3101_),
    .A(_3100_));
 sg13g2_nand2_1 _3982_ (.Y(_3102_),
    .A(_0185_),
    .B(_0184_));
 sg13g2_inv_1 _3983_ (.Y(_0000_),
    .A(_3102_));
 sg13g2_nand2_1 _3984_ (.Y(_3103_),
    .A(_3091_),
    .B(_3100_));
 sg13g2_and2_1 _3985_ (.A(_0002_),
    .B(_3103_),
    .X(_0001_));
 sg13g2_a21o_1 _3986_ (.A2(_3100_),
    .A1(_3087_),
    .B1(_0001_),
    .X(_0003_));
 sg13g2_nand2_1 _3987_ (.Y(_0004_),
    .A(_3101_),
    .B(_3103_));
 sg13g2_nand3_1 _3988_ (.B(_3091_),
    .C(_3100_),
    .A(_3075_),
    .Y(_0061_));
 sg13g2_nand2_1 _3989_ (.Y(_0062_),
    .A(_3087_),
    .B(_3094_));
 sg13g2_nor2b_1 _3990_ (.A(net822),
    .B_N(\r2[0] ),
    .Y(_3104_));
 sg13g2_nor2_1 _3991_ (.A(net798),
    .B(_3066_),
    .Y(_3105_));
 sg13g2_nand2b_2 _3992_ (.Y(_3106_),
    .B(net811),
    .A_N(_3066_));
 sg13g2_nor2_1 _3993_ (.A(_2397_),
    .B(net904),
    .Y(_3107_));
 sg13g2_a21oi_1 _3994_ (.A1(net866),
    .A2(_2590_),
    .Y(_3108_),
    .B1(_3107_));
 sg13g2_nor2_1 _3995_ (.A(net818),
    .B(net910),
    .Y(_3109_));
 sg13g2_nand2_1 _3996_ (.Y(_3110_),
    .A(net818),
    .B(net910));
 sg13g2_nand2b_1 _3997_ (.Y(_3111_),
    .B(_3110_),
    .A_N(_3109_));
 sg13g2_nor2_1 _3998_ (.A(net817),
    .B(\hvsync_gen.hpos[2] ),
    .Y(_3112_));
 sg13g2_nand2_1 _3999_ (.Y(_3113_),
    .A(net817),
    .B(net914));
 sg13g2_nand2b_1 _4000_ (.Y(_3114_),
    .B(_3113_),
    .A_N(_3112_));
 sg13g2_nor2_1 _4001_ (.A(_3111_),
    .B(_3114_),
    .Y(_3115_));
 sg13g2_nor2_1 _4002_ (.A(net880),
    .B(_2557_),
    .Y(_3116_));
 sg13g2_nand2_1 _4003_ (.Y(_3117_),
    .A(net880),
    .B(_2557_));
 sg13g2_nor2_1 _4004_ (.A(net889),
    .B(_2568_),
    .Y(_3118_));
 sg13g2_a21oi_1 _4005_ (.A1(_3117_),
    .A2(_3118_),
    .Y(_3119_),
    .B1(_3116_));
 sg13g2_a221oi_1 _4006_ (.B2(_3119_),
    .C1(_3109_),
    .B1(_3115_),
    .A1(_3110_),
    .Y(_3120_),
    .A2(_3112_));
 sg13g2_nor2_1 _4007_ (.A(net866),
    .B(_2590_),
    .Y(_3121_));
 sg13g2_xnor2_1 _4008_ (.Y(_3122_),
    .A(net866),
    .B(net908));
 sg13g2_o21ai_1 _4009_ (.B1(_3108_),
    .Y(_3123_),
    .A1(_3120_),
    .A2(_3121_));
 sg13g2_nor2_1 _4010_ (.A(net896),
    .B(_3053_),
    .Y(_3124_));
 sg13g2_nand2_2 _4011_ (.Y(_3125_),
    .A(_2633_),
    .B(net799));
 sg13g2_nor2_1 _4012_ (.A(net858),
    .B(_2601_),
    .Y(_3126_));
 sg13g2_nand2_1 _4013_ (.Y(_3127_),
    .A(_2397_),
    .B(net904));
 sg13g2_nor2b_1 _4014_ (.A(net900),
    .B_N(net898),
    .Y(_3128_));
 sg13g2_nor2_1 _4015_ (.A(_0033_),
    .B(_3126_),
    .Y(_3129_));
 sg13g2_nand4_1 _4016_ (.B(net795),
    .C(_3128_),
    .A(_3123_),
    .Y(_3130_),
    .D(_3129_));
 sg13g2_inv_2 _4017_ (.Y(_3131_),
    .A(net731));
 sg13g2_xnor2_1 _4018_ (.Y(_3132_),
    .A(net884),
    .B(\r2[0] ));
 sg13g2_nand2_1 _4019_ (.Y(_3133_),
    .A(_3057_),
    .B(_3128_));
 sg13g2_nor3_1 _4020_ (.A(_2622_),
    .B(net896),
    .C(_3133_),
    .Y(_3134_));
 sg13g2_nand3_1 _4021_ (.B(_3057_),
    .C(_3128_),
    .A(_3047_),
    .Y(_3135_));
 sg13g2_nor2_1 _4022_ (.A(net811),
    .B(net752),
    .Y(_3136_));
 sg13g2_nand2_2 _4023_ (.Y(_3137_),
    .A(net798),
    .B(net766));
 sg13g2_a21oi_1 _4024_ (.A1(_3104_),
    .A2(net732),
    .Y(_3138_),
    .B1(_3137_));
 sg13g2_o21ai_1 _4025_ (.B1(_3138_),
    .Y(_3139_),
    .A1(net732),
    .A2(_3132_));
 sg13g2_nand4_1 _4026_ (.B(net830),
    .C(net826),
    .A(net831),
    .Y(_3140_),
    .D(\hvsync_gen.vpos[8] ));
 sg13g2_nor2b_1 _4027_ (.A(\hvsync_gen.vpos[9] ),
    .B_N(_3140_),
    .Y(_3141_));
 sg13g2_and2_2 _4028_ (.A(_3053_),
    .B(_3141_),
    .X(_3142_));
 sg13g2_nand2_1 _4029_ (.Y(_3143_),
    .A(net811),
    .B(_3141_));
 sg13g2_and2_1 _4030_ (.A(net767),
    .B(_3141_),
    .X(_3144_));
 sg13g2_nor2_1 _4031_ (.A(net768),
    .B(_3143_),
    .Y(_3145_));
 sg13g2_nand2_1 _4032_ (.Y(_3146_),
    .A(net767),
    .B(_3142_));
 sg13g2_nor2_1 _4033_ (.A(net777),
    .B(net752),
    .Y(_3147_));
 sg13g2_nand2_2 _4034_ (.Y(_3148_),
    .A(net774),
    .B(net766));
 sg13g2_a21oi_1 _4035_ (.A1(net287),
    .A2(net750),
    .Y(_3149_),
    .B1(_3148_));
 sg13g2_a22oi_1 _4036_ (.Y(_3150_),
    .B1(_3139_),
    .B2(_3149_),
    .A2(net778),
    .A1(_3104_));
 sg13g2_nor2_2 _4037_ (.A(_3136_),
    .B(net749),
    .Y(_3151_));
 sg13g2_nand2_1 _4038_ (.Y(_3152_),
    .A(_3137_),
    .B(net748));
 sg13g2_o21ai_1 _4039_ (.B1(net928),
    .Y(_3153_),
    .A1(_3104_),
    .A2(_3152_));
 sg13g2_nor2_1 _4040_ (.A(_3150_),
    .B(_3153_),
    .Y(_0063_));
 sg13g2_nor2b_1 _4041_ (.A(net823),
    .B_N(\r2[1] ),
    .Y(_3154_));
 sg13g2_nand2_1 _4042_ (.Y(_3155_),
    .A(net778),
    .B(_3154_));
 sg13g2_nand2_1 _4043_ (.Y(_3156_),
    .A(net878),
    .B(\r2[1] ));
 sg13g2_xor2_1 _4044_ (.B(\r2[1] ),
    .A(net879),
    .X(_3157_));
 sg13g2_nand3_1 _4045_ (.B(\r2[0] ),
    .C(_3157_),
    .A(net884),
    .Y(_3158_));
 sg13g2_a21o_1 _4046_ (.A2(\r2[0] ),
    .A1(net884),
    .B1(_3157_),
    .X(_3159_));
 sg13g2_nand3_1 _4047_ (.B(_3158_),
    .C(_3159_),
    .A(net728),
    .Y(_3160_));
 sg13g2_a21oi_1 _4048_ (.A1(net733),
    .A2(_3154_),
    .Y(_3161_),
    .B1(_3137_));
 sg13g2_nand2_1 _4049_ (.Y(_3162_),
    .A(_3160_),
    .B(_3161_));
 sg13g2_nand2_2 _4050_ (.Y(_3163_),
    .A(net889),
    .B(_2568_));
 sg13g2_nor2b_2 _4051_ (.A(_3118_),
    .B_N(_3163_),
    .Y(_3164_));
 sg13g2_nand2b_2 _4052_ (.Y(_3165_),
    .B(_3163_),
    .A_N(_3118_));
 sg13g2_nor2_1 _4053_ (.A(_0023_),
    .B(_3164_),
    .Y(_3166_));
 sg13g2_xnor2_1 _4054_ (.Y(_3167_),
    .A(_0023_),
    .B(_3165_));
 sg13g2_xnor2_1 _4055_ (.Y(_3168_),
    .A(\r2[0] ),
    .B(_3167_));
 sg13g2_nor3_1 _4056_ (.A(net799),
    .B(_3144_),
    .C(_3154_),
    .Y(_3169_));
 sg13g2_a21oi_1 _4057_ (.A1(net750),
    .A2(_3168_),
    .Y(_3170_),
    .B1(_3169_));
 sg13g2_nand3_1 _4058_ (.B(_3162_),
    .C(_3170_),
    .A(net738),
    .Y(_3171_));
 sg13g2_a21oi_1 _4059_ (.A1(_3155_),
    .A2(_3171_),
    .Y(_0064_),
    .B1(net921));
 sg13g2_nor2b_1 _4060_ (.A(net823),
    .B_N(net267),
    .Y(_3172_));
 sg13g2_nor2_2 _4061_ (.A(net732),
    .B(_3137_),
    .Y(_3173_));
 sg13g2_nor2_1 _4062_ (.A(net750),
    .B(_3173_),
    .Y(_3174_));
 sg13g2_nand2_1 _4063_ (.Y(_3175_),
    .A(_3172_),
    .B(_3174_));
 sg13g2_a21oi_1 _4064_ (.A1(\r2[0] ),
    .A2(_3167_),
    .Y(_3176_),
    .B1(_3166_));
 sg13g2_nand2b_1 _4065_ (.Y(_3177_),
    .B(_3117_),
    .A_N(_3116_));
 sg13g2_xnor2_1 _4066_ (.Y(_3178_),
    .A(_3163_),
    .B(_3177_));
 sg13g2_xnor2_1 _4067_ (.Y(_3179_),
    .A(\r2[2] ),
    .B(net763));
 sg13g2_nor2_1 _4068_ (.A(_3176_),
    .B(_3179_),
    .Y(_3180_));
 sg13g2_xor2_1 _4069_ (.B(_3179_),
    .A(_3176_),
    .X(_3181_));
 sg13g2_nand2_1 _4070_ (.Y(_3182_),
    .A(net874),
    .B(\r2[2] ));
 sg13g2_xnor2_1 _4071_ (.Y(_3183_),
    .A(net874),
    .B(\r2[2] ));
 sg13g2_a21o_1 _4072_ (.A2(_3158_),
    .A1(_3156_),
    .B1(_3183_),
    .X(_3184_));
 sg13g2_nand3_1 _4073_ (.B(_3158_),
    .C(_3183_),
    .A(_3156_),
    .Y(_3185_));
 sg13g2_and2_1 _4074_ (.A(_3184_),
    .B(_3185_),
    .X(_3186_));
 sg13g2_a22oi_1 _4075_ (.Y(_3187_),
    .B1(_3186_),
    .B2(_3173_),
    .A2(_3181_),
    .A1(net750));
 sg13g2_nand2_1 _4076_ (.Y(_3188_),
    .A(_3175_),
    .B(_3187_));
 sg13g2_a22oi_1 _4077_ (.Y(_3189_),
    .B1(_3188_),
    .B2(net738),
    .A2(_3172_),
    .A1(net779));
 sg13g2_nor2_1 _4078_ (.A(net920),
    .B(_3189_),
    .Y(_0065_));
 sg13g2_nor2b_1 _4079_ (.A(net824),
    .B_N(\r2[3] ),
    .Y(_3190_));
 sg13g2_a21oi_2 _4080_ (.B1(_3116_),
    .Y(_3191_),
    .A2(_3163_),
    .A1(_3117_));
 sg13g2_inv_1 _4081_ (.Y(_3192_),
    .A(_3191_));
 sg13g2_xnor2_1 _4082_ (.Y(_3193_),
    .A(_3114_),
    .B(_3191_));
 sg13g2_inv_2 _4083_ (.Y(_3194_),
    .A(_3193_));
 sg13g2_nand2_1 _4084_ (.Y(_3195_),
    .A(\r2[3] ),
    .B(_3194_));
 sg13g2_xor2_1 _4085_ (.B(_3193_),
    .A(\r2[3] ),
    .X(_3196_));
 sg13g2_a21oi_1 _4086_ (.A1(_2959_),
    .A2(net763),
    .Y(_3197_),
    .B1(_3180_));
 sg13g2_or2_1 _4087_ (.X(_3198_),
    .B(_3197_),
    .A(_3196_));
 sg13g2_xnor2_1 _4088_ (.Y(_3199_),
    .A(_3196_),
    .B(_3197_));
 sg13g2_xnor2_1 _4089_ (.Y(_3200_),
    .A(net868),
    .B(\r2[3] ));
 sg13g2_a21oi_1 _4090_ (.A1(_3182_),
    .A2(_3184_),
    .Y(_3201_),
    .B1(_3200_));
 sg13g2_nand3_1 _4091_ (.B(_3184_),
    .C(_3200_),
    .A(_3182_),
    .Y(_3202_));
 sg13g2_nor2b_1 _4092_ (.A(_3201_),
    .B_N(_3202_),
    .Y(_3203_));
 sg13g2_a22oi_1 _4093_ (.Y(_3204_),
    .B1(_3203_),
    .B2(_3173_),
    .A2(_3190_),
    .A1(_3174_));
 sg13g2_o21ai_1 _4094_ (.B1(_3204_),
    .Y(_3205_),
    .A1(_3146_),
    .A2(_3199_));
 sg13g2_a22oi_1 _4095_ (.Y(_3206_),
    .B1(_3205_),
    .B2(net738),
    .A2(_3190_),
    .A1(net778));
 sg13g2_nor2_1 _4096_ (.A(net920),
    .B(_3206_),
    .Y(_0066_));
 sg13g2_nor2b_1 _4097_ (.A(net823),
    .B_N(net279),
    .Y(_3207_));
 sg13g2_o21ai_1 _4098_ (.B1(_3113_),
    .Y(_3208_),
    .A1(_3114_),
    .A2(_3191_));
 sg13g2_xnor2_1 _4099_ (.Y(_3209_),
    .A(_3111_),
    .B(_3208_));
 sg13g2_xnor2_1 _4100_ (.Y(_3210_),
    .A(\r2[4] ),
    .B(_3209_));
 sg13g2_nand3_1 _4101_ (.B(_3198_),
    .C(_3210_),
    .A(_3195_),
    .Y(_3211_));
 sg13g2_a21oi_1 _4102_ (.A1(_3195_),
    .A2(_3198_),
    .Y(_3212_),
    .B1(_3210_));
 sg13g2_nand3b_1 _4103_ (.B(net749),
    .C(_3211_),
    .Y(_3213_),
    .A_N(_3212_));
 sg13g2_xnor2_1 _4104_ (.Y(_3214_),
    .A(net862),
    .B(\r2[4] ));
 sg13g2_a21oi_1 _4105_ (.A1(net868),
    .A2(\r2[3] ),
    .Y(_3215_),
    .B1(_3201_));
 sg13g2_nor2_1 _4106_ (.A(_3214_),
    .B(_3215_),
    .Y(_3216_));
 sg13g2_and2_1 _4107_ (.A(_3214_),
    .B(_3215_),
    .X(_3217_));
 sg13g2_nor4_1 _4108_ (.A(net732),
    .B(_3137_),
    .C(_3216_),
    .D(_3217_),
    .Y(_3218_));
 sg13g2_a21oi_1 _4109_ (.A1(_3174_),
    .A2(_3207_),
    .Y(_3219_),
    .B1(_3218_));
 sg13g2_nand2_1 _4110_ (.Y(_3220_),
    .A(_3213_),
    .B(_3219_));
 sg13g2_a22oi_1 _4111_ (.Y(_3221_),
    .B1(_3220_),
    .B2(net738),
    .A2(_3207_),
    .A1(net779));
 sg13g2_nor2_1 _4112_ (.A(net921),
    .B(_3221_),
    .Y(_0067_));
 sg13g2_nor2b_1 _4113_ (.A(net823),
    .B_N(\r2[5] ),
    .Y(_3222_));
 sg13g2_a21o_1 _4114_ (.A2(_3209_),
    .A1(_2949_),
    .B1(_3212_),
    .X(_3223_));
 sg13g2_a21oi_1 _4115_ (.A1(_3115_),
    .A2(_3192_),
    .Y(_3224_),
    .B1(_3120_));
 sg13g2_inv_1 _4116_ (.Y(_3225_),
    .A(_3224_));
 sg13g2_xnor2_1 _4117_ (.Y(_3226_),
    .A(_3122_),
    .B(_3224_));
 sg13g2_nand2_1 _4118_ (.Y(_3227_),
    .A(\r2[5] ),
    .B(_3226_));
 sg13g2_xor2_1 _4119_ (.B(_3226_),
    .A(\r2[5] ),
    .X(_3228_));
 sg13g2_xnor2_1 _4120_ (.Y(_3229_),
    .A(_3223_),
    .B(_3228_));
 sg13g2_o21ai_1 _4121_ (.B1(net748),
    .Y(_3230_),
    .A1(_3136_),
    .A2(_3222_));
 sg13g2_o21ai_1 _4122_ (.B1(_3230_),
    .Y(_3231_),
    .A1(net748),
    .A2(_3229_));
 sg13g2_xnor2_1 _4123_ (.Y(_3232_),
    .A(net854),
    .B(\r2[5] ));
 sg13g2_a21oi_1 _4124_ (.A1(net862),
    .A2(\r2[4] ),
    .Y(_3233_),
    .B1(_3216_));
 sg13g2_nand2_1 _4125_ (.Y(_3234_),
    .A(_3232_),
    .B(_3233_));
 sg13g2_nor2_1 _4126_ (.A(_3232_),
    .B(_3233_),
    .Y(_3235_));
 sg13g2_nor2_1 _4127_ (.A(net732),
    .B(_3235_),
    .Y(_3236_));
 sg13g2_a22oi_1 _4128_ (.Y(_3237_),
    .B1(_3234_),
    .B2(_3236_),
    .A2(_3222_),
    .A1(net732));
 sg13g2_a21oi_1 _4129_ (.A1(_3136_),
    .A2(_3237_),
    .Y(_3238_),
    .B1(_3148_));
 sg13g2_a22oi_1 _4130_ (.Y(_3239_),
    .B1(_3231_),
    .B2(_3238_),
    .A2(_3222_),
    .A1(net778));
 sg13g2_nor2_1 _4131_ (.A(net921),
    .B(_3239_),
    .Y(_0068_));
 sg13g2_o21ai_1 _4132_ (.B1(_3223_),
    .Y(_3240_),
    .A1(\r2[5] ),
    .A2(_3226_));
 sg13g2_a21oi_1 _4133_ (.A1(_3122_),
    .A2(_3225_),
    .Y(_3241_),
    .B1(_3121_));
 sg13g2_nor2_1 _4134_ (.A(_3107_),
    .B(_3126_),
    .Y(_3242_));
 sg13g2_xnor2_1 _4135_ (.Y(_3243_),
    .A(_3241_),
    .B(_3242_));
 sg13g2_xnor2_1 _4136_ (.Y(_3244_),
    .A(\r2[6] ),
    .B(_3243_));
 sg13g2_nand3_1 _4137_ (.B(_3240_),
    .C(_3244_),
    .A(_3227_),
    .Y(_3245_));
 sg13g2_a21o_1 _4138_ (.A2(_3240_),
    .A1(_3227_),
    .B1(_3244_),
    .X(_3246_));
 sg13g2_nand2_1 _4139_ (.Y(_3247_),
    .A(_3066_),
    .B(_3144_));
 sg13g2_nand4_1 _4140_ (.B(_3144_),
    .C(_3245_),
    .A(_3066_),
    .Y(_3248_),
    .D(_3246_));
 sg13g2_nor2b_1 _4141_ (.A(net823),
    .B_N(\r2[6] ),
    .Y(_3249_));
 sg13g2_a21oi_1 _4142_ (.A1(_3247_),
    .A2(_3249_),
    .Y(_3250_),
    .B1(net799));
 sg13g2_a21oi_1 _4143_ (.A1(net854),
    .A2(\r2[5] ),
    .Y(_3251_),
    .B1(_3235_));
 sg13g2_nand2b_1 _4144_ (.Y(_3252_),
    .B(\r2[6] ),
    .A_N(_3251_));
 sg13g2_mux2_1 _4145_ (.A0(_3249_),
    .A1(_3252_),
    .S(_3131_),
    .X(_3253_));
 sg13g2_nand2b_1 _4146_ (.Y(_3254_),
    .B(_3251_),
    .A_N(net271));
 sg13g2_nand3_1 _4147_ (.B(_3253_),
    .C(_3254_),
    .A(net766),
    .Y(_3255_));
 sg13g2_nand2_1 _4148_ (.Y(_3256_),
    .A(net825),
    .B(net733));
 sg13g2_a221oi_1 _4149_ (.B2(net799),
    .C1(net920),
    .B1(_3255_),
    .A1(_3248_),
    .Y(_0069_),
    .A2(_3250_));
 sg13g2_nor2_1 _4150_ (.A(_2940_),
    .B(net822),
    .Y(_3257_));
 sg13g2_o21ai_1 _4151_ (.B1(_3127_),
    .Y(_3258_),
    .A1(_3107_),
    .A2(_3241_));
 sg13g2_nand2_1 _4152_ (.Y(_3259_),
    .A(net901),
    .B(_3258_));
 sg13g2_xnor2_1 _4153_ (.Y(_3260_),
    .A(_2611_),
    .B(_3258_));
 sg13g2_xnor2_1 _4154_ (.Y(_3261_),
    .A(\r2[7] ),
    .B(_3260_));
 sg13g2_nand2b_1 _4155_ (.Y(_3262_),
    .B(_3243_),
    .A_N(_0051_));
 sg13g2_a21oi_1 _4156_ (.A1(_3246_),
    .A2(_3262_),
    .Y(_3263_),
    .B1(_3261_));
 sg13g2_nand3_1 _4157_ (.B(_3261_),
    .C(_3262_),
    .A(_3246_),
    .Y(_3264_));
 sg13g2_nand2b_1 _4158_ (.Y(_3265_),
    .B(_3264_),
    .A_N(_3263_));
 sg13g2_o21ai_1 _4159_ (.B1(net737),
    .Y(_3266_),
    .A1(net736),
    .A2(_3257_));
 sg13g2_and2_1 _4160_ (.A(_2940_),
    .B(_3252_),
    .X(_3267_));
 sg13g2_nor2_1 _4161_ (.A(_2940_),
    .B(_3252_),
    .Y(_3268_));
 sg13g2_o21ai_1 _4162_ (.B1(net728),
    .Y(_3269_),
    .A1(_3267_),
    .A2(_3268_));
 sg13g2_a21oi_1 _4163_ (.A1(net732),
    .A2(_3257_),
    .Y(_3270_),
    .B1(_3137_));
 sg13g2_a221oi_1 _4164_ (.B2(_3270_),
    .C1(_3266_),
    .B1(_3269_),
    .A1(net749),
    .Y(_3271_),
    .A2(_3265_));
 sg13g2_a21oi_1 _4165_ (.A1(net778),
    .A2(_3257_),
    .Y(_3272_),
    .B1(_3271_));
 sg13g2_nor2_1 _4166_ (.A(net921),
    .B(_3272_),
    .Y(_0070_));
 sg13g2_nor2b_1 _4167_ (.A(net822),
    .B_N(net280),
    .Y(_3273_));
 sg13g2_a21oi_1 _4168_ (.A1(\r2[7] ),
    .A2(_3260_),
    .Y(_3274_),
    .B1(_3263_));
 sg13g2_nor2_1 _4169_ (.A(net897),
    .B(net815),
    .Y(_3275_));
 sg13g2_xor2_1 _4170_ (.B(_3259_),
    .A(net898),
    .X(_3276_));
 sg13g2_xnor2_1 _4171_ (.Y(_3277_),
    .A(\r2[8] ),
    .B(_3276_));
 sg13g2_nor2_1 _4172_ (.A(_3274_),
    .B(_3277_),
    .Y(_3278_));
 sg13g2_xnor2_1 _4173_ (.Y(_3279_),
    .A(_3274_),
    .B(_3277_));
 sg13g2_o21ai_1 _4174_ (.B1(net737),
    .Y(_3280_),
    .A1(net736),
    .A2(_3273_));
 sg13g2_o21ai_1 _4175_ (.B1(_3131_),
    .Y(_3281_),
    .A1(_0050_),
    .A2(_3267_));
 sg13g2_a21o_1 _4176_ (.A2(_3267_),
    .A1(_0050_),
    .B1(_3281_),
    .X(_3282_));
 sg13g2_a21oi_1 _4177_ (.A1(net732),
    .A2(_3273_),
    .Y(_3283_),
    .B1(_3137_));
 sg13g2_a221oi_1 _4178_ (.B2(_3283_),
    .C1(_3280_),
    .B1(_3282_),
    .A1(net750),
    .Y(_3284_),
    .A2(_3279_));
 sg13g2_a21oi_1 _4179_ (.A1(net777),
    .A2(_3273_),
    .Y(_3285_),
    .B1(_3284_));
 sg13g2_nor2_1 _4180_ (.A(net922),
    .B(net281),
    .Y(_0071_));
 sg13g2_nand2b_1 _4181_ (.Y(_3286_),
    .B(net917),
    .A_N(net822));
 sg13g2_a21oi_2 _4182_ (.B1(_3278_),
    .Y(_3287_),
    .A2(_3276_),
    .A1(_2930_));
 sg13g2_o21ai_1 _4183_ (.B1(_0022_),
    .Y(_3288_),
    .A1(net898),
    .A2(_3259_));
 sg13g2_nand2_1 _4184_ (.Y(_3289_),
    .A(net896),
    .B(_3288_));
 sg13g2_xnor2_1 _4185_ (.Y(_3290_),
    .A(_2633_),
    .B(_3288_));
 sg13g2_nand2_1 _4186_ (.Y(_3291_),
    .A(net917),
    .B(_3290_));
 sg13g2_nor2_1 _4187_ (.A(net917),
    .B(_3290_),
    .Y(_3292_));
 sg13g2_xor2_1 _4188_ (.B(_3290_),
    .A(net917),
    .X(_3293_));
 sg13g2_xnor2_1 _4189_ (.Y(_3294_),
    .A(_3287_),
    .B(_3293_));
 sg13g2_nand2_1 _4190_ (.Y(_3295_),
    .A(net917),
    .B(_3256_));
 sg13g2_mux2_1 _4191_ (.A0(net917),
    .A1(_3295_),
    .S(_3281_),
    .X(_3296_));
 sg13g2_a221oi_1 _4192_ (.B2(net798),
    .C1(_3148_),
    .B1(_3296_),
    .A1(_3151_),
    .Y(_3297_),
    .A2(_3286_));
 sg13g2_o21ai_1 _4193_ (.B1(_3297_),
    .Y(_3298_),
    .A1(net748),
    .A2(_3294_));
 sg13g2_o21ai_1 _4194_ (.B1(_3298_),
    .Y(_3299_),
    .A1(net775),
    .A2(_3286_));
 sg13g2_and2_1 _4195_ (.A(net925),
    .B(_3299_),
    .X(_0072_));
 sg13g2_nand2b_1 _4196_ (.Y(_3300_),
    .B(net284),
    .A_N(net821));
 sg13g2_a21oi_2 _4197_ (.B1(_3292_),
    .Y(_3301_),
    .A2(_3291_),
    .A1(_3287_));
 sg13g2_xnor2_1 _4198_ (.Y(_3302_),
    .A(_2622_),
    .B(_3289_));
 sg13g2_xor2_1 _4199_ (.B(_3302_),
    .A(\r2[10] ),
    .X(_3303_));
 sg13g2_xor2_1 _4200_ (.B(_3303_),
    .A(_3301_),
    .X(_3304_));
 sg13g2_nand2b_1 _4201_ (.Y(_3305_),
    .B(\r2[8] ),
    .A_N(net917));
 sg13g2_o21ai_1 _4202_ (.B1(_0025_),
    .Y(_3306_),
    .A1(_3267_),
    .A2(_3305_));
 sg13g2_nand2_1 _4203_ (.Y(_3307_),
    .A(net728),
    .B(_3306_));
 sg13g2_nand3_1 _4204_ (.B(_3256_),
    .C(_3307_),
    .A(\r2[10] ),
    .Y(_3308_));
 sg13g2_nor2_1 _4205_ (.A(\r2[10] ),
    .B(_3307_),
    .Y(_3309_));
 sg13g2_nor2_1 _4206_ (.A(net811),
    .B(_3309_),
    .Y(_3310_));
 sg13g2_a221oi_1 _4207_ (.B2(_3310_),
    .C1(_3148_),
    .B1(_3308_),
    .A1(_3151_),
    .Y(_3311_),
    .A2(_3300_));
 sg13g2_o21ai_1 _4208_ (.B1(_3311_),
    .Y(_3312_),
    .A1(net748),
    .A2(_3304_));
 sg13g2_o21ai_1 _4209_ (.B1(_3312_),
    .Y(_3313_),
    .A1(net774),
    .A2(_3300_));
 sg13g2_and2_1 _4210_ (.A(net928),
    .B(_3313_),
    .X(_0073_));
 sg13g2_nor2_1 _4211_ (.A(_2902_),
    .B(net820),
    .Y(_3314_));
 sg13g2_a22oi_1 _4212_ (.Y(_3315_),
    .B1(_3303_),
    .B2(_3301_),
    .A2(_3302_),
    .A1(_2921_));
 sg13g2_nor2_1 _4213_ (.A(\r2[11] ),
    .B(net718),
    .Y(_3316_));
 sg13g2_nand2_1 _4214_ (.Y(_3317_),
    .A(\r2[11] ),
    .B(net718));
 sg13g2_nand2b_1 _4215_ (.Y(_3318_),
    .B(_3317_),
    .A_N(_3316_));
 sg13g2_xnor2_1 _4216_ (.Y(_3319_),
    .A(_3315_),
    .B(_3318_));
 sg13g2_o21ai_1 _4217_ (.B1(net737),
    .Y(_3320_),
    .A1(net736),
    .A2(_3314_));
 sg13g2_and2_1 _4218_ (.A(\r2[10] ),
    .B(_3306_),
    .X(_3321_));
 sg13g2_a21oi_1 _4219_ (.A1(_0048_),
    .A2(_3321_),
    .Y(_3322_),
    .B1(net731));
 sg13g2_o21ai_1 _4220_ (.B1(_3322_),
    .Y(_3323_),
    .A1(net268),
    .A2(_3321_));
 sg13g2_o21ai_1 _4221_ (.B1(_3323_),
    .Y(_3324_),
    .A1(net728),
    .A2(_3314_));
 sg13g2_a221oi_1 _4222_ (.B2(net798),
    .C1(_3320_),
    .B1(_3324_),
    .A1(net749),
    .Y(_3325_),
    .A2(_3319_));
 sg13g2_a21oi_1 _4223_ (.A1(net777),
    .A2(_3314_),
    .Y(_3326_),
    .B1(_3325_));
 sg13g2_nor2_1 _4224_ (.A(net918),
    .B(net269),
    .Y(_0074_));
 sg13g2_or2_1 _4225_ (.X(_3327_),
    .B(_3316_),
    .A(_3315_));
 sg13g2_xnor2_1 _4226_ (.Y(_3328_),
    .A(\r2[12] ),
    .B(net717));
 sg13g2_nand3_1 _4227_ (.B(_3327_),
    .C(_3328_),
    .A(_3317_),
    .Y(_3329_));
 sg13g2_a21oi_1 _4228_ (.A1(_3317_),
    .A2(_3327_),
    .Y(_3330_),
    .B1(_3328_));
 sg13g2_nand3b_1 _4229_ (.B(net749),
    .C(_3329_),
    .Y(_3331_),
    .A_N(_3330_));
 sg13g2_nand2_1 _4230_ (.Y(_3332_),
    .A(\r2[11] ),
    .B(_3321_));
 sg13g2_xnor2_1 _4231_ (.Y(_3333_),
    .A(_2892_),
    .B(_3332_));
 sg13g2_nand2b_1 _4232_ (.Y(_3334_),
    .B(net226),
    .A_N(net820));
 sg13g2_a21oi_1 _4233_ (.A1(net730),
    .A2(_3334_),
    .Y(_3335_),
    .B1(net811));
 sg13g2_o21ai_1 _4234_ (.B1(_3335_),
    .Y(_3336_),
    .A1(net730),
    .A2(_3333_));
 sg13g2_o21ai_1 _4235_ (.B1(net737),
    .Y(_3337_),
    .A1(net736),
    .A2(_3334_));
 sg13g2_nor2b_1 _4236_ (.A(_3337_),
    .B_N(_3336_),
    .Y(_3338_));
 sg13g2_a221oi_1 _4237_ (.B2(_3331_),
    .C1(net918),
    .B1(_3338_),
    .A1(net777),
    .Y(_0075_),
    .A2(_3334_));
 sg13g2_nand2b_1 _4238_ (.Y(_3339_),
    .B(net249),
    .A_N(net820));
 sg13g2_or2_1 _4239_ (.X(_3340_),
    .B(_3339_),
    .A(net774));
 sg13g2_a21oi_2 _4240_ (.B1(_3330_),
    .Y(_3341_),
    .A2(net717),
    .A1(_2892_));
 sg13g2_nand2_1 _4241_ (.Y(_3342_),
    .A(\r2[13] ),
    .B(net717));
 sg13g2_nor2_1 _4242_ (.A(\r2[13] ),
    .B(net717),
    .Y(_3343_));
 sg13g2_xnor2_1 _4243_ (.Y(_3344_),
    .A(_2881_),
    .B(net717));
 sg13g2_a21oi_1 _4244_ (.A1(_3341_),
    .A2(_3344_),
    .Y(_3345_),
    .B1(net748));
 sg13g2_o21ai_1 _4245_ (.B1(_3345_),
    .Y(_3346_),
    .A1(_3341_),
    .A2(_3344_));
 sg13g2_nand3_1 _4246_ (.B(\r2[11] ),
    .C(_3321_),
    .A(\r2[12] ),
    .Y(_3347_));
 sg13g2_xnor2_1 _4247_ (.Y(_3348_),
    .A(_0046_),
    .B(_3347_));
 sg13g2_mux2_1 _4248_ (.A0(_3339_),
    .A1(_3348_),
    .S(net728),
    .X(_3349_));
 sg13g2_a221oi_1 _4249_ (.B2(net798),
    .C1(_3148_),
    .B1(_3349_),
    .A1(_3151_),
    .Y(_3350_),
    .A2(_3339_));
 sg13g2_nand2_1 _4250_ (.Y(_3351_),
    .A(_3346_),
    .B(_3350_));
 sg13g2_a21oi_1 _4251_ (.A1(_3340_),
    .A2(_3351_),
    .Y(_0076_),
    .B1(net918));
 sg13g2_nor2b_1 _4252_ (.A(net820),
    .B_N(net274),
    .Y(_3352_));
 sg13g2_o21ai_1 _4253_ (.B1(_3342_),
    .Y(_3353_),
    .A1(_3341_),
    .A2(_3343_));
 sg13g2_xor2_1 _4254_ (.B(net717),
    .A(\r2[14] ),
    .X(_3354_));
 sg13g2_xnor2_1 _4255_ (.Y(_3355_),
    .A(_3353_),
    .B(_3354_));
 sg13g2_a21oi_1 _4256_ (.A1(net730),
    .A2(_3352_),
    .Y(_3356_),
    .B1(_3137_));
 sg13g2_nor2_1 _4257_ (.A(_2881_),
    .B(_3347_),
    .Y(_3357_));
 sg13g2_xnor2_1 _4258_ (.Y(_3358_),
    .A(_0044_),
    .B(_3357_));
 sg13g2_nand2_1 _4259_ (.Y(_3359_),
    .A(net728),
    .B(_3358_));
 sg13g2_o21ai_1 _4260_ (.B1(net737),
    .Y(_3360_),
    .A1(net736),
    .A2(_3352_));
 sg13g2_a221oi_1 _4261_ (.B2(_3359_),
    .C1(_3360_),
    .B1(_3356_),
    .A1(net749),
    .Y(_3361_),
    .A2(_3355_));
 sg13g2_a21oi_1 _4262_ (.A1(net777),
    .A2(_3352_),
    .Y(_3362_),
    .B1(_3361_));
 sg13g2_nor2_1 _4263_ (.A(net918),
    .B(net275),
    .Y(_0077_));
 sg13g2_a22oi_1 _4264_ (.Y(_3363_),
    .B1(_3353_),
    .B2(_3354_),
    .A2(net717),
    .A1(_2861_));
 sg13g2_xor2_1 _4265_ (.B(net717),
    .A(\r2[15] ),
    .X(_3364_));
 sg13g2_nor2b_1 _4266_ (.A(_3363_),
    .B_N(_3364_),
    .Y(_3365_));
 sg13g2_nand2b_1 _4267_ (.Y(_3366_),
    .B(_3363_),
    .A_N(_3364_));
 sg13g2_nand3b_1 _4268_ (.B(_3366_),
    .C(net749),
    .Y(_3367_),
    .A_N(_3365_));
 sg13g2_nor4_1 _4269_ (.A(_0044_),
    .B(_2881_),
    .C(net731),
    .D(_3347_),
    .Y(_3368_));
 sg13g2_a21oi_1 _4270_ (.A1(net820),
    .A2(net730),
    .Y(_3369_),
    .B1(net811));
 sg13g2_xor2_1 _4271_ (.B(_3368_),
    .A(net238),
    .X(_3370_));
 sg13g2_nand2b_1 _4272_ (.Y(_3371_),
    .B(net238),
    .A_N(net820));
 sg13g2_o21ai_1 _4273_ (.B1(net737),
    .Y(_3372_),
    .A1(net736),
    .A2(_3371_));
 sg13g2_a21oi_1 _4274_ (.A1(_3369_),
    .A2(_3370_),
    .Y(_3373_),
    .B1(_3372_));
 sg13g2_a221oi_1 _4275_ (.B2(_3367_),
    .C1(net918),
    .B1(_3373_),
    .A1(net780),
    .Y(_0078_),
    .A2(_3371_));
 sg13g2_a21oi_1 _4276_ (.A1(_2851_),
    .A2(net718),
    .Y(_3374_),
    .B1(_3365_));
 sg13g2_xor2_1 _4277_ (.B(net718),
    .A(\r2[16] ),
    .X(_3375_));
 sg13g2_nand2b_2 _4278_ (.Y(_3376_),
    .B(_3375_),
    .A_N(_3374_));
 sg13g2_nand2b_1 _4279_ (.Y(_3377_),
    .B(_3374_),
    .A_N(_3375_));
 sg13g2_nand3_1 _4280_ (.B(_3376_),
    .C(_3377_),
    .A(net749),
    .Y(_3378_));
 sg13g2_and3_1 _4281_ (.X(_3379_),
    .A(\r2[15] ),
    .B(\r2[14] ),
    .C(_3357_));
 sg13g2_xnor2_1 _4282_ (.Y(_3380_),
    .A(_0026_),
    .B(_3379_));
 sg13g2_nand2b_1 _4283_ (.Y(_3381_),
    .B(net270),
    .A_N(net820));
 sg13g2_a21oi_1 _4284_ (.A1(net730),
    .A2(_3381_),
    .Y(_3382_),
    .B1(net811));
 sg13g2_o21ai_1 _4285_ (.B1(_3382_),
    .Y(_3383_),
    .A1(net730),
    .A2(_3380_));
 sg13g2_o21ai_1 _4286_ (.B1(_3383_),
    .Y(_3384_),
    .A1(net736),
    .A2(_3381_));
 sg13g2_nor2_1 _4287_ (.A(_3148_),
    .B(_3384_),
    .Y(_3385_));
 sg13g2_a221oi_1 _4288_ (.B2(_3378_),
    .C1(net918),
    .B1(_3385_),
    .A1(net780),
    .Y(_0079_),
    .A2(_3381_));
 sg13g2_nand2b_1 _4289_ (.Y(_3386_),
    .B(\r2[17] ),
    .A_N(net820));
 sg13g2_or2_1 _4290_ (.X(_3387_),
    .B(_3386_),
    .A(net774));
 sg13g2_nand2_1 _4291_ (.Y(_3388_),
    .A(_0026_),
    .B(net718));
 sg13g2_mux2_1 _4292_ (.A0(net718),
    .A1(_3388_),
    .S(_3376_),
    .X(_3389_));
 sg13g2_a21oi_1 _4293_ (.A1(\r2[17] ),
    .A2(_3389_),
    .Y(_3390_),
    .B1(net748));
 sg13g2_o21ai_1 _4294_ (.B1(_3390_),
    .Y(_3391_),
    .A1(\r2[17] ),
    .A2(_3389_));
 sg13g2_nand2_1 _4295_ (.Y(_3392_),
    .A(net730),
    .B(_3386_));
 sg13g2_nand2_1 _4296_ (.Y(_3393_),
    .A(\r2[16] ),
    .B(_3379_));
 sg13g2_xor2_1 _4297_ (.B(_3393_),
    .A(_0013_),
    .X(_3394_));
 sg13g2_o21ai_1 _4298_ (.B1(_3392_),
    .Y(_3395_),
    .A1(net730),
    .A2(_3394_));
 sg13g2_a22oi_1 _4299_ (.Y(_3396_),
    .B1(_3395_),
    .B2(net798),
    .A2(_3386_),
    .A1(_3151_));
 sg13g2_nand3_1 _4300_ (.B(_3391_),
    .C(_3396_),
    .A(net737),
    .Y(_3397_));
 sg13g2_a21oi_1 _4301_ (.A1(_3387_),
    .A2(_3397_),
    .Y(_0080_),
    .B1(net918));
 sg13g2_nor2b_1 _4302_ (.A(net819),
    .B_N(\r2[18] ),
    .Y(_3398_));
 sg13g2_o21ai_1 _4303_ (.B1(_0013_),
    .Y(_3399_),
    .A1(\r2[17] ),
    .A2(_0026_));
 sg13g2_mux2_1 _4304_ (.A0(_3376_),
    .A1(_3399_),
    .S(net718),
    .X(_3400_));
 sg13g2_nor2_1 _4305_ (.A(\r2[17] ),
    .B(_3376_),
    .Y(_3401_));
 sg13g2_nor2_1 _4306_ (.A(_3400_),
    .B(_3401_),
    .Y(_3402_));
 sg13g2_a21oi_1 _4307_ (.A1(net251),
    .A2(_3402_),
    .Y(_3403_),
    .B1(net748));
 sg13g2_o21ai_1 _4308_ (.B1(_3403_),
    .Y(_3404_),
    .A1(net251),
    .A2(_3402_));
 sg13g2_nand3_1 _4309_ (.B(\r2[17] ),
    .C(_3379_),
    .A(\r2[16] ),
    .Y(_3405_));
 sg13g2_xnor2_1 _4310_ (.Y(_3406_),
    .A(_0015_),
    .B(_3405_));
 sg13g2_nand2_1 _4311_ (.Y(_3407_),
    .A(net728),
    .B(_3406_));
 sg13g2_o21ai_1 _4312_ (.B1(_3407_),
    .Y(_3408_),
    .A1(net728),
    .A2(_3398_));
 sg13g2_o21ai_1 _4313_ (.B1(net737),
    .Y(_3409_),
    .A1(net736),
    .A2(_3398_));
 sg13g2_a21oi_1 _4314_ (.A1(net798),
    .A2(_3408_),
    .Y(_3410_),
    .B1(_3409_));
 sg13g2_a22oi_1 _4315_ (.Y(_3411_),
    .B1(_3404_),
    .B2(_3410_),
    .A2(_3398_),
    .A1(net777));
 sg13g2_nor2_1 _4316_ (.A(net918),
    .B(net252),
    .Y(_0081_));
 sg13g2_nand2_1 _4317_ (.Y(_0082_),
    .A(_3085_),
    .B(_3088_));
 sg13g2_xnor2_1 _4318_ (.Y(_3412_),
    .A(\title_r[12] ),
    .B(net899));
 sg13g2_xor2_1 _4319_ (.B(net899),
    .A(\title_r[9] ),
    .X(_3413_));
 sg13g2_nor2b_1 _4320_ (.A(net902),
    .B_N(\title_r[7] ),
    .Y(_3414_));
 sg13g2_xor2_1 _4321_ (.B(net902),
    .A(\title_r[7] ),
    .X(_3415_));
 sg13g2_nand2_1 _4322_ (.Y(_3416_),
    .A(\title_r[6] ),
    .B(net906));
 sg13g2_xnor2_1 _4323_ (.Y(_3417_),
    .A(\title_r[6] ),
    .B(net906));
 sg13g2_nand2_1 _4324_ (.Y(_3418_),
    .A(\title_r[5] ),
    .B(net909));
 sg13g2_xnor2_1 _4325_ (.Y(_3419_),
    .A(\title_r[5] ),
    .B(net909));
 sg13g2_nand2_1 _4326_ (.Y(_3420_),
    .A(\title_r[4] ),
    .B(net913));
 sg13g2_nand2_1 _4327_ (.Y(_3421_),
    .A(\title_r[3] ),
    .B(net914));
 sg13g2_xor2_1 _4328_ (.B(net914),
    .A(\title_r[3] ),
    .X(_3422_));
 sg13g2_and2_1 _4329_ (.A(\title_r[2] ),
    .B(\hvsync_gen.hpos[1] ),
    .X(_3423_));
 sg13g2_xnor2_1 _4330_ (.Y(_3424_),
    .A(\title_r[2] ),
    .B(net915));
 sg13g2_nor2_1 _4331_ (.A(\title_r[1] ),
    .B(\hvsync_gen.hpos[0] ),
    .Y(_3425_));
 sg13g2_a21oi_1 _4332_ (.A1(\title_r[1] ),
    .A2(\hvsync_gen.hpos[0] ),
    .Y(_3426_),
    .B1(\title_r[0] ));
 sg13g2_nor3_1 _4333_ (.A(_3424_),
    .B(_3425_),
    .C(_3426_),
    .Y(_3427_));
 sg13g2_o21ai_1 _4334_ (.B1(_3422_),
    .Y(_3428_),
    .A1(_3423_),
    .A2(_3427_));
 sg13g2_xnor2_1 _4335_ (.Y(_3429_),
    .A(\title_r[4] ),
    .B(net913));
 sg13g2_a21o_1 _4336_ (.A2(_3428_),
    .A1(_3421_),
    .B1(_3429_),
    .X(_3430_));
 sg13g2_a21o_1 _4337_ (.A2(_3430_),
    .A1(_3420_),
    .B1(_3419_),
    .X(_3431_));
 sg13g2_a21o_1 _4338_ (.A2(_3431_),
    .A1(_3418_),
    .B1(_3417_),
    .X(_3432_));
 sg13g2_a21oi_1 _4339_ (.A1(_3416_),
    .A2(_3432_),
    .Y(_3433_),
    .B1(_3415_));
 sg13g2_nand2_1 _4340_ (.Y(_3434_),
    .A(\title_r[8] ),
    .B(net815));
 sg13g2_xnor2_1 _4341_ (.Y(_3435_),
    .A(\title_r[8] ),
    .B(net902));
 sg13g2_o21ai_1 _4342_ (.B1(_3435_),
    .Y(_3436_),
    .A1(_3414_),
    .A2(_3433_));
 sg13g2_nor2_2 _4343_ (.A(_3413_),
    .B(_3436_),
    .Y(_3437_));
 sg13g2_xnor2_1 _4344_ (.Y(_3438_),
    .A(\title_r[10] ),
    .B(net899));
 sg13g2_xor2_1 _4345_ (.B(net899),
    .A(\title_r[11] ),
    .X(_3439_));
 sg13g2_inv_1 _4346_ (.Y(_3440_),
    .A(_3439_));
 sg13g2_nand3_1 _4347_ (.B(_3438_),
    .C(_3440_),
    .A(_3437_),
    .Y(_3441_));
 sg13g2_o21ai_1 _4348_ (.B1(_3434_),
    .Y(_3442_),
    .A1(_2367_),
    .A2(net899));
 sg13g2_o21ai_1 _4349_ (.B1(net815),
    .Y(_3443_),
    .A1(\title_r[11] ),
    .A2(\title_r[10] ));
 sg13g2_nand2_1 _4350_ (.Y(_3444_),
    .A(_3441_),
    .B(_3443_));
 sg13g2_nor2_1 _4351_ (.A(_3442_),
    .B(_3444_),
    .Y(_3445_));
 sg13g2_nor2b_1 _4352_ (.A(_3445_),
    .B_N(_3412_),
    .Y(_3446_));
 sg13g2_a21oi_1 _4353_ (.A1(\title_r[12] ),
    .A2(net815),
    .Y(_3447_),
    .B1(_3446_));
 sg13g2_xor2_1 _4354_ (.B(net899),
    .A(\title_r[13] ),
    .X(_3448_));
 sg13g2_o21ai_1 _4355_ (.B1(net764),
    .Y(_3449_),
    .A1(_3447_),
    .A2(_3448_));
 sg13g2_a21oi_1 _4356_ (.A1(_3447_),
    .A2(_3448_),
    .Y(_3450_),
    .B1(_3449_));
 sg13g2_nand2_1 _4357_ (.Y(_3451_),
    .A(\title_r[12] ),
    .B(net828));
 sg13g2_nor2b_1 _4358_ (.A(\title_r[11] ),
    .B_N(net828),
    .Y(_3452_));
 sg13g2_xnor2_1 _4359_ (.Y(_3453_),
    .A(\title_r[12] ),
    .B(net828));
 sg13g2_nor2_1 _4360_ (.A(_3452_),
    .B(_3453_),
    .Y(_3454_));
 sg13g2_a21oi_1 _4361_ (.A1(\title_r[12] ),
    .A2(_3452_),
    .Y(_3455_),
    .B1(_3454_));
 sg13g2_nand2_1 _4362_ (.Y(_3456_),
    .A(\title_r[6] ),
    .B(\hvsync_gen.vpos[5] ));
 sg13g2_nor2b_1 _4363_ (.A(\title_r[7] ),
    .B_N(net829),
    .Y(_3457_));
 sg13g2_xnor2_1 _4364_ (.Y(_3458_),
    .A(\title_r[7] ),
    .B(net828));
 sg13g2_nor2_1 _4365_ (.A(_3456_),
    .B(_3458_),
    .Y(_3459_));
 sg13g2_xor2_1 _4366_ (.B(\hvsync_gen.vpos[5] ),
    .A(\title_r[6] ),
    .X(_3460_));
 sg13g2_nand3_1 _4367_ (.B(net834),
    .C(_3460_),
    .A(\title_r[5] ),
    .Y(_3461_));
 sg13g2_xnor2_1 _4368_ (.Y(_3462_),
    .A(\title_r[5] ),
    .B(net834));
 sg13g2_nand2_1 _4369_ (.Y(_3463_),
    .A(\title_r[4] ),
    .B(net836));
 sg13g2_nor2_1 _4370_ (.A(_3462_),
    .B(_3463_),
    .Y(_3464_));
 sg13g2_xor2_1 _4371_ (.B(net836),
    .A(\title_r[4] ),
    .X(_3465_));
 sg13g2_nand3_1 _4372_ (.B(\hvsync_gen.vpos[2] ),
    .C(_3465_),
    .A(\title_r[3] ),
    .Y(_3466_));
 sg13g2_xnor2_1 _4373_ (.Y(_3467_),
    .A(\title_r[3] ),
    .B(\hvsync_gen.vpos[2] ));
 sg13g2_nand2_1 _4374_ (.Y(_3468_),
    .A(\title_r[2] ),
    .B(net839));
 sg13g2_nor2_1 _4375_ (.A(_3467_),
    .B(_3468_),
    .Y(_3469_));
 sg13g2_xnor2_1 _4376_ (.Y(_3470_),
    .A(\title_r[2] ),
    .B(net839));
 sg13g2_nor2_1 _4377_ (.A(\title_r[0] ),
    .B(net841),
    .Y(_3471_));
 sg13g2_a21oi_1 _4378_ (.A1(\title_r[0] ),
    .A2(net841),
    .Y(_3472_),
    .B1(\title_r[1] ));
 sg13g2_or3_1 _4379_ (.A(_3470_),
    .B(_3471_),
    .C(_3472_),
    .X(_3473_));
 sg13g2_xnor2_1 _4380_ (.Y(_3474_),
    .A(_3467_),
    .B(_3468_));
 sg13g2_nor2_1 _4381_ (.A(_3473_),
    .B(_3474_),
    .Y(_3475_));
 sg13g2_a21o_1 _4382_ (.A2(\hvsync_gen.vpos[2] ),
    .A1(\title_r[3] ),
    .B1(_3465_),
    .X(_3476_));
 sg13g2_and2_1 _4383_ (.A(_3466_),
    .B(_3476_),
    .X(_3477_));
 sg13g2_o21ai_1 _4384_ (.B1(_3477_),
    .Y(_3478_),
    .A1(_3469_),
    .A2(_3475_));
 sg13g2_xnor2_1 _4385_ (.Y(_3479_),
    .A(_3462_),
    .B(_3463_));
 sg13g2_a21oi_1 _4386_ (.A1(_3466_),
    .A2(_3478_),
    .Y(_3480_),
    .B1(_3479_));
 sg13g2_a21o_1 _4387_ (.A2(net834),
    .A1(\title_r[5] ),
    .B1(_3460_),
    .X(_3481_));
 sg13g2_and2_1 _4388_ (.A(_3461_),
    .B(_3481_),
    .X(_3482_));
 sg13g2_o21ai_1 _4389_ (.B1(_3482_),
    .Y(_3483_),
    .A1(_3464_),
    .A2(_3480_));
 sg13g2_xnor2_1 _4390_ (.Y(_3484_),
    .A(_3456_),
    .B(_3458_));
 sg13g2_a21oi_1 _4391_ (.A1(_3461_),
    .A2(_3483_),
    .Y(_3485_),
    .B1(_3484_));
 sg13g2_nor2_2 _4392_ (.A(_3459_),
    .B(_3485_),
    .Y(_3486_));
 sg13g2_nor2b_1 _4393_ (.A(\title_r[10] ),
    .B_N(net828),
    .Y(_3487_));
 sg13g2_xnor2_1 _4394_ (.Y(_3488_),
    .A(\title_r[11] ),
    .B(net828));
 sg13g2_nor2_1 _4395_ (.A(_3487_),
    .B(_3488_),
    .Y(_3489_));
 sg13g2_a21o_1 _4396_ (.A2(_3487_),
    .A1(\title_r[11] ),
    .B1(_3489_),
    .X(_3490_));
 sg13g2_nor2b_1 _4397_ (.A(\title_r[9] ),
    .B_N(net829),
    .Y(_3491_));
 sg13g2_xnor2_1 _4398_ (.Y(_3492_),
    .A(\title_r[10] ),
    .B(net829));
 sg13g2_nor2_1 _4399_ (.A(_3491_),
    .B(_3492_),
    .Y(_3493_));
 sg13g2_nor2b_1 _4400_ (.A(\title_r[8] ),
    .B_N(net829),
    .Y(_3494_));
 sg13g2_xnor2_1 _4401_ (.Y(_3495_),
    .A(\title_r[9] ),
    .B(net828));
 sg13g2_nor2_1 _4402_ (.A(_3494_),
    .B(_3495_),
    .Y(_3496_));
 sg13g2_a21oi_1 _4403_ (.A1(\title_r[9] ),
    .A2(_3494_),
    .Y(_3497_),
    .B1(_3496_));
 sg13g2_xnor2_1 _4404_ (.Y(_3498_),
    .A(\title_r[8] ),
    .B(net828));
 sg13g2_nor2_1 _4405_ (.A(_3457_),
    .B(_3498_),
    .Y(_3499_));
 sg13g2_nand2_1 _4406_ (.Y(_3500_),
    .A(_3497_),
    .B(_3499_));
 sg13g2_nand2b_1 _4407_ (.Y(_3501_),
    .B(_3500_),
    .A_N(_3496_));
 sg13g2_a21oi_1 _4408_ (.A1(\title_r[10] ),
    .A2(_3491_),
    .Y(_3502_),
    .B1(_3493_));
 sg13g2_a21oi_1 _4409_ (.A1(_3501_),
    .A2(_3502_),
    .Y(_3503_),
    .B1(_3493_));
 sg13g2_nor2_1 _4410_ (.A(_3490_),
    .B(_3503_),
    .Y(_3504_));
 sg13g2_nor2_1 _4411_ (.A(_3489_),
    .B(_3504_),
    .Y(_3505_));
 sg13g2_o21ai_1 _4412_ (.B1(_3505_),
    .Y(_3506_),
    .A1(\title_r[11] ),
    .A2(_3486_));
 sg13g2_a21oi_1 _4413_ (.A1(_3455_),
    .A2(_3506_),
    .Y(_3507_),
    .B1(_3454_));
 sg13g2_xnor2_1 _4414_ (.Y(_3508_),
    .A(_2550_),
    .B(_3451_));
 sg13g2_xnor2_1 _4415_ (.Y(_3509_),
    .A(_3507_),
    .B(_3508_));
 sg13g2_a21oi_1 _4416_ (.A1(net751),
    .A2(_3509_),
    .Y(_3510_),
    .B1(_3450_));
 sg13g2_nor3_1 _4417_ (.A(net832),
    .B(net833),
    .C(_3142_),
    .Y(_3511_));
 sg13g2_nand3_1 _4418_ (.B(_3064_),
    .C(_3511_),
    .A(net237),
    .Y(_3512_));
 sg13g2_mux2_1 _4419_ (.A0(_2550_),
    .A1(_3510_),
    .S(net793),
    .X(_3513_));
 sg13g2_a21oi_1 _4420_ (.A1(_3512_),
    .A2(_3513_),
    .Y(_0083_),
    .B1(net924));
 sg13g2_nand2_2 _4421_ (.Y(_3514_),
    .A(net930),
    .B(_3142_));
 sg13g2_nor2b_1 _4422_ (.A(\frame_counter[7] ),
    .B_N(net850),
    .Y(_3515_));
 sg13g2_nor2b_2 _4423_ (.A(net851),
    .B_N(_3515_),
    .Y(_3516_));
 sg13g2_nand2b_1 _4424_ (.Y(_3517_),
    .B(_3515_),
    .A_N(net851));
 sg13g2_nor2b_2 _4425_ (.A(\frame_counter[8] ),
    .B_N(net852),
    .Y(_3518_));
 sg13g2_nand2_2 _4426_ (.Y(_3519_),
    .A(_0034_),
    .B(_3518_));
 sg13g2_nand2b_1 _4427_ (.Y(_3520_),
    .B(net850),
    .A_N(net851));
 sg13g2_and2_1 _4428_ (.A(net851),
    .B(net852),
    .X(_3521_));
 sg13g2_and2_1 _4429_ (.A(net850),
    .B(_3521_),
    .X(_3522_));
 sg13g2_a21o_2 _4430_ (.A2(_0017_),
    .A1(net852),
    .B1(_3515_),
    .X(_3523_));
 sg13g2_nor2_2 _4431_ (.A(_2388_),
    .B(net852),
    .Y(_3524_));
 sg13g2_and2_2 _4432_ (.A(\frame_counter[8] ),
    .B(_3524_),
    .X(_3525_));
 sg13g2_nand2_2 _4433_ (.Y(_3526_),
    .A(net851),
    .B(_3524_));
 sg13g2_nand2_2 _4434_ (.Y(_3527_),
    .A(net873),
    .B(net817));
 sg13g2_nor2_2 _4435_ (.A(_3526_),
    .B(_3527_),
    .Y(_3528_));
 sg13g2_nand2_1 _4436_ (.Y(_3529_),
    .A(\envelopeA[0] ),
    .B(_3528_));
 sg13g2_nand2_1 _4437_ (.Y(_3530_),
    .A(net816),
    .B(net839));
 sg13g2_xnor2_1 _4438_ (.Y(_3531_),
    .A(net889),
    .B(net839));
 sg13g2_nand3_1 _4439_ (.B(_3528_),
    .C(_3531_),
    .A(net892),
    .Y(_3532_));
 sg13g2_a21o_1 _4440_ (.A2(_3528_),
    .A1(net892),
    .B1(_3531_),
    .X(_3533_));
 sg13g2_nand2_1 _4441_ (.Y(_3534_),
    .A(_3532_),
    .B(_3533_));
 sg13g2_a21oi_1 _4442_ (.A1(_0057_),
    .A2(_3529_),
    .Y(_3535_),
    .B1(_3534_));
 sg13g2_nor2_1 _4443_ (.A(_3519_),
    .B(_3527_),
    .Y(_3536_));
 sg13g2_nor3_1 _4444_ (.A(_2456_),
    .B(_3519_),
    .C(_3527_),
    .Y(_3537_));
 sg13g2_nand3_1 _4445_ (.B(_3529_),
    .C(_3534_),
    .A(_0057_),
    .Y(_3538_));
 sg13g2_nor2b_1 _4446_ (.A(_3535_),
    .B_N(_3538_),
    .Y(_3539_));
 sg13g2_a21oi_1 _4447_ (.A1(_3537_),
    .A2(_3538_),
    .Y(_3540_),
    .B1(_3535_));
 sg13g2_nand2_1 _4448_ (.Y(_3541_),
    .A(net889),
    .B(_3536_));
 sg13g2_and2_1 _4449_ (.A(_3530_),
    .B(_3532_),
    .X(_3542_));
 sg13g2_xnor2_1 _4450_ (.Y(_3543_),
    .A(net883),
    .B(net837));
 sg13g2_and3_1 _4451_ (.X(_3544_),
    .A(_0012_),
    .B(_3528_),
    .C(_3543_));
 sg13g2_a21oi_1 _4452_ (.A1(_0012_),
    .A2(_3528_),
    .Y(_3545_),
    .B1(_3543_));
 sg13g2_or2_1 _4453_ (.X(_3546_),
    .B(_3545_),
    .A(_3544_));
 sg13g2_or2_1 _4454_ (.X(_3547_),
    .B(_3546_),
    .A(_3542_));
 sg13g2_xor2_1 _4455_ (.B(_3546_),
    .A(_3542_),
    .X(_3548_));
 sg13g2_nand2b_1 _4456_ (.Y(_3549_),
    .B(_3548_),
    .A_N(_3541_));
 sg13g2_xor2_1 _4457_ (.B(_3548_),
    .A(_3541_),
    .X(_3550_));
 sg13g2_nor2_1 _4458_ (.A(_3540_),
    .B(_3550_),
    .Y(_3551_));
 sg13g2_xnor2_1 _4459_ (.Y(_3552_),
    .A(_3537_),
    .B(_3539_));
 sg13g2_xor2_1 _4460_ (.B(_3529_),
    .A(net840),
    .X(_3553_));
 sg13g2_and2_1 _4461_ (.A(frame_counter_frac),
    .B(_3536_),
    .X(_3554_));
 sg13g2_xnor2_1 _4462_ (.Y(_3555_),
    .A(net813),
    .B(_3553_));
 sg13g2_a22oi_1 _4463_ (.Y(_3556_),
    .B1(_3554_),
    .B2(_3555_),
    .A2(_3553_),
    .A1(_2456_));
 sg13g2_nor2_1 _4464_ (.A(_3552_),
    .B(_3556_),
    .Y(_3557_));
 sg13g2_xor2_1 _4465_ (.B(_3550_),
    .A(_3540_),
    .X(_3558_));
 sg13g2_a21oi_1 _4466_ (.A1(_3557_),
    .A2(_3558_),
    .Y(_3559_),
    .B1(_3551_));
 sg13g2_and2_1 _4467_ (.A(_0053_),
    .B(_3536_),
    .X(_3560_));
 sg13g2_a21oi_1 _4468_ (.A1(_2437_),
    .A2(net837),
    .Y(_3561_),
    .B1(_3544_));
 sg13g2_nand2_1 _4469_ (.Y(_3562_),
    .A(_0053_),
    .B(_3528_));
 sg13g2_xor2_1 _4470_ (.B(net836),
    .A(net875),
    .X(_3563_));
 sg13g2_xnor2_1 _4471_ (.Y(_3564_),
    .A(_3562_),
    .B(_3563_));
 sg13g2_nor2_1 _4472_ (.A(_3561_),
    .B(_3564_),
    .Y(_3565_));
 sg13g2_xnor2_1 _4473_ (.Y(_3566_),
    .A(_3561_),
    .B(_3564_));
 sg13g2_inv_1 _4474_ (.Y(_3567_),
    .A(_3566_));
 sg13g2_xor2_1 _4475_ (.B(_3566_),
    .A(net762),
    .X(_3568_));
 sg13g2_a21oi_1 _4476_ (.A1(_3547_),
    .A2(_3549_),
    .Y(_3569_),
    .B1(_3568_));
 sg13g2_nand3_1 _4477_ (.B(_3549_),
    .C(_3568_),
    .A(_3547_),
    .Y(_3570_));
 sg13g2_nor2b_1 _4478_ (.A(_3569_),
    .B_N(_3570_),
    .Y(_3571_));
 sg13g2_nand2b_1 _4479_ (.Y(_3572_),
    .B(_3571_),
    .A_N(_3559_));
 sg13g2_xnor2_1 _4480_ (.Y(_3573_),
    .A(_3559_),
    .B(_3571_));
 sg13g2_and2_1 _4481_ (.A(net791),
    .B(_3573_),
    .X(_3574_));
 sg13g2_a21oi_2 _4482_ (.B1(_3525_),
    .Y(_3575_),
    .A2(_3518_),
    .A1(\frame_counter[9] ));
 sg13g2_a21o_1 _4483_ (.A2(_3518_),
    .A1(\frame_counter[9] ),
    .B1(_3525_),
    .X(_3576_));
 sg13g2_nand2_1 _4484_ (.Y(_3577_),
    .A(net863),
    .B(net869));
 sg13g2_xnor2_1 _4485_ (.Y(_3578_),
    .A(net853),
    .B(_3577_));
 sg13g2_xnor2_1 _4486_ (.Y(_3579_),
    .A(_2695_),
    .B(_3577_));
 sg13g2_nor2_2 _4487_ (.A(net862),
    .B(net867),
    .Y(_3580_));
 sg13g2_xor2_1 _4488_ (.B(net869),
    .A(net863),
    .X(_3581_));
 sg13g2_xnor2_1 _4489_ (.Y(_3582_),
    .A(net863),
    .B(net869));
 sg13g2_nor3_1 _4490_ (.A(net854),
    .B(net862),
    .C(net867),
    .Y(_3583_));
 sg13g2_nand2_2 _4491_ (.Y(_3584_),
    .A(_2397_),
    .B(_3580_));
 sg13g2_nor2_1 _4492_ (.A(_0038_),
    .B(_3584_),
    .Y(_3585_));
 sg13g2_nand2_1 _4493_ (.Y(_3586_),
    .A(_2789_),
    .B(net805));
 sg13g2_xnor2_1 _4494_ (.Y(_3587_),
    .A(_2789_),
    .B(net805));
 sg13g2_nor2_1 _4495_ (.A(_0039_),
    .B(net805),
    .Y(_3588_));
 sg13g2_xnor2_1 _4496_ (.Y(_3589_),
    .A(_3580_),
    .B(net854));
 sg13g2_a21oi_2 _4497_ (.B1(_3588_),
    .Y(_3590_),
    .A2(_3589_),
    .A1(_2820_));
 sg13g2_xnor2_1 _4498_ (.Y(_3591_),
    .A(_3580_),
    .B(net853));
 sg13g2_xnor2_1 _4499_ (.Y(_3592_),
    .A(_0040_),
    .B(_3591_));
 sg13g2_inv_1 _4500_ (.Y(_3593_),
    .A(_3592_));
 sg13g2_xnor2_1 _4501_ (.Y(_3594_),
    .A(_0039_),
    .B(net805));
 sg13g2_or2_1 _4502_ (.X(_3595_),
    .B(_3594_),
    .A(_3592_));
 sg13g2_nand2b_1 _4503_ (.Y(_3596_),
    .B(net874),
    .A_N(net846));
 sg13g2_nand2b_1 _4504_ (.Y(_3597_),
    .B(net848),
    .A_N(net884));
 sg13g2_nor2b_1 _4505_ (.A(\r1[1] ),
    .B_N(net893),
    .Y(_3598_));
 sg13g2_nor2b_1 _4506_ (.A(net848),
    .B_N(net884),
    .Y(_3599_));
 sg13g2_xnor2_1 _4507_ (.Y(_3600_),
    .A(net884),
    .B(net848));
 sg13g2_o21ai_1 _4508_ (.B1(_3597_),
    .Y(_3601_),
    .A1(_3599_),
    .A2(_3598_));
 sg13g2_nor2b_1 _4509_ (.A(net878),
    .B_N(net847),
    .Y(_3602_));
 sg13g2_nand2b_1 _4510_ (.Y(_3603_),
    .B(net878),
    .A_N(net847));
 sg13g2_xor2_1 _4511_ (.B(net847),
    .A(net878),
    .X(_3604_));
 sg13g2_nor2b_1 _4512_ (.A(net874),
    .B_N(net846),
    .Y(_3605_));
 sg13g2_xor2_1 _4513_ (.B(net846),
    .A(net874),
    .X(_3606_));
 sg13g2_nor2_1 _4514_ (.A(_3604_),
    .B(_3606_),
    .Y(_3607_));
 sg13g2_a221oi_1 _4515_ (.B2(_3607_),
    .C1(_3605_),
    .B1(_3601_),
    .A1(_3596_),
    .Y(_3608_),
    .A2(_3602_));
 sg13g2_and2_1 _4516_ (.A(net867),
    .B(\r1[5] ),
    .X(_3609_));
 sg13g2_nand2_1 _4517_ (.Y(_3610_),
    .A(net867),
    .B(net845));
 sg13g2_xnor2_1 _4518_ (.Y(_3611_),
    .A(net867),
    .B(net845));
 sg13g2_xnor2_1 _4519_ (.Y(_3612_),
    .A(\r1[6] ),
    .B(net807));
 sg13g2_nand2b_1 _4520_ (.Y(_3613_),
    .B(_3612_),
    .A_N(_3611_));
 sg13g2_or2_1 _4521_ (.X(_3614_),
    .B(_3613_),
    .A(net152));
 sg13g2_a22oi_1 _4522_ (.Y(_3615_),
    .B1(_3609_),
    .B2(_3612_),
    .A2(net810),
    .A1(_2831_));
 sg13g2_and2_1 _4523_ (.A(_3590_),
    .B(_3615_),
    .X(_3616_));
 sg13g2_a22oi_1 _4524_ (.Y(_3617_),
    .B1(_3614_),
    .B2(_3616_),
    .A2(_3595_),
    .A1(_3590_));
 sg13g2_a221oi_1 _4525_ (.B2(_3616_),
    .C1(_3587_),
    .B1(_3614_),
    .A1(_3595_),
    .Y(_3618_),
    .A2(_3590_));
 sg13g2_xor2_1 _4526_ (.B(_3617_),
    .A(_3587_),
    .X(_0186_));
 sg13g2_nand2b_1 _4527_ (.Y(_0187_),
    .B(_0186_),
    .A_N(\r2[10] ));
 sg13g2_nand3b_1 _4528_ (.B(_0037_),
    .C(_3586_),
    .Y(_0188_),
    .A_N(_3618_));
 sg13g2_o21ai_1 _4529_ (.B1(_2799_),
    .Y(_0189_),
    .A1(_3585_),
    .A2(_3618_));
 sg13g2_nand3_1 _4530_ (.B(_0188_),
    .C(_0189_),
    .A(_2911_),
    .Y(_0190_));
 sg13g2_a21o_1 _4531_ (.A2(_0189_),
    .A1(_0188_),
    .B1(_2911_),
    .X(_0191_));
 sg13g2_a21oi_1 _4532_ (.A1(_0190_),
    .A2(_0191_),
    .Y(_0192_),
    .B1(_0187_));
 sg13g2_and3_1 _4533_ (.X(_0193_),
    .A(_0187_),
    .B(_0190_),
    .C(_0191_));
 sg13g2_nand3_1 _4534_ (.B(_0190_),
    .C(_0191_),
    .A(_0187_),
    .Y(_0194_));
 sg13g2_nor2_1 _4535_ (.A(_0192_),
    .B(_0193_),
    .Y(_0195_));
 sg13g2_inv_1 _4536_ (.Y(_0196_),
    .A(_0195_));
 sg13g2_o21ai_1 _4537_ (.B1(_3615_),
    .Y(_0197_),
    .A1(net153),
    .A2(_3613_));
 sg13g2_a22oi_1 _4538_ (.Y(_0198_),
    .B1(_3593_),
    .B2(_0197_),
    .A2(_3589_),
    .A1(_2820_));
 sg13g2_xnor2_1 _4539_ (.Y(_0199_),
    .A(_3594_),
    .B(_0198_));
 sg13g2_nand2b_1 _4540_ (.Y(_0200_),
    .B(\r2[9] ),
    .A_N(_0199_));
 sg13g2_xnor2_1 _4541_ (.Y(_0201_),
    .A(_2921_),
    .B(_0186_));
 sg13g2_nor2_1 _4542_ (.A(_0200_),
    .B(_0201_),
    .Y(_0202_));
 sg13g2_or2_1 _4543_ (.X(_0203_),
    .B(_0201_),
    .A(_0200_));
 sg13g2_xnor2_1 _4544_ (.Y(_0204_),
    .A(_0200_),
    .B(_0201_));
 sg13g2_xnor2_1 _4545_ (.Y(_0205_),
    .A(_3593_),
    .B(_0197_));
 sg13g2_nand2_2 _4546_ (.Y(_0206_),
    .A(_0050_),
    .B(_0205_));
 sg13g2_xnor2_1 _4547_ (.Y(_0207_),
    .A(net917),
    .B(_0199_));
 sg13g2_nor2_1 _4548_ (.A(_0206_),
    .B(_0207_),
    .Y(_0208_));
 sg13g2_o21ai_1 _4549_ (.B1(_3610_),
    .Y(_0209_),
    .A1(net152),
    .A2(_3611_));
 sg13g2_xor2_1 _4550_ (.B(_0209_),
    .A(_3612_),
    .X(_0210_));
 sg13g2_nand2_1 _4551_ (.Y(_0211_),
    .A(\r2[7] ),
    .B(_0210_));
 sg13g2_xor2_1 _4552_ (.B(_0205_),
    .A(\r2[8] ),
    .X(_0212_));
 sg13g2_nor2b_1 _4553_ (.A(_0211_),
    .B_N(_0212_),
    .Y(_0213_));
 sg13g2_nand2b_1 _4554_ (.Y(_0214_),
    .B(_0212_),
    .A_N(_0211_));
 sg13g2_a21oi_1 _4555_ (.A1(_0206_),
    .A2(_0207_),
    .Y(_0215_),
    .B1(_0213_));
 sg13g2_nor2_1 _4556_ (.A(_0208_),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_inv_1 _4557_ (.Y(_0217_),
    .A(_0216_));
 sg13g2_xor2_1 _4558_ (.B(_0207_),
    .A(_0206_),
    .X(_0218_));
 sg13g2_xnor2_1 _4559_ (.Y(_0219_),
    .A(_0206_),
    .B(_0207_));
 sg13g2_xnor2_1 _4560_ (.Y(_0220_),
    .A(_0211_),
    .B(_0212_));
 sg13g2_xnor2_1 _4561_ (.Y(_0221_),
    .A(net152),
    .B(_3611_));
 sg13g2_xnor2_1 _4562_ (.Y(_0222_),
    .A(\r2[6] ),
    .B(_0221_));
 sg13g2_nor2_1 _4563_ (.A(_0051_),
    .B(_0221_),
    .Y(_0223_));
 sg13g2_a21oi_1 _4564_ (.A1(net853),
    .A2(_0222_),
    .Y(_0224_),
    .B1(_0223_));
 sg13g2_xor2_1 _4565_ (.B(_0210_),
    .A(\r2[7] ),
    .X(_0225_));
 sg13g2_nor2b_1 _4566_ (.A(_0224_),
    .B_N(_0225_),
    .Y(_0226_));
 sg13g2_nand2b_2 _4567_ (.Y(_0227_),
    .B(_0224_),
    .A_N(_0225_));
 sg13g2_xnor2_1 _4568_ (.Y(_0228_),
    .A(_2695_),
    .B(_0222_));
 sg13g2_a21oi_1 _4569_ (.A1(_3601_),
    .A2(_3603_),
    .Y(_0229_),
    .B1(_3602_));
 sg13g2_xor2_1 _4570_ (.B(_0229_),
    .A(_3606_),
    .X(_0230_));
 sg13g2_and2_1 _4571_ (.A(\r2[5] ),
    .B(_0230_),
    .X(_0231_));
 sg13g2_xor2_1 _4572_ (.B(_0230_),
    .A(\r2[5] ),
    .X(_0232_));
 sg13g2_a21oi_1 _4573_ (.A1(net861),
    .A2(_0232_),
    .Y(_0233_),
    .B1(_0231_));
 sg13g2_nand2b_1 _4574_ (.Y(_0234_),
    .B(_0228_),
    .A_N(_0233_));
 sg13g2_xnor2_1 _4575_ (.Y(_0235_),
    .A(_0228_),
    .B(_0233_));
 sg13g2_inv_1 _4576_ (.Y(_0236_),
    .A(_0235_));
 sg13g2_xnor2_1 _4577_ (.Y(_0237_),
    .A(_3601_),
    .B(_3604_));
 sg13g2_xnor2_1 _4578_ (.Y(_0238_),
    .A(\r2[4] ),
    .B(_0237_));
 sg13g2_nor2_1 _4579_ (.A(_2767_),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_a21oi_2 _4580_ (.B1(_0239_),
    .Y(_0240_),
    .A2(_0237_),
    .A1(_2949_));
 sg13g2_xnor2_1 _4581_ (.Y(_0241_),
    .A(net861),
    .B(_0232_));
 sg13g2_nor2_1 _4582_ (.A(_0240_),
    .B(_0241_),
    .Y(_0242_));
 sg13g2_xnor2_1 _4583_ (.Y(_0243_),
    .A(_2767_),
    .B(_0238_));
 sg13g2_xnor2_1 _4584_ (.Y(_0244_),
    .A(_3598_),
    .B(_3600_));
 sg13g2_and2_1 _4585_ (.A(\r2[3] ),
    .B(_0244_),
    .X(_0245_));
 sg13g2_xor2_1 _4586_ (.B(_0244_),
    .A(\r2[3] ),
    .X(_0246_));
 sg13g2_a21oi_1 _4587_ (.A1(_0032_),
    .A2(_0246_),
    .Y(_0247_),
    .B1(_0245_));
 sg13g2_or2_1 _4588_ (.X(_0248_),
    .B(_0247_),
    .A(_0243_));
 sg13g2_xnor2_1 _4589_ (.Y(_0249_),
    .A(_0243_),
    .B(_0247_));
 sg13g2_xor2_1 _4590_ (.B(\r1[1] ),
    .A(net893),
    .X(_0250_));
 sg13g2_nand2_1 _4591_ (.Y(_0251_),
    .A(\r2[2] ),
    .B(_0250_));
 sg13g2_xnor2_1 _4592_ (.Y(_0252_),
    .A(_2959_),
    .B(_0250_));
 sg13g2_nand2b_1 _4593_ (.Y(_0253_),
    .B(_0053_),
    .A_N(_0252_));
 sg13g2_xnor2_1 _4594_ (.Y(_0254_),
    .A(_0032_),
    .B(_0246_));
 sg13g2_a21oi_1 _4595_ (.A1(_0251_),
    .A2(_0253_),
    .Y(_0255_),
    .B1(_0254_));
 sg13g2_nand3_1 _4596_ (.B(_0253_),
    .C(_0254_),
    .A(_0251_),
    .Y(_0256_));
 sg13g2_xnor2_1 _4597_ (.Y(_0257_),
    .A(_0053_),
    .B(_0252_));
 sg13g2_nor2_1 _4598_ (.A(\r2[1] ),
    .B(\r1[0] ),
    .Y(_0258_));
 sg13g2_xor2_1 _4599_ (.B(\r1[0] ),
    .A(\r2[1] ),
    .X(_0259_));
 sg13g2_a21oi_2 _4600_ (.B1(_0258_),
    .Y(_0260_),
    .A2(_0259_),
    .A1(net885));
 sg13g2_nor2_1 _4601_ (.A(_0257_),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_inv_1 _4602_ (.Y(_0262_),
    .A(_0261_));
 sg13g2_o21ai_1 _4603_ (.B1(_0256_),
    .Y(_0263_),
    .A1(_0255_),
    .A2(_0262_));
 sg13g2_o21ai_1 _4604_ (.B1(_0248_),
    .Y(_0264_),
    .A1(_0263_),
    .A2(_0249_));
 sg13g2_xor2_1 _4605_ (.B(_0241_),
    .A(_0240_),
    .X(_0265_));
 sg13g2_a21oi_2 _4606_ (.B1(_0242_),
    .Y(_0266_),
    .A2(_0265_),
    .A1(_0264_));
 sg13g2_o21ai_1 _4607_ (.B1(_0234_),
    .Y(_0267_),
    .A1(_0236_),
    .A2(_0266_));
 sg13g2_nor2b_1 _4608_ (.A(_0226_),
    .B_N(_0234_),
    .Y(_0268_));
 sg13g2_o21ai_1 _4609_ (.B1(_0268_),
    .Y(_0269_),
    .A1(_0266_),
    .A2(_0236_));
 sg13g2_and3_1 _4610_ (.X(_0270_),
    .A(_0220_),
    .B(_0269_),
    .C(_0227_));
 sg13g2_nand3_1 _4611_ (.B(_0227_),
    .C(_0269_),
    .A(_0220_),
    .Y(_0271_));
 sg13g2_nand4_1 _4612_ (.B(_0220_),
    .C(_0227_),
    .A(_0269_),
    .Y(_0272_),
    .D(_0218_));
 sg13g2_a21oi_1 _4613_ (.A1(_0217_),
    .A2(_0272_),
    .Y(_0273_),
    .B1(_0204_));
 sg13g2_nand3b_1 _4614_ (.B(_0195_),
    .C(_0203_),
    .Y(_0274_),
    .A_N(_0273_));
 sg13g2_o21ai_1 _4615_ (.B1(_0196_),
    .Y(_0275_),
    .A1(_0202_),
    .A2(_0273_));
 sg13g2_nand2_2 _4616_ (.Y(_0276_),
    .A(_0274_),
    .B(_0275_));
 sg13g2_nor2_1 _4617_ (.A(net885),
    .B(net893),
    .Y(_0277_));
 sg13g2_xor2_1 _4618_ (.B(net893),
    .A(net884),
    .X(_0278_));
 sg13g2_xnor2_1 _4619_ (.Y(_0279_),
    .A(net884),
    .B(net893));
 sg13g2_a21oi_2 _4620_ (.B1(net802),
    .Y(_0280_),
    .A2(_0275_),
    .A1(_0274_));
 sg13g2_and3_1 _4621_ (.X(_0281_),
    .A(_0204_),
    .B(_0217_),
    .C(_0272_));
 sg13g2_or2_2 _4622_ (.X(_0282_),
    .B(_0281_),
    .A(_0273_));
 sg13g2_nor2_1 _4623_ (.A(net891),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_a21oi_1 _4624_ (.A1(_0274_),
    .A2(_0275_),
    .Y(_0284_),
    .B1(net891));
 sg13g2_nor2_1 _4625_ (.A(net802),
    .B(_0282_),
    .Y(_0285_));
 sg13g2_nand2_1 _4626_ (.Y(_0286_),
    .A(_0280_),
    .B(_0283_));
 sg13g2_nor3_2 _4627_ (.A(_0213_),
    .B(_0218_),
    .C(_0270_),
    .Y(_0287_));
 sg13g2_a21oi_2 _4628_ (.B1(_0219_),
    .Y(_0288_),
    .A2(_0271_),
    .A1(_0214_));
 sg13g2_nor2_2 _4629_ (.A(_0287_),
    .B(_0288_),
    .Y(_0289_));
 sg13g2_nor3_2 _4630_ (.A(net878),
    .B(net885),
    .C(net894),
    .Y(_0290_));
 sg13g2_xnor2_1 _4631_ (.Y(_0291_),
    .A(net879),
    .B(_0277_));
 sg13g2_xnor2_1 _4632_ (.Y(_0292_),
    .A(_2437_),
    .B(_0277_));
 sg13g2_nand2_1 _4633_ (.Y(_0293_),
    .A(_0289_),
    .B(net787));
 sg13g2_xnor2_1 _4634_ (.Y(_0294_),
    .A(_0284_),
    .B(_0285_));
 sg13g2_o21ai_1 _4635_ (.B1(_0286_),
    .Y(_0295_),
    .A1(_0293_),
    .A2(_0294_));
 sg13g2_nor2_1 _4636_ (.A(_0282_),
    .B(_0292_),
    .Y(_0296_));
 sg13g2_nor3_2 _4637_ (.A(_0192_),
    .B(_0193_),
    .C(_0204_),
    .Y(_0297_));
 sg13g2_and2_1 _4638_ (.A(_0218_),
    .B(_0220_),
    .X(_0298_));
 sg13g2_nand4_1 _4639_ (.B(_0269_),
    .C(_0227_),
    .A(_0297_),
    .Y(_0299_),
    .D(_0298_));
 sg13g2_a21oi_1 _4640_ (.A1(_0194_),
    .A2(_0203_),
    .Y(_0300_),
    .B1(_0192_));
 sg13g2_a21oi_2 _4641_ (.B1(_0300_),
    .Y(_0301_),
    .A2(_0297_),
    .A1(_0216_));
 sg13g2_nand3_1 _4642_ (.B(_0188_),
    .C(_0189_),
    .A(_2902_),
    .Y(_0302_));
 sg13g2_nand2_1 _4643_ (.Y(_0303_),
    .A(_0037_),
    .B(_3586_));
 sg13g2_a21o_2 _4644_ (.A2(_3618_),
    .A1(_2778_),
    .B1(_0303_),
    .X(_0304_));
 sg13g2_nor2_1 _4645_ (.A(net843),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_xor2_1 _4646_ (.B(_0304_),
    .A(net844),
    .X(_0306_));
 sg13g2_xnor2_1 _4647_ (.Y(_0307_),
    .A(_0047_),
    .B(_0306_));
 sg13g2_nand2_1 _4648_ (.Y(_0308_),
    .A(_0302_),
    .B(_0307_));
 sg13g2_xnor2_1 _4649_ (.Y(_0309_),
    .A(_0302_),
    .B(_0307_));
 sg13g2_a21o_1 _4650_ (.A2(_0301_),
    .A1(_0299_),
    .B1(_0309_),
    .X(_0310_));
 sg13g2_nand3_1 _4651_ (.B(_0301_),
    .C(_0309_),
    .A(_0299_),
    .Y(_0311_));
 sg13g2_and2_1 _4652_ (.A(_0310_),
    .B(_0311_),
    .X(_0312_));
 sg13g2_nand2_1 _4653_ (.Y(_0313_),
    .A(net804),
    .B(net719));
 sg13g2_and2_1 _4654_ (.A(net814),
    .B(net719),
    .X(_0314_));
 sg13g2_and2_1 _4655_ (.A(_0280_),
    .B(_0314_),
    .X(_0315_));
 sg13g2_xor2_1 _4656_ (.B(_0314_),
    .A(_0280_),
    .X(_0316_));
 sg13g2_xnor2_1 _4657_ (.Y(_0317_),
    .A(_0296_),
    .B(_0316_));
 sg13g2_nor2b_1 _4658_ (.A(_0317_),
    .B_N(_0295_),
    .Y(_0318_));
 sg13g2_nand2b_1 _4659_ (.Y(_0319_),
    .B(_0317_),
    .A_N(_0295_));
 sg13g2_xor2_1 _4660_ (.B(_0317_),
    .A(_0295_),
    .X(_0320_));
 sg13g2_and2_1 _4661_ (.A(_2427_),
    .B(_0290_),
    .X(_0321_));
 sg13g2_nand2_2 _4662_ (.Y(_0322_),
    .A(_2416_),
    .B(_0321_));
 sg13g2_nor2_2 _4663_ (.A(net863),
    .B(_0322_),
    .Y(_0323_));
 sg13g2_xnor2_1 _4664_ (.Y(_0324_),
    .A(_2407_),
    .B(_0322_));
 sg13g2_xnor2_1 _4665_ (.Y(_0325_),
    .A(net863),
    .B(_0322_));
 sg13g2_nand2b_1 _4666_ (.Y(_0326_),
    .B(_0227_),
    .A_N(_0226_));
 sg13g2_xnor2_1 _4667_ (.Y(_0327_),
    .A(_0267_),
    .B(_0326_));
 sg13g2_nand2_1 _4668_ (.Y(_0328_),
    .A(net757),
    .B(net726));
 sg13g2_inv_1 _4669_ (.Y(_0329_),
    .A(_0328_));
 sg13g2_xnor2_1 _4670_ (.Y(_0330_),
    .A(net869),
    .B(_0321_));
 sg13g2_xnor2_1 _4671_ (.Y(_0331_),
    .A(_2416_),
    .B(_0321_));
 sg13g2_nand2_1 _4672_ (.Y(_0332_),
    .A(_0289_),
    .B(net772));
 sg13g2_xnor2_1 _4673_ (.Y(_0333_),
    .A(net875),
    .B(_0290_));
 sg13g2_xnor2_1 _4674_ (.Y(_0334_),
    .A(_2427_),
    .B(_0290_));
 sg13g2_a21oi_2 _4675_ (.B1(_0220_),
    .Y(_0335_),
    .A2(_0269_),
    .A1(_0227_));
 sg13g2_or2_1 _4676_ (.X(_0336_),
    .B(_0335_),
    .A(_0270_));
 sg13g2_nand2_1 _4677_ (.Y(_0337_),
    .A(_0289_),
    .B(net785));
 sg13g2_or2_1 _4678_ (.X(_0338_),
    .B(net725),
    .A(_0331_));
 sg13g2_nor2_1 _4679_ (.A(_0337_),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_xor2_1 _4680_ (.B(_0338_),
    .A(_0337_),
    .X(_0340_));
 sg13g2_xnor2_1 _4681_ (.Y(_0341_),
    .A(_0328_),
    .B(_0340_));
 sg13g2_a21oi_1 _4682_ (.A1(_0319_),
    .A2(_0341_),
    .Y(_0342_),
    .B1(_0318_));
 sg13g2_or2_1 _4683_ (.X(_0343_),
    .B(_0336_),
    .A(_0325_));
 sg13g2_nor2_1 _4684_ (.A(_0282_),
    .B(_0331_),
    .Y(_0344_));
 sg13g2_nand2b_1 _4685_ (.Y(_0345_),
    .B(_0344_),
    .A_N(_0337_));
 sg13g2_o21ai_1 _4686_ (.B1(_0332_),
    .Y(_0346_),
    .A1(_0282_),
    .A2(net784));
 sg13g2_nand2_1 _4687_ (.Y(_0347_),
    .A(_0345_),
    .B(_0346_));
 sg13g2_xor2_1 _4688_ (.B(_0347_),
    .A(_0343_),
    .X(_0348_));
 sg13g2_a21oi_1 _4689_ (.A1(_0296_),
    .A2(_0316_),
    .Y(_0349_),
    .B1(_0315_));
 sg13g2_nand2_1 _4690_ (.Y(_0350_),
    .A(net716),
    .B(net788));
 sg13g2_nor2b_1 _4691_ (.A(\r2[12] ),
    .B_N(_0306_),
    .Y(_0351_));
 sg13g2_or3_1 _4692_ (.A(net844),
    .B(_2871_),
    .C(_0304_),
    .X(_0352_));
 sg13g2_o21ai_1 _4693_ (.B1(_2871_),
    .Y(_0353_),
    .A1(net844),
    .A2(_0304_));
 sg13g2_nand3_1 _4694_ (.B(_0352_),
    .C(_0353_),
    .A(_0046_),
    .Y(_0354_));
 sg13g2_a21o_1 _4695_ (.A2(_0353_),
    .A1(_0352_),
    .B1(_0046_),
    .X(_0355_));
 sg13g2_nand3_1 _4696_ (.B(_0354_),
    .C(_0355_),
    .A(_0351_),
    .Y(_0356_));
 sg13g2_a21o_1 _4697_ (.A2(_0355_),
    .A1(_0354_),
    .B1(_0351_),
    .X(_0357_));
 sg13g2_and2_1 _4698_ (.A(_0356_),
    .B(_0357_),
    .X(_0358_));
 sg13g2_inv_1 _4699_ (.Y(_0359_),
    .A(_0358_));
 sg13g2_a21oi_2 _4700_ (.B1(_0359_),
    .Y(_0360_),
    .A2(_0310_),
    .A1(_0308_));
 sg13g2_and3_2 _4701_ (.X(_0361_),
    .A(_0308_),
    .B(_0310_),
    .C(_0359_));
 sg13g2_nor2_2 _4702_ (.A(_0360_),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_nor3_2 _4703_ (.A(net802),
    .B(_0360_),
    .C(_0361_),
    .Y(_0363_));
 sg13g2_nor3_1 _4704_ (.A(net890),
    .B(_0360_),
    .C(_0361_),
    .Y(_0364_));
 sg13g2_nand2_1 _4705_ (.Y(_0365_),
    .A(_0314_),
    .B(_0363_));
 sg13g2_xor2_1 _4706_ (.B(_0364_),
    .A(_0313_),
    .X(_0366_));
 sg13g2_xnor2_1 _4707_ (.Y(_0367_),
    .A(_0350_),
    .B(_0366_));
 sg13g2_nor2_1 _4708_ (.A(_0349_),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_xor2_1 _4709_ (.B(_0367_),
    .A(_0349_),
    .X(_0369_));
 sg13g2_xnor2_1 _4710_ (.Y(_0370_),
    .A(_0348_),
    .B(_0369_));
 sg13g2_nor2_1 _4711_ (.A(_0342_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_xor2_1 _4712_ (.B(_0370_),
    .A(_0342_),
    .X(_0372_));
 sg13g2_xnor2_1 _4713_ (.Y(_0373_),
    .A(_0235_),
    .B(_0266_));
 sg13g2_nor3_2 _4714_ (.A(net863),
    .B(_2695_),
    .C(_0322_),
    .Y(_0374_));
 sg13g2_nand2_2 _4715_ (.Y(_0375_),
    .A(net853),
    .B(_0323_));
 sg13g2_nand2_1 _4716_ (.Y(_0376_),
    .A(net727),
    .B(net755));
 sg13g2_xor2_1 _4717_ (.B(net862),
    .A(net854),
    .X(_0377_));
 sg13g2_xnor2_1 _4718_ (.Y(_0378_),
    .A(net858),
    .B(net866));
 sg13g2_xnor2_1 _4719_ (.Y(_0379_),
    .A(\center_x[5] ),
    .B(_0323_));
 sg13g2_xnor2_1 _4720_ (.Y(_0380_),
    .A(_2397_),
    .B(_0323_));
 sg13g2_xnor2_1 _4721_ (.Y(_0381_),
    .A(net157),
    .B(_0265_));
 sg13g2_nor2_1 _4722_ (.A(_0380_),
    .B(_0381_),
    .Y(_0382_));
 sg13g2_nand2_1 _4723_ (.Y(_0383_),
    .A(net727),
    .B(net747));
 sg13g2_nor2_2 _4724_ (.A(_0375_),
    .B(_0381_),
    .Y(_0384_));
 sg13g2_nand3_1 _4725_ (.B(net747),
    .C(_0384_),
    .A(net727),
    .Y(_0385_));
 sg13g2_inv_1 _4726_ (.Y(_0386_),
    .A(_0385_));
 sg13g2_a21oi_1 _4727_ (.A1(_0329_),
    .A2(_0340_),
    .Y(_0387_),
    .B1(_0339_));
 sg13g2_nand2_1 _4728_ (.Y(_0388_),
    .A(net726),
    .B(net755));
 sg13g2_nand2_1 _4729_ (.Y(_0389_),
    .A(net726),
    .B(net747));
 sg13g2_or2_1 _4730_ (.X(_0390_),
    .B(_0389_),
    .A(_0376_));
 sg13g2_xor2_1 _4731_ (.B(_0389_),
    .A(_0376_),
    .X(_0391_));
 sg13g2_nor2b_1 _4732_ (.A(_0387_),
    .B_N(_0391_),
    .Y(_0392_));
 sg13g2_xnor2_1 _4733_ (.Y(_0393_),
    .A(_0387_),
    .B(_0391_));
 sg13g2_xnor2_1 _4734_ (.Y(_0394_),
    .A(_0385_),
    .B(_0393_));
 sg13g2_a21oi_1 _4735_ (.A1(_0372_),
    .A2(_0394_),
    .Y(_0395_),
    .B1(_0371_));
 sg13g2_o21ai_1 _4736_ (.B1(_0345_),
    .Y(_0396_),
    .A1(_0343_),
    .A2(_0347_));
 sg13g2_o21ai_1 _4737_ (.B1(_0388_),
    .Y(_0397_),
    .A1(_0336_),
    .A2(_0380_));
 sg13g2_nor2_1 _4738_ (.A(net725),
    .B(_0375_),
    .Y(_0398_));
 sg13g2_or3_1 _4739_ (.A(net725),
    .B(_0380_),
    .C(_0388_),
    .X(_0399_));
 sg13g2_nand2_1 _4740_ (.Y(_0400_),
    .A(_0397_),
    .B(_0399_));
 sg13g2_nand2b_1 _4741_ (.Y(_0401_),
    .B(_0396_),
    .A_N(_0400_));
 sg13g2_xor2_1 _4742_ (.B(_0400_),
    .A(_0396_),
    .X(_0402_));
 sg13g2_xnor2_1 _4743_ (.Y(_0403_),
    .A(_0390_),
    .B(_0402_));
 sg13g2_inv_1 _4744_ (.Y(_0404_),
    .A(_0403_));
 sg13g2_a21oi_1 _4745_ (.A1(_0348_),
    .A2(_0369_),
    .Y(_0405_),
    .B1(_0368_));
 sg13g2_o21ai_1 _4746_ (.B1(_0365_),
    .Y(_0406_),
    .A1(_0350_),
    .A2(_0366_));
 sg13g2_and2_1 _4747_ (.A(net788),
    .B(net719),
    .X(_0407_));
 sg13g2_and3_1 _4748_ (.X(_0408_),
    .A(_2881_),
    .B(_0352_),
    .C(_0353_));
 sg13g2_or2_1 _4749_ (.X(_0409_),
    .B(\r1[12] ),
    .A(\r1[13] ));
 sg13g2_nand2_1 _4750_ (.Y(_0410_),
    .A(net842),
    .B(\r1[12] ));
 sg13g2_nand2_1 _4751_ (.Y(_0411_),
    .A(_0409_),
    .B(_0410_));
 sg13g2_mux2_1 _4752_ (.A0(net842),
    .A1(_0411_),
    .S(_0305_),
    .X(_0412_));
 sg13g2_xnor2_1 _4753_ (.Y(_0413_),
    .A(_2861_),
    .B(_0412_));
 sg13g2_nor2b_1 _4754_ (.A(_0408_),
    .B_N(_0413_),
    .Y(_0414_));
 sg13g2_inv_1 _4755_ (.Y(_0415_),
    .A(_0414_));
 sg13g2_xnor2_1 _4756_ (.Y(_0416_),
    .A(_0408_),
    .B(_0413_));
 sg13g2_xor2_1 _4757_ (.B(_0413_),
    .A(_0408_),
    .X(_0417_));
 sg13g2_nand3b_1 _4758_ (.B(_0356_),
    .C(_0357_),
    .Y(_0418_),
    .A_N(_0309_));
 sg13g2_a21oi_2 _4759_ (.B1(_0418_),
    .Y(_0419_),
    .A2(_0301_),
    .A1(_0299_));
 sg13g2_a21o_1 _4760_ (.A2(_0301_),
    .A1(_0299_),
    .B1(_0418_),
    .X(_0420_));
 sg13g2_nand2_1 _4761_ (.Y(_0421_),
    .A(_0308_),
    .B(_0357_));
 sg13g2_and2_1 _4762_ (.A(_0356_),
    .B(_0421_),
    .X(_0422_));
 sg13g2_nand2_1 _4763_ (.Y(_0423_),
    .A(_0356_),
    .B(_0421_));
 sg13g2_a21oi_2 _4764_ (.B1(_0417_),
    .Y(_0424_),
    .A2(_0423_),
    .A1(_0420_));
 sg13g2_o21ai_1 _4765_ (.B1(_0416_),
    .Y(_0425_),
    .A1(_0419_),
    .A2(_0422_));
 sg13g2_nor3_2 _4766_ (.A(_0416_),
    .B(_0419_),
    .C(_0422_),
    .Y(_0426_));
 sg13g2_nor2_2 _4767_ (.A(_0424_),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_nand2_1 _4768_ (.Y(_0428_),
    .A(_0278_),
    .B(net714));
 sg13g2_nor3_2 _4769_ (.A(net890),
    .B(_0424_),
    .C(_0426_),
    .Y(_0429_));
 sg13g2_and2_1 _4770_ (.A(_0363_),
    .B(_0429_),
    .X(_0430_));
 sg13g2_xor2_1 _4771_ (.B(_0429_),
    .A(_0363_),
    .X(_0431_));
 sg13g2_xor2_1 _4772_ (.B(_0431_),
    .A(_0407_),
    .X(_0432_));
 sg13g2_xnor2_1 _4773_ (.Y(_0433_),
    .A(_0406_),
    .B(_0432_));
 sg13g2_nand2_1 _4774_ (.Y(_0434_),
    .A(_0289_),
    .B(net757));
 sg13g2_a21oi_2 _4775_ (.B1(net784),
    .Y(_0435_),
    .A2(_0275_),
    .A1(_0274_));
 sg13g2_nand2_1 _4776_ (.Y(_0436_),
    .A(_0344_),
    .B(_0435_));
 sg13g2_xnor2_1 _4777_ (.Y(_0437_),
    .A(_0344_),
    .B(_0435_));
 sg13g2_xor2_1 _4778_ (.B(_0437_),
    .A(_0434_),
    .X(_0438_));
 sg13g2_nor2b_1 _4779_ (.A(_0433_),
    .B_N(_0438_),
    .Y(_0439_));
 sg13g2_xor2_1 _4780_ (.B(_0438_),
    .A(_0433_),
    .X(_0440_));
 sg13g2_nor2_1 _4781_ (.A(_0405_),
    .B(_0440_),
    .Y(_0441_));
 sg13g2_xor2_1 _4782_ (.B(_0440_),
    .A(_0405_),
    .X(_0442_));
 sg13g2_xnor2_1 _4783_ (.Y(_0443_),
    .A(_0403_),
    .B(_0442_));
 sg13g2_nor2b_1 _4784_ (.A(_0395_),
    .B_N(_0443_),
    .Y(_0444_));
 sg13g2_a21oi_1 _4785_ (.A1(_0386_),
    .A2(_0393_),
    .Y(_0445_),
    .B1(_0392_));
 sg13g2_xnor2_1 _4786_ (.Y(_0446_),
    .A(_0395_),
    .B(_0443_));
 sg13g2_nor2b_1 _4787_ (.A(_0445_),
    .B_N(_0446_),
    .Y(_0447_));
 sg13g2_nor2_1 _4788_ (.A(_0444_),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_or2_1 _4789_ (.X(_0449_),
    .B(_0447_),
    .A(_0444_));
 sg13g2_o21ai_1 _4790_ (.B1(_0401_),
    .Y(_0450_),
    .A1(_0390_),
    .A2(_0402_));
 sg13g2_a21oi_1 _4791_ (.A1(_0404_),
    .A2(_0442_),
    .Y(_0451_),
    .B1(_0441_));
 sg13g2_o21ai_1 _4792_ (.B1(_0436_),
    .Y(_0452_),
    .A1(_0434_),
    .A2(_0437_));
 sg13g2_nand2_1 _4793_ (.Y(_0453_),
    .A(_0289_),
    .B(net747));
 sg13g2_nand2_1 _4794_ (.Y(_0454_),
    .A(_0289_),
    .B(net755));
 sg13g2_nor3_1 _4795_ (.A(net725),
    .B(_0375_),
    .C(_0453_),
    .Y(_0455_));
 sg13g2_xnor2_1 _4796_ (.Y(_0456_),
    .A(_0398_),
    .B(_0453_));
 sg13g2_xnor2_1 _4797_ (.Y(_0457_),
    .A(_0452_),
    .B(_0456_));
 sg13g2_xnor2_1 _4798_ (.Y(_0458_),
    .A(_0399_),
    .B(_0457_));
 sg13g2_a21oi_2 _4799_ (.B1(_0439_),
    .Y(_0459_),
    .A2(_0432_),
    .A1(_0406_));
 sg13g2_nor2_1 _4800_ (.A(_0282_),
    .B(_0325_),
    .Y(_0460_));
 sg13g2_and2_1 _4801_ (.A(net719),
    .B(_0330_),
    .X(_0461_));
 sg13g2_a22oi_1 _4802_ (.Y(_0462_),
    .B1(net786),
    .B2(net719),
    .A2(net772),
    .A1(net716));
 sg13g2_a21oi_1 _4803_ (.A1(_0435_),
    .A2(_0461_),
    .Y(_0463_),
    .B1(_0462_));
 sg13g2_xor2_1 _4804_ (.B(_0463_),
    .A(_0460_),
    .X(_0464_));
 sg13g2_a21oi_1 _4805_ (.A1(_0407_),
    .A2(_0431_),
    .Y(_0465_),
    .B1(_0430_));
 sg13g2_nand2_1 _4806_ (.Y(_0466_),
    .A(net788),
    .B(net715));
 sg13g2_inv_1 _4807_ (.Y(_0467_),
    .A(_0466_));
 sg13g2_nor2_1 _4808_ (.A(\r2[14] ),
    .B(_0412_),
    .Y(_0468_));
 sg13g2_nor3_1 _4809_ (.A(net843),
    .B(_0304_),
    .C(_0409_),
    .Y(_0469_));
 sg13g2_xnor2_1 _4810_ (.Y(_0470_),
    .A(_0042_),
    .B(_0469_));
 sg13g2_xnor2_1 _4811_ (.Y(_0471_),
    .A(_0043_),
    .B(_0470_));
 sg13g2_nor2_1 _4812_ (.A(_0468_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_xnor2_1 _4813_ (.Y(_0473_),
    .A(_0468_),
    .B(_0471_));
 sg13g2_inv_1 _4814_ (.Y(_0474_),
    .A(_0473_));
 sg13g2_nor3_2 _4815_ (.A(_0414_),
    .B(_0424_),
    .C(_0473_),
    .Y(_0475_));
 sg13g2_a21oi_2 _4816_ (.B1(_0474_),
    .Y(_0476_),
    .A2(_0425_),
    .A1(_0415_));
 sg13g2_or2_2 _4817_ (.X(_0477_),
    .B(_0476_),
    .A(_0475_));
 sg13g2_o21ai_1 _4818_ (.B1(net893),
    .Y(_0478_),
    .A1(_0475_),
    .A2(_0476_));
 sg13g2_nor2_1 _4819_ (.A(_0428_),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_xor2_1 _4820_ (.B(_0478_),
    .A(_0428_),
    .X(_0480_));
 sg13g2_xnor2_1 _4821_ (.Y(_0481_),
    .A(_0467_),
    .B(_0480_));
 sg13g2_nor2_1 _4822_ (.A(_0465_),
    .B(_0481_),
    .Y(_0482_));
 sg13g2_xor2_1 _4823_ (.B(_0481_),
    .A(_0465_),
    .X(_0483_));
 sg13g2_xor2_1 _4824_ (.B(_0483_),
    .A(_0464_),
    .X(_0484_));
 sg13g2_nand2b_1 _4825_ (.Y(_0485_),
    .B(_0484_),
    .A_N(_0459_));
 sg13g2_nor2b_1 _4826_ (.A(_0484_),
    .B_N(_0459_),
    .Y(_0486_));
 sg13g2_xnor2_1 _4827_ (.Y(_0487_),
    .A(_0459_),
    .B(_0484_));
 sg13g2_xnor2_1 _4828_ (.Y(_0488_),
    .A(_0458_),
    .B(_0487_));
 sg13g2_nor2b_1 _4829_ (.A(_0451_),
    .B_N(_0488_),
    .Y(_0489_));
 sg13g2_xnor2_1 _4830_ (.Y(_0490_),
    .A(_0451_),
    .B(_0488_));
 sg13g2_xor2_1 _4831_ (.B(_0490_),
    .A(_0450_),
    .X(_0491_));
 sg13g2_nor2_1 _4832_ (.A(_0449_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_nand2b_1 _4833_ (.Y(_0493_),
    .B(_0448_),
    .A_N(_0491_));
 sg13g2_xnor2_1 _4834_ (.Y(_0494_),
    .A(_0448_),
    .B(_0491_));
 sg13g2_xor2_1 _4835_ (.B(_0446_),
    .A(_0445_),
    .X(_0495_));
 sg13g2_nor3_1 _4836_ (.A(net890),
    .B(_0287_),
    .C(_0288_),
    .Y(_0496_));
 sg13g2_nor3_2 _4837_ (.A(net802),
    .B(_0287_),
    .C(_0288_),
    .Y(_0497_));
 sg13g2_nand2_1 _4838_ (.Y(_0498_),
    .A(_0283_),
    .B(_0497_));
 sg13g2_or2_1 _4839_ (.X(_0499_),
    .B(net725),
    .A(_0292_));
 sg13g2_xnor2_1 _4840_ (.Y(_0500_),
    .A(_0283_),
    .B(_0497_));
 sg13g2_o21ai_1 _4841_ (.B1(_0498_),
    .Y(_0501_),
    .A1(_0499_),
    .A2(_0500_));
 sg13g2_xor2_1 _4842_ (.B(_0294_),
    .A(_0293_),
    .X(_0502_));
 sg13g2_nand2_1 _4843_ (.Y(_0503_),
    .A(_0501_),
    .B(_0502_));
 sg13g2_nand2_1 _4844_ (.Y(_0504_),
    .A(net757),
    .B(net727));
 sg13g2_inv_1 _4845_ (.Y(_0505_),
    .A(_0504_));
 sg13g2_nand2_1 _4846_ (.Y(_0506_),
    .A(net726),
    .B(net785));
 sg13g2_nand2_1 _4847_ (.Y(_0507_),
    .A(_0327_),
    .B(net771));
 sg13g2_nor2_1 _4848_ (.A(_0338_),
    .B(_0506_),
    .Y(_0508_));
 sg13g2_o21ai_1 _4849_ (.B1(_0507_),
    .Y(_0509_),
    .A1(net784),
    .A2(net725));
 sg13g2_nor2b_1 _4850_ (.A(_0508_),
    .B_N(_0509_),
    .Y(_0510_));
 sg13g2_xnor2_1 _4851_ (.Y(_0511_),
    .A(_0504_),
    .B(_0510_));
 sg13g2_inv_1 _4852_ (.Y(_0512_),
    .A(_0511_));
 sg13g2_xnor2_1 _4853_ (.Y(_0513_),
    .A(_0501_),
    .B(_0502_));
 sg13g2_o21ai_1 _4854_ (.B1(_0503_),
    .Y(_0514_),
    .A1(_0512_),
    .A2(_0513_));
 sg13g2_xnor2_1 _4855_ (.Y(_0515_),
    .A(_0320_),
    .B(_0341_));
 sg13g2_nand2_1 _4856_ (.Y(_0516_),
    .A(_0514_),
    .B(_0515_));
 sg13g2_a21oi_1 _4857_ (.A1(_0505_),
    .A2(_0509_),
    .Y(_0517_),
    .B1(_0508_));
 sg13g2_xnor2_1 _4858_ (.Y(_0518_),
    .A(_0383_),
    .B(_0384_));
 sg13g2_nand2b_1 _4859_ (.Y(_0519_),
    .B(_0518_),
    .A_N(_0517_));
 sg13g2_xnor2_1 _4860_ (.Y(_0520_),
    .A(_0517_),
    .B(_0518_));
 sg13g2_xnor2_1 _4861_ (.Y(_0521_),
    .A(_0249_),
    .B(_0263_));
 sg13g2_nor2_2 _4862_ (.A(_0380_),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_nand3_1 _4863_ (.B(_0520_),
    .C(_0522_),
    .A(_0384_),
    .Y(_0523_));
 sg13g2_a21o_1 _4864_ (.A2(_0522_),
    .A1(_0384_),
    .B1(_0520_),
    .X(_0524_));
 sg13g2_nor2_1 _4865_ (.A(_0375_),
    .B(_0521_),
    .Y(_0525_));
 sg13g2_nand2_1 _4866_ (.Y(_0526_),
    .A(_0523_),
    .B(_0524_));
 sg13g2_xnor2_1 _4867_ (.Y(_0527_),
    .A(_0514_),
    .B(_0515_));
 sg13g2_o21ai_1 _4868_ (.B1(_0516_),
    .Y(_0528_),
    .A1(_0526_),
    .A2(_0527_));
 sg13g2_xnor2_1 _4869_ (.Y(_0529_),
    .A(_0372_),
    .B(_0394_));
 sg13g2_nor2b_1 _4870_ (.A(_0529_),
    .B_N(_0528_),
    .Y(_0530_));
 sg13g2_inv_1 _4871_ (.Y(_0531_),
    .A(_0530_));
 sg13g2_and2_1 _4872_ (.A(_0519_),
    .B(_0523_),
    .X(_0532_));
 sg13g2_xor2_1 _4873_ (.B(_0529_),
    .A(_0528_),
    .X(_0533_));
 sg13g2_or2_1 _4874_ (.X(_0534_),
    .B(_0533_),
    .A(_0532_));
 sg13g2_a21oi_1 _4875_ (.A1(_0531_),
    .A2(_0534_),
    .Y(_0535_),
    .B1(_0495_));
 sg13g2_inv_1 _4876_ (.Y(_0536_),
    .A(_0535_));
 sg13g2_nand3_1 _4877_ (.B(_0531_),
    .C(_0534_),
    .A(_0495_),
    .Y(_0537_));
 sg13g2_nor2b_1 _4878_ (.A(_0535_),
    .B_N(_0537_),
    .Y(_0538_));
 sg13g2_inv_1 _4879_ (.Y(_0539_),
    .A(_0538_));
 sg13g2_nor3_2 _4880_ (.A(net890),
    .B(_0270_),
    .C(_0335_),
    .Y(_0540_));
 sg13g2_nor2_1 _4881_ (.A(net802),
    .B(net725),
    .Y(_0541_));
 sg13g2_nand2_1 _4882_ (.Y(_0542_),
    .A(net787),
    .B(net726));
 sg13g2_inv_1 _4883_ (.Y(_0543_),
    .A(_0542_));
 sg13g2_xor2_1 _4884_ (.B(_0541_),
    .A(_0496_),
    .X(_0544_));
 sg13g2_a22oi_1 _4885_ (.Y(_0545_),
    .B1(_0543_),
    .B2(_0544_),
    .A2(_0540_),
    .A1(_0497_));
 sg13g2_xor2_1 _4886_ (.B(_0500_),
    .A(_0499_),
    .X(_0546_));
 sg13g2_nor2b_1 _4887_ (.A(_0545_),
    .B_N(_0546_),
    .Y(_0547_));
 sg13g2_or2_1 _4888_ (.X(_0548_),
    .B(_0381_),
    .A(_0325_));
 sg13g2_inv_1 _4889_ (.Y(_0549_),
    .A(_0548_));
 sg13g2_nand2_1 _4890_ (.Y(_0550_),
    .A(net785),
    .B(_0373_));
 sg13g2_and2_1 _4891_ (.A(net771),
    .B(net727),
    .X(_0551_));
 sg13g2_nor2_1 _4892_ (.A(_0507_),
    .B(_0550_),
    .Y(_0552_));
 sg13g2_xnor2_1 _4893_ (.Y(_0553_),
    .A(_0506_),
    .B(_0551_));
 sg13g2_xnor2_1 _4894_ (.Y(_0554_),
    .A(_0548_),
    .B(_0553_));
 sg13g2_xnor2_1 _4895_ (.Y(_0555_),
    .A(_0545_),
    .B(_0546_));
 sg13g2_a21o_1 _4896_ (.A2(_0555_),
    .A1(_0554_),
    .B1(_0547_),
    .X(_0556_));
 sg13g2_xnor2_1 _4897_ (.Y(_0557_),
    .A(_0512_),
    .B(_0513_));
 sg13g2_nand2b_1 _4898_ (.Y(_0558_),
    .B(_0556_),
    .A_N(_0557_));
 sg13g2_a21oi_1 _4899_ (.A1(_0549_),
    .A2(_0553_),
    .Y(_0559_),
    .B1(_0552_));
 sg13g2_xor2_1 _4900_ (.B(_0525_),
    .A(_0382_),
    .X(_0560_));
 sg13g2_inv_1 _4901_ (.Y(_0561_),
    .A(_0560_));
 sg13g2_xnor2_1 _4902_ (.Y(_0562_),
    .A(_0559_),
    .B(_0560_));
 sg13g2_nand2b_1 _4903_ (.Y(_0563_),
    .B(_0256_),
    .A_N(_0255_));
 sg13g2_xnor2_1 _4904_ (.Y(_0564_),
    .A(_0262_),
    .B(_0563_));
 sg13g2_and2_1 _4905_ (.A(net747),
    .B(net729),
    .X(_0565_));
 sg13g2_nand3_1 _4906_ (.B(_0562_),
    .C(_0565_),
    .A(_0525_),
    .Y(_0566_));
 sg13g2_a21o_1 _4907_ (.A2(_0565_),
    .A1(_0525_),
    .B1(_0562_),
    .X(_0567_));
 sg13g2_and2_1 _4908_ (.A(net755),
    .B(net729),
    .X(_0568_));
 sg13g2_nand2_1 _4909_ (.Y(_0569_),
    .A(_0566_),
    .B(_0567_));
 sg13g2_xor2_1 _4910_ (.B(_0557_),
    .A(_0556_),
    .X(_0570_));
 sg13g2_o21ai_1 _4911_ (.B1(_0558_),
    .Y(_0571_),
    .A1(_0569_),
    .A2(_0570_));
 sg13g2_xor2_1 _4912_ (.B(_0527_),
    .A(_0526_),
    .X(_0572_));
 sg13g2_nand2_1 _4913_ (.Y(_0573_),
    .A(_0571_),
    .B(_0572_));
 sg13g2_o21ai_1 _4914_ (.B1(_0566_),
    .Y(_0574_),
    .A1(_0559_),
    .A2(_0561_));
 sg13g2_xnor2_1 _4915_ (.Y(_0575_),
    .A(_0571_),
    .B(_0572_));
 sg13g2_nand2b_1 _4916_ (.Y(_0576_),
    .B(_0574_),
    .A_N(_0575_));
 sg13g2_xnor2_1 _4917_ (.Y(_0577_),
    .A(_0532_),
    .B(_0533_));
 sg13g2_nand3_1 _4918_ (.B(_0576_),
    .C(_0577_),
    .A(_0573_),
    .Y(_0578_));
 sg13g2_a21o_1 _4919_ (.A2(_0576_),
    .A1(_0573_),
    .B1(_0577_),
    .X(_0579_));
 sg13g2_xor2_1 _4920_ (.B(_0575_),
    .A(_0574_),
    .X(_0580_));
 sg13g2_nand2_1 _4921_ (.Y(_0581_),
    .A(net804),
    .B(net726));
 sg13g2_nor3_1 _4922_ (.A(net891),
    .B(net725),
    .C(_0581_),
    .Y(_0582_));
 sg13g2_nand2_1 _4923_ (.Y(_0583_),
    .A(net787),
    .B(net727));
 sg13g2_inv_1 _4924_ (.Y(_0584_),
    .A(_0583_));
 sg13g2_xnor2_1 _4925_ (.Y(_0585_),
    .A(_0540_),
    .B(_0581_));
 sg13g2_a21oi_1 _4926_ (.A1(_0584_),
    .A2(_0585_),
    .Y(_0586_),
    .B1(_0582_));
 sg13g2_xnor2_1 _4927_ (.Y(_0587_),
    .A(_0543_),
    .B(_0544_));
 sg13g2_nor2_1 _4928_ (.A(_0586_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_nor2_1 _4929_ (.A(_0325_),
    .B(_0521_),
    .Y(_0589_));
 sg13g2_nor2_1 _4930_ (.A(net784),
    .B(_0381_),
    .Y(_0590_));
 sg13g2_nor2_1 _4931_ (.A(_0331_),
    .B(_0381_),
    .Y(_0591_));
 sg13g2_and2_1 _4932_ (.A(_0551_),
    .B(_0590_),
    .X(_0592_));
 sg13g2_xnor2_1 _4933_ (.Y(_0593_),
    .A(_0550_),
    .B(_0591_));
 sg13g2_xor2_1 _4934_ (.B(_0593_),
    .A(_0589_),
    .X(_0594_));
 sg13g2_xor2_1 _4935_ (.B(_0587_),
    .A(_0586_),
    .X(_0595_));
 sg13g2_a21oi_1 _4936_ (.A1(_0594_),
    .A2(_0595_),
    .Y(_0596_),
    .B1(_0588_));
 sg13g2_xnor2_1 _4937_ (.Y(_0597_),
    .A(_0554_),
    .B(_0555_));
 sg13g2_nor2_1 _4938_ (.A(_0596_),
    .B(_0597_),
    .Y(_0598_));
 sg13g2_xor2_1 _4939_ (.B(_0260_),
    .A(_0257_),
    .X(_0599_));
 sg13g2_xnor2_1 _4940_ (.Y(_0600_),
    .A(_0257_),
    .B(_0260_));
 sg13g2_nor2_1 _4941_ (.A(_0380_),
    .B(_0599_),
    .Y(_0601_));
 sg13g2_nor2_1 _4942_ (.A(_0375_),
    .B(_0599_),
    .Y(_0602_));
 sg13g2_nand2_1 _4943_ (.Y(_0603_),
    .A(_0565_),
    .B(_0602_));
 sg13g2_a21o_1 _4944_ (.A2(_0593_),
    .A1(_0589_),
    .B1(_0592_),
    .X(_0604_));
 sg13g2_xnor2_1 _4945_ (.Y(_0605_),
    .A(_0522_),
    .B(_0568_));
 sg13g2_nand2b_1 _4946_ (.Y(_0606_),
    .B(_0604_),
    .A_N(_0605_));
 sg13g2_xor2_1 _4947_ (.B(_0605_),
    .A(_0604_),
    .X(_0607_));
 sg13g2_xor2_1 _4948_ (.B(_0607_),
    .A(_0603_),
    .X(_0608_));
 sg13g2_xor2_1 _4949_ (.B(_0597_),
    .A(_0596_),
    .X(_0609_));
 sg13g2_a21oi_1 _4950_ (.A1(_0608_),
    .A2(_0609_),
    .Y(_0610_),
    .B1(_0598_));
 sg13g2_xor2_1 _4951_ (.B(_0570_),
    .A(_0569_),
    .X(_0611_));
 sg13g2_nor2b_1 _4952_ (.A(_0610_),
    .B_N(_0611_),
    .Y(_0612_));
 sg13g2_o21ai_1 _4953_ (.B1(_0606_),
    .Y(_0613_),
    .A1(_0603_),
    .A2(_0607_));
 sg13g2_xnor2_1 _4954_ (.Y(_0614_),
    .A(_0610_),
    .B(_0611_));
 sg13g2_a21oi_1 _4955_ (.A1(_0613_),
    .A2(_0614_),
    .Y(_0615_),
    .B1(_0612_));
 sg13g2_nor2_1 _4956_ (.A(_0580_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_nand2_1 _4957_ (.Y(_0617_),
    .A(_0578_),
    .B(_0616_));
 sg13g2_nand2_1 _4958_ (.Y(_0618_),
    .A(_0579_),
    .B(_0617_));
 sg13g2_nand2_1 _4959_ (.Y(_0619_),
    .A(net814),
    .B(net727));
 sg13g2_and2_1 _4960_ (.A(net804),
    .B(net727),
    .X(_0620_));
 sg13g2_nor2_1 _4961_ (.A(_0581_),
    .B(_0619_),
    .Y(_0621_));
 sg13g2_nand3_1 _4962_ (.B(net726),
    .C(_0620_),
    .A(net814),
    .Y(_0622_));
 sg13g2_nor2_1 _4963_ (.A(_0292_),
    .B(_0381_),
    .Y(_0623_));
 sg13g2_a21o_1 _4964_ (.A2(net726),
    .A1(net814),
    .B1(_0620_),
    .X(_0624_));
 sg13g2_and3_1 _4965_ (.X(_0625_),
    .A(_0622_),
    .B(_0623_),
    .C(_0624_));
 sg13g2_nor2_1 _4966_ (.A(_0621_),
    .B(_0625_),
    .Y(_0626_));
 sg13g2_xnor2_1 _4967_ (.Y(_0627_),
    .A(_0584_),
    .B(_0585_));
 sg13g2_nor2_1 _4968_ (.A(_0626_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nand2_1 _4969_ (.Y(_0629_),
    .A(net757),
    .B(net729));
 sg13g2_nor2_1 _4970_ (.A(net784),
    .B(_0521_),
    .Y(_0630_));
 sg13g2_nor2_1 _4971_ (.A(_0331_),
    .B(_0521_),
    .Y(_0631_));
 sg13g2_nand2_1 _4972_ (.Y(_0632_),
    .A(_0591_),
    .B(_0630_));
 sg13g2_nor2_1 _4973_ (.A(_0590_),
    .B(_0631_),
    .Y(_0633_));
 sg13g2_a21oi_1 _4974_ (.A1(_0591_),
    .A2(_0630_),
    .Y(_0634_),
    .B1(_0633_));
 sg13g2_xnor2_1 _4975_ (.Y(_0635_),
    .A(_0629_),
    .B(_0634_));
 sg13g2_xor2_1 _4976_ (.B(_0627_),
    .A(_0626_),
    .X(_0636_));
 sg13g2_a21oi_1 _4977_ (.A1(_0635_),
    .A2(_0636_),
    .Y(_0637_),
    .B1(_0628_));
 sg13g2_xor2_1 _4978_ (.B(_0595_),
    .A(_0594_),
    .X(_0638_));
 sg13g2_nor2b_1 _4979_ (.A(_0637_),
    .B_N(_0638_),
    .Y(_0639_));
 sg13g2_o21ai_1 _4980_ (.B1(_0632_),
    .Y(_0640_),
    .A1(_0629_),
    .A2(_0633_));
 sg13g2_xor2_1 _4981_ (.B(_0602_),
    .A(_0565_),
    .X(_0641_));
 sg13g2_nand2_1 _4982_ (.Y(_0642_),
    .A(_0640_),
    .B(_0641_));
 sg13g2_xnor2_1 _4983_ (.Y(_0643_),
    .A(_0640_),
    .B(_0641_));
 sg13g2_xnor2_1 _4984_ (.Y(_0644_),
    .A(net885),
    .B(_0259_));
 sg13g2_nand2_1 _4985_ (.Y(_0645_),
    .A(net755),
    .B(net783));
 sg13g2_nand3_1 _4986_ (.B(_0601_),
    .C(_0644_),
    .A(net755),
    .Y(_0646_));
 sg13g2_xor2_1 _4987_ (.B(_0646_),
    .A(_0643_),
    .X(_0647_));
 sg13g2_xnor2_1 _4988_ (.Y(_0648_),
    .A(_0637_),
    .B(_0638_));
 sg13g2_a21oi_1 _4989_ (.A1(_0647_),
    .A2(_0648_),
    .Y(_0649_),
    .B1(_0639_));
 sg13g2_xnor2_1 _4990_ (.Y(_0650_),
    .A(_0608_),
    .B(_0609_));
 sg13g2_nor2_1 _4991_ (.A(_0649_),
    .B(_0650_),
    .Y(_0651_));
 sg13g2_o21ai_1 _4992_ (.B1(_0642_),
    .Y(_0652_),
    .A1(_0643_),
    .A2(_0646_));
 sg13g2_xor2_1 _4993_ (.B(_0650_),
    .A(_0649_),
    .X(_0653_));
 sg13g2_a21oi_1 _4994_ (.A1(_0652_),
    .A2(_0653_),
    .Y(_0654_),
    .B1(_0651_));
 sg13g2_xnor2_1 _4995_ (.Y(_0655_),
    .A(_0613_),
    .B(_0614_));
 sg13g2_or2_1 _4996_ (.X(_0656_),
    .B(_0655_),
    .A(_0654_));
 sg13g2_nor2_1 _4997_ (.A(net890),
    .B(_0381_),
    .Y(_0657_));
 sg13g2_nor2_1 _4998_ (.A(net802),
    .B(_0381_),
    .Y(_0658_));
 sg13g2_nor2_1 _4999_ (.A(_0292_),
    .B(_0521_),
    .Y(_0659_));
 sg13g2_xnor2_1 _5000_ (.Y(_0660_),
    .A(_0619_),
    .B(_0658_));
 sg13g2_a22oi_1 _5001_ (.Y(_0661_),
    .B1(_0659_),
    .B2(_0660_),
    .A2(_0657_),
    .A1(_0620_));
 sg13g2_a21oi_1 _5002_ (.A1(_0622_),
    .A2(_0624_),
    .Y(_0662_),
    .B1(_0623_));
 sg13g2_nor3_1 _5003_ (.A(_0625_),
    .B(_0661_),
    .C(_0662_),
    .Y(_0663_));
 sg13g2_nand2_1 _5004_ (.Y(_0664_),
    .A(net757),
    .B(_0600_));
 sg13g2_and2_1 _5005_ (.A(net785),
    .B(_0564_),
    .X(_0665_));
 sg13g2_a21oi_1 _5006_ (.A1(net771),
    .A2(net729),
    .Y(_0666_),
    .B1(_0630_));
 sg13g2_a21o_1 _5007_ (.A2(_0665_),
    .A1(_0631_),
    .B1(_0666_),
    .X(_0667_));
 sg13g2_nor2_1 _5008_ (.A(_0664_),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_xor2_1 _5009_ (.B(_0667_),
    .A(_0664_),
    .X(_0669_));
 sg13g2_o21ai_1 _5010_ (.B1(_0661_),
    .Y(_0670_),
    .A1(_0625_),
    .A2(_0662_));
 sg13g2_nor2b_1 _5011_ (.A(_0663_),
    .B_N(_0670_),
    .Y(_0671_));
 sg13g2_a21oi_2 _5012_ (.B1(_0663_),
    .Y(_0672_),
    .A2(_0670_),
    .A1(_0669_));
 sg13g2_xnor2_1 _5013_ (.Y(_0673_),
    .A(_0635_),
    .B(_0636_));
 sg13g2_nor2_1 _5014_ (.A(_0672_),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_a21oi_2 _5015_ (.B1(_0668_),
    .Y(_0675_),
    .A2(_0665_),
    .A1(_0631_));
 sg13g2_xnor2_1 _5016_ (.Y(_0676_),
    .A(_0601_),
    .B(_0645_));
 sg13g2_nor2b_1 _5017_ (.A(_0675_),
    .B_N(_0676_),
    .Y(_0677_));
 sg13g2_xnor2_1 _5018_ (.Y(_0678_),
    .A(_0675_),
    .B(_0676_));
 sg13g2_xor2_1 _5019_ (.B(_3132_),
    .A(_0012_),
    .X(_0679_));
 sg13g2_nand2_1 _5020_ (.Y(_0680_),
    .A(net747),
    .B(net782));
 sg13g2_and4_1 _5021_ (.A(net755),
    .B(net747),
    .C(net783),
    .D(net782),
    .X(_0681_));
 sg13g2_xnor2_1 _5022_ (.Y(_0682_),
    .A(_0678_),
    .B(_0681_));
 sg13g2_inv_1 _5023_ (.Y(_0683_),
    .A(_0682_));
 sg13g2_xor2_1 _5024_ (.B(_0673_),
    .A(_0672_),
    .X(_0684_));
 sg13g2_a21oi_1 _5025_ (.A1(_0683_),
    .A2(_0684_),
    .Y(_0685_),
    .B1(_0674_));
 sg13g2_xnor2_1 _5026_ (.Y(_0686_),
    .A(_0647_),
    .B(_0648_));
 sg13g2_nor2_1 _5027_ (.A(_0685_),
    .B(_0686_),
    .Y(_0687_));
 sg13g2_a21oi_1 _5028_ (.A1(_0678_),
    .A2(_0681_),
    .Y(_0688_),
    .B1(_0677_));
 sg13g2_inv_1 _5029_ (.Y(_0689_),
    .A(_0688_));
 sg13g2_xor2_1 _5030_ (.B(_0686_),
    .A(_0685_),
    .X(_0690_));
 sg13g2_a21oi_1 _5031_ (.A1(_0689_),
    .A2(_0690_),
    .Y(_0691_),
    .B1(_0687_));
 sg13g2_xnor2_1 _5032_ (.Y(_0692_),
    .A(_0652_),
    .B(_0653_));
 sg13g2_nor2_1 _5033_ (.A(_0691_),
    .B(_0692_),
    .Y(_0693_));
 sg13g2_nor2_1 _5034_ (.A(net890),
    .B(_0521_),
    .Y(_0694_));
 sg13g2_nor2_1 _5035_ (.A(net802),
    .B(_0521_),
    .Y(_0695_));
 sg13g2_nand2_1 _5036_ (.Y(_0696_),
    .A(net787),
    .B(net729));
 sg13g2_inv_1 _5037_ (.Y(_0697_),
    .A(_0696_));
 sg13g2_xor2_1 _5038_ (.B(_0695_),
    .A(_0657_),
    .X(_0698_));
 sg13g2_a22oi_1 _5039_ (.Y(_0699_),
    .B1(_0697_),
    .B2(_0698_),
    .A2(_0694_),
    .A1(_0658_));
 sg13g2_xnor2_1 _5040_ (.Y(_0700_),
    .A(_0659_),
    .B(_0660_));
 sg13g2_nor2_1 _5041_ (.A(_0699_),
    .B(_0700_),
    .Y(_0701_));
 sg13g2_nand2_1 _5042_ (.Y(_0702_),
    .A(net757),
    .B(_0644_));
 sg13g2_nor2_1 _5043_ (.A(net784),
    .B(_0599_),
    .Y(_0703_));
 sg13g2_nand2_1 _5044_ (.Y(_0704_),
    .A(net771),
    .B(_0600_));
 sg13g2_nand3_1 _5045_ (.B(net729),
    .C(_0703_),
    .A(net771),
    .Y(_0705_));
 sg13g2_xnor2_1 _5046_ (.Y(_0706_),
    .A(_0665_),
    .B(_0704_));
 sg13g2_nand2b_1 _5047_ (.Y(_0707_),
    .B(_0706_),
    .A_N(_0702_));
 sg13g2_xnor2_1 _5048_ (.Y(_0708_),
    .A(_0702_),
    .B(_0706_));
 sg13g2_xor2_1 _5049_ (.B(_0700_),
    .A(_0699_),
    .X(_0709_));
 sg13g2_a21oi_2 _5050_ (.B1(_0701_),
    .Y(_0710_),
    .A2(_0709_),
    .A1(_0708_));
 sg13g2_xnor2_1 _5051_ (.Y(_0711_),
    .A(_0669_),
    .B(_0671_));
 sg13g2_nor2_1 _5052_ (.A(_0710_),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_nand2_1 _5053_ (.Y(_0713_),
    .A(_0705_),
    .B(_0707_));
 sg13g2_a22oi_1 _5054_ (.Y(_0714_),
    .B1(net782),
    .B2(net755),
    .A2(net783),
    .A1(net747));
 sg13g2_or2_1 _5055_ (.X(_0715_),
    .B(_0714_),
    .A(_0681_));
 sg13g2_a21oi_1 _5056_ (.A1(_0705_),
    .A2(_0707_),
    .Y(_0716_),
    .B1(_0715_));
 sg13g2_xnor2_1 _5057_ (.Y(_0717_),
    .A(_0713_),
    .B(_0715_));
 sg13g2_nand2_1 _5058_ (.Y(_0718_),
    .A(_0710_),
    .B(_0711_));
 sg13g2_xnor2_1 _5059_ (.Y(_0719_),
    .A(_0710_),
    .B(_0711_));
 sg13g2_a21oi_1 _5060_ (.A1(_0717_),
    .A2(_0718_),
    .Y(_0720_),
    .B1(_0712_));
 sg13g2_xnor2_1 _5061_ (.Y(_0721_),
    .A(_0682_),
    .B(_0684_));
 sg13g2_nand2b_1 _5062_ (.Y(_0722_),
    .B(_0721_),
    .A_N(_0720_));
 sg13g2_xnor2_1 _5063_ (.Y(_0723_),
    .A(_0720_),
    .B(_0721_));
 sg13g2_nand2_1 _5064_ (.Y(_0724_),
    .A(_0716_),
    .B(_0723_));
 sg13g2_and2_1 _5065_ (.A(_0722_),
    .B(_0724_),
    .X(_0725_));
 sg13g2_xnor2_1 _5066_ (.Y(_0726_),
    .A(_0688_),
    .B(_0690_));
 sg13g2_nand2b_1 _5067_ (.Y(_0727_),
    .B(_0726_),
    .A_N(_0725_));
 sg13g2_xor2_1 _5068_ (.B(_0726_),
    .A(_0725_),
    .X(_0728_));
 sg13g2_xnor2_1 _5069_ (.Y(_0729_),
    .A(_0716_),
    .B(_0723_));
 sg13g2_xnor2_1 _5070_ (.Y(_0730_),
    .A(_0717_),
    .B(_0719_));
 sg13g2_and2_1 _5071_ (.A(net814),
    .B(net729),
    .X(_0731_));
 sg13g2_nand2_1 _5072_ (.Y(_0732_),
    .A(net787),
    .B(_0600_));
 sg13g2_a21oi_1 _5073_ (.A1(net804),
    .A2(net729),
    .Y(_0733_),
    .B1(_0694_));
 sg13g2_a21o_1 _5074_ (.A2(_0731_),
    .A1(_0695_),
    .B1(_0733_),
    .X(_0734_));
 sg13g2_nor2_1 _5075_ (.A(_0732_),
    .B(_0734_),
    .Y(_0735_));
 sg13g2_a21oi_1 _5076_ (.A1(_0695_),
    .A2(_0731_),
    .Y(_0736_),
    .B1(_0735_));
 sg13g2_xnor2_1 _5077_ (.Y(_0737_),
    .A(_0697_),
    .B(_0698_));
 sg13g2_nor2_1 _5078_ (.A(_0736_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_nand2_1 _5079_ (.Y(_0739_),
    .A(net757),
    .B(_0679_));
 sg13g2_nand2_1 _5080_ (.Y(_0740_),
    .A(net771),
    .B(net783));
 sg13g2_nand3_1 _5081_ (.B(net783),
    .C(_0703_),
    .A(net771),
    .Y(_0741_));
 sg13g2_xor2_1 _5082_ (.B(_0740_),
    .A(_0703_),
    .X(_0742_));
 sg13g2_xor2_1 _5083_ (.B(_0742_),
    .A(_0739_),
    .X(_0743_));
 sg13g2_xor2_1 _5084_ (.B(_0737_),
    .A(_0736_),
    .X(_0744_));
 sg13g2_a21oi_1 _5085_ (.A1(_0743_),
    .A2(_0744_),
    .Y(_0745_),
    .B1(_0738_));
 sg13g2_xnor2_1 _5086_ (.Y(_0746_),
    .A(_0708_),
    .B(_0709_));
 sg13g2_nor2_1 _5087_ (.A(_0745_),
    .B(_0746_),
    .Y(_0747_));
 sg13g2_o21ai_1 _5088_ (.B1(_0741_),
    .Y(_0748_),
    .A1(_0739_),
    .A2(_0742_));
 sg13g2_nand2b_1 _5089_ (.Y(_0749_),
    .B(_0748_),
    .A_N(_0680_));
 sg13g2_inv_1 _5090_ (.Y(_0750_),
    .A(_0749_));
 sg13g2_xnor2_1 _5091_ (.Y(_0751_),
    .A(_0680_),
    .B(_0748_));
 sg13g2_xor2_1 _5092_ (.B(_0746_),
    .A(_0745_),
    .X(_0752_));
 sg13g2_a21oi_1 _5093_ (.A1(_0751_),
    .A2(_0752_),
    .Y(_0753_),
    .B1(_0747_));
 sg13g2_nand2b_1 _5094_ (.Y(_0754_),
    .B(_0730_),
    .A_N(_0753_));
 sg13g2_xnor2_1 _5095_ (.Y(_0755_),
    .A(_0730_),
    .B(_0753_));
 sg13g2_nand2_1 _5096_ (.Y(_0756_),
    .A(net785),
    .B(net782));
 sg13g2_or2_1 _5097_ (.X(_0757_),
    .B(_0756_),
    .A(_0740_));
 sg13g2_inv_1 _5098_ (.Y(_0758_),
    .A(_0757_));
 sg13g2_xnor2_1 _5099_ (.Y(_0759_),
    .A(_0743_),
    .B(_0744_));
 sg13g2_nor2_1 _5100_ (.A(net890),
    .B(_0599_),
    .Y(_0760_));
 sg13g2_nor2_1 _5101_ (.A(net802),
    .B(_0599_),
    .Y(_0761_));
 sg13g2_nand2_1 _5102_ (.Y(_0762_),
    .A(net787),
    .B(net783));
 sg13g2_xnor2_1 _5103_ (.Y(_0763_),
    .A(_0731_),
    .B(_0761_));
 sg13g2_nor2_1 _5104_ (.A(_0762_),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_a21oi_1 _5105_ (.A1(_0731_),
    .A2(_0761_),
    .Y(_0765_),
    .B1(_0764_));
 sg13g2_xor2_1 _5106_ (.B(_0734_),
    .A(_0732_),
    .X(_0766_));
 sg13g2_nor2b_1 _5107_ (.A(_0765_),
    .B_N(_0766_),
    .Y(_0767_));
 sg13g2_a22oi_1 _5108_ (.Y(_0768_),
    .B1(net782),
    .B2(net771),
    .A2(net783),
    .A1(net785));
 sg13g2_nor2_1 _5109_ (.A(_0758_),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_xnor2_1 _5110_ (.Y(_0770_),
    .A(_0765_),
    .B(_0766_));
 sg13g2_a21oi_1 _5111_ (.A1(_0769_),
    .A2(_0770_),
    .Y(_0771_),
    .B1(_0767_));
 sg13g2_nor2_1 _5112_ (.A(_0759_),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_xnor2_1 _5113_ (.Y(_0773_),
    .A(_0759_),
    .B(_0771_));
 sg13g2_and2_1 _5114_ (.A(net804),
    .B(net783),
    .X(_0774_));
 sg13g2_xor2_1 _5115_ (.B(_0774_),
    .A(_0760_),
    .X(_0775_));
 sg13g2_and3_1 _5116_ (.X(_0776_),
    .A(net787),
    .B(net782),
    .C(_0775_));
 sg13g2_a21oi_1 _5117_ (.A1(_0760_),
    .A2(_0774_),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_xnor2_1 _5118_ (.Y(_0778_),
    .A(_0762_),
    .B(_0763_));
 sg13g2_nor2_1 _5119_ (.A(_0777_),
    .B(_0778_),
    .Y(_0779_));
 sg13g2_and2_1 _5120_ (.A(_0777_),
    .B(_0778_),
    .X(_0780_));
 sg13g2_o21ai_1 _5121_ (.B1(_0756_),
    .Y(_0781_),
    .A1(_0779_),
    .A2(_0780_));
 sg13g2_a21oi_1 _5122_ (.A1(net787),
    .A2(net782),
    .Y(_0782_),
    .B1(_0775_));
 sg13g2_nor3_1 _5123_ (.A(net890),
    .B(_0776_),
    .C(_0782_),
    .Y(_0783_));
 sg13g2_and4_1 _5124_ (.A(net782),
    .B(_0774_),
    .C(_0781_),
    .D(_0783_),
    .X(_0784_));
 sg13g2_nor2_1 _5125_ (.A(_0756_),
    .B(_0780_),
    .Y(_0785_));
 sg13g2_or3_1 _5126_ (.A(_0779_),
    .B(_0784_),
    .C(_0785_),
    .X(_0786_));
 sg13g2_xor2_1 _5127_ (.B(_0770_),
    .A(_0769_),
    .X(_0787_));
 sg13g2_a22oi_1 _5128_ (.Y(_0788_),
    .B1(_0786_),
    .B2(_0787_),
    .A2(_0784_),
    .A1(_0779_));
 sg13g2_a21oi_1 _5129_ (.A1(_0757_),
    .A2(_0773_),
    .Y(_0789_),
    .B1(_0788_));
 sg13g2_nor2_1 _5130_ (.A(_0757_),
    .B(_0773_),
    .Y(_0790_));
 sg13g2_nor3_1 _5131_ (.A(_0772_),
    .B(_0789_),
    .C(_0790_),
    .Y(_0791_));
 sg13g2_xor2_1 _5132_ (.B(_0752_),
    .A(_0751_),
    .X(_0792_));
 sg13g2_a21oi_1 _5133_ (.A1(_0772_),
    .A2(_0789_),
    .Y(_0793_),
    .B1(_0792_));
 sg13g2_nor2_1 _5134_ (.A(_0791_),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_o21ai_1 _5135_ (.B1(_0794_),
    .Y(_0795_),
    .A1(_0750_),
    .A2(_0755_));
 sg13g2_nand2_1 _5136_ (.Y(_0796_),
    .A(_0750_),
    .B(_0755_));
 sg13g2_a21oi_1 _5137_ (.A1(_0729_),
    .A2(_0795_),
    .Y(_0797_),
    .B1(_0754_));
 sg13g2_a21oi_1 _5138_ (.A1(_0795_),
    .A2(_0796_),
    .Y(_0798_),
    .B1(_0729_));
 sg13g2_nor2_1 _5139_ (.A(_0797_),
    .B(_0798_),
    .Y(_0799_));
 sg13g2_o21ai_1 _5140_ (.B1(_0727_),
    .Y(_0800_),
    .A1(_0799_),
    .A2(_0728_));
 sg13g2_xor2_1 _5141_ (.B(_0692_),
    .A(_0691_),
    .X(_0801_));
 sg13g2_a21oi_2 _5142_ (.B1(_0693_),
    .Y(_0802_),
    .A2(_0801_),
    .A1(_0800_));
 sg13g2_xor2_1 _5143_ (.B(_0655_),
    .A(_0654_),
    .X(_0803_));
 sg13g2_inv_1 _5144_ (.Y(_0804_),
    .A(_0803_));
 sg13g2_o21ai_1 _5145_ (.B1(_0656_),
    .Y(_0805_),
    .A1(_0804_),
    .A2(_0802_));
 sg13g2_nand2_1 _5146_ (.Y(_0806_),
    .A(_0578_),
    .B(_0579_));
 sg13g2_xor2_1 _5147_ (.B(_0615_),
    .A(_0580_),
    .X(_0807_));
 sg13g2_nor2b_1 _5148_ (.A(_0806_),
    .B_N(_0807_),
    .Y(_0808_));
 sg13g2_a21oi_1 _5149_ (.A1(_0805_),
    .A2(_0808_),
    .Y(_0809_),
    .B1(_0618_));
 sg13g2_o21ai_1 _5150_ (.B1(_0536_),
    .Y(_0810_),
    .A1(_0539_),
    .A2(_0809_));
 sg13g2_xnor2_1 _5151_ (.Y(_0811_),
    .A(_0494_),
    .B(_0810_));
 sg13g2_xnor2_1 _5152_ (.Y(_0812_),
    .A(_0538_),
    .B(_0809_));
 sg13g2_nand2_1 _5153_ (.Y(_0813_),
    .A(_3582_),
    .B(_0812_));
 sg13g2_o21ai_1 _5154_ (.B1(_0813_),
    .Y(_0814_),
    .A1(_3582_),
    .A2(_0811_));
 sg13g2_nor2_2 _5155_ (.A(_2416_),
    .B(_3096_),
    .Y(_0815_));
 sg13g2_nand2_2 _5156_ (.Y(_0816_),
    .A(net869),
    .B(net797));
 sg13g2_a21oi_1 _5157_ (.A1(_0805_),
    .A2(_0807_),
    .Y(_0817_),
    .B1(_0616_));
 sg13g2_xor2_1 _5158_ (.B(_0817_),
    .A(_0806_),
    .X(_0818_));
 sg13g2_xnor2_1 _5159_ (.Y(_0819_),
    .A(_0805_),
    .B(_0807_));
 sg13g2_nor2_1 _5160_ (.A(net809),
    .B(_0819_),
    .Y(_0820_));
 sg13g2_a21oi_2 _5161_ (.B1(_0820_),
    .Y(_0821_),
    .A2(_0818_),
    .A1(net808));
 sg13g2_o21ai_1 _5162_ (.B1(_0816_),
    .Y(_0822_),
    .A1(net790),
    .A2(_0821_));
 sg13g2_a21oi_1 _5163_ (.A1(net789),
    .A2(_0814_),
    .Y(_0823_),
    .B1(_0822_));
 sg13g2_a22oi_1 _5164_ (.Y(_0824_),
    .B1(_0463_),
    .B2(_0460_),
    .A2(_0461_),
    .A1(_0435_));
 sg13g2_nor2_1 _5165_ (.A(_0282_),
    .B(_0380_),
    .Y(_0825_));
 sg13g2_nor2_1 _5166_ (.A(_0282_),
    .B(_0375_),
    .Y(_0826_));
 sg13g2_nand2b_1 _5167_ (.Y(_0827_),
    .B(_0825_),
    .A_N(_0454_));
 sg13g2_xor2_1 _5168_ (.B(_0825_),
    .A(_0454_),
    .X(_0828_));
 sg13g2_nor2_1 _5169_ (.A(_0824_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_xor2_1 _5170_ (.B(_0828_),
    .A(_0824_),
    .X(_0830_));
 sg13g2_a21oi_1 _5171_ (.A1(_0455_),
    .A2(_0830_),
    .Y(_0831_),
    .B1(_0829_));
 sg13g2_a21oi_2 _5172_ (.B1(_0482_),
    .Y(_0832_),
    .A2(_0483_),
    .A1(_0464_));
 sg13g2_nand2_1 _5173_ (.Y(_0833_),
    .A(net716),
    .B(net758));
 sg13g2_nand2_1 _5174_ (.Y(_0834_),
    .A(net786),
    .B(net715));
 sg13g2_nand3_1 _5175_ (.B(net715),
    .C(_0461_),
    .A(net786),
    .Y(_0835_));
 sg13g2_xor2_1 _5176_ (.B(_0834_),
    .A(_0461_),
    .X(_0836_));
 sg13g2_xor2_1 _5177_ (.B(_0836_),
    .A(_0833_),
    .X(_0837_));
 sg13g2_a21oi_1 _5178_ (.A1(_0467_),
    .A2(_0480_),
    .Y(_0838_),
    .B1(_0479_));
 sg13g2_nand2_1 _5179_ (.Y(_0839_),
    .A(net788),
    .B(net714));
 sg13g2_nor4_2 _5180_ (.A(\r1[14] ),
    .B(net843),
    .C(_0304_),
    .Y(_0840_),
    .D(_0409_));
 sg13g2_xnor2_1 _5181_ (.Y(_0841_),
    .A(_0036_),
    .B(_0840_));
 sg13g2_nor2_1 _5182_ (.A(\r2[16] ),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_xor2_1 _5183_ (.B(_0841_),
    .A(\r2[16] ),
    .X(_0843_));
 sg13g2_nor2_1 _5184_ (.A(\r2[15] ),
    .B(_0470_),
    .Y(_0844_));
 sg13g2_nor2_1 _5185_ (.A(_0843_),
    .B(_0844_),
    .Y(_0845_));
 sg13g2_or2_2 _5186_ (.X(_0846_),
    .B(_0844_),
    .A(_0843_));
 sg13g2_xnor2_1 _5187_ (.Y(_0847_),
    .A(_0843_),
    .B(_0844_));
 sg13g2_nor2_1 _5188_ (.A(_0417_),
    .B(_0473_),
    .Y(_0848_));
 sg13g2_o21ai_1 _5189_ (.B1(_0848_),
    .Y(_0849_),
    .A1(_0419_),
    .A2(_0422_));
 sg13g2_a21oi_1 _5190_ (.A1(_0414_),
    .A2(_0474_),
    .Y(_0850_),
    .B1(_0472_));
 sg13g2_a21o_2 _5191_ (.A2(_0850_),
    .A1(_0849_),
    .B1(_0847_),
    .X(_0851_));
 sg13g2_nand3_1 _5192_ (.B(_0849_),
    .C(_0850_),
    .A(_0847_),
    .Y(_0852_));
 sg13g2_nand2_2 _5193_ (.Y(_0853_),
    .A(_0851_),
    .B(_0852_));
 sg13g2_and3_1 _5194_ (.X(_0854_),
    .A(net814),
    .B(_0851_),
    .C(_0852_));
 sg13g2_o21ai_1 _5195_ (.B1(_0278_),
    .Y(_0855_),
    .A1(_0475_),
    .A2(_0476_));
 sg13g2_nand3_1 _5196_ (.B(net713),
    .C(_0854_),
    .A(net804),
    .Y(_0856_));
 sg13g2_xor2_1 _5197_ (.B(_0855_),
    .A(_0854_),
    .X(_0857_));
 sg13g2_xor2_1 _5198_ (.B(_0857_),
    .A(_0839_),
    .X(_0858_));
 sg13g2_nor2b_1 _5199_ (.A(_0838_),
    .B_N(_0858_),
    .Y(_0859_));
 sg13g2_xnor2_1 _5200_ (.Y(_0860_),
    .A(_0838_),
    .B(_0858_));
 sg13g2_xnor2_1 _5201_ (.Y(_0861_),
    .A(_0837_),
    .B(_0860_));
 sg13g2_xnor2_1 _5202_ (.Y(_0862_),
    .A(_0455_),
    .B(_0830_));
 sg13g2_xor2_1 _5203_ (.B(_0861_),
    .A(_0832_),
    .X(_0863_));
 sg13g2_nand2b_1 _5204_ (.Y(_0864_),
    .B(_0863_),
    .A_N(_0862_));
 sg13g2_o21ai_1 _5205_ (.B1(_0864_),
    .Y(_0865_),
    .A1(_0832_),
    .A2(_0861_));
 sg13g2_o21ai_1 _5206_ (.B1(_0835_),
    .Y(_0866_),
    .A1(_0833_),
    .A2(_0836_));
 sg13g2_nand3_1 _5207_ (.B(net746),
    .C(_0826_),
    .A(net716),
    .Y(_0867_));
 sg13g2_a21o_1 _5208_ (.A2(net746),
    .A1(net716),
    .B1(_0826_),
    .X(_0868_));
 sg13g2_nand2_1 _5209_ (.Y(_0869_),
    .A(_0867_),
    .B(_0868_));
 sg13g2_nand2b_1 _5210_ (.Y(_0870_),
    .B(_0866_),
    .A_N(_0869_));
 sg13g2_xor2_1 _5211_ (.B(_0869_),
    .A(_0866_),
    .X(_0871_));
 sg13g2_xor2_1 _5212_ (.B(_0871_),
    .A(_0827_),
    .X(_0872_));
 sg13g2_a21oi_1 _5213_ (.A1(_0837_),
    .A2(_0860_),
    .Y(_0873_),
    .B1(_0859_));
 sg13g2_and2_1 _5214_ (.A(net719),
    .B(net758),
    .X(_0874_));
 sg13g2_nand2_1 _5215_ (.Y(_0875_),
    .A(net772),
    .B(net714));
 sg13g2_nand2_1 _5216_ (.Y(_0876_),
    .A(net786),
    .B(net714));
 sg13g2_nor2_1 _5217_ (.A(_0834_),
    .B(_0875_),
    .Y(_0877_));
 sg13g2_a22oi_1 _5218_ (.Y(_0878_),
    .B1(net714),
    .B2(net786),
    .A2(net715),
    .A1(net772));
 sg13g2_nor2_1 _5219_ (.A(_0877_),
    .B(_0878_),
    .Y(_0879_));
 sg13g2_xnor2_1 _5220_ (.Y(_0880_),
    .A(_0874_),
    .B(_0879_));
 sg13g2_o21ai_1 _5221_ (.B1(_0856_),
    .Y(_0881_),
    .A1(_0839_),
    .A2(_0857_));
 sg13g2_nand2_1 _5222_ (.Y(_0882_),
    .A(net788),
    .B(net713));
 sg13g2_nor2b_1 _5223_ (.A(\r1[15] ),
    .B_N(_0840_),
    .Y(_0883_));
 sg13g2_xnor2_1 _5224_ (.Y(_0884_),
    .A(_0014_),
    .B(_0883_));
 sg13g2_xor2_1 _5225_ (.B(_0884_),
    .A(_0013_),
    .X(_0885_));
 sg13g2_nor2b_1 _5226_ (.A(_0842_),
    .B_N(_0885_),
    .Y(_0886_));
 sg13g2_xnor2_1 _5227_ (.Y(_0887_),
    .A(_0842_),
    .B(_0885_));
 sg13g2_nand3_1 _5228_ (.B(_0851_),
    .C(_0887_),
    .A(_0846_),
    .Y(_0888_));
 sg13g2_a21o_1 _5229_ (.A2(_0851_),
    .A1(_0846_),
    .B1(_0887_),
    .X(_0889_));
 sg13g2_nand2_2 _5230_ (.Y(_0890_),
    .A(_0888_),
    .B(_0889_));
 sg13g2_and2_1 _5231_ (.A(_0888_),
    .B(_0889_),
    .X(_0891_));
 sg13g2_a21oi_1 _5232_ (.A1(_0888_),
    .A2(_0889_),
    .Y(_0892_),
    .B1(net803));
 sg13g2_a21oi_1 _5233_ (.A1(_0888_),
    .A2(_0889_),
    .Y(_0893_),
    .B1(net891));
 sg13g2_nor2_1 _5234_ (.A(net803),
    .B(_0853_),
    .Y(_0894_));
 sg13g2_nand2_1 _5235_ (.Y(_0895_),
    .A(_0854_),
    .B(_0892_));
 sg13g2_xnor2_1 _5236_ (.Y(_0896_),
    .A(_0893_),
    .B(_0894_));
 sg13g2_xor2_1 _5237_ (.B(_0896_),
    .A(_0882_),
    .X(_0897_));
 sg13g2_nand2_1 _5238_ (.Y(_0898_),
    .A(_0881_),
    .B(_0897_));
 sg13g2_xnor2_1 _5239_ (.Y(_0899_),
    .A(_0881_),
    .B(_0897_));
 sg13g2_xor2_1 _5240_ (.B(_0899_),
    .A(_0880_),
    .X(_0900_));
 sg13g2_nor2b_1 _5241_ (.A(_0873_),
    .B_N(_0900_),
    .Y(_0901_));
 sg13g2_xnor2_1 _5242_ (.Y(_0902_),
    .A(_0873_),
    .B(_0900_));
 sg13g2_xnor2_1 _5243_ (.Y(_0903_),
    .A(_0872_),
    .B(_0902_));
 sg13g2_nor2b_1 _5244_ (.A(_0903_),
    .B_N(_0865_),
    .Y(_0904_));
 sg13g2_xor2_1 _5245_ (.B(_0903_),
    .A(_0865_),
    .X(_0905_));
 sg13g2_nor2_1 _5246_ (.A(_0831_),
    .B(_0905_),
    .Y(_0906_));
 sg13g2_xor2_1 _5247_ (.B(_0905_),
    .A(_0831_),
    .X(_0907_));
 sg13g2_o21ai_1 _5248_ (.B1(_0485_),
    .Y(_0908_),
    .A1(_0458_),
    .A2(_0486_));
 sg13g2_xnor2_1 _5249_ (.Y(_0909_),
    .A(_0862_),
    .B(_0863_));
 sg13g2_nor2_1 _5250_ (.A(_0399_),
    .B(_0457_),
    .Y(_0910_));
 sg13g2_a21oi_1 _5251_ (.A1(_0452_),
    .A2(_0456_),
    .Y(_0911_),
    .B1(_0910_));
 sg13g2_xnor2_1 _5252_ (.Y(_0912_),
    .A(_0908_),
    .B(_0909_));
 sg13g2_nor2_1 _5253_ (.A(_0911_),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_a21oi_2 _5254_ (.B1(_0913_),
    .Y(_0914_),
    .A2(_0909_),
    .A1(_0908_));
 sg13g2_nand2b_1 _5255_ (.Y(_0915_),
    .B(_0914_),
    .A_N(_0907_));
 sg13g2_nor2b_1 _5256_ (.A(_0914_),
    .B_N(_0907_),
    .Y(_0916_));
 sg13g2_xnor2_1 _5257_ (.Y(_0917_),
    .A(_0907_),
    .B(_0914_));
 sg13g2_xor2_1 _5258_ (.B(_0912_),
    .A(_0911_),
    .X(_0918_));
 sg13g2_a21o_1 _5259_ (.A2(_0490_),
    .A1(_0450_),
    .B1(_0489_),
    .X(_0919_));
 sg13g2_and2_1 _5260_ (.A(_0918_),
    .B(_0919_),
    .X(_0920_));
 sg13g2_a21o_1 _5261_ (.A2(_0491_),
    .A1(_0449_),
    .B1(_0535_),
    .X(_0921_));
 sg13g2_a221oi_1 _5262_ (.B2(_0493_),
    .C1(_0618_),
    .B1(_0921_),
    .A1(_0808_),
    .Y(_0922_),
    .A2(_0805_));
 sg13g2_a21oi_1 _5263_ (.A1(_0449_),
    .A2(_0491_),
    .Y(_0923_),
    .B1(_0537_));
 sg13g2_nor2_1 _5264_ (.A(_0492_),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_nor2b_1 _5265_ (.A(_0922_),
    .B_N(_0924_),
    .Y(_0925_));
 sg13g2_xor2_1 _5266_ (.B(_0919_),
    .A(_0918_),
    .X(_0926_));
 sg13g2_a21oi_1 _5267_ (.A1(_0925_),
    .A2(_0926_),
    .Y(_0927_),
    .B1(_0920_));
 sg13g2_xnor2_1 _5268_ (.Y(_0928_),
    .A(_0917_),
    .B(_0927_));
 sg13g2_xnor2_1 _5269_ (.Y(_0929_),
    .A(_0925_),
    .B(_0926_));
 sg13g2_nor2_1 _5270_ (.A(net808),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_a21oi_1 _5271_ (.A1(net808),
    .A2(_0928_),
    .Y(_0931_),
    .B1(_0930_));
 sg13g2_nand2_1 _5272_ (.Y(_0932_),
    .A(_3578_),
    .B(_0931_));
 sg13g2_a21oi_1 _5273_ (.A1(_0872_),
    .A2(_0902_),
    .Y(_0933_),
    .B1(_0901_));
 sg13g2_a21oi_1 _5274_ (.A1(_0874_),
    .A2(_0879_),
    .Y(_0934_),
    .B1(_0877_));
 sg13g2_a22oi_1 _5275_ (.Y(_0935_),
    .B1(net746),
    .B2(net719),
    .A2(net756),
    .A1(net716));
 sg13g2_nand2_1 _5276_ (.Y(_0936_),
    .A(net720),
    .B(net756));
 sg13g2_nand4_1 _5277_ (.B(net719),
    .C(net756),
    .A(net716),
    .Y(_0937_),
    .D(net746));
 sg13g2_inv_1 _5278_ (.Y(_0938_),
    .A(_0937_));
 sg13g2_nand2b_1 _5279_ (.Y(_0939_),
    .B(_0937_),
    .A_N(_0935_));
 sg13g2_nor2_1 _5280_ (.A(_0934_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_xor2_1 _5281_ (.B(_0939_),
    .A(_0934_),
    .X(_0941_));
 sg13g2_nor2b_1 _5282_ (.A(_0867_),
    .B_N(_0941_),
    .Y(_0942_));
 sg13g2_xor2_1 _5283_ (.B(_0941_),
    .A(_0867_),
    .X(_0943_));
 sg13g2_o21ai_1 _5284_ (.B1(_0898_),
    .Y(_0944_),
    .A1(_0880_),
    .A2(_0899_));
 sg13g2_nand2_1 _5285_ (.Y(_0945_),
    .A(net758),
    .B(net715));
 sg13g2_nand2_1 _5286_ (.Y(_0946_),
    .A(net772),
    .B(net713));
 sg13g2_nand2_1 _5287_ (.Y(_0947_),
    .A(net785),
    .B(net713));
 sg13g2_nor2_1 _5288_ (.A(_0876_),
    .B(_0946_),
    .Y(_0948_));
 sg13g2_xor2_1 _5289_ (.B(_0947_),
    .A(_0875_),
    .X(_0949_));
 sg13g2_nor2b_1 _5290_ (.A(_0945_),
    .B_N(_0949_),
    .Y(_0950_));
 sg13g2_xor2_1 _5291_ (.B(_0949_),
    .A(_0945_),
    .X(_0951_));
 sg13g2_o21ai_1 _5292_ (.B1(_0895_),
    .Y(_0952_),
    .A1(_0882_),
    .A2(_0896_));
 sg13g2_nor2_1 _5293_ (.A(_0292_),
    .B(_0853_),
    .Y(_0953_));
 sg13g2_nand2b_1 _5294_ (.Y(_0954_),
    .B(_0887_),
    .A_N(_0847_));
 sg13g2_a21oi_1 _5295_ (.A1(_0849_),
    .A2(_0850_),
    .Y(_0955_),
    .B1(_0954_));
 sg13g2_a21oi_1 _5296_ (.A1(_0845_),
    .A2(_0887_),
    .Y(_0956_),
    .B1(_0886_));
 sg13g2_inv_1 _5297_ (.Y(_0957_),
    .A(_0956_));
 sg13g2_nor2_1 _5298_ (.A(\r2[17] ),
    .B(_0884_),
    .Y(_0958_));
 sg13g2_and2_1 _5299_ (.A(_2979_),
    .B(_0883_),
    .X(_0959_));
 sg13g2_and2_1 _5300_ (.A(_2998_),
    .B(_0959_),
    .X(_0960_));
 sg13g2_xnor2_1 _5301_ (.Y(_0961_),
    .A(_0016_),
    .B(_0959_));
 sg13g2_xnor2_1 _5302_ (.Y(_0962_),
    .A(_0015_),
    .B(_0961_));
 sg13g2_or2_2 _5303_ (.X(_0963_),
    .B(_0962_),
    .A(_0958_));
 sg13g2_xor2_1 _5304_ (.B(_0962_),
    .A(_0958_),
    .X(_0964_));
 sg13g2_o21ai_1 _5305_ (.B1(_0964_),
    .Y(_0965_),
    .A1(_0957_),
    .A2(_0955_));
 sg13g2_or3_2 _5306_ (.A(_0955_),
    .B(_0957_),
    .C(_0964_),
    .X(_0966_));
 sg13g2_nand2_2 _5307_ (.Y(_0967_),
    .A(net151),
    .B(_0966_));
 sg13g2_nor2_1 _5308_ (.A(net803),
    .B(_0967_),
    .Y(_0968_));
 sg13g2_nand3_1 _5309_ (.B(net151),
    .C(_0966_),
    .A(net814),
    .Y(_0969_));
 sg13g2_xnor2_1 _5310_ (.Y(_0970_),
    .A(_0892_),
    .B(_0969_));
 sg13g2_xnor2_1 _5311_ (.Y(_0971_),
    .A(_0953_),
    .B(_0970_));
 sg13g2_nor2b_1 _5312_ (.A(_0971_),
    .B_N(_0952_),
    .Y(_0972_));
 sg13g2_xor2_1 _5313_ (.B(_0971_),
    .A(_0952_),
    .X(_0973_));
 sg13g2_nor2_1 _5314_ (.A(_0951_),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_xor2_1 _5315_ (.B(_0973_),
    .A(_0951_),
    .X(_0975_));
 sg13g2_nand2_1 _5316_ (.Y(_0976_),
    .A(_0944_),
    .B(_0975_));
 sg13g2_xnor2_1 _5317_ (.Y(_0977_),
    .A(_0944_),
    .B(_0975_));
 sg13g2_xnor2_1 _5318_ (.Y(_0978_),
    .A(_0943_),
    .B(_0977_));
 sg13g2_nor2_1 _5319_ (.A(_0933_),
    .B(_0978_),
    .Y(_0979_));
 sg13g2_o21ai_1 _5320_ (.B1(_0870_),
    .Y(_0980_),
    .A1(_0827_),
    .A2(_0871_));
 sg13g2_xor2_1 _5321_ (.B(_0978_),
    .A(_0933_),
    .X(_0981_));
 sg13g2_a21o_1 _5322_ (.A2(_0981_),
    .A1(_0980_),
    .B1(_0979_),
    .X(_0982_));
 sg13g2_inv_1 _5323_ (.Y(_0983_),
    .A(_0982_));
 sg13g2_nor2_2 _5324_ (.A(_0940_),
    .B(_0942_),
    .Y(_0984_));
 sg13g2_o21ai_1 _5325_ (.B1(_0976_),
    .Y(_0985_),
    .A1(_0943_),
    .A2(_0977_));
 sg13g2_nor2_1 _5326_ (.A(_0948_),
    .B(_0950_),
    .Y(_0986_));
 sg13g2_nand2_1 _5327_ (.Y(_0987_),
    .A(net715),
    .B(net746));
 sg13g2_or2_1 _5328_ (.X(_0988_),
    .B(_0987_),
    .A(_0936_));
 sg13g2_xnor2_1 _5329_ (.Y(_0989_),
    .A(_0936_),
    .B(_0987_));
 sg13g2_nor2_1 _5330_ (.A(_0986_),
    .B(_0989_),
    .Y(_0990_));
 sg13g2_xor2_1 _5331_ (.B(_0989_),
    .A(_0986_),
    .X(_0991_));
 sg13g2_xnor2_1 _5332_ (.Y(_0992_),
    .A(_0937_),
    .B(_0991_));
 sg13g2_nor2_1 _5333_ (.A(_0972_),
    .B(_0974_),
    .Y(_0993_));
 sg13g2_nand2_1 _5334_ (.Y(_0994_),
    .A(net758),
    .B(net714));
 sg13g2_nor2_1 _5335_ (.A(_0331_),
    .B(_0853_),
    .Y(_0995_));
 sg13g2_nand2b_1 _5336_ (.Y(_0996_),
    .B(_0995_),
    .A_N(_0947_));
 sg13g2_o21ai_1 _5337_ (.B1(_0946_),
    .Y(_0997_),
    .A1(_0334_),
    .A2(_0853_));
 sg13g2_and2_1 _5338_ (.A(_0996_),
    .B(_0997_),
    .X(_0998_));
 sg13g2_nand2b_1 _5339_ (.Y(_0999_),
    .B(_0998_),
    .A_N(_0994_));
 sg13g2_xnor2_1 _5340_ (.Y(_1000_),
    .A(_0994_),
    .B(_0998_));
 sg13g2_a22oi_1 _5341_ (.Y(_1001_),
    .B1(_0970_),
    .B2(_0953_),
    .A2(_0968_),
    .A1(_0893_));
 sg13g2_nand2_1 _5342_ (.Y(_1002_),
    .A(net788),
    .B(_0890_));
 sg13g2_inv_1 _5343_ (.Y(_1003_),
    .A(_1002_));
 sg13g2_o21ai_1 _5344_ (.B1(\r2[18] ),
    .Y(_1004_),
    .A1(_2998_),
    .A2(_0959_));
 sg13g2_o21ai_1 _5345_ (.B1(_1004_),
    .Y(_1005_),
    .A1(\r2[18] ),
    .A2(_0960_));
 sg13g2_xor2_1 _5346_ (.B(_1005_),
    .A(_0015_),
    .X(_1006_));
 sg13g2_a21o_1 _5347_ (.A2(net151),
    .A1(_0963_),
    .B1(_1006_),
    .X(_1007_));
 sg13g2_nand3_1 _5348_ (.B(net151),
    .C(_1006_),
    .A(_0963_),
    .Y(_1008_));
 sg13g2_nand2_1 _5349_ (.Y(_1009_),
    .A(_1007_),
    .B(_1008_));
 sg13g2_nand3_1 _5350_ (.B(_1007_),
    .C(_1008_),
    .A(net804),
    .Y(_1010_));
 sg13g2_and3_1 _5351_ (.X(_1011_),
    .A(net814),
    .B(_1007_),
    .C(_1008_));
 sg13g2_nor2_1 _5352_ (.A(_0969_),
    .B(_1010_),
    .Y(_1012_));
 sg13g2_xor2_1 _5353_ (.B(_1011_),
    .A(_0968_),
    .X(_1013_));
 sg13g2_xnor2_1 _5354_ (.Y(_1014_),
    .A(_1003_),
    .B(_1013_));
 sg13g2_nor2_1 _5355_ (.A(_1001_),
    .B(_1014_),
    .Y(_1015_));
 sg13g2_xor2_1 _5356_ (.B(_1014_),
    .A(_1001_),
    .X(_1016_));
 sg13g2_xnor2_1 _5357_ (.Y(_1017_),
    .A(_1000_),
    .B(_1016_));
 sg13g2_nor2_1 _5358_ (.A(_0993_),
    .B(_1017_),
    .Y(_1018_));
 sg13g2_xor2_1 _5359_ (.B(_1017_),
    .A(_0993_),
    .X(_1019_));
 sg13g2_xnor2_1 _5360_ (.Y(_1020_),
    .A(_0992_),
    .B(_1019_));
 sg13g2_nand2b_1 _5361_ (.Y(_1021_),
    .B(_0985_),
    .A_N(_1020_));
 sg13g2_xor2_1 _5362_ (.B(_1020_),
    .A(_0985_),
    .X(_1022_));
 sg13g2_xor2_1 _5363_ (.B(_1022_),
    .A(_0984_),
    .X(_1023_));
 sg13g2_xnor2_1 _5364_ (.Y(_1024_),
    .A(_0984_),
    .B(_1022_));
 sg13g2_nor2_1 _5365_ (.A(_0982_),
    .B(_1023_),
    .Y(_1025_));
 sg13g2_nand2_1 _5366_ (.Y(_1026_),
    .A(_0982_),
    .B(_1023_));
 sg13g2_nor2b_1 _5367_ (.A(_1025_),
    .B_N(_1026_),
    .Y(_1027_));
 sg13g2_xor2_1 _5368_ (.B(_0981_),
    .A(_0980_),
    .X(_1028_));
 sg13g2_o21ai_1 _5369_ (.B1(_1028_),
    .Y(_1029_),
    .A1(_0904_),
    .A2(_0906_));
 sg13g2_nor3_1 _5370_ (.A(_0904_),
    .B(_0906_),
    .C(_1028_),
    .Y(_1030_));
 sg13g2_inv_1 _5371_ (.Y(_1031_),
    .A(_1030_));
 sg13g2_nand2_1 _5372_ (.Y(_1032_),
    .A(_1029_),
    .B(_1031_));
 sg13g2_and2_1 _5373_ (.A(_0917_),
    .B(_0926_),
    .X(_1033_));
 sg13g2_nand3b_1 _5374_ (.B(_0924_),
    .C(_1033_),
    .Y(_1034_),
    .A_N(_0922_));
 sg13g2_a21oi_1 _5375_ (.A1(_0915_),
    .A2(_0920_),
    .Y(_1035_),
    .B1(_0916_));
 sg13g2_and2_1 _5376_ (.A(_1034_),
    .B(_1035_),
    .X(_1036_));
 sg13g2_o21ai_1 _5377_ (.B1(_1029_),
    .Y(_1037_),
    .A1(_1032_),
    .A2(_1036_));
 sg13g2_xor2_1 _5378_ (.B(_1037_),
    .A(_1027_),
    .X(_1038_));
 sg13g2_xor2_1 _5379_ (.B(_1036_),
    .A(_1032_),
    .X(_1039_));
 sg13g2_mux2_1 _5380_ (.A0(_1038_),
    .A1(_1039_),
    .S(net807),
    .X(_1040_));
 sg13g2_o21ai_1 _5381_ (.B1(_0932_),
    .Y(_1041_),
    .A1(_3578_),
    .A2(_1040_));
 sg13g2_a21oi_2 _5382_ (.B1(_0823_),
    .Y(_1042_),
    .A2(_1041_),
    .A1(_0815_));
 sg13g2_a21o_2 _5383_ (.A2(_1041_),
    .A1(net781),
    .B1(_0823_),
    .X(_1043_));
 sg13g2_mux2_1 _5384_ (.A0(_0812_),
    .A1(_0818_),
    .S(net807),
    .X(_1044_));
 sg13g2_xnor2_1 _5385_ (.Y(_1045_),
    .A(_0802_),
    .B(_0803_));
 sg13g2_nand2_1 _5386_ (.Y(_1046_),
    .A(net807),
    .B(_1045_));
 sg13g2_o21ai_1 _5387_ (.B1(_1046_),
    .Y(_1047_),
    .A1(net807),
    .A2(_0819_));
 sg13g2_mux2_1 _5388_ (.A0(_0811_),
    .A1(_0929_),
    .S(net808),
    .X(_1048_));
 sg13g2_mux2_1 _5389_ (.A0(_0928_),
    .A1(_1039_),
    .S(_3581_),
    .X(_1049_));
 sg13g2_nor2_1 _5390_ (.A(net790),
    .B(_1048_),
    .Y(_1050_));
 sg13g2_a21o_1 _5391_ (.A2(_1049_),
    .A1(net789),
    .B1(_1050_),
    .X(_1051_));
 sg13g2_nor2_1 _5392_ (.A(net789),
    .B(_1047_),
    .Y(_1052_));
 sg13g2_o21ai_1 _5393_ (.B1(_0816_),
    .Y(_1053_),
    .A1(_3578_),
    .A2(_1044_));
 sg13g2_nor2_1 _5394_ (.A(_1052_),
    .B(_1053_),
    .Y(_1054_));
 sg13g2_a21oi_2 _5395_ (.B1(_1054_),
    .Y(_1055_),
    .A2(_1051_),
    .A1(net781));
 sg13g2_or2_1 _5396_ (.X(_1056_),
    .B(_1055_),
    .A(_1043_));
 sg13g2_a21o_1 _5397_ (.A2(_1024_),
    .A1(_0983_),
    .B1(_1029_),
    .X(_1057_));
 sg13g2_and3_1 _5398_ (.X(_1058_),
    .A(_1026_),
    .B(_1035_),
    .C(_1057_));
 sg13g2_nand2_1 _5399_ (.Y(_1059_),
    .A(_1034_),
    .B(_1058_));
 sg13g2_nand2b_1 _5400_ (.Y(_1060_),
    .B(_1031_),
    .A_N(_1025_));
 sg13g2_nand2_1 _5401_ (.Y(_1061_),
    .A(_1026_),
    .B(_1060_));
 sg13g2_a21oi_1 _5402_ (.A1(_0938_),
    .A2(_0991_),
    .Y(_1062_),
    .B1(_0990_));
 sg13g2_a21oi_1 _5403_ (.A1(_0992_),
    .A2(_1019_),
    .Y(_1063_),
    .B1(_1018_));
 sg13g2_nand2_1 _5404_ (.Y(_1064_),
    .A(_0996_),
    .B(_0999_));
 sg13g2_a22oi_1 _5405_ (.Y(_1065_),
    .B1(_0379_),
    .B2(_0427_),
    .A2(net756),
    .A1(net715));
 sg13g2_nand2_1 _5406_ (.Y(_1066_),
    .A(net756),
    .B(_0427_));
 sg13g2_nand4_1 _5407_ (.B(net756),
    .C(net746),
    .A(_0362_),
    .Y(_1067_),
    .D(_0427_));
 sg13g2_nand2b_1 _5408_ (.Y(_1068_),
    .B(_1067_),
    .A_N(_1065_));
 sg13g2_nand2b_1 _5409_ (.Y(_1069_),
    .B(_1064_),
    .A_N(_1068_));
 sg13g2_xor2_1 _5410_ (.B(_1068_),
    .A(_1064_),
    .X(_1070_));
 sg13g2_xor2_1 _5411_ (.B(_1070_),
    .A(_0988_),
    .X(_1071_));
 sg13g2_a21oi_1 _5412_ (.A1(_1000_),
    .A2(_1016_),
    .Y(_1072_),
    .B1(_1015_));
 sg13g2_nand2_1 _5413_ (.Y(_1073_),
    .A(net758),
    .B(_0477_));
 sg13g2_nand2_1 _5414_ (.Y(_1074_),
    .A(net772),
    .B(_0890_));
 sg13g2_nor2_1 _5415_ (.A(_0334_),
    .B(_0891_),
    .Y(_1075_));
 sg13g2_nand2_1 _5416_ (.Y(_1076_),
    .A(_0995_),
    .B(_1075_));
 sg13g2_xnor2_1 _5417_ (.Y(_1077_),
    .A(_0995_),
    .B(_1075_));
 sg13g2_xor2_1 _5418_ (.B(_1077_),
    .A(_1073_),
    .X(_1078_));
 sg13g2_a21oi_1 _5419_ (.A1(_1003_),
    .A2(_1013_),
    .Y(_1079_),
    .B1(_1012_));
 sg13g2_a21oi_1 _5420_ (.A1(net891),
    .A2(net803),
    .Y(_1080_),
    .B1(_1009_));
 sg13g2_mux2_1 _5421_ (.A0(net891),
    .A1(_1011_),
    .S(_1010_),
    .X(_1081_));
 sg13g2_nor2_1 _5422_ (.A(_0292_),
    .B(_0967_),
    .Y(_1082_));
 sg13g2_xnor2_1 _5423_ (.Y(_1083_),
    .A(_1081_),
    .B(_1082_));
 sg13g2_nor2_1 _5424_ (.A(_1079_),
    .B(_1083_),
    .Y(_1084_));
 sg13g2_xor2_1 _5425_ (.B(_1083_),
    .A(_1079_),
    .X(_1085_));
 sg13g2_xnor2_1 _5426_ (.Y(_1086_),
    .A(_1078_),
    .B(_1085_));
 sg13g2_nor2_1 _5427_ (.A(_1072_),
    .B(_1086_),
    .Y(_1087_));
 sg13g2_xor2_1 _5428_ (.B(_1086_),
    .A(_1072_),
    .X(_1088_));
 sg13g2_xnor2_1 _5429_ (.Y(_1089_),
    .A(_1071_),
    .B(_1088_));
 sg13g2_nor2_1 _5430_ (.A(_1063_),
    .B(_1089_),
    .Y(_1090_));
 sg13g2_xor2_1 _5431_ (.B(_1089_),
    .A(_1063_),
    .X(_1091_));
 sg13g2_nand2b_1 _5432_ (.Y(_1092_),
    .B(_1091_),
    .A_N(_1062_));
 sg13g2_xnor2_1 _5433_ (.Y(_1093_),
    .A(_1062_),
    .B(_1091_));
 sg13g2_o21ai_1 _5434_ (.B1(_1021_),
    .Y(_1094_),
    .A1(_0984_),
    .A2(_1022_));
 sg13g2_and2_1 _5435_ (.A(_1093_),
    .B(_1094_),
    .X(_1095_));
 sg13g2_inv_1 _5436_ (.Y(_1096_),
    .A(_1095_));
 sg13g2_or2_1 _5437_ (.X(_1097_),
    .B(_1094_),
    .A(_1093_));
 sg13g2_nand2b_1 _5438_ (.Y(_1098_),
    .B(_1097_),
    .A_N(_1095_));
 sg13g2_a221oi_1 _5439_ (.B2(_1026_),
    .C1(_1098_),
    .B1(_1060_),
    .A1(_1058_),
    .Y(_1099_),
    .A2(_1034_));
 sg13g2_a22oi_1 _5440_ (.Y(_1100_),
    .B1(_1096_),
    .B2(_1097_),
    .A2(_1061_),
    .A1(_1059_));
 sg13g2_nor2_1 _5441_ (.A(_1099_),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_nor2b_1 _5442_ (.A(_1090_),
    .B_N(_1092_),
    .Y(_1102_));
 sg13g2_o21ai_1 _5443_ (.B1(_1069_),
    .Y(_1103_),
    .A1(_0988_),
    .A2(_1070_));
 sg13g2_a21oi_1 _5444_ (.A1(_1071_),
    .A2(_1088_),
    .Y(_1104_),
    .B1(_1087_));
 sg13g2_o21ai_1 _5445_ (.B1(_1076_),
    .Y(_1105_),
    .A1(_1073_),
    .A2(_1077_));
 sg13g2_nand2_2 _5446_ (.Y(_1106_),
    .A(net746),
    .B(net713));
 sg13g2_nand2_1 _5447_ (.Y(_1107_),
    .A(net756),
    .B(net713));
 sg13g2_or2_1 _5448_ (.X(_1108_),
    .B(_1106_),
    .A(_1066_));
 sg13g2_xor2_1 _5449_ (.B(_1106_),
    .A(_1066_),
    .X(_1109_));
 sg13g2_xnor2_1 _5450_ (.Y(_1110_),
    .A(_1105_),
    .B(_1109_));
 sg13g2_xnor2_1 _5451_ (.Y(_1111_),
    .A(_1067_),
    .B(_1110_));
 sg13g2_a21oi_2 _5452_ (.B1(_1084_),
    .Y(_1112_),
    .A2(_1085_),
    .A1(_1078_));
 sg13g2_nor2_1 _5453_ (.A(_0325_),
    .B(_0853_),
    .Y(_1113_));
 sg13g2_nor2_2 _5454_ (.A(_0331_),
    .B(_0967_),
    .Y(_1114_));
 sg13g2_nand2_1 _5455_ (.Y(_1115_),
    .A(_1075_),
    .B(_1114_));
 sg13g2_o21ai_1 _5456_ (.B1(_1074_),
    .Y(_1116_),
    .A1(net784),
    .A2(_0967_));
 sg13g2_and2_1 _5457_ (.A(_1115_),
    .B(_1116_),
    .X(_1117_));
 sg13g2_nand2_1 _5458_ (.Y(_1118_),
    .A(_1113_),
    .B(_1117_));
 sg13g2_xnor2_1 _5459_ (.Y(_1119_),
    .A(_1113_),
    .B(_1117_));
 sg13g2_inv_1 _5460_ (.Y(_1120_),
    .A(_1119_));
 sg13g2_nor3_2 _5461_ (.A(\center_x[1] ),
    .B(net891),
    .C(_1010_),
    .Y(_1121_));
 sg13g2_nand3_1 _5462_ (.B(_1007_),
    .C(_1008_),
    .A(net788),
    .Y(_1122_));
 sg13g2_a22oi_1 _5463_ (.Y(_1123_),
    .B1(_1081_),
    .B2(_1082_),
    .A2(_1011_),
    .A1(net804));
 sg13g2_xor2_1 _5464_ (.B(_1122_),
    .A(_1081_),
    .X(_1124_));
 sg13g2_a21oi_2 _5465_ (.B1(_1121_),
    .Y(_1125_),
    .A2(_1124_),
    .A1(_1123_));
 sg13g2_xnor2_1 _5466_ (.Y(_1126_),
    .A(_1119_),
    .B(_1125_));
 sg13g2_nand2b_1 _5467_ (.Y(_1127_),
    .B(_1126_),
    .A_N(_1112_));
 sg13g2_xnor2_1 _5468_ (.Y(_1128_),
    .A(_1112_),
    .B(_1126_));
 sg13g2_nand2b_1 _5469_ (.Y(_1129_),
    .B(_1128_),
    .A_N(_1111_));
 sg13g2_xnor2_1 _5470_ (.Y(_1130_),
    .A(_1111_),
    .B(_1128_));
 sg13g2_nor2b_1 _5471_ (.A(_1104_),
    .B_N(_1130_),
    .Y(_1131_));
 sg13g2_xnor2_1 _5472_ (.Y(_1132_),
    .A(_1104_),
    .B(_1130_));
 sg13g2_xnor2_1 _5473_ (.Y(_1133_),
    .A(_1103_),
    .B(_1132_));
 sg13g2_nand2_1 _5474_ (.Y(_1134_),
    .A(_1102_),
    .B(_1133_));
 sg13g2_xnor2_1 _5475_ (.Y(_1135_),
    .A(_1102_),
    .B(_1133_));
 sg13g2_nor2_1 _5476_ (.A(_1095_),
    .B(_1099_),
    .Y(_1136_));
 sg13g2_xnor2_1 _5477_ (.Y(_1137_),
    .A(_1135_),
    .B(_1136_));
 sg13g2_xor2_1 _5478_ (.B(_1136_),
    .A(_1135_),
    .X(_1138_));
 sg13g2_mux2_1 _5479_ (.A0(_1101_),
    .A1(_1138_),
    .S(net809),
    .X(_1139_));
 sg13g2_a221oi_1 _5480_ (.B2(net790),
    .C1(_0816_),
    .B1(_1139_),
    .A1(_2695_),
    .Y(_1140_),
    .A2(_1040_));
 sg13g2_nor2_1 _5481_ (.A(net789),
    .B(_0814_),
    .Y(_1141_));
 sg13g2_a21oi_1 _5482_ (.A1(net789),
    .A2(_0931_),
    .Y(_1142_),
    .B1(_1141_));
 sg13g2_nor2_1 _5483_ (.A(net781),
    .B(_1142_),
    .Y(_1143_));
 sg13g2_nor2_2 _5484_ (.A(_1140_),
    .B(_1143_),
    .Y(_1144_));
 sg13g2_or2_2 _5485_ (.X(_1145_),
    .B(_1143_),
    .A(_1140_));
 sg13g2_xnor2_1 _5486_ (.Y(_1146_),
    .A(_0800_),
    .B(_0801_));
 sg13g2_nand2_1 _5487_ (.Y(_1147_),
    .A(net790),
    .B(_1047_));
 sg13g2_xor2_1 _5488_ (.B(_0799_),
    .A(_0728_),
    .X(_1148_));
 sg13g2_o21ai_1 _5489_ (.B1(_3578_),
    .Y(_1149_),
    .A1(net808),
    .A2(_1148_));
 sg13g2_a21oi_1 _5490_ (.A1(net808),
    .A2(_1146_),
    .Y(_1150_),
    .B1(_1149_));
 sg13g2_nor2_1 _5491_ (.A(net789),
    .B(_1044_),
    .Y(_1151_));
 sg13g2_a21oi_1 _5492_ (.A1(net789),
    .A2(_1048_),
    .Y(_1152_),
    .B1(_1151_));
 sg13g2_a21o_1 _5493_ (.A2(_1048_),
    .A1(net789),
    .B1(_1151_),
    .X(_1153_));
 sg13g2_nor2_1 _5494_ (.A(net781),
    .B(_1150_),
    .Y(_1154_));
 sg13g2_nand2_1 _5495_ (.Y(_1155_),
    .A(_1147_),
    .B(_1154_));
 sg13g2_o21ai_1 _5496_ (.B1(_1155_),
    .Y(_1156_),
    .A1(_0816_),
    .A2(_1152_));
 sg13g2_a22oi_1 _5497_ (.Y(_1157_),
    .B1(_1154_),
    .B2(_1147_),
    .A2(_1153_),
    .A1(net781));
 sg13g2_nand2_1 _5498_ (.Y(_1158_),
    .A(_1144_),
    .B(net709));
 sg13g2_mux2_1 _5499_ (.A0(_1038_),
    .A1(_1101_),
    .S(net809),
    .X(_1159_));
 sg13g2_mux4_1 _5500_ (.S0(net790),
    .A0(_0928_),
    .A1(_1038_),
    .A2(_1039_),
    .A3(_1101_),
    .S1(net809),
    .X(_1160_));
 sg13g2_mux2_2 _5501_ (.A0(_1152_),
    .A1(_1160_),
    .S(net781),
    .X(_1161_));
 sg13g2_inv_2 _5502_ (.Y(_1162_),
    .A(_1161_));
 sg13g2_o21ai_1 _5503_ (.B1(_3578_),
    .Y(_1163_),
    .A1(net808),
    .A2(_1146_));
 sg13g2_a21oi_1 _5504_ (.A1(net808),
    .A2(_1045_),
    .Y(_1164_),
    .B1(_1163_));
 sg13g2_a221oi_1 _5505_ (.B2(_0821_),
    .C1(_1164_),
    .B1(net790),
    .A1(net869),
    .Y(_1165_),
    .A2(net797));
 sg13g2_a21oi_2 _5506_ (.B1(_1165_),
    .Y(_1166_),
    .A2(_1142_),
    .A1(net781));
 sg13g2_nor2b_1 _5507_ (.A(_1166_),
    .B_N(_1161_),
    .Y(_1167_));
 sg13g2_or3_2 _5508_ (.A(_1140_),
    .B(_1143_),
    .C(_1166_),
    .X(_1168_));
 sg13g2_nand2_1 _5509_ (.Y(_1169_),
    .A(net709),
    .B(_1161_));
 sg13g2_or2_1 _5510_ (.X(_1170_),
    .B(_1169_),
    .A(_1168_));
 sg13g2_a21oi_1 _5511_ (.A1(_1144_),
    .A2(net709),
    .Y(_1171_),
    .B1(_1167_));
 sg13g2_xnor2_1 _5512_ (.Y(_1172_),
    .A(_1158_),
    .B(_1167_));
 sg13g2_xnor2_1 _5513_ (.Y(_1173_),
    .A(_1056_),
    .B(_1172_));
 sg13g2_o21ai_1 _5514_ (.B1(_1170_),
    .Y(_1174_),
    .A1(_1056_),
    .A2(_1171_));
 sg13g2_nand2b_2 _5515_ (.Y(_1175_),
    .B(_1161_),
    .A_N(_1055_));
 sg13g2_inv_1 _5516_ (.Y(_1176_),
    .A(_1175_));
 sg13g2_nor2_2 _5517_ (.A(net781),
    .B(_1051_),
    .Y(_1177_));
 sg13g2_o21ai_1 _5518_ (.B1(_1096_),
    .Y(_1178_),
    .A1(_1102_),
    .A2(_1133_));
 sg13g2_o21ai_1 _5519_ (.B1(_1134_),
    .Y(_1179_),
    .A1(_1178_),
    .A2(_1099_));
 sg13g2_a21oi_1 _5520_ (.A1(_1103_),
    .A2(_1132_),
    .Y(_1180_),
    .B1(_1131_));
 sg13g2_nor2_1 _5521_ (.A(_1067_),
    .B(_1110_),
    .Y(_1181_));
 sg13g2_a21oi_1 _5522_ (.A1(_1105_),
    .A2(_1109_),
    .Y(_1182_),
    .B1(_1181_));
 sg13g2_nand2_1 _5523_ (.Y(_1183_),
    .A(_1127_),
    .B(_1129_));
 sg13g2_nor2_1 _5524_ (.A(_0380_),
    .B(_0853_),
    .Y(_1184_));
 sg13g2_xor2_1 _5525_ (.B(_1184_),
    .A(_1107_),
    .X(_1185_));
 sg13g2_a21oi_1 _5526_ (.A1(_1115_),
    .A2(_1118_),
    .Y(_1186_),
    .B1(_1185_));
 sg13g2_nand3_1 _5527_ (.B(_1118_),
    .C(_1185_),
    .A(_1115_),
    .Y(_1187_));
 sg13g2_nand2b_1 _5528_ (.Y(_1188_),
    .B(_1187_),
    .A_N(_1186_));
 sg13g2_xnor2_1 _5529_ (.Y(_1189_),
    .A(_1108_),
    .B(_1188_));
 sg13g2_a21oi_1 _5530_ (.A1(_1120_),
    .A2(_1125_),
    .Y(_1190_),
    .B1(_1121_));
 sg13g2_nand2b_1 _5531_ (.Y(_1191_),
    .B(_1122_),
    .A_N(_1080_));
 sg13g2_nor2b_1 _5532_ (.A(_1121_),
    .B_N(_1191_),
    .Y(_1192_));
 sg13g2_nand2_1 _5533_ (.Y(_1193_),
    .A(net757),
    .B(_0890_));
 sg13g2_nor2_1 _5534_ (.A(net784),
    .B(_1009_),
    .Y(_1194_));
 sg13g2_xor2_1 _5535_ (.B(_1194_),
    .A(_1114_),
    .X(_1195_));
 sg13g2_nor2b_1 _5536_ (.A(_1193_),
    .B_N(_1195_),
    .Y(_1196_));
 sg13g2_xnor2_1 _5537_ (.Y(_1197_),
    .A(_1193_),
    .B(_1195_));
 sg13g2_xnor2_1 _5538_ (.Y(_1198_),
    .A(_1192_),
    .B(_1197_));
 sg13g2_xor2_1 _5539_ (.B(_1198_),
    .A(_1190_),
    .X(_1199_));
 sg13g2_nand2b_1 _5540_ (.Y(_1200_),
    .B(_1199_),
    .A_N(_1189_));
 sg13g2_xnor2_1 _5541_ (.Y(_1201_),
    .A(_1189_),
    .B(_1199_));
 sg13g2_nand2_1 _5542_ (.Y(_1202_),
    .A(_1183_),
    .B(_1201_));
 sg13g2_xnor2_1 _5543_ (.Y(_1203_),
    .A(_1183_),
    .B(_1201_));
 sg13g2_xor2_1 _5544_ (.B(_1203_),
    .A(_1182_),
    .X(_1204_));
 sg13g2_nand2b_1 _5545_ (.Y(_1205_),
    .B(_1204_),
    .A_N(_1180_));
 sg13g2_xnor2_1 _5546_ (.Y(_1206_),
    .A(_1180_),
    .B(_1204_));
 sg13g2_inv_1 _5547_ (.Y(_1207_),
    .A(_1206_));
 sg13g2_xnor2_1 _5548_ (.Y(_1208_),
    .A(_1179_),
    .B(_1206_));
 sg13g2_nand2b_1 _5549_ (.Y(_1209_),
    .B(net809),
    .A_N(_1208_));
 sg13g2_a21oi_1 _5550_ (.A1(net807),
    .A2(_1137_),
    .Y(_1210_),
    .B1(_3578_));
 sg13g2_a221oi_1 _5551_ (.B2(_1209_),
    .C1(_0816_),
    .B1(_1210_),
    .A1(_2695_),
    .Y(_1211_),
    .A2(_1159_));
 sg13g2_or2_1 _5552_ (.X(_1212_),
    .B(_1211_),
    .A(_1177_));
 sg13g2_nor3_2 _5553_ (.A(_1166_),
    .B(_1177_),
    .C(net156),
    .Y(_1213_));
 sg13g2_inv_1 _5554_ (.Y(_1214_),
    .A(_1213_));
 sg13g2_nor3_2 _5555_ (.A(_1156_),
    .B(_1177_),
    .C(_1211_),
    .Y(_1215_));
 sg13g2_nor2_1 _5556_ (.A(_1158_),
    .B(_1214_),
    .Y(_1216_));
 sg13g2_xnor2_1 _5557_ (.Y(_1217_),
    .A(_1168_),
    .B(_1215_));
 sg13g2_xnor2_1 _5558_ (.Y(_1218_),
    .A(_1175_),
    .B(_1217_));
 sg13g2_nand2_1 _5559_ (.Y(_1219_),
    .A(_1174_),
    .B(_1218_));
 sg13g2_xnor2_1 _5560_ (.Y(_1220_),
    .A(_1174_),
    .B(_1218_));
 sg13g2_nor2_1 _5561_ (.A(_1043_),
    .B(_1162_),
    .Y(_1221_));
 sg13g2_xnor2_1 _5562_ (.Y(_1222_),
    .A(_1042_),
    .B(_1175_));
 sg13g2_nand2b_1 _5563_ (.Y(_1223_),
    .B(_1222_),
    .A_N(_1168_));
 sg13g2_xor2_1 _5564_ (.B(_1222_),
    .A(_1168_),
    .X(_1224_));
 sg13g2_xor2_1 _5565_ (.B(_1224_),
    .A(_1220_),
    .X(_1225_));
 sg13g2_nand2_1 _5566_ (.Y(_1226_),
    .A(_1173_),
    .B(_1225_));
 sg13g2_nand2_1 _5567_ (.Y(_1227_),
    .A(_1174_),
    .B(_1215_));
 sg13g2_xnor2_1 _5568_ (.Y(_1228_),
    .A(_1174_),
    .B(_1215_));
 sg13g2_nor2_1 _5569_ (.A(_1173_),
    .B(_1225_),
    .Y(_1229_));
 sg13g2_o21ai_1 _5570_ (.B1(_1226_),
    .Y(_1230_),
    .A1(_1228_),
    .A2(_1229_));
 sg13g2_o21ai_1 _5571_ (.B1(_1219_),
    .Y(_1231_),
    .A1(_1220_),
    .A2(_1224_));
 sg13g2_o21ai_1 _5572_ (.B1(_1205_),
    .Y(_1232_),
    .A1(_1179_),
    .A2(_1207_));
 sg13g2_o21ai_1 _5573_ (.B1(_1202_),
    .Y(_1233_),
    .A1(_1182_),
    .A2(_1203_));
 sg13g2_o21ai_1 _5574_ (.B1(_1200_),
    .Y(_1234_),
    .A1(_1190_),
    .A2(_1198_));
 sg13g2_nor2_1 _5575_ (.A(_1108_),
    .B(_1188_),
    .Y(_1235_));
 sg13g2_nor2_1 _5576_ (.A(_1186_),
    .B(_1235_),
    .Y(_1236_));
 sg13g2_xnor2_1 _5577_ (.Y(_1237_),
    .A(net772),
    .B(net785));
 sg13g2_nor2_1 _5578_ (.A(_1009_),
    .B(_1237_),
    .Y(_1238_));
 sg13g2_nand2_1 _5579_ (.Y(_1239_),
    .A(net746),
    .B(_0890_));
 sg13g2_nand4_1 _5580_ (.B(_0851_),
    .C(_0852_),
    .A(net756),
    .Y(_1240_),
    .D(_1106_));
 sg13g2_o21ai_1 _5581_ (.B1(_1240_),
    .Y(_1241_),
    .A1(_0325_),
    .A2(_0967_));
 sg13g2_xnor2_1 _5582_ (.Y(_1242_),
    .A(_1239_),
    .B(_1241_));
 sg13g2_xnor2_1 _5583_ (.Y(_1243_),
    .A(_1238_),
    .B(_1242_));
 sg13g2_xnor2_1 _5584_ (.Y(_1244_),
    .A(_1236_),
    .B(_1243_));
 sg13g2_a21oi_1 _5585_ (.A1(_1114_),
    .A2(_1194_),
    .Y(_1245_),
    .B1(_1196_));
 sg13g2_nand2b_1 _5586_ (.Y(_1246_),
    .B(_1197_),
    .A_N(_1121_));
 sg13g2_nand2_1 _5587_ (.Y(_1247_),
    .A(_1191_),
    .B(_1246_));
 sg13g2_xor2_1 _5588_ (.B(_1247_),
    .A(_1245_),
    .X(_1248_));
 sg13g2_xnor2_1 _5589_ (.Y(_1249_),
    .A(_1244_),
    .B(_1248_));
 sg13g2_xnor2_1 _5590_ (.Y(_1250_),
    .A(_1234_),
    .B(_1249_));
 sg13g2_xnor2_1 _5591_ (.Y(_1251_),
    .A(_1233_),
    .B(_1250_));
 sg13g2_xnor2_1 _5592_ (.Y(_1252_),
    .A(_1232_),
    .B(_1251_));
 sg13g2_o21ai_1 _5593_ (.B1(net790),
    .Y(_1253_),
    .A1(net809),
    .A2(_1208_));
 sg13g2_a21o_1 _5594_ (.A2(_1252_),
    .A1(net809),
    .B1(_1253_),
    .X(_1254_));
 sg13g2_a21oi_1 _5595_ (.A1(_2695_),
    .A2(_1139_),
    .Y(_1255_),
    .B1(_0816_));
 sg13g2_a22oi_1 _5596_ (.Y(_1256_),
    .B1(_1254_),
    .B2(_1255_),
    .A2(_1041_),
    .A1(_0816_));
 sg13g2_inv_1 _5597_ (.Y(_1257_),
    .A(net706));
 sg13g2_nand2_1 _5598_ (.Y(_1258_),
    .A(net709),
    .B(net706));
 sg13g2_a21oi_1 _5599_ (.A1(net709),
    .A2(net706),
    .Y(_1259_),
    .B1(_1213_));
 sg13g2_nand2b_2 _5600_ (.Y(_1260_),
    .B(net706),
    .A_N(_1166_));
 sg13g2_nand3_1 _5601_ (.B(_1213_),
    .C(net706),
    .A(net709),
    .Y(_1261_));
 sg13g2_nand2b_1 _5602_ (.Y(_1262_),
    .B(_1261_),
    .A_N(_1259_));
 sg13g2_a21oi_1 _5603_ (.A1(_1176_),
    .A2(_1217_),
    .Y(_1263_),
    .B1(_1216_));
 sg13g2_xor2_1 _5604_ (.B(_1263_),
    .A(_1262_),
    .X(_1264_));
 sg13g2_and2_1 _5605_ (.A(_1231_),
    .B(_1264_),
    .X(_1265_));
 sg13g2_xor2_1 _5606_ (.B(_1264_),
    .A(_1231_),
    .X(_1266_));
 sg13g2_o21ai_1 _5607_ (.B1(_1223_),
    .Y(_1267_),
    .A1(_1043_),
    .A2(_1175_));
 sg13g2_xnor2_1 _5608_ (.Y(_1268_),
    .A(_1214_),
    .B(_1267_));
 sg13g2_nor2b_1 _5609_ (.A(_1258_),
    .B_N(_1268_),
    .Y(_1269_));
 sg13g2_xnor2_1 _5610_ (.Y(_1270_),
    .A(_1258_),
    .B(_1268_));
 sg13g2_xnor2_1 _5611_ (.Y(_1271_),
    .A(_1266_),
    .B(_1270_));
 sg13g2_nand2b_1 _5612_ (.Y(_1272_),
    .B(_1230_),
    .A_N(_1271_));
 sg13g2_xor2_1 _5613_ (.B(_1271_),
    .A(_1230_),
    .X(_1273_));
 sg13g2_o21ai_1 _5614_ (.B1(_1272_),
    .Y(_1274_),
    .A1(_1227_),
    .A2(_1273_));
 sg13g2_a21o_1 _5615_ (.A2(_1267_),
    .A1(_1213_),
    .B1(_1269_),
    .X(_1275_));
 sg13g2_a21oi_2 _5616_ (.B1(_1265_),
    .Y(_1276_),
    .A2(_1270_),
    .A1(_1266_));
 sg13g2_nor2_1 _5617_ (.A(_1055_),
    .B(net707),
    .Y(_1277_));
 sg13g2_nand2b_2 _5618_ (.Y(_1278_),
    .B(net706),
    .A_N(_1055_));
 sg13g2_xnor2_1 _5619_ (.Y(_1279_),
    .A(_1260_),
    .B(_1277_));
 sg13g2_nand2b_1 _5620_ (.Y(_1280_),
    .B(_1144_),
    .A_N(_1055_));
 sg13g2_a21oi_1 _5621_ (.A1(_1261_),
    .A2(_1280_),
    .Y(_1281_),
    .B1(_1259_));
 sg13g2_nand2_1 _5622_ (.Y(_1282_),
    .A(_1279_),
    .B(_1281_));
 sg13g2_xnor2_1 _5623_ (.Y(_1283_),
    .A(_1279_),
    .B(_1281_));
 sg13g2_xnor2_1 _5624_ (.Y(_1284_),
    .A(_1283_),
    .B(_1162_));
 sg13g2_mux2_1 _5625_ (.A0(_1263_),
    .A1(_1280_),
    .S(_1262_),
    .X(_1285_));
 sg13g2_nor2_1 _5626_ (.A(_1284_),
    .B(_1285_),
    .Y(_1286_));
 sg13g2_xor2_1 _5627_ (.B(_1284_),
    .A(_1285_),
    .X(_1287_));
 sg13g2_nor2_1 _5628_ (.A(_1162_),
    .B(net707),
    .Y(_1288_));
 sg13g2_nor2_1 _5629_ (.A(_1043_),
    .B(net707),
    .Y(_1289_));
 sg13g2_inv_1 _5630_ (.Y(_1290_),
    .A(_1289_));
 sg13g2_nand2_1 _5631_ (.Y(_1291_),
    .A(_1176_),
    .B(_1289_));
 sg13g2_o21ai_1 _5632_ (.B1(_1291_),
    .Y(_1292_),
    .A1(_1221_),
    .A2(_1277_));
 sg13g2_xor2_1 _5633_ (.B(_1292_),
    .A(_1260_),
    .X(_1293_));
 sg13g2_xnor2_1 _5634_ (.Y(_1294_),
    .A(_1287_),
    .B(_1293_));
 sg13g2_xor2_1 _5635_ (.B(_1276_),
    .A(_1294_),
    .X(_1295_));
 sg13g2_nand2_1 _5636_ (.Y(_1296_),
    .A(_1275_),
    .B(_1295_));
 sg13g2_xnor2_1 _5637_ (.Y(_1297_),
    .A(_1275_),
    .B(_1295_));
 sg13g2_nor2b_1 _5638_ (.A(_1297_),
    .B_N(_1274_),
    .Y(_1298_));
 sg13g2_or2_1 _5639_ (.X(_1299_),
    .B(_1166_),
    .A(_1043_));
 sg13g2_nor2_1 _5640_ (.A(_1169_),
    .B(_1299_),
    .Y(_1300_));
 sg13g2_and2_1 _5641_ (.A(_1169_),
    .B(_1299_),
    .X(_1301_));
 sg13g2_or2_1 _5642_ (.X(_1302_),
    .B(_1166_),
    .A(_1055_));
 sg13g2_nor2_1 _5643_ (.A(_1301_),
    .B(_1302_),
    .Y(_1303_));
 sg13g2_nor2_1 _5644_ (.A(_1300_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_xnor2_1 _5645_ (.Y(_1305_),
    .A(_1043_),
    .B(_1173_));
 sg13g2_nand2b_1 _5646_ (.Y(_1306_),
    .B(_1305_),
    .A_N(_1304_));
 sg13g2_xor2_1 _5647_ (.B(_1305_),
    .A(_1304_),
    .X(_1307_));
 sg13g2_nand2b_2 _5648_ (.Y(_1308_),
    .B(net709),
    .A_N(_1056_));
 sg13g2_nor2_1 _5649_ (.A(_1300_),
    .B(_1301_),
    .Y(_1309_));
 sg13g2_xor2_1 _5650_ (.B(_1309_),
    .A(_1302_),
    .X(_1310_));
 sg13g2_or2_1 _5651_ (.X(_1311_),
    .B(_1310_),
    .A(_1308_));
 sg13g2_o21ai_1 _5652_ (.B1(_1306_),
    .Y(_1312_),
    .A1(_1307_),
    .A2(_1311_));
 sg13g2_xor2_1 _5653_ (.B(_1273_),
    .A(_1227_),
    .X(_1313_));
 sg13g2_and2_1 _5654_ (.A(_1312_),
    .B(_1313_),
    .X(_1314_));
 sg13g2_nand2b_1 _5655_ (.Y(_1315_),
    .B(_1297_),
    .A_N(_1274_));
 sg13g2_xor2_1 _5656_ (.B(_1297_),
    .A(_1274_),
    .X(_1316_));
 sg13g2_a21oi_1 _5657_ (.A1(_1314_),
    .A2(_1315_),
    .Y(_1317_),
    .B1(_1298_));
 sg13g2_o21ai_1 _5658_ (.B1(_1296_),
    .Y(_1318_),
    .A1(_1276_),
    .A2(_1294_));
 sg13g2_o21ai_1 _5659_ (.B1(_1291_),
    .Y(_1319_),
    .A1(_1260_),
    .A2(_1292_));
 sg13g2_a21oi_1 _5660_ (.A1(_1287_),
    .A2(_1293_),
    .Y(_1320_),
    .B1(_1286_));
 sg13g2_o21ai_1 _5661_ (.B1(_1282_),
    .Y(_1321_),
    .A1(_1162_),
    .A2(_1283_));
 sg13g2_nor2_1 _5662_ (.A(_1213_),
    .B(_1278_),
    .Y(_1322_));
 sg13g2_xnor2_1 _5663_ (.Y(_1323_),
    .A(_1289_),
    .B(_1322_));
 sg13g2_nand2b_1 _5664_ (.Y(_1324_),
    .B(_1321_),
    .A_N(_1323_));
 sg13g2_xor2_1 _5665_ (.B(_1323_),
    .A(_1321_),
    .X(_1325_));
 sg13g2_nor2_1 _5666_ (.A(_1145_),
    .B(net707),
    .Y(_1326_));
 sg13g2_xnor2_1 _5667_ (.Y(_1327_),
    .A(_1145_),
    .B(net707));
 sg13g2_or2_1 _5668_ (.X(_1328_),
    .B(_1327_),
    .A(_1043_));
 sg13g2_nor2_1 _5669_ (.A(_1278_),
    .B(_1328_),
    .Y(_1329_));
 sg13g2_xor2_1 _5670_ (.B(_1328_),
    .A(_1278_),
    .X(_1330_));
 sg13g2_inv_1 _5671_ (.Y(_1331_),
    .A(_1330_));
 sg13g2_xnor2_1 _5672_ (.Y(_1332_),
    .A(_1325_),
    .B(_1331_));
 sg13g2_or2_1 _5673_ (.X(_1333_),
    .B(_1332_),
    .A(_1320_));
 sg13g2_xor2_1 _5674_ (.B(_1332_),
    .A(_1320_),
    .X(_1334_));
 sg13g2_nand2_1 _5675_ (.Y(_1335_),
    .A(_1319_),
    .B(_1334_));
 sg13g2_xnor2_1 _5676_ (.Y(_1336_),
    .A(_1319_),
    .B(_1334_));
 sg13g2_inv_1 _5677_ (.Y(_1337_),
    .A(_1336_));
 sg13g2_nor2_1 _5678_ (.A(_1318_),
    .B(_1337_),
    .Y(_1338_));
 sg13g2_xnor2_1 _5679_ (.Y(_1339_),
    .A(_1318_),
    .B(_1336_));
 sg13g2_xnor2_1 _5680_ (.Y(_1340_),
    .A(_1317_),
    .B(_1339_));
 sg13g2_nand2_1 _5681_ (.Y(_1341_),
    .A(net886),
    .B(_1340_));
 sg13g2_xnor2_1 _5682_ (.Y(_1342_),
    .A(_1314_),
    .B(_1316_));
 sg13g2_and2_1 _5683_ (.A(net812),
    .B(_1342_),
    .X(_1343_));
 sg13g2_and3_1 _5684_ (.X(_1344_),
    .A(net887),
    .B(_1340_),
    .C(_1343_));
 sg13g2_xor2_1 _5685_ (.B(_1313_),
    .A(_1312_),
    .X(_1345_));
 sg13g2_nand2_1 _5686_ (.Y(_1346_),
    .A(net881),
    .B(_1345_));
 sg13g2_a22oi_1 _5687_ (.Y(_1347_),
    .B1(_1342_),
    .B2(net887),
    .A2(_1340_),
    .A1(net812));
 sg13g2_or3_1 _5688_ (.A(_1344_),
    .B(_1346_),
    .C(_1347_),
    .X(_1348_));
 sg13g2_nand2b_1 _5689_ (.Y(_1349_),
    .B(_1348_),
    .A_N(_1344_));
 sg13g2_nand2_1 _5690_ (.Y(_1350_),
    .A(net881),
    .B(_1342_));
 sg13g2_inv_1 _5691_ (.Y(_1351_),
    .A(_1350_));
 sg13g2_a21oi_2 _5692_ (.B1(_1329_),
    .Y(_1352_),
    .A2(_1326_),
    .A1(_1042_));
 sg13g2_o21ai_1 _5693_ (.B1(_1324_),
    .Y(_1353_),
    .A1(_1325_),
    .A2(_1331_));
 sg13g2_nand2_1 _5694_ (.Y(_1354_),
    .A(_1042_),
    .B(net706));
 sg13g2_nor2_1 _5695_ (.A(_1162_),
    .B(_1327_),
    .Y(_1355_));
 sg13g2_nand2_1 _5696_ (.Y(_1356_),
    .A(_1161_),
    .B(net706));
 sg13g2_xnor2_1 _5697_ (.Y(_1357_),
    .A(_1354_),
    .B(_1355_));
 sg13g2_a21oi_1 _5698_ (.A1(_1214_),
    .A2(_1290_),
    .Y(_1358_),
    .B1(_1278_));
 sg13g2_nand2b_2 _5699_ (.Y(_1359_),
    .B(_1256_),
    .A_N(net708));
 sg13g2_nor3_1 _5700_ (.A(_1162_),
    .B(net707),
    .C(_1354_),
    .Y(_1360_));
 sg13g2_xor2_1 _5701_ (.B(_1354_),
    .A(_1288_),
    .X(_1361_));
 sg13g2_nor2_1 _5702_ (.A(_1145_),
    .B(_1361_),
    .Y(_1362_));
 sg13g2_xnor2_1 _5703_ (.Y(_1363_),
    .A(_1144_),
    .B(_1361_));
 sg13g2_and2_1 _5704_ (.A(_1358_),
    .B(_1363_),
    .X(_1364_));
 sg13g2_xor2_1 _5705_ (.B(_1363_),
    .A(_1358_),
    .X(_1365_));
 sg13g2_xnor2_1 _5706_ (.Y(_1366_),
    .A(_1357_),
    .B(_1365_));
 sg13g2_nor2b_1 _5707_ (.A(_1366_),
    .B_N(_1353_),
    .Y(_1367_));
 sg13g2_xnor2_1 _5708_ (.Y(_1368_),
    .A(_1353_),
    .B(_1366_));
 sg13g2_nor2b_1 _5709_ (.A(_1352_),
    .B_N(_1368_),
    .Y(_1369_));
 sg13g2_xor2_1 _5710_ (.B(_1368_),
    .A(_1352_),
    .X(_1370_));
 sg13g2_a21oi_1 _5711_ (.A1(_1333_),
    .A2(_1335_),
    .Y(_1371_),
    .B1(_1370_));
 sg13g2_inv_1 _5712_ (.Y(_1372_),
    .A(_1371_));
 sg13g2_nand3_1 _5713_ (.B(_1335_),
    .C(_1370_),
    .A(_1333_),
    .Y(_1373_));
 sg13g2_nand2b_1 _5714_ (.Y(_1374_),
    .B(_1373_),
    .A_N(_1371_));
 sg13g2_a221oi_1 _5715_ (.B2(_1337_),
    .C1(_1298_),
    .B1(_1318_),
    .A1(_1315_),
    .Y(_1375_),
    .A2(_1314_));
 sg13g2_or3_2 _5716_ (.A(_1338_),
    .B(_1375_),
    .C(_1374_),
    .X(_1376_));
 sg13g2_o21ai_1 _5717_ (.B1(_1374_),
    .Y(_1377_),
    .A1(_1338_),
    .A2(net158));
 sg13g2_and2_2 _5718_ (.A(_1376_),
    .B(_1377_),
    .X(_1378_));
 sg13g2_and2_1 _5719_ (.A(net886),
    .B(_1378_),
    .X(_1379_));
 sg13g2_nand3_1 _5720_ (.B(_1376_),
    .C(_1377_),
    .A(net812),
    .Y(_1380_));
 sg13g2_nor2_1 _5721_ (.A(_1341_),
    .B(_1380_),
    .Y(_1381_));
 sg13g2_xor2_1 _5722_ (.B(_1380_),
    .A(_1341_),
    .X(_1382_));
 sg13g2_xnor2_1 _5723_ (.Y(_1383_),
    .A(_1350_),
    .B(_1382_));
 sg13g2_nand2_1 _5724_ (.Y(_1384_),
    .A(_1349_),
    .B(_1383_));
 sg13g2_xor2_1 _5725_ (.B(_1310_),
    .A(_1308_),
    .X(_1385_));
 sg13g2_nand2_1 _5726_ (.Y(_1386_),
    .A(net865),
    .B(_1385_));
 sg13g2_xor2_1 _5727_ (.B(_1311_),
    .A(_1307_),
    .X(_1387_));
 sg13g2_nand2_1 _5728_ (.Y(_1388_),
    .A(net876),
    .B(_1387_));
 sg13g2_nand2_1 _5729_ (.Y(_1389_),
    .A(net876),
    .B(_1345_));
 sg13g2_nand2_1 _5730_ (.Y(_1390_),
    .A(net871),
    .B(_1387_));
 sg13g2_xor2_1 _5731_ (.B(_1390_),
    .A(_1389_),
    .X(_1391_));
 sg13g2_nand2b_1 _5732_ (.Y(_1392_),
    .B(_1391_),
    .A_N(_1386_));
 sg13g2_xor2_1 _5733_ (.B(_1391_),
    .A(_1386_),
    .X(_1393_));
 sg13g2_xnor2_1 _5734_ (.Y(_1394_),
    .A(_1349_),
    .B(_1383_));
 sg13g2_o21ai_1 _5735_ (.B1(_1384_),
    .Y(_1395_),
    .A1(_1393_),
    .A2(_1394_));
 sg13g2_nand2_1 _5736_ (.Y(_1396_),
    .A(net865),
    .B(_1387_));
 sg13g2_inv_1 _5737_ (.Y(_1397_),
    .A(_1396_));
 sg13g2_nand2_1 _5738_ (.Y(_1398_),
    .A(net870),
    .B(_1342_));
 sg13g2_nor2_1 _5739_ (.A(_1389_),
    .B(_1398_),
    .Y(_1399_));
 sg13g2_a22oi_1 _5740_ (.Y(_1400_),
    .B1(_1345_),
    .B2(net870),
    .A2(_1342_),
    .A1(net876));
 sg13g2_nor2_1 _5741_ (.A(_1399_),
    .B(_1400_),
    .Y(_1401_));
 sg13g2_xnor2_1 _5742_ (.Y(_1402_),
    .A(_1396_),
    .B(_1401_));
 sg13g2_a21oi_1 _5743_ (.A1(_1351_),
    .A2(_1382_),
    .Y(_1403_),
    .B1(_1381_));
 sg13g2_nand2_1 _5744_ (.Y(_1404_),
    .A(net881),
    .B(_1340_));
 sg13g2_nor2_2 _5745_ (.A(_1367_),
    .B(_1369_),
    .Y(_1405_));
 sg13g2_nand2_1 _5746_ (.Y(_1406_),
    .A(_1161_),
    .B(_1326_));
 sg13g2_o21ai_1 _5747_ (.B1(_1406_),
    .Y(_1407_),
    .A1(_1328_),
    .A2(_1356_));
 sg13g2_nor2_1 _5748_ (.A(_1360_),
    .B(_1362_),
    .Y(_1408_));
 sg13g2_a21oi_1 _5749_ (.A1(_1357_),
    .A2(_1365_),
    .Y(_1409_),
    .B1(_1364_));
 sg13g2_nor2_1 _5750_ (.A(_1408_),
    .B(_1409_),
    .Y(_1410_));
 sg13g2_xor2_1 _5751_ (.B(_1409_),
    .A(_1408_),
    .X(_1411_));
 sg13g2_xnor2_1 _5752_ (.Y(_1412_),
    .A(_1407_),
    .B(_1411_));
 sg13g2_nor2_1 _5753_ (.A(_1405_),
    .B(_1412_),
    .Y(_1413_));
 sg13g2_xnor2_1 _5754_ (.Y(_1414_),
    .A(_1405_),
    .B(_1412_));
 sg13g2_a21oi_2 _5755_ (.B1(_1414_),
    .Y(_1415_),
    .A2(_1376_),
    .A1(_1372_));
 sg13g2_and3_1 _5756_ (.X(_1416_),
    .A(_1372_),
    .B(_1376_),
    .C(_1414_));
 sg13g2_nor2_2 _5757_ (.A(_1415_),
    .B(_1416_),
    .Y(_1417_));
 sg13g2_nor3_2 _5758_ (.A(net892),
    .B(_1415_),
    .C(_1416_),
    .Y(_1418_));
 sg13g2_xor2_1 _5759_ (.B(_1418_),
    .A(_1379_),
    .X(_1419_));
 sg13g2_nor2b_1 _5760_ (.A(_1404_),
    .B_N(_1419_),
    .Y(_1420_));
 sg13g2_xnor2_1 _5761_ (.Y(_1421_),
    .A(_1404_),
    .B(_1419_));
 sg13g2_nor2b_1 _5762_ (.A(_1403_),
    .B_N(_1421_),
    .Y(_1422_));
 sg13g2_xnor2_1 _5763_ (.Y(_1423_),
    .A(_1403_),
    .B(_1421_));
 sg13g2_xnor2_1 _5764_ (.Y(_1424_),
    .A(_1402_),
    .B(_1423_));
 sg13g2_nand2b_1 _5765_ (.Y(_1425_),
    .B(_1395_),
    .A_N(_1424_));
 sg13g2_o21ai_1 _5766_ (.B1(_1392_),
    .Y(_1426_),
    .A1(_1389_),
    .A2(_1390_));
 sg13g2_xor2_1 _5767_ (.B(_1424_),
    .A(_1395_),
    .X(_1427_));
 sg13g2_nand2b_1 _5768_ (.Y(_1428_),
    .B(_1426_),
    .A_N(_1427_));
 sg13g2_nand2_1 _5769_ (.Y(_1429_),
    .A(_1425_),
    .B(_1428_));
 sg13g2_a21oi_1 _5770_ (.A1(_1397_),
    .A2(_1401_),
    .Y(_1430_),
    .B1(_1399_));
 sg13g2_a21o_1 _5771_ (.A2(_1423_),
    .A1(_1402_),
    .B1(_1422_),
    .X(_1431_));
 sg13g2_a21o_1 _5772_ (.A2(_1418_),
    .A1(_1379_),
    .B1(_1420_),
    .X(_1432_));
 sg13g2_and2_1 _5773_ (.A(net881),
    .B(_1378_),
    .X(_1433_));
 sg13g2_nor2_1 _5774_ (.A(_1257_),
    .B(_1406_),
    .Y(_1434_));
 sg13g2_nor2_1 _5775_ (.A(net707),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_nor2b_1 _5776_ (.A(_1326_),
    .B_N(_1356_),
    .Y(_1436_));
 sg13g2_nor3_2 _5777_ (.A(net708),
    .B(_1434_),
    .C(_1436_),
    .Y(_1437_));
 sg13g2_a21oi_1 _5778_ (.A1(net707),
    .A2(_1356_),
    .Y(_1438_),
    .B1(_1437_));
 sg13g2_a21oi_1 _5779_ (.A1(_1407_),
    .A2(_1411_),
    .Y(_1439_),
    .B1(_1410_));
 sg13g2_nor2b_1 _5780_ (.A(_1439_),
    .B_N(_1438_),
    .Y(_1440_));
 sg13g2_xnor2_1 _5781_ (.Y(_1441_),
    .A(_1438_),
    .B(_1439_));
 sg13g2_inv_1 _5782_ (.Y(_1442_),
    .A(_1441_));
 sg13g2_nor2_1 _5783_ (.A(_1371_),
    .B(_1413_),
    .Y(_1443_));
 sg13g2_a22oi_1 _5784_ (.Y(_1444_),
    .B1(_1443_),
    .B2(_1376_),
    .A2(_1412_),
    .A1(_1405_));
 sg13g2_a221oi_1 _5785_ (.B2(_1376_),
    .C1(_1442_),
    .B1(_1443_),
    .A1(_1405_),
    .Y(_1445_),
    .A2(_1412_));
 sg13g2_xnor2_1 _5786_ (.Y(_1446_),
    .A(_1442_),
    .B(_1444_));
 sg13g2_nand2_1 _5787_ (.Y(_1447_),
    .A(net886),
    .B(_1446_));
 sg13g2_and3_1 _5788_ (.X(_1448_),
    .A(net886),
    .B(_1418_),
    .C(_1446_));
 sg13g2_a22oi_1 _5789_ (.Y(_1449_),
    .B1(_1446_),
    .B2(net812),
    .A2(_1417_),
    .A1(net886));
 sg13g2_nor2_1 _5790_ (.A(_1448_),
    .B(_1449_),
    .Y(_1450_));
 sg13g2_xor2_1 _5791_ (.B(_1450_),
    .A(_1433_),
    .X(_1451_));
 sg13g2_nand2_1 _5792_ (.Y(_1452_),
    .A(_1432_),
    .B(_1451_));
 sg13g2_xnor2_1 _5793_ (.Y(_1453_),
    .A(_1432_),
    .B(_1451_));
 sg13g2_nand2_1 _5794_ (.Y(_1454_),
    .A(net864),
    .B(_1345_));
 sg13g2_nand2_1 _5795_ (.Y(_1455_),
    .A(net876),
    .B(_1340_));
 sg13g2_xor2_1 _5796_ (.B(_1455_),
    .A(_1398_),
    .X(_1456_));
 sg13g2_nand2b_1 _5797_ (.Y(_1457_),
    .B(_1456_),
    .A_N(_1454_));
 sg13g2_xor2_1 _5798_ (.B(_1456_),
    .A(_1454_),
    .X(_1458_));
 sg13g2_xor2_1 _5799_ (.B(_1458_),
    .A(_1453_),
    .X(_1459_));
 sg13g2_nand2_1 _5800_ (.Y(_1460_),
    .A(_1431_),
    .B(_1459_));
 sg13g2_xnor2_1 _5801_ (.Y(_1461_),
    .A(_1431_),
    .B(_1459_));
 sg13g2_xnor2_1 _5802_ (.Y(_1462_),
    .A(_1430_),
    .B(_1461_));
 sg13g2_nand2b_1 _5803_ (.Y(_1463_),
    .B(_1429_),
    .A_N(_1462_));
 sg13g2_nand2_1 _5804_ (.Y(_1464_),
    .A(net856),
    .B(_1387_));
 sg13g2_xnor2_1 _5805_ (.Y(_1465_),
    .A(_1429_),
    .B(_1462_));
 sg13g2_nand2b_1 _5806_ (.Y(_1466_),
    .B(_1465_),
    .A_N(_1464_));
 sg13g2_nand2_1 _5807_ (.Y(_1467_),
    .A(net856),
    .B(_1345_));
 sg13g2_o21ai_1 _5808_ (.B1(_1460_),
    .Y(_1468_),
    .A1(_1430_),
    .A2(_1461_));
 sg13g2_o21ai_1 _5809_ (.B1(_1457_),
    .Y(_1469_),
    .A1(_1398_),
    .A2(_1455_));
 sg13g2_o21ai_1 _5810_ (.B1(_1452_),
    .Y(_1470_),
    .A1(_1453_),
    .A2(_1458_));
 sg13g2_nand2_1 _5811_ (.Y(_1471_),
    .A(net864),
    .B(_1342_));
 sg13g2_inv_1 _5812_ (.Y(_1472_),
    .A(_1471_));
 sg13g2_nand2_1 _5813_ (.Y(_1473_),
    .A(net870),
    .B(_1378_));
 sg13g2_nor2_1 _5814_ (.A(_1455_),
    .B(_1473_),
    .Y(_1474_));
 sg13g2_a22oi_1 _5815_ (.Y(_1475_),
    .B1(_1378_),
    .B2(net876),
    .A2(_1340_),
    .A1(net870));
 sg13g2_nor2_1 _5816_ (.A(_1474_),
    .B(_1475_),
    .Y(_1476_));
 sg13g2_xnor2_1 _5817_ (.Y(_1477_),
    .A(_1471_),
    .B(_1476_));
 sg13g2_a21oi_1 _5818_ (.A1(_1433_),
    .A2(_1450_),
    .Y(_1478_),
    .B1(_1448_));
 sg13g2_nand2_1 _5819_ (.Y(_1479_),
    .A(net882),
    .B(_1417_));
 sg13g2_nor3_1 _5820_ (.A(_1145_),
    .B(_1257_),
    .C(_1288_),
    .Y(_1480_));
 sg13g2_and2_1 _5821_ (.A(_1437_),
    .B(_1480_),
    .X(_1481_));
 sg13g2_xor2_1 _5822_ (.B(_1480_),
    .A(_1437_),
    .X(_1482_));
 sg13g2_or3_1 _5823_ (.A(_1440_),
    .B(_1445_),
    .C(_1482_),
    .X(_1483_));
 sg13g2_o21ai_1 _5824_ (.B1(_1482_),
    .Y(_1484_),
    .A1(_1440_),
    .A2(_1445_));
 sg13g2_and2_2 _5825_ (.A(_1483_),
    .B(_1484_),
    .X(_1485_));
 sg13g2_nand3_1 _5826_ (.B(_1483_),
    .C(_1484_),
    .A(net886),
    .Y(_1486_));
 sg13g2_nand3_1 _5827_ (.B(_1483_),
    .C(_1484_),
    .A(net812),
    .Y(_1487_));
 sg13g2_or2_1 _5828_ (.X(_1488_),
    .B(_1487_),
    .A(_1447_));
 sg13g2_and2_1 _5829_ (.A(_1447_),
    .B(_1487_),
    .X(_1489_));
 sg13g2_xor2_1 _5830_ (.B(_1487_),
    .A(_1447_),
    .X(_1490_));
 sg13g2_xnor2_1 _5831_ (.Y(_1491_),
    .A(_1479_),
    .B(_1490_));
 sg13g2_nor2b_1 _5832_ (.A(_1478_),
    .B_N(_1491_),
    .Y(_1492_));
 sg13g2_xnor2_1 _5833_ (.Y(_1493_),
    .A(_1478_),
    .B(_1491_));
 sg13g2_xnor2_1 _5834_ (.Y(_1494_),
    .A(_1477_),
    .B(_1493_));
 sg13g2_nor2b_1 _5835_ (.A(_1494_),
    .B_N(_1470_),
    .Y(_1495_));
 sg13g2_xnor2_1 _5836_ (.Y(_1496_),
    .A(_1470_),
    .B(_1494_));
 sg13g2_xnor2_1 _5837_ (.Y(_1497_),
    .A(_1469_),
    .B(_1496_));
 sg13g2_nor2b_1 _5838_ (.A(_1497_),
    .B_N(_1468_),
    .Y(_1498_));
 sg13g2_xor2_1 _5839_ (.B(_1497_),
    .A(_1468_),
    .X(_1499_));
 sg13g2_nor2_1 _5840_ (.A(_1467_),
    .B(_1499_),
    .Y(_1500_));
 sg13g2_xnor2_1 _5841_ (.Y(_1501_),
    .A(_1467_),
    .B(_1499_));
 sg13g2_a21o_1 _5842_ (.A2(_1466_),
    .A1(_1463_),
    .B1(_1501_),
    .X(_1502_));
 sg13g2_nand3_1 _5843_ (.B(_1466_),
    .C(_1501_),
    .A(_1463_),
    .Y(_1503_));
 sg13g2_nand2_1 _5844_ (.Y(_1504_),
    .A(net812),
    .B(_1345_));
 sg13g2_nand2_1 _5845_ (.Y(_1505_),
    .A(net886),
    .B(_1345_));
 sg13g2_inv_1 _5846_ (.Y(_1506_),
    .A(_1505_));
 sg13g2_and2_1 _5847_ (.A(_1343_),
    .B(_1506_),
    .X(_1507_));
 sg13g2_nand2_1 _5848_ (.Y(_1508_),
    .A(net881),
    .B(_1387_));
 sg13g2_inv_1 _5849_ (.Y(_1509_),
    .A(_1508_));
 sg13g2_xnor2_1 _5850_ (.Y(_1510_),
    .A(_1343_),
    .B(_1505_));
 sg13g2_a21o_1 _5851_ (.A2(_1510_),
    .A1(_1509_),
    .B1(_1507_),
    .X(_1511_));
 sg13g2_o21ai_1 _5852_ (.B1(_1346_),
    .Y(_1512_),
    .A1(_1344_),
    .A2(_1347_));
 sg13g2_nand3_1 _5853_ (.B(_1511_),
    .C(_1512_),
    .A(_1348_),
    .Y(_1513_));
 sg13g2_o21ai_1 _5854_ (.B1(_1055_),
    .Y(_1514_),
    .A1(_1043_),
    .A2(_1156_));
 sg13g2_nor2_1 _5855_ (.A(net709),
    .B(_1166_),
    .Y(_1515_));
 sg13g2_nand2_2 _5856_ (.Y(_1516_),
    .A(_1308_),
    .B(_1514_));
 sg13g2_nor2_2 _5857_ (.A(net705),
    .B(_1516_),
    .Y(_1517_));
 sg13g2_nand2_1 _5858_ (.Y(_1518_),
    .A(net865),
    .B(_1517_));
 sg13g2_nand2_1 _5859_ (.Y(_1519_),
    .A(net877),
    .B(_1385_));
 sg13g2_nand2_1 _5860_ (.Y(_1520_),
    .A(net870),
    .B(_1385_));
 sg13g2_xor2_1 _5861_ (.B(_1520_),
    .A(_1388_),
    .X(_1521_));
 sg13g2_nand2b_1 _5862_ (.Y(_1522_),
    .B(_1521_),
    .A_N(_1518_));
 sg13g2_xnor2_1 _5863_ (.Y(_1523_),
    .A(_1518_),
    .B(_1521_));
 sg13g2_a21o_1 _5864_ (.A2(_1512_),
    .A1(_1348_),
    .B1(_1511_),
    .X(_1524_));
 sg13g2_nand3_1 _5865_ (.B(_1523_),
    .C(_1524_),
    .A(_1513_),
    .Y(_1525_));
 sg13g2_nand2_1 _5866_ (.Y(_1526_),
    .A(_1513_),
    .B(_1525_));
 sg13g2_xor2_1 _5867_ (.B(_1394_),
    .A(_1393_),
    .X(_1527_));
 sg13g2_nand2_1 _5868_ (.Y(_1528_),
    .A(_1526_),
    .B(_1527_));
 sg13g2_o21ai_1 _5869_ (.B1(_1522_),
    .Y(_1529_),
    .A1(_1388_),
    .A2(_1520_));
 sg13g2_inv_1 _5870_ (.Y(_1530_),
    .A(_1529_));
 sg13g2_xnor2_1 _5871_ (.Y(_1531_),
    .A(_1526_),
    .B(_1527_));
 sg13g2_o21ai_1 _5872_ (.B1(_1528_),
    .Y(_1532_),
    .A1(_1530_),
    .A2(_1531_));
 sg13g2_xor2_1 _5873_ (.B(_1427_),
    .A(_1426_),
    .X(_1533_));
 sg13g2_nand2b_1 _5874_ (.Y(_1534_),
    .B(_1532_),
    .A_N(_1533_));
 sg13g2_nand2_1 _5875_ (.Y(_1535_),
    .A(net856),
    .B(_1385_));
 sg13g2_xor2_1 _5876_ (.B(_1533_),
    .A(_1532_),
    .X(_1536_));
 sg13g2_o21ai_1 _5877_ (.B1(_1534_),
    .Y(_1537_),
    .A1(_1535_),
    .A2(_1536_));
 sg13g2_xnor2_1 _5878_ (.Y(_1538_),
    .A(_1464_),
    .B(_1465_));
 sg13g2_nor2_1 _5879_ (.A(_1537_),
    .B(_1538_),
    .Y(_1539_));
 sg13g2_xnor2_1 _5880_ (.Y(_1540_),
    .A(_1535_),
    .B(_1536_));
 sg13g2_nand2_1 _5881_ (.Y(_1541_),
    .A(net856),
    .B(_1517_));
 sg13g2_and2_1 _5882_ (.A(net813),
    .B(_1387_),
    .X(_1542_));
 sg13g2_nand2_1 _5883_ (.Y(_1543_),
    .A(net886),
    .B(_1387_));
 sg13g2_nand2_1 _5884_ (.Y(_1544_),
    .A(net881),
    .B(_1385_));
 sg13g2_xnor2_1 _5885_ (.Y(_1545_),
    .A(_1504_),
    .B(_1543_));
 sg13g2_nor2_1 _5886_ (.A(_1544_),
    .B(_1545_),
    .Y(_1546_));
 sg13g2_a21oi_1 _5887_ (.A1(_1506_),
    .A2(_1542_),
    .Y(_1547_),
    .B1(_1546_));
 sg13g2_xnor2_1 _5888_ (.Y(_1548_),
    .A(_1508_),
    .B(_1510_));
 sg13g2_nor2b_1 _5889_ (.A(_1547_),
    .B_N(_1548_),
    .Y(_1549_));
 sg13g2_xnor2_1 _5890_ (.Y(_1550_),
    .A(_1055_),
    .B(_1166_));
 sg13g2_nor2_2 _5891_ (.A(_1156_),
    .B(_1550_),
    .Y(_1551_));
 sg13g2_nor3_2 _5892_ (.A(_2407_),
    .B(_1156_),
    .C(_1550_),
    .Y(_1552_));
 sg13g2_nor3_2 _5893_ (.A(_2427_),
    .B(_1515_),
    .C(_1516_),
    .Y(_1553_));
 sg13g2_nand2_1 _5894_ (.Y(_1554_),
    .A(net870),
    .B(_1517_));
 sg13g2_nor2_1 _5895_ (.A(_1519_),
    .B(_1554_),
    .Y(_1555_));
 sg13g2_xor2_1 _5896_ (.B(_1554_),
    .A(_1519_),
    .X(_1556_));
 sg13g2_xnor2_1 _5897_ (.Y(_1557_),
    .A(_1552_),
    .B(_1556_));
 sg13g2_inv_1 _5898_ (.Y(_1558_),
    .A(_1557_));
 sg13g2_xnor2_1 _5899_ (.Y(_1559_),
    .A(_1547_),
    .B(_1548_));
 sg13g2_a21o_1 _5900_ (.A2(_1559_),
    .A1(_1558_),
    .B1(_1549_),
    .X(_1560_));
 sg13g2_a21o_1 _5901_ (.A2(_1524_),
    .A1(_1513_),
    .B1(_1523_),
    .X(_1561_));
 sg13g2_nand3_1 _5902_ (.B(_1560_),
    .C(_1561_),
    .A(_1525_),
    .Y(_1562_));
 sg13g2_a21oi_1 _5903_ (.A1(_1552_),
    .A2(_1556_),
    .Y(_1563_),
    .B1(_1555_));
 sg13g2_inv_1 _5904_ (.Y(_1564_),
    .A(_1563_));
 sg13g2_a21o_1 _5905_ (.A2(_1561_),
    .A1(_1525_),
    .B1(_1560_),
    .X(_1565_));
 sg13g2_nand3_1 _5906_ (.B(_1564_),
    .C(_1565_),
    .A(_1562_),
    .Y(_1566_));
 sg13g2_nand2_1 _5907_ (.Y(_1567_),
    .A(_1562_),
    .B(_1566_));
 sg13g2_xnor2_1 _5908_ (.Y(_1568_),
    .A(_1530_),
    .B(_1531_));
 sg13g2_nor2b_1 _5909_ (.A(_1568_),
    .B_N(_1567_),
    .Y(_1569_));
 sg13g2_xor2_1 _5910_ (.B(_1568_),
    .A(_1567_),
    .X(_1570_));
 sg13g2_nor2_1 _5911_ (.A(_1541_),
    .B(_1570_),
    .Y(_1571_));
 sg13g2_xnor2_1 _5912_ (.Y(_1572_),
    .A(_1541_),
    .B(_1570_));
 sg13g2_and2_1 _5913_ (.A(net887),
    .B(_1385_),
    .X(_1573_));
 sg13g2_nand2_1 _5914_ (.Y(_1574_),
    .A(net881),
    .B(_1517_));
 sg13g2_xnor2_1 _5915_ (.Y(_1575_),
    .A(_1542_),
    .B(_1573_));
 sg13g2_nor2_1 _5916_ (.A(_1574_),
    .B(_1575_),
    .Y(_1576_));
 sg13g2_a21oi_1 _5917_ (.A1(_1542_),
    .A2(_1573_),
    .Y(_1577_),
    .B1(_1576_));
 sg13g2_xnor2_1 _5918_ (.Y(_1578_),
    .A(_1544_),
    .B(_1545_));
 sg13g2_nor2_1 _5919_ (.A(_1577_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_nand2_1 _5920_ (.Y(_1580_),
    .A(net865),
    .B(net705));
 sg13g2_nand3_1 _5921_ (.B(_1551_),
    .C(_1553_),
    .A(net872),
    .Y(_1581_));
 sg13g2_inv_1 _5922_ (.Y(_1582_),
    .A(_1581_));
 sg13g2_a21oi_1 _5923_ (.A1(net872),
    .A2(_1551_),
    .Y(_1583_),
    .B1(_1553_));
 sg13g2_o21ai_1 _5924_ (.B1(_1580_),
    .Y(_1584_),
    .A1(_1582_),
    .A2(_1583_));
 sg13g2_xor2_1 _5925_ (.B(_1578_),
    .A(_1577_),
    .X(_1585_));
 sg13g2_a21oi_1 _5926_ (.A1(_1584_),
    .A2(_1585_),
    .Y(_1586_),
    .B1(_1579_));
 sg13g2_xnor2_1 _5927_ (.Y(_1587_),
    .A(_1557_),
    .B(_1559_));
 sg13g2_nor2b_1 _5928_ (.A(_1586_),
    .B_N(_1587_),
    .Y(_1588_));
 sg13g2_xnor2_1 _5929_ (.Y(_1589_),
    .A(_1586_),
    .B(_1587_));
 sg13g2_a21o_1 _5930_ (.A2(_1589_),
    .A1(_1582_),
    .B1(_1588_),
    .X(_1590_));
 sg13g2_a21o_1 _5931_ (.A2(_1565_),
    .A1(_1562_),
    .B1(_1564_),
    .X(_1591_));
 sg13g2_and2_1 _5932_ (.A(_1566_),
    .B(_1591_),
    .X(_1592_));
 sg13g2_and3_1 _5933_ (.X(_1593_),
    .A(_1566_),
    .B(_1590_),
    .C(_1591_));
 sg13g2_nand2_1 _5934_ (.Y(_1594_),
    .A(net857),
    .B(net710));
 sg13g2_nand2_1 _5935_ (.Y(_1595_),
    .A(net855),
    .B(_1551_));
 sg13g2_a21oi_1 _5936_ (.A1(_1566_),
    .A2(_1591_),
    .Y(_1596_),
    .B1(_1590_));
 sg13g2_nor3_1 _5937_ (.A(_1593_),
    .B(_1595_),
    .C(_1596_),
    .Y(_1597_));
 sg13g2_or3_1 _5938_ (.A(_1593_),
    .B(_1595_),
    .C(_1596_),
    .X(_1598_));
 sg13g2_o21ai_1 _5939_ (.B1(_1595_),
    .Y(_1599_),
    .A1(_1593_),
    .A2(_1596_));
 sg13g2_xnor2_1 _5940_ (.Y(_1600_),
    .A(_1581_),
    .B(_1589_));
 sg13g2_xnor2_1 _5941_ (.Y(_1601_),
    .A(_1584_),
    .B(_1585_));
 sg13g2_nor3_2 _5942_ (.A(net892),
    .B(net705),
    .C(_1516_),
    .Y(_1602_));
 sg13g2_nand2_1 _5943_ (.Y(_1603_),
    .A(net881),
    .B(_1551_));
 sg13g2_a22oi_1 _5944_ (.Y(_1604_),
    .B1(_1517_),
    .B2(net887),
    .A2(_1385_),
    .A1(net812));
 sg13g2_a21o_1 _5945_ (.A2(_1602_),
    .A1(_1573_),
    .B1(_1604_),
    .X(_1605_));
 sg13g2_nor2_1 _5946_ (.A(_1603_),
    .B(_1605_),
    .Y(_1606_));
 sg13g2_a21oi_1 _5947_ (.A1(_1573_),
    .A2(_1602_),
    .Y(_1607_),
    .B1(_1606_));
 sg13g2_xor2_1 _5948_ (.B(_1575_),
    .A(_1574_),
    .X(_1608_));
 sg13g2_nor2b_1 _5949_ (.A(_1607_),
    .B_N(_1608_),
    .Y(_1609_));
 sg13g2_nand2_1 _5950_ (.Y(_1610_),
    .A(net872),
    .B(net705));
 sg13g2_nand2_1 _5951_ (.Y(_1611_),
    .A(net877),
    .B(net710));
 sg13g2_o21ai_1 _5952_ (.B1(_1610_),
    .Y(_1612_),
    .A1(_1550_),
    .A2(_1611_));
 sg13g2_xnor2_1 _5953_ (.Y(_1613_),
    .A(_1607_),
    .B(_1608_));
 sg13g2_a21o_1 _5954_ (.A2(_1613_),
    .A1(_1612_),
    .B1(_1609_),
    .X(_1614_));
 sg13g2_nor2b_1 _5955_ (.A(_1601_),
    .B_N(_1614_),
    .Y(_1615_));
 sg13g2_xor2_1 _5956_ (.B(_1614_),
    .A(_1601_),
    .X(_1616_));
 sg13g2_nand3_1 _5957_ (.B(_1551_),
    .C(_1602_),
    .A(net887),
    .Y(_1617_));
 sg13g2_inv_1 _5958_ (.Y(_1618_),
    .A(_1617_));
 sg13g2_xor2_1 _5959_ (.B(_1605_),
    .A(_1603_),
    .X(_1619_));
 sg13g2_a22oi_1 _5960_ (.Y(_1620_),
    .B1(net705),
    .B2(net877),
    .A2(net710),
    .A1(net865));
 sg13g2_xnor2_1 _5961_ (.Y(_1621_),
    .A(_1618_),
    .B(_1619_));
 sg13g2_nor2_1 _5962_ (.A(_1620_),
    .B(_1621_),
    .Y(_1622_));
 sg13g2_a21oi_1 _5963_ (.A1(_1618_),
    .A2(_1619_),
    .Y(_1623_),
    .B1(_1622_));
 sg13g2_xnor2_1 _5964_ (.Y(_1624_),
    .A(_1612_),
    .B(_1613_));
 sg13g2_nor2_1 _5965_ (.A(_1623_),
    .B(_1624_),
    .Y(_1625_));
 sg13g2_a21o_1 _5966_ (.A2(_1551_),
    .A1(net887),
    .B1(_1602_),
    .X(_1626_));
 sg13g2_a22oi_1 _5967_ (.Y(_1627_),
    .B1(_1617_),
    .B2(_1626_),
    .A2(net705),
    .A1(net883));
 sg13g2_nor3_1 _5968_ (.A(net818),
    .B(_1156_),
    .C(_1627_),
    .Y(_1628_));
 sg13g2_nand4_1 _5969_ (.B(net813),
    .C(net710),
    .A(net877),
    .Y(_1629_),
    .D(_1551_));
 sg13g2_a21oi_1 _5970_ (.A1(net818),
    .A2(_1627_),
    .Y(_1630_),
    .B1(_1629_));
 sg13g2_nor2_1 _5971_ (.A(_1628_),
    .B(_1630_),
    .Y(_1631_));
 sg13g2_xnor2_1 _5972_ (.Y(_1632_),
    .A(_1620_),
    .B(_1621_));
 sg13g2_nor3_1 _5973_ (.A(_1594_),
    .B(_1631_),
    .C(_1632_),
    .Y(_1633_));
 sg13g2_nand2_1 _5974_ (.Y(_1634_),
    .A(_1625_),
    .B(_1633_));
 sg13g2_o21ai_1 _5975_ (.B1(_1594_),
    .Y(_1635_),
    .A1(_1631_),
    .A2(_1632_));
 sg13g2_nand3b_1 _5976_ (.B(_1623_),
    .C(_1624_),
    .Y(_1636_),
    .A_N(_1633_));
 sg13g2_o21ai_1 _5977_ (.B1(_1636_),
    .Y(_1637_),
    .A1(_1625_),
    .A2(_1635_));
 sg13g2_a21oi_1 _5978_ (.A1(_1616_),
    .A2(_1634_),
    .Y(_1638_),
    .B1(_1637_));
 sg13g2_nand3_1 _5979_ (.B(net705),
    .C(_1638_),
    .A(net857),
    .Y(_1639_));
 sg13g2_nor2_1 _5980_ (.A(_1600_),
    .B(_1615_),
    .Y(_1640_));
 sg13g2_a221oi_1 _5981_ (.B2(_1615_),
    .C1(_1638_),
    .B1(_1600_),
    .A1(net857),
    .Y(_1641_),
    .A2(net705));
 sg13g2_a21oi_1 _5982_ (.A1(_1639_),
    .A2(_1640_),
    .Y(_1642_),
    .B1(_1641_));
 sg13g2_nand4_1 _5983_ (.B(_1598_),
    .C(_1599_),
    .A(_1593_),
    .Y(_1643_),
    .D(_1642_));
 sg13g2_a221oi_1 _5984_ (.B2(_1642_),
    .C1(_1597_),
    .B1(_1599_),
    .A1(_1590_),
    .Y(_1644_),
    .A2(_1592_));
 sg13g2_a21o_1 _5985_ (.A2(_1643_),
    .A1(_1572_),
    .B1(_1644_),
    .X(_1645_));
 sg13g2_nor2_1 _5986_ (.A(_1569_),
    .B(_1571_),
    .Y(_1646_));
 sg13g2_nand2_1 _5987_ (.Y(_1647_),
    .A(_1540_),
    .B(_1646_));
 sg13g2_o21ai_1 _5988_ (.B1(_1645_),
    .Y(_1648_),
    .A1(_1540_),
    .A2(_1646_));
 sg13g2_a22oi_1 _5989_ (.Y(_1649_),
    .B1(_1647_),
    .B2(_1648_),
    .A2(_1538_),
    .A1(_1537_));
 sg13g2_or2_1 _5990_ (.X(_1650_),
    .B(_1649_),
    .A(_1539_));
 sg13g2_o21ai_1 _5991_ (.B1(_1502_),
    .Y(_1651_),
    .A1(_1539_),
    .A2(_1649_));
 sg13g2_a21oi_1 _5992_ (.A1(_1469_),
    .A2(_1496_),
    .Y(_1652_),
    .B1(_1495_));
 sg13g2_a21oi_1 _5993_ (.A1(_1472_),
    .A2(_1476_),
    .Y(_1653_),
    .B1(_1474_));
 sg13g2_a21oi_2 _5994_ (.B1(_1492_),
    .Y(_1654_),
    .A2(_1493_),
    .A1(_1477_));
 sg13g2_o21ai_1 _5995_ (.B1(_1488_),
    .Y(_1655_),
    .A1(_1479_),
    .A2(_1489_));
 sg13g2_nand2_1 _5996_ (.Y(_1656_),
    .A(net882),
    .B(_1446_));
 sg13g2_nand2_1 _5997_ (.Y(_1657_),
    .A(_1441_),
    .B(_1482_));
 sg13g2_a221oi_1 _5998_ (.B2(_1376_),
    .C1(_1657_),
    .B1(_1443_),
    .A1(_1405_),
    .Y(_1658_),
    .A2(_1412_));
 sg13g2_a21oi_1 _5999_ (.A1(_1440_),
    .A2(_1482_),
    .Y(_1659_),
    .B1(_1481_));
 sg13g2_inv_1 _6000_ (.Y(_1660_),
    .A(_1659_));
 sg13g2_nor2_1 _6001_ (.A(_1257_),
    .B(_1435_),
    .Y(_1661_));
 sg13g2_o21ai_1 _6002_ (.B1(_1661_),
    .Y(_1662_),
    .A1(_1660_),
    .A2(_1658_));
 sg13g2_or3_1 _6003_ (.A(_1658_),
    .B(_1660_),
    .C(_1661_),
    .X(_1663_));
 sg13g2_and2_1 _6004_ (.A(net704),
    .B(_1663_),
    .X(_1664_));
 sg13g2_nand2_1 _6005_ (.Y(_1665_),
    .A(net704),
    .B(_1663_));
 sg13g2_nand3_1 _6006_ (.B(_1662_),
    .C(_1663_),
    .A(net888),
    .Y(_1666_));
 sg13g2_nand3_1 _6007_ (.B(net704),
    .C(_1663_),
    .A(net812),
    .Y(_1667_));
 sg13g2_or2_1 _6008_ (.X(_1668_),
    .B(_1666_),
    .A(_1487_));
 sg13g2_xnor2_1 _6009_ (.Y(_1669_),
    .A(_1486_),
    .B(_1667_));
 sg13g2_xor2_1 _6010_ (.B(_1669_),
    .A(_1656_),
    .X(_1670_));
 sg13g2_and2_1 _6011_ (.A(_1655_),
    .B(_1670_),
    .X(_1671_));
 sg13g2_or2_1 _6012_ (.X(_1672_),
    .B(_1670_),
    .A(_1655_));
 sg13g2_xnor2_1 _6013_ (.Y(_1673_),
    .A(_1655_),
    .B(_1670_));
 sg13g2_nand2_1 _6014_ (.Y(_1674_),
    .A(net864),
    .B(_1340_));
 sg13g2_nand2_1 _6015_ (.Y(_1675_),
    .A(net870),
    .B(_1417_));
 sg13g2_nand2_1 _6016_ (.Y(_1676_),
    .A(net876),
    .B(_1417_));
 sg13g2_xor2_1 _6017_ (.B(_1676_),
    .A(_1473_),
    .X(_1677_));
 sg13g2_nand2b_1 _6018_ (.Y(_1678_),
    .B(_1677_),
    .A_N(_1674_));
 sg13g2_xnor2_1 _6019_ (.Y(_1679_),
    .A(_1674_),
    .B(_1677_));
 sg13g2_xnor2_1 _6020_ (.Y(_1680_),
    .A(_1673_),
    .B(_1679_));
 sg13g2_nand2b_1 _6021_ (.Y(_1681_),
    .B(_1680_),
    .A_N(_1654_));
 sg13g2_nor2b_1 _6022_ (.A(_1680_),
    .B_N(_1654_),
    .Y(_1682_));
 sg13g2_xnor2_1 _6023_ (.Y(_1683_),
    .A(_1654_),
    .B(_1680_));
 sg13g2_xnor2_1 _6024_ (.Y(_1684_),
    .A(_1653_),
    .B(_1683_));
 sg13g2_nor2b_1 _6025_ (.A(_1652_),
    .B_N(_1684_),
    .Y(_1685_));
 sg13g2_nand2_1 _6026_ (.Y(_1686_),
    .A(net856),
    .B(_1342_));
 sg13g2_inv_1 _6027_ (.Y(_1687_),
    .A(_1686_));
 sg13g2_xnor2_1 _6028_ (.Y(_1688_),
    .A(_1652_),
    .B(_1684_));
 sg13g2_a21oi_1 _6029_ (.A1(_1687_),
    .A2(_1688_),
    .Y(_1689_),
    .B1(_1685_));
 sg13g2_nand2_1 _6030_ (.Y(_1690_),
    .A(net855),
    .B(_1340_));
 sg13g2_o21ai_1 _6031_ (.B1(_1681_),
    .Y(_1691_),
    .A1(_1653_),
    .A2(_1682_));
 sg13g2_o21ai_1 _6032_ (.B1(_1678_),
    .Y(_1692_),
    .A1(_1473_),
    .A2(_1676_));
 sg13g2_a21oi_1 _6033_ (.A1(_1672_),
    .A2(_1679_),
    .Y(_1693_),
    .B1(_1671_));
 sg13g2_nand2_1 _6034_ (.Y(_1694_),
    .A(net864),
    .B(_1378_));
 sg13g2_nand2_1 _6035_ (.Y(_1695_),
    .A(net870),
    .B(_1446_));
 sg13g2_nand2_1 _6036_ (.Y(_1696_),
    .A(net876),
    .B(_1446_));
 sg13g2_xor2_1 _6037_ (.B(_1696_),
    .A(_1675_),
    .X(_1697_));
 sg13g2_nand2b_1 _6038_ (.Y(_1698_),
    .B(_1697_),
    .A_N(_1694_));
 sg13g2_xnor2_1 _6039_ (.Y(_1699_),
    .A(_1694_),
    .B(_1697_));
 sg13g2_inv_1 _6040_ (.Y(_1700_),
    .A(_1699_));
 sg13g2_o21ai_1 _6041_ (.B1(_1668_),
    .Y(_1701_),
    .A1(_1669_),
    .A2(_1656_));
 sg13g2_nand2_1 _6042_ (.Y(_1702_),
    .A(net882),
    .B(_1485_));
 sg13g2_nand2_1 _6043_ (.Y(_1703_),
    .A(_1359_),
    .B(net704));
 sg13g2_a21oi_1 _6044_ (.A1(_1359_),
    .A2(net704),
    .Y(_1704_),
    .B1(_2445_));
 sg13g2_a21oi_2 _6045_ (.B1(net892),
    .Y(_1705_),
    .A2(_1662_),
    .A1(_1359_));
 sg13g2_nand2b_1 _6046_ (.Y(_1706_),
    .B(_1705_),
    .A_N(_1666_));
 sg13g2_a21oi_1 _6047_ (.A1(net888),
    .A2(_1664_),
    .Y(_1707_),
    .B1(_1705_));
 sg13g2_xnor2_1 _6048_ (.Y(_1708_),
    .A(_1666_),
    .B(_1705_));
 sg13g2_xnor2_1 _6049_ (.Y(_1709_),
    .A(_1702_),
    .B(_1708_));
 sg13g2_xnor2_1 _6050_ (.Y(_1710_),
    .A(_1701_),
    .B(_1709_));
 sg13g2_nor2_1 _6051_ (.A(_1700_),
    .B(_1710_),
    .Y(_1711_));
 sg13g2_xnor2_1 _6052_ (.Y(_1712_),
    .A(_1700_),
    .B(_1710_));
 sg13g2_nor2_1 _6053_ (.A(_1693_),
    .B(_1712_),
    .Y(_1713_));
 sg13g2_xor2_1 _6054_ (.B(_1693_),
    .A(_1712_),
    .X(_1714_));
 sg13g2_xnor2_1 _6055_ (.Y(_1715_),
    .A(_1692_),
    .B(_1714_));
 sg13g2_nand2b_1 _6056_ (.Y(_1716_),
    .B(_1691_),
    .A_N(_1715_));
 sg13g2_xor2_1 _6057_ (.B(_1715_),
    .A(_1691_),
    .X(_1717_));
 sg13g2_xor2_1 _6058_ (.B(_1717_),
    .A(_1690_),
    .X(_1718_));
 sg13g2_nand2b_1 _6059_ (.Y(_1719_),
    .B(_1718_),
    .A_N(_1689_));
 sg13g2_nor2b_1 _6060_ (.A(_1718_),
    .B_N(_1689_),
    .Y(_1720_));
 sg13g2_inv_1 _6061_ (.Y(_1721_),
    .A(_1720_));
 sg13g2_xnor2_1 _6062_ (.Y(_1722_),
    .A(_1689_),
    .B(_1718_));
 sg13g2_nand2_1 _6063_ (.Y(_1723_),
    .A(_1719_),
    .B(_1721_));
 sg13g2_xnor2_1 _6064_ (.Y(_1724_),
    .A(_1686_),
    .B(_1688_));
 sg13g2_nor2_1 _6065_ (.A(_1498_),
    .B(_1500_),
    .Y(_1725_));
 sg13g2_o21ai_1 _6066_ (.B1(_1724_),
    .Y(_1726_),
    .A1(_1498_),
    .A2(_1500_));
 sg13g2_inv_1 _6067_ (.Y(_1727_),
    .A(_1726_));
 sg13g2_xnor2_1 _6068_ (.Y(_1728_),
    .A(_1724_),
    .B(_1725_));
 sg13g2_nand4_1 _6069_ (.B(_1651_),
    .C(_1503_),
    .A(_1722_),
    .Y(_1729_),
    .D(_1728_));
 sg13g2_a21o_1 _6070_ (.A2(_1726_),
    .A1(_1719_),
    .B1(_1720_),
    .X(_1730_));
 sg13g2_o21ai_1 _6071_ (.B1(_1716_),
    .Y(_1731_),
    .A1(_1690_),
    .A2(_1717_));
 sg13g2_nand2_1 _6072_ (.Y(_1732_),
    .A(net855),
    .B(_1378_));
 sg13g2_a21oi_1 _6073_ (.A1(_1692_),
    .A2(_1714_),
    .Y(_1733_),
    .B1(_1713_));
 sg13g2_o21ai_1 _6074_ (.B1(_1698_),
    .Y(_1734_),
    .A1(_1675_),
    .A2(_1696_));
 sg13g2_a21oi_1 _6075_ (.A1(_1701_),
    .A2(_1709_),
    .Y(_1735_),
    .B1(_1711_));
 sg13g2_nand2_1 _6076_ (.Y(_1736_),
    .A(net864),
    .B(_1417_));
 sg13g2_nand2_1 _6077_ (.Y(_1737_),
    .A(net871),
    .B(_1485_));
 sg13g2_nand2_1 _6078_ (.Y(_1738_),
    .A(net876),
    .B(_1485_));
 sg13g2_xor2_1 _6079_ (.B(_1738_),
    .A(_1695_),
    .X(_1739_));
 sg13g2_nand2b_1 _6080_ (.Y(_1740_),
    .B(_1739_),
    .A_N(_1736_));
 sg13g2_xor2_1 _6081_ (.B(_1739_),
    .A(_1736_),
    .X(_1741_));
 sg13g2_o21ai_1 _6082_ (.B1(_1706_),
    .Y(_1742_),
    .A1(_1702_),
    .A2(_1707_));
 sg13g2_nor2_1 _6083_ (.A(_2437_),
    .B(_1665_),
    .Y(_1743_));
 sg13g2_nand2_1 _6084_ (.Y(_1744_),
    .A(_1704_),
    .B(_1743_));
 sg13g2_xnor2_1 _6085_ (.Y(_1745_),
    .A(_1704_),
    .B(_1743_));
 sg13g2_nor2b_1 _6086_ (.A(_1745_),
    .B_N(_1742_),
    .Y(_1746_));
 sg13g2_xor2_1 _6087_ (.B(_1745_),
    .A(_1742_),
    .X(_1747_));
 sg13g2_nor2_1 _6088_ (.A(_1741_),
    .B(_1747_),
    .Y(_1748_));
 sg13g2_xnor2_1 _6089_ (.Y(_1749_),
    .A(_1741_),
    .B(_1747_));
 sg13g2_nor2_1 _6090_ (.A(_1735_),
    .B(_1749_),
    .Y(_1750_));
 sg13g2_xor2_1 _6091_ (.B(_1749_),
    .A(_1735_),
    .X(_1751_));
 sg13g2_xnor2_1 _6092_ (.Y(_1752_),
    .A(_1734_),
    .B(_1751_));
 sg13g2_nor2_1 _6093_ (.A(_1733_),
    .B(_1752_),
    .Y(_1753_));
 sg13g2_xor2_1 _6094_ (.B(_1752_),
    .A(_1733_),
    .X(_1754_));
 sg13g2_nor2b_1 _6095_ (.A(_1732_),
    .B_N(_1754_),
    .Y(_1755_));
 sg13g2_xnor2_1 _6096_ (.Y(_1756_),
    .A(_1732_),
    .B(_1754_));
 sg13g2_nand2_1 _6097_ (.Y(_1757_),
    .A(_1731_),
    .B(_1756_));
 sg13g2_xnor2_1 _6098_ (.Y(_1758_),
    .A(_1731_),
    .B(_1756_));
 sg13g2_a21o_1 _6099_ (.A2(_1730_),
    .A1(_1729_),
    .B1(_1758_),
    .X(_1759_));
 sg13g2_nand3_1 _6100_ (.B(_1730_),
    .C(_1758_),
    .A(_1729_),
    .Y(_1760_));
 sg13g2_and2_1 _6101_ (.A(_1759_),
    .B(_1760_),
    .X(_1761_));
 sg13g2_nand2_1 _6102_ (.Y(_1762_),
    .A(net855),
    .B(_1446_));
 sg13g2_nor2_1 _6103_ (.A(_1746_),
    .B(_1748_),
    .Y(_1763_));
 sg13g2_nor2_1 _6104_ (.A(_0053_),
    .B(_1744_),
    .Y(_1764_));
 sg13g2_a21oi_1 _6105_ (.A1(_1359_),
    .A2(net704),
    .Y(_1765_),
    .B1(_0053_));
 sg13g2_mux2_1 _6106_ (.A0(_0053_),
    .A1(_1765_),
    .S(_1744_),
    .X(_1766_));
 sg13g2_nand2_1 _6107_ (.Y(_1767_),
    .A(net864),
    .B(_1446_));
 sg13g2_nand2b_1 _6108_ (.Y(_1768_),
    .B(_1664_),
    .A_N(_0032_));
 sg13g2_xor2_1 _6109_ (.B(_1768_),
    .A(_1737_),
    .X(_1769_));
 sg13g2_nand2b_1 _6110_ (.Y(_1770_),
    .B(_1769_),
    .A_N(_1767_));
 sg13g2_xnor2_1 _6111_ (.Y(_1771_),
    .A(_1767_),
    .B(_1769_));
 sg13g2_xnor2_1 _6112_ (.Y(_1772_),
    .A(_1766_),
    .B(_1771_));
 sg13g2_nor2_1 _6113_ (.A(_1763_),
    .B(_1772_),
    .Y(_1773_));
 sg13g2_o21ai_1 _6114_ (.B1(_1740_),
    .Y(_1774_),
    .A1(_1695_),
    .A2(_1738_));
 sg13g2_xor2_1 _6115_ (.B(_1772_),
    .A(_1763_),
    .X(_1775_));
 sg13g2_a21oi_1 _6116_ (.A1(_1774_),
    .A2(_1775_),
    .Y(_1776_),
    .B1(_1773_));
 sg13g2_o21ai_1 _6117_ (.B1(_1770_),
    .Y(_1777_),
    .A1(_1737_),
    .A2(_1768_));
 sg13g2_a21oi_1 _6118_ (.A1(_1766_),
    .A2(_1771_),
    .Y(_1778_),
    .B1(_1764_));
 sg13g2_nand2_1 _6119_ (.Y(_1779_),
    .A(net864),
    .B(_1485_));
 sg13g2_nor2_2 _6120_ (.A(net818),
    .B(_1665_),
    .Y(_1780_));
 sg13g2_a21oi_1 _6121_ (.A1(_1359_),
    .A2(net704),
    .Y(_1781_),
    .B1(_0032_));
 sg13g2_nand2_1 _6122_ (.Y(_1782_),
    .A(_1780_),
    .B(_1781_));
 sg13g2_xor2_1 _6123_ (.B(_1781_),
    .A(_1780_),
    .X(_1783_));
 sg13g2_nand2b_1 _6124_ (.Y(_1784_),
    .B(_1783_),
    .A_N(_1779_));
 sg13g2_xnor2_1 _6125_ (.Y(_1785_),
    .A(_1779_),
    .B(_1783_));
 sg13g2_nand2b_1 _6126_ (.Y(_1786_),
    .B(_1785_),
    .A_N(_1778_));
 sg13g2_xnor2_1 _6127_ (.Y(_1787_),
    .A(_1778_),
    .B(_1785_));
 sg13g2_nand2_1 _6128_ (.Y(_1788_),
    .A(_1777_),
    .B(_1787_));
 sg13g2_xnor2_1 _6129_ (.Y(_1789_),
    .A(_1777_),
    .B(_1787_));
 sg13g2_or2_1 _6130_ (.X(_1790_),
    .B(_1789_),
    .A(_1776_));
 sg13g2_xor2_1 _6131_ (.B(_1789_),
    .A(_1776_),
    .X(_1791_));
 sg13g2_nand2b_1 _6132_ (.Y(_1792_),
    .B(_1791_),
    .A_N(_1762_));
 sg13g2_xnor2_1 _6133_ (.Y(_1793_),
    .A(_1762_),
    .B(_1791_));
 sg13g2_a21oi_1 _6134_ (.A1(_1734_),
    .A2(_1751_),
    .Y(_1794_),
    .B1(_1750_));
 sg13g2_xnor2_1 _6135_ (.Y(_1795_),
    .A(_1774_),
    .B(_1775_));
 sg13g2_nand2_1 _6136_ (.Y(_1796_),
    .A(net855),
    .B(_1417_));
 sg13g2_xor2_1 _6137_ (.B(_1795_),
    .A(_1794_),
    .X(_1797_));
 sg13g2_nand2b_1 _6138_ (.Y(_1798_),
    .B(_1797_),
    .A_N(_1796_));
 sg13g2_o21ai_1 _6139_ (.B1(_1798_),
    .Y(_1799_),
    .A1(_1794_),
    .A2(_1795_));
 sg13g2_nand2_1 _6140_ (.Y(_1800_),
    .A(_1793_),
    .B(_1799_));
 sg13g2_xor2_1 _6141_ (.B(_1799_),
    .A(_1793_),
    .X(_1801_));
 sg13g2_nor2_1 _6142_ (.A(_1753_),
    .B(_1755_),
    .Y(_1802_));
 sg13g2_xnor2_1 _6143_ (.Y(_1803_),
    .A(_1796_),
    .B(_1797_));
 sg13g2_nor2b_1 _6144_ (.A(_1802_),
    .B_N(_1803_),
    .Y(_1804_));
 sg13g2_xnor2_1 _6145_ (.Y(_1805_),
    .A(_1802_),
    .B(_1803_));
 sg13g2_inv_1 _6146_ (.Y(_1806_),
    .A(_1805_));
 sg13g2_a21oi_2 _6147_ (.B1(_1806_),
    .Y(_1807_),
    .A2(_1759_),
    .A1(_1757_));
 sg13g2_o21ai_1 _6148_ (.B1(_1801_),
    .Y(_1808_),
    .A1(_1807_),
    .A2(_1804_));
 sg13g2_or3_1 _6149_ (.A(_1801_),
    .B(_1804_),
    .C(_1807_),
    .X(_1809_));
 sg13g2_a21o_1 _6150_ (.A2(_1809_),
    .A1(_1808_),
    .B1(net759),
    .X(_1810_));
 sg13g2_or2_1 _6151_ (.X(_1811_),
    .B(_1761_),
    .A(_3575_));
 sg13g2_nand3_1 _6152_ (.B(_1810_),
    .C(_1811_),
    .A(_3574_),
    .Y(_1812_));
 sg13g2_nor2_1 _6153_ (.A(net866),
    .B(_3193_),
    .Y(_1813_));
 sg13g2_nand3_1 _6154_ (.B(net800),
    .C(_1813_),
    .A(_3178_),
    .Y(_1814_));
 sg13g2_a21o_1 _6155_ (.A2(net800),
    .A1(net763),
    .B1(_1813_),
    .X(_1815_));
 sg13g2_a22oi_1 _6156_ (.Y(_1816_),
    .B1(_1814_),
    .B2(_1815_),
    .A2(_3165_),
    .A1(net796));
 sg13g2_nand2_1 _6157_ (.Y(_1817_),
    .A(net860),
    .B(net763));
 sg13g2_nand4_1 _6158_ (.B(_3165_),
    .C(net763),
    .A(net859),
    .Y(_1818_),
    .D(net800));
 sg13g2_or2_1 _6159_ (.X(_1819_),
    .B(_1818_),
    .A(_1816_));
 sg13g2_nand2_1 _6160_ (.Y(_1820_),
    .A(net796),
    .B(net763));
 sg13g2_nand2_1 _6161_ (.Y(_1821_),
    .A(net860),
    .B(_3209_));
 sg13g2_nor2_1 _6162_ (.A(_3193_),
    .B(_0378_),
    .Y(_1822_));
 sg13g2_nand3_1 _6163_ (.B(_3209_),
    .C(_1822_),
    .A(net859),
    .Y(_1823_));
 sg13g2_xor2_1 _6164_ (.B(_1822_),
    .A(_1821_),
    .X(_1824_));
 sg13g2_xnor2_1 _6165_ (.Y(_1825_),
    .A(_1820_),
    .B(_1824_));
 sg13g2_xnor2_1 _6166_ (.Y(_1826_),
    .A(_1814_),
    .B(_1825_));
 sg13g2_nor2_1 _6167_ (.A(_1819_),
    .B(_1826_),
    .Y(_1827_));
 sg13g2_inv_1 _6168_ (.Y(_1828_),
    .A(_1827_));
 sg13g2_nor3_2 _6169_ (.A(_2388_),
    .B(net851),
    .C(net852),
    .Y(_1829_));
 sg13g2_nor2_1 _6170_ (.A(_3516_),
    .B(_1829_),
    .Y(_1830_));
 sg13g2_or2_2 _6171_ (.X(_1831_),
    .B(_1829_),
    .A(_3516_));
 sg13g2_a21oi_1 _6172_ (.A1(_1819_),
    .A2(_1826_),
    .Y(_1832_),
    .B1(net770));
 sg13g2_nand2_2 _6173_ (.Y(_1833_),
    .A(_1828_),
    .B(_1832_));
 sg13g2_a21o_1 _6174_ (.A2(_1811_),
    .A1(_1810_),
    .B1(_3574_),
    .X(_1834_));
 sg13g2_and3_1 _6175_ (.X(_1835_),
    .A(_1812_),
    .B(_1833_),
    .C(_1834_));
 sg13g2_nand3_1 _6176_ (.B(_1833_),
    .C(_1834_),
    .A(_1812_),
    .Y(_1836_));
 sg13g2_nand2_1 _6177_ (.Y(_1837_),
    .A(_1812_),
    .B(_1836_));
 sg13g2_o21ai_1 _6178_ (.B1(_1828_),
    .Y(_1838_),
    .A1(_1814_),
    .A2(_1825_));
 sg13g2_nor2_1 _6179_ (.A(_3096_),
    .B(_3193_),
    .Y(_1839_));
 sg13g2_nand2_1 _6180_ (.Y(_1840_),
    .A(_3226_),
    .B(net801));
 sg13g2_nor2_1 _6181_ (.A(_1821_),
    .B(_1840_),
    .Y(_1841_));
 sg13g2_a22oi_1 _6182_ (.Y(_1842_),
    .B1(net801),
    .B2(_3209_),
    .A2(_3226_),
    .A1(net860));
 sg13g2_nor2_1 _6183_ (.A(_1841_),
    .B(_1842_),
    .Y(_1843_));
 sg13g2_xnor2_1 _6184_ (.Y(_1844_),
    .A(_1839_),
    .B(_1843_));
 sg13g2_o21ai_1 _6185_ (.B1(_1823_),
    .Y(_1845_),
    .A1(_1820_),
    .A2(_1824_));
 sg13g2_nand2b_1 _6186_ (.Y(_1846_),
    .B(_1845_),
    .A_N(_1844_));
 sg13g2_xnor2_1 _6187_ (.Y(_1847_),
    .A(_1844_),
    .B(_1845_));
 sg13g2_nand2_1 _6188_ (.Y(_1848_),
    .A(_1838_),
    .B(_1847_));
 sg13g2_o21ai_1 _6189_ (.B1(_1831_),
    .Y(_1849_),
    .A1(_1838_),
    .A2(_1847_));
 sg13g2_nor2b_2 _6190_ (.A(_1849_),
    .B_N(_1848_),
    .Y(_1850_));
 sg13g2_nand2b_1 _6191_ (.Y(_1851_),
    .B(_3572_),
    .A_N(_3569_));
 sg13g2_a21oi_1 _6192_ (.A1(net762),
    .A2(_3567_),
    .Y(_1852_),
    .B1(_3565_));
 sg13g2_nand2_1 _6193_ (.Y(_1853_),
    .A(net868),
    .B(net834));
 sg13g2_xor2_1 _6194_ (.B(net833),
    .A(net873),
    .X(_1854_));
 sg13g2_a22oi_1 _6195_ (.Y(_1855_),
    .B1(_0053_),
    .B2(_3528_),
    .A2(net836),
    .A1(net817));
 sg13g2_nand2b_1 _6196_ (.Y(_1856_),
    .B(_1854_),
    .A_N(_1855_));
 sg13g2_xnor2_1 _6197_ (.Y(_1857_),
    .A(_1854_),
    .B(_1855_));
 sg13g2_nand2_1 _6198_ (.Y(_1858_),
    .A(net762),
    .B(_1857_));
 sg13g2_xnor2_1 _6199_ (.Y(_1859_),
    .A(net762),
    .B(_1857_));
 sg13g2_nor2_1 _6200_ (.A(_1852_),
    .B(_1859_),
    .Y(_1860_));
 sg13g2_xor2_1 _6201_ (.B(_1859_),
    .A(_1852_),
    .X(_1861_));
 sg13g2_xor2_1 _6202_ (.B(_1861_),
    .A(_1851_),
    .X(_1862_));
 sg13g2_nand2_1 _6203_ (.Y(_1863_),
    .A(net791),
    .B(_1862_));
 sg13g2_and3_1 _6204_ (.X(_1864_),
    .A(_1757_),
    .B(_1759_),
    .C(_1806_));
 sg13g2_or3_1 _6205_ (.A(_3575_),
    .B(_1807_),
    .C(_1864_),
    .X(_1865_));
 sg13g2_nand2_1 _6206_ (.Y(_1866_),
    .A(net855),
    .B(_1485_));
 sg13g2_a21oi_1 _6207_ (.A1(_1359_),
    .A2(net704),
    .Y(_1867_),
    .B1(_2407_));
 sg13g2_nand2_1 _6208_ (.Y(_1868_),
    .A(_1780_),
    .B(_1867_));
 sg13g2_a22oi_1 _6209_ (.Y(_1869_),
    .B1(_1703_),
    .B2(net871),
    .A2(_1664_),
    .A1(net864));
 sg13g2_a21o_1 _6210_ (.A2(_1867_),
    .A1(_1780_),
    .B1(_1869_),
    .X(_1870_));
 sg13g2_a21oi_2 _6211_ (.B1(_1870_),
    .Y(_1871_),
    .A2(_1784_),
    .A1(_1782_));
 sg13g2_nand3_1 _6212_ (.B(_1784_),
    .C(_1870_),
    .A(_1782_),
    .Y(_1872_));
 sg13g2_nand2b_1 _6213_ (.Y(_1873_),
    .B(_1872_),
    .A_N(_1871_));
 sg13g2_and2_1 _6214_ (.A(_1786_),
    .B(_1788_),
    .X(_1874_));
 sg13g2_nor2_1 _6215_ (.A(_1873_),
    .B(_1874_),
    .Y(_1875_));
 sg13g2_xnor2_1 _6216_ (.Y(_1876_),
    .A(_1873_),
    .B(_1874_));
 sg13g2_nor2_1 _6217_ (.A(_1866_),
    .B(_1876_),
    .Y(_1877_));
 sg13g2_xnor2_1 _6218_ (.Y(_1878_),
    .A(_1866_),
    .B(_1876_));
 sg13g2_a21oi_2 _6219_ (.B1(_1878_),
    .Y(_1879_),
    .A2(_1792_),
    .A1(_1790_));
 sg13g2_nand3_1 _6220_ (.B(_1792_),
    .C(_1878_),
    .A(_1790_),
    .Y(_1880_));
 sg13g2_nor2b_1 _6221_ (.A(_1879_),
    .B_N(_1880_),
    .Y(_1881_));
 sg13g2_inv_1 _6222_ (.Y(_1882_),
    .A(_1881_));
 sg13g2_and3_1 _6223_ (.X(_1883_),
    .A(_1800_),
    .B(_1808_),
    .C(_1881_));
 sg13g2_a21oi_1 _6224_ (.A1(_1800_),
    .A2(_1808_),
    .Y(_1884_),
    .B1(_1881_));
 sg13g2_nor2_1 _6225_ (.A(_1800_),
    .B(_1882_),
    .Y(_1885_));
 sg13g2_or2_1 _6226_ (.X(_1886_),
    .B(_1884_),
    .A(_1883_));
 sg13g2_o21ai_1 _6227_ (.B1(net760),
    .Y(_1887_),
    .A1(_1883_),
    .A2(_1884_));
 sg13g2_a21oi_1 _6228_ (.A1(_1865_),
    .A2(_1887_),
    .Y(_1888_),
    .B1(_1863_));
 sg13g2_and3_1 _6229_ (.X(_1889_),
    .A(_1863_),
    .B(_1865_),
    .C(_1887_));
 sg13g2_or3_1 _6230_ (.A(_1850_),
    .B(_1888_),
    .C(_1889_),
    .X(_1890_));
 sg13g2_o21ai_1 _6231_ (.B1(_1850_),
    .Y(_1891_),
    .A1(_1888_),
    .A2(_1889_));
 sg13g2_nand3_1 _6232_ (.B(_1890_),
    .C(_1891_),
    .A(_1837_),
    .Y(_1892_));
 sg13g2_xnor2_1 _6233_ (.Y(_1893_),
    .A(_3557_),
    .B(_3558_));
 sg13g2_inv_1 _6234_ (.Y(_1894_),
    .A(_1893_));
 sg13g2_xnor2_1 _6235_ (.Y(_1895_),
    .A(_3552_),
    .B(_3556_));
 sg13g2_inv_2 _6236_ (.Y(_1896_),
    .A(_1895_));
 sg13g2_nand2_1 _6237_ (.Y(_1897_),
    .A(net800),
    .B(_1896_));
 sg13g2_nor3_1 _6238_ (.A(net866),
    .B(_1893_),
    .C(_1897_),
    .Y(_1898_));
 sg13g2_inv_1 _6239_ (.Y(_1899_),
    .A(_1898_));
 sg13g2_nor2_1 _6240_ (.A(_3096_),
    .B(_1895_),
    .Y(_1900_));
 sg13g2_nand2_1 _6241_ (.Y(_1901_),
    .A(net859),
    .B(_3573_));
 sg13g2_nor2_1 _6242_ (.A(_0378_),
    .B(_1893_),
    .Y(_1902_));
 sg13g2_nor2b_1 _6243_ (.A(_1901_),
    .B_N(_1902_),
    .Y(_1903_));
 sg13g2_xnor2_1 _6244_ (.Y(_1904_),
    .A(_1901_),
    .B(_1902_));
 sg13g2_xnor2_1 _6245_ (.Y(_1905_),
    .A(_1900_),
    .B(_1904_));
 sg13g2_and2_1 _6246_ (.A(net859),
    .B(_1896_),
    .X(_1906_));
 sg13g2_xor2_1 _6247_ (.B(_3555_),
    .A(_3554_),
    .X(_1907_));
 sg13g2_inv_1 _6248_ (.Y(_1908_),
    .A(_1907_));
 sg13g2_nand3_1 _6249_ (.B(_1906_),
    .C(_1907_),
    .A(net800),
    .Y(_1909_));
 sg13g2_inv_1 _6250_ (.Y(_1910_),
    .A(_1909_));
 sg13g2_o21ai_1 _6251_ (.B1(_1897_),
    .Y(_1911_),
    .A1(net866),
    .A2(_1893_));
 sg13g2_a22oi_1 _6252_ (.Y(_1912_),
    .B1(_1911_),
    .B2(_1899_),
    .A2(_1907_),
    .A1(net796));
 sg13g2_nand2b_1 _6253_ (.Y(_1913_),
    .B(_1910_),
    .A_N(_1912_));
 sg13g2_xnor2_1 _6254_ (.Y(_1914_),
    .A(_1899_),
    .B(_1905_));
 sg13g2_or2_1 _6255_ (.X(_1915_),
    .B(_1914_),
    .A(_1913_));
 sg13g2_o21ai_1 _6256_ (.B1(_1915_),
    .Y(_1916_),
    .A1(_1899_),
    .A2(_1905_));
 sg13g2_nor2_1 _6257_ (.A(_3096_),
    .B(_1893_),
    .Y(_1917_));
 sg13g2_nand2_1 _6258_ (.Y(_1918_),
    .A(net800),
    .B(_1862_));
 sg13g2_nand2_1 _6259_ (.Y(_1919_),
    .A(net859),
    .B(_1862_));
 sg13g2_nand2_1 _6260_ (.Y(_1920_),
    .A(_3573_),
    .B(net800));
 sg13g2_xor2_1 _6261_ (.B(_1920_),
    .A(_1919_),
    .X(_1921_));
 sg13g2_nand2_1 _6262_ (.Y(_1922_),
    .A(_1917_),
    .B(_1921_));
 sg13g2_xnor2_1 _6263_ (.Y(_1923_),
    .A(_1917_),
    .B(_1921_));
 sg13g2_a21o_1 _6264_ (.A2(_1904_),
    .A1(_1900_),
    .B1(_1903_),
    .X(_1924_));
 sg13g2_nor2b_1 _6265_ (.A(_1923_),
    .B_N(_1924_),
    .Y(_1925_));
 sg13g2_xnor2_1 _6266_ (.Y(_1926_),
    .A(_1923_),
    .B(_1924_));
 sg13g2_nor2_1 _6267_ (.A(_1916_),
    .B(_1926_),
    .Y(_1927_));
 sg13g2_and2_1 _6268_ (.A(_1916_),
    .B(_1926_),
    .X(_1928_));
 sg13g2_nor3_2 _6269_ (.A(net770),
    .B(_1927_),
    .C(_1928_),
    .Y(_1929_));
 sg13g2_a21o_1 _6270_ (.A2(_1891_),
    .A1(_1890_),
    .B1(_1837_),
    .X(_1930_));
 sg13g2_nand3_1 _6271_ (.B(_1929_),
    .C(_1930_),
    .A(_1892_),
    .Y(_1931_));
 sg13g2_nand2_1 _6272_ (.Y(_1932_),
    .A(_1892_),
    .B(_1931_));
 sg13g2_or2_1 _6273_ (.X(_1933_),
    .B(_1928_),
    .A(_1925_));
 sg13g2_nand2_1 _6274_ (.Y(_1934_),
    .A(net796),
    .B(_3573_));
 sg13g2_a21oi_1 _6275_ (.A1(_1851_),
    .A2(_1861_),
    .Y(_1935_),
    .B1(_1860_));
 sg13g2_and2_1 _6276_ (.A(_1856_),
    .B(_1858_),
    .X(_1936_));
 sg13g2_nand2_1 _6277_ (.Y(_1937_),
    .A(net831),
    .B(net810));
 sg13g2_xnor2_1 _6278_ (.Y(_1938_),
    .A(net832),
    .B(net810));
 sg13g2_or2_1 _6279_ (.X(_1939_),
    .B(_1938_),
    .A(_1853_));
 sg13g2_xor2_1 _6280_ (.B(_1938_),
    .A(_1853_),
    .X(_1940_));
 sg13g2_nand2_1 _6281_ (.Y(_1941_),
    .A(net762),
    .B(_1940_));
 sg13g2_xnor2_1 _6282_ (.Y(_1942_),
    .A(net761),
    .B(_1940_));
 sg13g2_or2_1 _6283_ (.X(_1943_),
    .B(_1942_),
    .A(_1936_));
 sg13g2_xnor2_1 _6284_ (.Y(_1944_),
    .A(_1936_),
    .B(_1942_));
 sg13g2_xor2_1 _6285_ (.B(_1944_),
    .A(_1935_),
    .X(_1945_));
 sg13g2_nand2_1 _6286_ (.Y(_1946_),
    .A(net801),
    .B(_1945_));
 sg13g2_nand2_1 _6287_ (.Y(_1947_),
    .A(net859),
    .B(_1945_));
 sg13g2_xor2_1 _6288_ (.B(_1947_),
    .A(_1918_),
    .X(_1948_));
 sg13g2_nand2b_1 _6289_ (.Y(_1949_),
    .B(_1948_),
    .A_N(_1934_));
 sg13g2_xnor2_1 _6290_ (.Y(_1950_),
    .A(_1934_),
    .B(_1948_));
 sg13g2_o21ai_1 _6291_ (.B1(_1922_),
    .Y(_1951_),
    .A1(_1919_),
    .A2(_1920_));
 sg13g2_xor2_1 _6292_ (.B(_1951_),
    .A(_1950_),
    .X(_1952_));
 sg13g2_and2_1 _6293_ (.A(_1933_),
    .B(_1952_),
    .X(_1953_));
 sg13g2_nor2_1 _6294_ (.A(net770),
    .B(_1953_),
    .Y(_1954_));
 sg13g2_o21ai_1 _6295_ (.B1(_1954_),
    .Y(_1955_),
    .A1(_1933_),
    .A2(_1952_));
 sg13g2_inv_1 _6296_ (.Y(_1956_),
    .A(_1955_));
 sg13g2_nor2b_1 _6297_ (.A(_1888_),
    .B_N(_1890_),
    .Y(_1957_));
 sg13g2_nand2_1 _6298_ (.Y(_1958_),
    .A(net796),
    .B(_3209_));
 sg13g2_nand2_1 _6299_ (.Y(_1959_),
    .A(_3243_),
    .B(net801));
 sg13g2_nand2_1 _6300_ (.Y(_1960_),
    .A(net860),
    .B(_3243_));
 sg13g2_or2_1 _6301_ (.X(_1961_),
    .B(_1960_),
    .A(_1840_));
 sg13g2_xnor2_1 _6302_ (.Y(_1962_),
    .A(_1840_),
    .B(_1960_));
 sg13g2_xnor2_1 _6303_ (.Y(_1963_),
    .A(_1958_),
    .B(_1962_));
 sg13g2_a21oi_1 _6304_ (.A1(_1839_),
    .A2(_1843_),
    .Y(_1964_),
    .B1(_1841_));
 sg13g2_nor2_1 _6305_ (.A(_1963_),
    .B(_1964_),
    .Y(_1965_));
 sg13g2_xnor2_1 _6306_ (.Y(_1966_),
    .A(_1963_),
    .B(_1964_));
 sg13g2_and3_1 _6307_ (.X(_1967_),
    .A(_1846_),
    .B(_1848_),
    .C(_1966_));
 sg13g2_a21oi_1 _6308_ (.A1(_1846_),
    .A2(_1848_),
    .Y(_1968_),
    .B1(_1966_));
 sg13g2_nor3_2 _6309_ (.A(net770),
    .B(_1967_),
    .C(_1968_),
    .Y(_1969_));
 sg13g2_nand2_1 _6310_ (.Y(_1970_),
    .A(_3523_),
    .B(_1945_));
 sg13g2_nor2_1 _6311_ (.A(_1879_),
    .B(_1885_),
    .Y(_1971_));
 sg13g2_o21ai_1 _6312_ (.B1(_1971_),
    .Y(_1972_),
    .A1(_1882_),
    .A2(_1808_));
 sg13g2_nor2_1 _6313_ (.A(_1875_),
    .B(_1877_),
    .Y(_1973_));
 sg13g2_nand2_1 _6314_ (.Y(_1974_),
    .A(net855),
    .B(_1664_));
 sg13g2_o21ai_1 _6315_ (.B1(_1867_),
    .Y(_1975_),
    .A1(net818),
    .A2(_1665_));
 sg13g2_inv_1 _6316_ (.Y(_1976_),
    .A(_1975_));
 sg13g2_xnor2_1 _6317_ (.Y(_1977_),
    .A(_1871_),
    .B(_1976_));
 sg13g2_nor2_1 _6318_ (.A(_1974_),
    .B(_1977_),
    .Y(_1978_));
 sg13g2_xor2_1 _6319_ (.B(_1977_),
    .A(_1974_),
    .X(_1979_));
 sg13g2_o21ai_1 _6320_ (.B1(_1979_),
    .Y(_1980_),
    .A1(_1875_),
    .A2(_1877_));
 sg13g2_inv_1 _6321_ (.Y(_1981_),
    .A(_1980_));
 sg13g2_xnor2_1 _6322_ (.Y(_1982_),
    .A(_1973_),
    .B(_1979_));
 sg13g2_xnor2_1 _6323_ (.Y(_1983_),
    .A(_1972_),
    .B(_1982_));
 sg13g2_a21oi_1 _6324_ (.A1(_1808_),
    .A2(_1809_),
    .Y(_1984_),
    .B1(net760));
 sg13g2_a21o_1 _6325_ (.A2(_1983_),
    .A1(net760),
    .B1(_1984_),
    .X(_1985_));
 sg13g2_or2_1 _6326_ (.X(_1986_),
    .B(_1985_),
    .A(_1970_));
 sg13g2_xnor2_1 _6327_ (.Y(_1987_),
    .A(_1970_),
    .B(_1985_));
 sg13g2_xnor2_1 _6328_ (.Y(_1988_),
    .A(_1969_),
    .B(_1987_));
 sg13g2_nor2_1 _6329_ (.A(_1957_),
    .B(_1988_),
    .Y(_1989_));
 sg13g2_xor2_1 _6330_ (.B(_1988_),
    .A(_1957_),
    .X(_1990_));
 sg13g2_xnor2_1 _6331_ (.Y(_1991_),
    .A(_1955_),
    .B(_1990_));
 sg13g2_and2_1 _6332_ (.A(_1932_),
    .B(_1991_),
    .X(_1992_));
 sg13g2_nand2_1 _6333_ (.Y(_1993_),
    .A(_3260_),
    .B(net791));
 sg13g2_xor2_1 _6334_ (.B(_1932_),
    .A(_1991_),
    .X(_1994_));
 sg13g2_a21o_1 _6335_ (.A2(_1994_),
    .A1(_1993_),
    .B1(_1992_),
    .X(_1995_));
 sg13g2_and2_1 _6336_ (.A(_3276_),
    .B(net791),
    .X(_1996_));
 sg13g2_a21o_1 _6337_ (.A2(_1990_),
    .A1(_1956_),
    .B1(_1989_),
    .X(_1997_));
 sg13g2_a21o_1 _6338_ (.A2(_1951_),
    .A1(_1950_),
    .B1(_1953_),
    .X(_1998_));
 sg13g2_nand2_1 _6339_ (.Y(_1999_),
    .A(net796),
    .B(_1862_));
 sg13g2_o21ai_1 _6340_ (.B1(_1943_),
    .Y(_2000_),
    .A1(_1935_),
    .A2(_1944_));
 sg13g2_xnor2_1 _6341_ (.Y(_2001_),
    .A(_0024_),
    .B(net148));
 sg13g2_nor2_1 _6342_ (.A(_1937_),
    .B(_2001_),
    .Y(_2002_));
 sg13g2_xor2_1 _6343_ (.B(_2001_),
    .A(_1937_),
    .X(_2003_));
 sg13g2_xnor2_1 _6344_ (.Y(_2004_),
    .A(net761),
    .B(_2003_));
 sg13g2_a21oi_1 _6345_ (.A1(_1939_),
    .A2(_1941_),
    .Y(_2005_),
    .B1(_2004_));
 sg13g2_nand3_1 _6346_ (.B(_1941_),
    .C(_2004_),
    .A(_1939_),
    .Y(_2006_));
 sg13g2_nor2b_1 _6347_ (.A(_2005_),
    .B_N(_2006_),
    .Y(_2007_));
 sg13g2_xor2_1 _6348_ (.B(_2007_),
    .A(_2000_),
    .X(_2008_));
 sg13g2_nand2_1 _6349_ (.Y(_2009_),
    .A(net859),
    .B(_2008_));
 sg13g2_or2_1 _6350_ (.X(_2010_),
    .B(_2009_),
    .A(_1946_));
 sg13g2_xnor2_1 _6351_ (.Y(_2011_),
    .A(_1946_),
    .B(_2009_));
 sg13g2_xnor2_1 _6352_ (.Y(_2012_),
    .A(_1999_),
    .B(_2011_));
 sg13g2_o21ai_1 _6353_ (.B1(_1949_),
    .Y(_2013_),
    .A1(_1918_),
    .A2(_1947_));
 sg13g2_nor2b_1 _6354_ (.A(_2012_),
    .B_N(_2013_),
    .Y(_2014_));
 sg13g2_xnor2_1 _6355_ (.Y(_2015_),
    .A(_2012_),
    .B(_2013_));
 sg13g2_and2_1 _6356_ (.A(_1998_),
    .B(_2015_),
    .X(_2016_));
 sg13g2_o21ai_1 _6357_ (.B1(_1831_),
    .Y(_2017_),
    .A1(_1998_),
    .A2(_2015_));
 sg13g2_nor2_2 _6358_ (.A(_2016_),
    .B(_2017_),
    .Y(_2018_));
 sg13g2_o21ai_1 _6359_ (.B1(_1986_),
    .Y(_2019_),
    .A1(_1969_),
    .A2(_1987_));
 sg13g2_nor2_1 _6360_ (.A(_1965_),
    .B(_1968_),
    .Y(_2020_));
 sg13g2_nand2_1 _6361_ (.Y(_2021_),
    .A(net796),
    .B(_3226_));
 sg13g2_nand2_1 _6362_ (.Y(_2022_),
    .A(net860),
    .B(_3260_));
 sg13g2_or2_1 _6363_ (.X(_2023_),
    .B(_2022_),
    .A(_1959_));
 sg13g2_xnor2_1 _6364_ (.Y(_2024_),
    .A(_1959_),
    .B(_2022_));
 sg13g2_xnor2_1 _6365_ (.Y(_2025_),
    .A(_2021_),
    .B(_2024_));
 sg13g2_o21ai_1 _6366_ (.B1(_1961_),
    .Y(_2026_),
    .A1(_1958_),
    .A2(_1962_));
 sg13g2_nand2b_1 _6367_ (.Y(_2027_),
    .B(_2026_),
    .A_N(_2025_));
 sg13g2_xor2_1 _6368_ (.B(_2026_),
    .A(_2025_),
    .X(_2028_));
 sg13g2_or2_1 _6369_ (.X(_2029_),
    .B(_2028_),
    .A(_2020_));
 sg13g2_a21oi_1 _6370_ (.A1(_2020_),
    .A2(_2028_),
    .Y(_2030_),
    .B1(net770));
 sg13g2_nand2_2 _6371_ (.Y(_2031_),
    .A(_2029_),
    .B(_2030_));
 sg13g2_and2_1 _6372_ (.A(_3523_),
    .B(_2008_),
    .X(_2032_));
 sg13g2_inv_1 _6373_ (.Y(_2033_),
    .A(_2032_));
 sg13g2_nand2_1 _6374_ (.Y(_2034_),
    .A(net855),
    .B(_1703_));
 sg13g2_nor2_2 _6375_ (.A(_2397_),
    .B(_1868_),
    .Y(_2035_));
 sg13g2_a21oi_2 _6376_ (.B1(_2035_),
    .Y(_2036_),
    .A2(_2034_),
    .A1(_1868_));
 sg13g2_a21oi_2 _6377_ (.B1(_1978_),
    .Y(_2037_),
    .A2(_1976_),
    .A1(_1871_));
 sg13g2_nor2b_1 _6378_ (.A(_2037_),
    .B_N(_2036_),
    .Y(_2038_));
 sg13g2_xor2_1 _6379_ (.B(_2037_),
    .A(_2036_),
    .X(_2039_));
 sg13g2_inv_1 _6380_ (.Y(_2040_),
    .A(_2039_));
 sg13g2_a21o_1 _6381_ (.A2(_1982_),
    .A1(_1972_),
    .B1(_1981_),
    .X(_2041_));
 sg13g2_nand2b_1 _6382_ (.Y(_2042_),
    .B(_2039_),
    .A_N(_2041_));
 sg13g2_and2_1 _6383_ (.A(_2040_),
    .B(_2041_),
    .X(_2043_));
 sg13g2_a21oi_1 _6384_ (.A1(_2040_),
    .A2(_2041_),
    .Y(_2044_),
    .B1(net759));
 sg13g2_xnor2_1 _6385_ (.Y(_2045_),
    .A(_2040_),
    .B(_2041_));
 sg13g2_nor2_1 _6386_ (.A(net760),
    .B(_1886_),
    .Y(_2046_));
 sg13g2_a21oi_2 _6387_ (.B1(_2046_),
    .Y(_2047_),
    .A2(_2045_),
    .A1(net760));
 sg13g2_nand2_1 _6388_ (.Y(_2048_),
    .A(_2032_),
    .B(_2047_));
 sg13g2_a221oi_1 _6389_ (.B2(_2044_),
    .C1(_2033_),
    .B1(_2042_),
    .A1(net759),
    .Y(_2049_),
    .A2(_1886_));
 sg13g2_a221oi_1 _6390_ (.B2(net760),
    .C1(_2046_),
    .B1(_2045_),
    .A1(net791),
    .Y(_2050_),
    .A2(_2008_));
 sg13g2_o21ai_1 _6391_ (.B1(_2031_),
    .Y(_2051_),
    .A1(_2049_),
    .A2(_2050_));
 sg13g2_or3_1 _6392_ (.A(_2031_),
    .B(_2049_),
    .C(_2050_),
    .X(_2052_));
 sg13g2_nand3_1 _6393_ (.B(_2051_),
    .C(_2052_),
    .A(_2019_),
    .Y(_2053_));
 sg13g2_a21o_1 _6394_ (.A2(_2052_),
    .A1(_2051_),
    .B1(_2019_),
    .X(_2054_));
 sg13g2_nand3_1 _6395_ (.B(_2053_),
    .C(_2054_),
    .A(_2018_),
    .Y(_2055_));
 sg13g2_a21o_1 _6396_ (.A2(_2054_),
    .A1(_2053_),
    .B1(_2018_),
    .X(_2056_));
 sg13g2_and3_1 _6397_ (.X(_2057_),
    .A(_1997_),
    .B(_2055_),
    .C(_2056_));
 sg13g2_a21oi_1 _6398_ (.A1(_2055_),
    .A2(_2056_),
    .Y(_2058_),
    .B1(_1997_));
 sg13g2_or3_1 _6399_ (.A(_1996_),
    .B(_2057_),
    .C(_2058_),
    .X(_2059_));
 sg13g2_o21ai_1 _6400_ (.B1(_1996_),
    .Y(_2060_),
    .A1(_2057_),
    .A2(_2058_));
 sg13g2_and3_1 _6401_ (.X(_2061_),
    .A(_1995_),
    .B(_2059_),
    .C(_2060_));
 sg13g2_nand3_1 _6402_ (.B(_2059_),
    .C(_2060_),
    .A(_1995_),
    .Y(_2062_));
 sg13g2_nor2b_1 _6403_ (.A(_1893_),
    .B_N(net792),
    .Y(_2063_));
 sg13g2_and3_1 _6404_ (.X(_2064_),
    .A(_1503_),
    .B(_1651_),
    .C(_1728_));
 sg13g2_nand3b_1 _6405_ (.B(_1722_),
    .C(_1726_),
    .Y(_2065_),
    .A_N(_2064_));
 sg13g2_o21ai_1 _6406_ (.B1(_1723_),
    .Y(_2066_),
    .A1(_1727_),
    .A2(_2064_));
 sg13g2_o21ai_1 _6407_ (.B1(net760),
    .Y(_2067_),
    .A1(_1807_),
    .A2(_1864_));
 sg13g2_nand3_1 _6408_ (.B(_2065_),
    .C(_2066_),
    .A(net759),
    .Y(_2068_));
 sg13g2_and3_1 _6409_ (.X(_2069_),
    .A(_2063_),
    .B(_2067_),
    .C(_2068_));
 sg13g2_nand3_1 _6410_ (.B(_2067_),
    .C(_2068_),
    .A(_2063_),
    .Y(_2070_));
 sg13g2_a21oi_1 _6411_ (.A1(_1816_),
    .A2(_1818_),
    .Y(_2071_),
    .B1(_1830_));
 sg13g2_nand2_2 _6412_ (.Y(_2072_),
    .A(_1819_),
    .B(_2071_));
 sg13g2_a21o_1 _6413_ (.A2(_2068_),
    .A1(_2067_),
    .B1(_2063_),
    .X(_2073_));
 sg13g2_nand3_1 _6414_ (.B(_2072_),
    .C(_2073_),
    .A(_2070_),
    .Y(_2074_));
 sg13g2_a21oi_1 _6415_ (.A1(_2072_),
    .A2(_2073_),
    .Y(_2075_),
    .B1(_2069_));
 sg13g2_a21oi_1 _6416_ (.A1(_1812_),
    .A2(_1834_),
    .Y(_2076_),
    .B1(_1833_));
 sg13g2_a21o_1 _6417_ (.A2(_1834_),
    .A1(_1812_),
    .B1(_1833_),
    .X(_2077_));
 sg13g2_nor3_1 _6418_ (.A(_1835_),
    .B(_2075_),
    .C(_2076_),
    .Y(_2078_));
 sg13g2_or3_1 _6419_ (.A(_1835_),
    .B(_2075_),
    .C(_2076_),
    .X(_2079_));
 sg13g2_a21oi_1 _6420_ (.A1(_1913_),
    .A2(_1914_),
    .Y(_2080_),
    .B1(net770));
 sg13g2_and2_1 _6421_ (.A(_1915_),
    .B(_2080_),
    .X(_2081_));
 sg13g2_inv_1 _6422_ (.Y(_2082_),
    .A(_2081_));
 sg13g2_a221oi_1 _6423_ (.B2(_1836_),
    .C1(_2069_),
    .B1(_2077_),
    .A1(_2072_),
    .Y(_2083_),
    .A2(_2073_));
 sg13g2_o21ai_1 _6424_ (.B1(_2075_),
    .Y(_2084_),
    .A1(_1835_),
    .A2(_2076_));
 sg13g2_nor3_1 _6425_ (.A(_2078_),
    .B(_2082_),
    .C(_2083_),
    .Y(_2085_));
 sg13g2_nand3_1 _6426_ (.B(_2081_),
    .C(_2084_),
    .A(_2079_),
    .Y(_2086_));
 sg13g2_nand2_1 _6427_ (.Y(_2087_),
    .A(_2079_),
    .B(_2086_));
 sg13g2_a21o_1 _6428_ (.A2(_1930_),
    .A1(_1892_),
    .B1(_1929_),
    .X(_2088_));
 sg13g2_nand3_1 _6429_ (.B(_2087_),
    .C(_2088_),
    .A(_1931_),
    .Y(_2089_));
 sg13g2_and2_1 _6430_ (.A(_3243_),
    .B(net791),
    .X(_2090_));
 sg13g2_nand2_1 _6431_ (.Y(_2091_),
    .A(_3243_),
    .B(net791));
 sg13g2_a21oi_1 _6432_ (.A1(_1931_),
    .A2(_2088_),
    .Y(_2092_),
    .B1(_2087_));
 sg13g2_a21o_1 _6433_ (.A2(_2088_),
    .A1(_1931_),
    .B1(_2087_),
    .X(_2093_));
 sg13g2_and3_1 _6434_ (.X(_2094_),
    .A(_2089_),
    .B(_2091_),
    .C(_2093_));
 sg13g2_o21ai_1 _6435_ (.B1(_2089_),
    .Y(_2095_),
    .A1(_2090_),
    .A2(_2092_));
 sg13g2_xor2_1 _6436_ (.B(_1994_),
    .A(_1993_),
    .X(_2096_));
 sg13g2_nor2_1 _6437_ (.A(_2095_),
    .B(_2096_),
    .Y(_2097_));
 sg13g2_nand2_1 _6438_ (.Y(_2098_),
    .A(net792),
    .B(_1896_));
 sg13g2_a21oi_1 _6439_ (.A1(_1503_),
    .A2(_1651_),
    .Y(_2099_),
    .B1(_1728_));
 sg13g2_o21ai_1 _6440_ (.B1(net759),
    .Y(_2100_),
    .A1(_2064_),
    .A2(_2099_));
 sg13g2_o21ai_1 _6441_ (.B1(_2100_),
    .Y(_2101_),
    .A1(_3576_),
    .A2(_1761_));
 sg13g2_and2_1 _6442_ (.A(_2098_),
    .B(_2101_),
    .X(_2102_));
 sg13g2_inv_1 _6443_ (.Y(_2103_),
    .A(_2102_));
 sg13g2_xnor2_1 _6444_ (.Y(_2104_),
    .A(_2098_),
    .B(_2101_));
 sg13g2_inv_1 _6445_ (.Y(_2105_),
    .A(_2104_));
 sg13g2_nand2_1 _6446_ (.Y(_2106_),
    .A(net792),
    .B(_1907_));
 sg13g2_and3_2 _6447_ (.X(_2107_),
    .A(net760),
    .B(_2065_),
    .C(_2066_));
 sg13g2_nand2_1 _6448_ (.Y(_2108_),
    .A(_1502_),
    .B(_1503_));
 sg13g2_xnor2_1 _6449_ (.Y(_2109_),
    .A(_1650_),
    .B(_2108_));
 sg13g2_nand2_1 _6450_ (.Y(_2110_),
    .A(net759),
    .B(_2109_));
 sg13g2_inv_2 _6451_ (.Y(_2111_),
    .A(_2110_));
 sg13g2_nor3_1 _6452_ (.A(_2106_),
    .B(_2107_),
    .C(_2111_),
    .Y(_2112_));
 sg13g2_nand3_1 _6453_ (.B(_3165_),
    .C(_1831_),
    .A(net859),
    .Y(_2113_));
 sg13g2_o21ai_1 _6454_ (.B1(_2106_),
    .Y(_2114_),
    .A1(_2107_),
    .A2(_2111_));
 sg13g2_nor2b_1 _6455_ (.A(_2112_),
    .B_N(_2114_),
    .Y(_2115_));
 sg13g2_and2_1 _6456_ (.A(_2113_),
    .B(_2115_),
    .X(_2116_));
 sg13g2_a21oi_1 _6457_ (.A1(_2113_),
    .A2(_2114_),
    .Y(_2117_),
    .B1(_2112_));
 sg13g2_a21oi_1 _6458_ (.A1(net800),
    .A2(_1907_),
    .Y(_2118_),
    .B1(_1906_));
 sg13g2_nor3_1 _6459_ (.A(net770),
    .B(_1910_),
    .C(_2118_),
    .Y(_2119_));
 sg13g2_xnor2_1 _6460_ (.Y(_2120_),
    .A(_2104_),
    .B(_2117_));
 sg13g2_nand2_1 _6461_ (.Y(_2121_),
    .A(_2119_),
    .B(_2120_));
 sg13g2_o21ai_1 _6462_ (.B1(_2121_),
    .Y(_2122_),
    .A1(_2105_),
    .A2(_2117_));
 sg13g2_nand2_1 _6463_ (.Y(_2123_),
    .A(_1831_),
    .B(_1913_));
 sg13g2_a21oi_2 _6464_ (.B1(_2123_),
    .Y(_2124_),
    .A2(_1912_),
    .A1(_1909_));
 sg13g2_inv_1 _6465_ (.Y(_2125_),
    .A(_2124_));
 sg13g2_a21o_1 _6466_ (.A2(_2073_),
    .A1(_2070_),
    .B1(_2072_),
    .X(_2126_));
 sg13g2_and3_1 _6467_ (.X(_2127_),
    .A(_2074_),
    .B(_2103_),
    .C(_2126_));
 sg13g2_nand3_1 _6468_ (.B(_2103_),
    .C(_2126_),
    .A(_2074_),
    .Y(_2128_));
 sg13g2_a21oi_1 _6469_ (.A1(_2074_),
    .A2(_2126_),
    .Y(_2129_),
    .B1(_2103_));
 sg13g2_nand3b_1 _6470_ (.B(_2124_),
    .C(_2128_),
    .Y(_2130_),
    .A_N(_2129_));
 sg13g2_o21ai_1 _6471_ (.B1(_2125_),
    .Y(_2131_),
    .A1(_2127_),
    .A2(_2129_));
 sg13g2_nand3_1 _6472_ (.B(_2130_),
    .C(_2131_),
    .A(_2122_),
    .Y(_2132_));
 sg13g2_nand2_1 _6473_ (.Y(_2133_),
    .A(_3209_),
    .B(net792));
 sg13g2_inv_1 _6474_ (.Y(_2134_),
    .A(_2133_));
 sg13g2_a21oi_1 _6475_ (.A1(_2130_),
    .A2(_2131_),
    .Y(_2135_),
    .B1(_2122_));
 sg13g2_a21o_1 _6476_ (.A2(_2131_),
    .A1(_2130_),
    .B1(_2122_),
    .X(_2136_));
 sg13g2_and3_1 _6477_ (.X(_2137_),
    .A(_2132_),
    .B(_2133_),
    .C(_2136_));
 sg13g2_o21ai_1 _6478_ (.B1(_2132_),
    .Y(_2138_),
    .A1(_2134_),
    .A2(_2135_));
 sg13g2_nand2_1 _6479_ (.Y(_2139_),
    .A(_3226_),
    .B(net792));
 sg13g2_inv_1 _6480_ (.Y(_2140_),
    .A(_2139_));
 sg13g2_and2_1 _6481_ (.A(_2128_),
    .B(_2130_),
    .X(_2141_));
 sg13g2_nand2_1 _6482_ (.Y(_2142_),
    .A(_2128_),
    .B(_2130_));
 sg13g2_a21oi_1 _6483_ (.A1(_2079_),
    .A2(_2084_),
    .Y(_2143_),
    .B1(_2081_));
 sg13g2_o21ai_1 _6484_ (.B1(_2082_),
    .Y(_2144_),
    .A1(_2078_),
    .A2(_2083_));
 sg13g2_nor3_1 _6485_ (.A(_2085_),
    .B(_2141_),
    .C(_2143_),
    .Y(_2145_));
 sg13g2_nand3_1 _6486_ (.B(_2142_),
    .C(_2144_),
    .A(_2086_),
    .Y(_2146_));
 sg13g2_a21oi_1 _6487_ (.A1(_2086_),
    .A2(_2144_),
    .Y(_2147_),
    .B1(_2142_));
 sg13g2_o21ai_1 _6488_ (.B1(_2141_),
    .Y(_2148_),
    .A1(_2085_),
    .A2(_2143_));
 sg13g2_nor3_1 _6489_ (.A(_2140_),
    .B(_2145_),
    .C(_2147_),
    .Y(_2149_));
 sg13g2_nand3_1 _6490_ (.B(_2146_),
    .C(_2148_),
    .A(_2139_),
    .Y(_2150_));
 sg13g2_a21oi_1 _6491_ (.A1(_2146_),
    .A2(_2148_),
    .Y(_2151_),
    .B1(_2139_));
 sg13g2_o21ai_1 _6492_ (.B1(_2140_),
    .Y(_2152_),
    .A1(_2145_),
    .A2(_2147_));
 sg13g2_nand3_1 _6493_ (.B(_2150_),
    .C(_2152_),
    .A(_2138_),
    .Y(_2153_));
 sg13g2_a21oi_1 _6494_ (.A1(_2132_),
    .A2(_2136_),
    .Y(_2154_),
    .B1(_2133_));
 sg13g2_o21ai_1 _6495_ (.B1(_1817_),
    .Y(_2155_),
    .A1(_3164_),
    .A2(_0378_));
 sg13g2_nand3_1 _6496_ (.B(_1831_),
    .C(_2155_),
    .A(_1818_),
    .Y(_2156_));
 sg13g2_inv_1 _6497_ (.Y(_2157_),
    .A(_2156_));
 sg13g2_nor2_1 _6498_ (.A(_2113_),
    .B(_2115_),
    .Y(_2158_));
 sg13g2_nor2_1 _6499_ (.A(_2116_),
    .B(_2158_),
    .Y(_2159_));
 sg13g2_nor3_1 _6500_ (.A(_2116_),
    .B(_2157_),
    .C(_2158_),
    .Y(_2160_));
 sg13g2_nor3_2 _6501_ (.A(net862),
    .B(net770),
    .C(_1908_),
    .Y(_2161_));
 sg13g2_o21ai_1 _6502_ (.B1(_2157_),
    .Y(_2162_),
    .A1(_2116_),
    .A2(_2158_));
 sg13g2_nand2b_1 _6503_ (.Y(_2163_),
    .B(_2162_),
    .A_N(_2160_));
 sg13g2_a21oi_1 _6504_ (.A1(_2161_),
    .A2(_2162_),
    .Y(_2164_),
    .B1(_2160_));
 sg13g2_xnor2_1 _6505_ (.Y(_2165_),
    .A(_2119_),
    .B(_2120_));
 sg13g2_nor2_1 _6506_ (.A(_2164_),
    .B(_2165_),
    .Y(_2166_));
 sg13g2_nand2_1 _6507_ (.Y(_2167_),
    .A(_3194_),
    .B(net792));
 sg13g2_xor2_1 _6508_ (.B(_2165_),
    .A(_2164_),
    .X(_2168_));
 sg13g2_a21oi_2 _6509_ (.B1(_2166_),
    .Y(_2169_),
    .A2(_2168_),
    .A1(_2167_));
 sg13g2_nor3_1 _6510_ (.A(_2137_),
    .B(_2154_),
    .C(_2169_),
    .Y(_2170_));
 sg13g2_xnor2_1 _6511_ (.Y(_2171_),
    .A(_2161_),
    .B(_2163_));
 sg13g2_nand2_1 _6512_ (.Y(_2172_),
    .A(_2156_),
    .B(_2171_));
 sg13g2_nand2_1 _6513_ (.Y(_2173_),
    .A(net763),
    .B(net792));
 sg13g2_xor2_1 _6514_ (.B(_2161_),
    .A(_2159_),
    .X(_2174_));
 sg13g2_nand2_1 _6515_ (.Y(_2175_),
    .A(_2173_),
    .B(_2174_));
 sg13g2_xnor2_1 _6516_ (.Y(_2176_),
    .A(_2167_),
    .B(_2168_));
 sg13g2_a21oi_2 _6517_ (.B1(_2176_),
    .Y(_2177_),
    .A2(_2175_),
    .A1(_2172_));
 sg13g2_o21ai_1 _6518_ (.B1(_2169_),
    .Y(_2178_),
    .A1(_2137_),
    .A2(_2154_));
 sg13g2_nor2b_1 _6519_ (.A(_2170_),
    .B_N(_2178_),
    .Y(_2179_));
 sg13g2_a21oi_2 _6520_ (.B1(_2170_),
    .Y(_2180_),
    .A2(_2178_),
    .A1(_2177_));
 sg13g2_a21oi_1 _6521_ (.A1(_2150_),
    .A2(_2152_),
    .Y(_2181_),
    .B1(_2138_));
 sg13g2_nor3_1 _6522_ (.A(_2138_),
    .B(_2149_),
    .C(_2151_),
    .Y(_2182_));
 sg13g2_o21ai_1 _6523_ (.B1(_2138_),
    .Y(_2183_),
    .A1(_2149_),
    .A2(_2151_));
 sg13g2_nand2b_1 _6524_ (.Y(_2184_),
    .B(_2183_),
    .A_N(_2182_));
 sg13g2_o21ai_1 _6525_ (.B1(_2153_),
    .Y(_2185_),
    .A1(_2180_),
    .A2(_2181_));
 sg13g2_a21oi_1 _6526_ (.A1(_2089_),
    .A2(_2093_),
    .Y(_2186_),
    .B1(_2091_));
 sg13g2_nor2_1 _6527_ (.A(_2145_),
    .B(_2149_),
    .Y(_2187_));
 sg13g2_nor3_1 _6528_ (.A(_2094_),
    .B(_2186_),
    .C(_2187_),
    .Y(_2188_));
 sg13g2_or3_1 _6529_ (.A(_2094_),
    .B(_2186_),
    .C(_2187_),
    .X(_2189_));
 sg13g2_o21ai_1 _6530_ (.B1(_2187_),
    .Y(_2190_),
    .A1(_2094_),
    .A2(_2186_));
 sg13g2_and3_1 _6531_ (.X(_2191_),
    .A(_2185_),
    .B(_2189_),
    .C(_2190_));
 sg13g2_a221oi_1 _6532_ (.B2(_2190_),
    .C1(_2188_),
    .B1(_2185_),
    .A1(_2095_),
    .Y(_2192_),
    .A2(_2096_));
 sg13g2_nor2_1 _6533_ (.A(_2097_),
    .B(_2192_),
    .Y(_2193_));
 sg13g2_a21oi_1 _6534_ (.A1(_2059_),
    .A2(_2060_),
    .Y(_2194_),
    .B1(_1995_));
 sg13g2_or2_1 _6535_ (.X(_2195_),
    .B(_2194_),
    .A(_2061_));
 sg13g2_or4_1 _6536_ (.A(_2061_),
    .B(_2097_),
    .C(_2192_),
    .D(_2194_),
    .X(_2196_));
 sg13g2_nor2b_1 _6537_ (.A(_2057_),
    .B_N(_2059_),
    .Y(_2197_));
 sg13g2_nand2_1 _6538_ (.Y(_2198_),
    .A(_3290_),
    .B(net791));
 sg13g2_nand2_1 _6539_ (.Y(_2199_),
    .A(_2053_),
    .B(_2055_));
 sg13g2_nand2_1 _6540_ (.Y(_2200_),
    .A(_2048_),
    .B(_2051_));
 sg13g2_nor4_1 _6541_ (.A(net759),
    .B(_2035_),
    .C(_2038_),
    .D(_2043_),
    .Y(_2201_));
 sg13g2_a21oi_1 _6542_ (.A1(net759),
    .A2(_1983_),
    .Y(_2202_),
    .B1(_2201_));
 sg13g2_a21oi_1 _6543_ (.A1(_2000_),
    .A2(_2007_),
    .Y(_2203_),
    .B1(_2005_));
 sg13g2_a21oi_1 _6544_ (.A1(net761),
    .A2(_2003_),
    .Y(_2204_),
    .B1(_2002_));
 sg13g2_nand2_1 _6545_ (.Y(_2205_),
    .A(net830),
    .B(net155));
 sg13g2_a21oi_1 _6546_ (.A1(net830),
    .A2(net154),
    .Y(_2206_),
    .B1(net806));
 sg13g2_xnor2_1 _6547_ (.Y(_2207_),
    .A(net826),
    .B(_2206_));
 sg13g2_nand2b_1 _6548_ (.Y(_2208_),
    .B(net761),
    .A_N(_2207_));
 sg13g2_xnor2_1 _6549_ (.Y(_2209_),
    .A(net761),
    .B(_2207_));
 sg13g2_inv_1 _6550_ (.Y(_2210_),
    .A(_2209_));
 sg13g2_xnor2_1 _6551_ (.Y(_2211_),
    .A(_2204_),
    .B(_2209_));
 sg13g2_nand2b_1 _6552_ (.Y(_2212_),
    .B(_2211_),
    .A_N(_2203_));
 sg13g2_xnor2_1 _6553_ (.Y(_2213_),
    .A(_2203_),
    .B(_2211_));
 sg13g2_nand2_1 _6554_ (.Y(_2214_),
    .A(net792),
    .B(_2213_));
 sg13g2_o21ai_1 _6555_ (.B1(_2023_),
    .Y(_2215_),
    .A1(_2021_),
    .A2(_2024_));
 sg13g2_nand2_1 _6556_ (.Y(_2216_),
    .A(_2407_),
    .B(_3276_));
 sg13g2_a22oi_1 _6557_ (.Y(_2217_),
    .B1(_3260_),
    .B2(net801),
    .A2(_3243_),
    .A1(net796));
 sg13g2_xnor2_1 _6558_ (.Y(_2218_),
    .A(_2216_),
    .B(_2217_));
 sg13g2_xor2_1 _6559_ (.B(_2218_),
    .A(_2215_),
    .X(_2219_));
 sg13g2_a21o_1 _6560_ (.A2(_2029_),
    .A1(_2027_),
    .B1(_2219_),
    .X(_2220_));
 sg13g2_nand3_1 _6561_ (.B(_2029_),
    .C(_2219_),
    .A(_2027_),
    .Y(_2221_));
 sg13g2_nand3_1 _6562_ (.B(_2220_),
    .C(_2221_),
    .A(_1831_),
    .Y(_2222_));
 sg13g2_xnor2_1 _6563_ (.Y(_2223_),
    .A(_2214_),
    .B(_2222_));
 sg13g2_o21ai_1 _6564_ (.B1(_2010_),
    .Y(_2224_),
    .A1(_1999_),
    .A2(_2011_));
 sg13g2_nand2_1 _6565_ (.Y(_2225_),
    .A(_2407_),
    .B(_2213_));
 sg13g2_a22oi_1 _6566_ (.Y(_2226_),
    .B1(_2008_),
    .B2(net801),
    .A2(_1945_),
    .A1(net797));
 sg13g2_xnor2_1 _6567_ (.Y(_2227_),
    .A(_2225_),
    .B(_2226_));
 sg13g2_xnor2_1 _6568_ (.Y(_2228_),
    .A(_2224_),
    .B(_2227_));
 sg13g2_o21ai_1 _6569_ (.B1(_2228_),
    .Y(_2229_),
    .A1(_2014_),
    .A2(_2016_));
 sg13g2_or3_1 _6570_ (.A(_2014_),
    .B(_2016_),
    .C(_2228_),
    .X(_2230_));
 sg13g2_nand3_1 _6571_ (.B(_2229_),
    .C(_2230_),
    .A(_1831_),
    .Y(_2231_));
 sg13g2_xnor2_1 _6572_ (.Y(_2232_),
    .A(_2223_),
    .B(_2231_));
 sg13g2_xnor2_1 _6573_ (.Y(_2233_),
    .A(_2202_),
    .B(_2232_));
 sg13g2_xnor2_1 _6574_ (.Y(_2234_),
    .A(_2200_),
    .B(_2233_));
 sg13g2_xnor2_1 _6575_ (.Y(_2235_),
    .A(_2199_),
    .B(_2234_));
 sg13g2_xor2_1 _6576_ (.B(_2235_),
    .A(_2198_),
    .X(_2236_));
 sg13g2_xnor2_1 _6577_ (.Y(_2237_),
    .A(_2197_),
    .B(_2236_));
 sg13g2_a21o_1 _6578_ (.A2(_2196_),
    .A1(_2062_),
    .B1(_2237_),
    .X(_2238_));
 sg13g2_nand3_1 _6579_ (.B(_2196_),
    .C(_2237_),
    .A(_2062_),
    .Y(_2239_));
 sg13g2_a21oi_1 _6580_ (.A1(_2388_),
    .A2(_3518_),
    .Y(_2240_),
    .B1(_3525_));
 sg13g2_a21o_2 _6581_ (.A2(_3518_),
    .A1(_2388_),
    .B1(_3525_),
    .X(_2241_));
 sg13g2_nand3_1 _6582_ (.B(_2239_),
    .C(_2240_),
    .A(_2238_),
    .Y(_2242_));
 sg13g2_nand2_1 _6583_ (.Y(_2243_),
    .A(net830),
    .B(_3260_));
 sg13g2_nand2_1 _6584_ (.Y(_2244_),
    .A(_0890_),
    .B(_2243_));
 sg13g2_xnor2_1 _6585_ (.Y(_2245_),
    .A(_0891_),
    .B(_2243_));
 sg13g2_nand2_1 _6586_ (.Y(_2246_),
    .A(net832),
    .B(_3243_));
 sg13g2_nor2b_1 _6587_ (.A(_0853_),
    .B_N(_2246_),
    .Y(_2247_));
 sg13g2_xor2_1 _6588_ (.B(_2246_),
    .A(_0853_),
    .X(_2248_));
 sg13g2_nand2_1 _6589_ (.Y(_2249_),
    .A(net833),
    .B(_3226_));
 sg13g2_nand2_1 _6590_ (.Y(_2250_),
    .A(net836),
    .B(_3209_));
 sg13g2_nand2_1 _6591_ (.Y(_2251_),
    .A(net714),
    .B(_2250_));
 sg13g2_xnor2_1 _6592_ (.Y(_2252_),
    .A(net714),
    .B(_2250_));
 sg13g2_nand2_1 _6593_ (.Y(_2253_),
    .A(net837),
    .B(_3194_));
 sg13g2_nand2_1 _6594_ (.Y(_2254_),
    .A(_0362_),
    .B(_2253_));
 sg13g2_nand2_1 _6595_ (.Y(_2255_),
    .A(net838),
    .B(net763));
 sg13g2_nand2_1 _6596_ (.Y(_2256_),
    .A(net720),
    .B(_2255_));
 sg13g2_nor2_1 _6597_ (.A(net720),
    .B(_2255_),
    .Y(_2257_));
 sg13g2_xor2_1 _6598_ (.B(_2255_),
    .A(net720),
    .X(_2258_));
 sg13g2_nor3_2 _6599_ (.A(_0057_),
    .B(_3164_),
    .C(_0276_),
    .Y(_2259_));
 sg13g2_o21ai_1 _6600_ (.B1(_2256_),
    .Y(_2260_),
    .A1(_2257_),
    .A2(_2259_));
 sg13g2_xnor2_1 _6601_ (.Y(_2261_),
    .A(net715),
    .B(_2253_));
 sg13g2_nand2b_1 _6602_ (.Y(_2262_),
    .B(_2260_),
    .A_N(_2261_));
 sg13g2_nand2_1 _6603_ (.Y(_2263_),
    .A(_2254_),
    .B(_2262_));
 sg13g2_nand2b_1 _6604_ (.Y(_2264_),
    .B(_2263_),
    .A_N(_2252_));
 sg13g2_xnor2_1 _6605_ (.Y(_2265_),
    .A(net713),
    .B(_2249_));
 sg13g2_a21oi_1 _6606_ (.A1(_2251_),
    .A2(_2264_),
    .Y(_2266_),
    .B1(_2265_));
 sg13g2_a21oi_1 _6607_ (.A1(net713),
    .A2(_2249_),
    .Y(_2267_),
    .B1(_2266_));
 sg13g2_nor2_1 _6608_ (.A(_2248_),
    .B(_2267_),
    .Y(_2268_));
 sg13g2_o21ai_1 _6609_ (.B1(_2245_),
    .Y(_2269_),
    .A1(_2247_),
    .A2(_2268_));
 sg13g2_nand2_1 _6610_ (.Y(_2270_),
    .A(_2244_),
    .B(_2269_));
 sg13g2_a21oi_1 _6611_ (.A1(_0967_),
    .A2(_2270_),
    .Y(_2271_),
    .B1(net754));
 sg13g2_o21ai_1 _6612_ (.B1(_2271_),
    .Y(_2272_),
    .A1(_0967_),
    .A2(_2270_));
 sg13g2_or3_1 _6613_ (.A(_2245_),
    .B(_2247_),
    .C(_2268_),
    .X(_2273_));
 sg13g2_nand2_2 _6614_ (.Y(_2274_),
    .A(_2269_),
    .B(_2273_));
 sg13g2_nor2_1 _6615_ (.A(_2240_),
    .B(_2274_),
    .Y(_2275_));
 sg13g2_xnor2_1 _6616_ (.Y(_2276_),
    .A(_2193_),
    .B(_2195_));
 sg13g2_a21oi_2 _6617_ (.B1(_2275_),
    .Y(_2277_),
    .A2(_2276_),
    .A1(net754));
 sg13g2_nand3_1 _6618_ (.B(_2272_),
    .C(_2277_),
    .A(_2242_),
    .Y(_2278_));
 sg13g2_and2_1 _6619_ (.A(_3522_),
    .B(_2278_),
    .X(_2279_));
 sg13g2_xnor2_1 _6620_ (.Y(_2280_),
    .A(_2248_),
    .B(_2267_));
 sg13g2_and2_1 _6621_ (.A(_2241_),
    .B(_2280_),
    .X(_2281_));
 sg13g2_xnor2_1 _6622_ (.Y(_2282_),
    .A(_2095_),
    .B(_2096_));
 sg13g2_a21oi_1 _6623_ (.A1(_2185_),
    .A2(_2190_),
    .Y(_2283_),
    .B1(_2188_));
 sg13g2_xnor2_1 _6624_ (.Y(_2284_),
    .A(_2282_),
    .B(_2283_));
 sg13g2_a21oi_2 _6625_ (.B1(_2281_),
    .Y(_2285_),
    .A2(_2284_),
    .A1(net754));
 sg13g2_inv_1 _6626_ (.Y(_2286_),
    .A(_2285_));
 sg13g2_nand3_1 _6627_ (.B(_2264_),
    .C(_2265_),
    .A(_2251_),
    .Y(_2287_));
 sg13g2_nor2_2 _6628_ (.A(net754),
    .B(_2266_),
    .Y(_2288_));
 sg13g2_a21oi_1 _6629_ (.A1(_2189_),
    .A2(_2190_),
    .Y(_2289_),
    .B1(_2185_));
 sg13g2_nor3_1 _6630_ (.A(_2191_),
    .B(_2241_),
    .C(_2289_),
    .Y(_2290_));
 sg13g2_a21o_2 _6631_ (.A2(_2288_),
    .A1(_2287_),
    .B1(_2290_),
    .X(_2291_));
 sg13g2_inv_1 _6632_ (.Y(_2292_),
    .A(_2291_));
 sg13g2_nand2_1 _6633_ (.Y(_2293_),
    .A(_2285_),
    .B(_2291_));
 sg13g2_nor2_1 _6634_ (.A(_2277_),
    .B(_2293_),
    .Y(_2294_));
 sg13g2_nand2_1 _6635_ (.Y(_2295_),
    .A(_1829_),
    .B(_2294_));
 sg13g2_nand2_1 _6636_ (.Y(_2296_),
    .A(_2601_),
    .B(\title_r_pixels_in_scanline[5] ));
 sg13g2_nand2_1 _6637_ (.Y(_2297_),
    .A(net905),
    .B(\title_r_pixels_in_scanline[5] ));
 sg13g2_nor2_1 _6638_ (.A(net905),
    .B(\title_r_pixels_in_scanline[5] ),
    .Y(_2298_));
 sg13g2_xor2_1 _6639_ (.B(\title_r_pixels_in_scanline[5] ),
    .A(net905),
    .X(_2299_));
 sg13g2_nand2b_1 _6640_ (.Y(_2300_),
    .B(\title_r_pixels_in_scanline[3] ),
    .A_N(net912));
 sg13g2_nand2_1 _6641_ (.Y(_2301_),
    .A(net915),
    .B(\title_r_pixels_in_scanline[1] ));
 sg13g2_nor2_1 _6642_ (.A(net915),
    .B(\title_r_pixels_in_scanline[1] ),
    .Y(_2302_));
 sg13g2_xor2_1 _6643_ (.B(\title_r_pixels_in_scanline[1] ),
    .A(net915),
    .X(_2303_));
 sg13g2_a21oi_1 _6644_ (.A1(net916),
    .A2(_3007_),
    .Y(_2304_),
    .B1(_2303_));
 sg13g2_a221oi_1 _6645_ (.B2(_2557_),
    .C1(_2304_),
    .B1(\title_r_pixels_in_scanline[1] ),
    .A1(_2579_),
    .Y(_2305_),
    .A2(\title_r_pixels_in_scanline[2] ));
 sg13g2_xnor2_1 _6646_ (.Y(_2306_),
    .A(net912),
    .B(\title_r_pixels_in_scanline[3] ));
 sg13g2_o21ai_1 _6647_ (.B1(_2306_),
    .Y(_2307_),
    .A1(_2579_),
    .A2(\title_r_pixels_in_scanline[2] ));
 sg13g2_or2_1 _6648_ (.X(_2308_),
    .B(_2307_),
    .A(_2305_));
 sg13g2_xor2_1 _6649_ (.B(\title_r_pixels_in_scanline[4] ),
    .A(net908),
    .X(_2309_));
 sg13g2_a21oi_1 _6650_ (.A1(_2300_),
    .A2(_2308_),
    .Y(_2310_),
    .B1(_2309_));
 sg13g2_a21oi_1 _6651_ (.A1(_2590_),
    .A2(\title_r_pixels_in_scanline[4] ),
    .Y(_2311_),
    .B1(_2310_));
 sg13g2_o21ai_1 _6652_ (.B1(_2296_),
    .Y(_2312_),
    .A1(_2299_),
    .A2(_2311_));
 sg13g2_xor2_1 _6653_ (.B(\title_r_pixels_in_scanline[2] ),
    .A(net914),
    .X(_2313_));
 sg13g2_nor2_1 _6654_ (.A(net916),
    .B(\title_r_pixels_in_scanline[0] ),
    .Y(_2314_));
 sg13g2_xor2_1 _6655_ (.B(\title_r_pixels_in_scanline[0] ),
    .A(net916),
    .X(_2315_));
 sg13g2_nor3_1 _6656_ (.A(_2303_),
    .B(_2313_),
    .C(_2315_),
    .Y(_2316_));
 sg13g2_nand2_1 _6657_ (.Y(_2317_),
    .A(_0019_),
    .B(_2306_));
 sg13g2_nor3_1 _6658_ (.A(_2299_),
    .B(_2309_),
    .C(_2317_),
    .Y(_2318_));
 sg13g2_nor3_2 _6659_ (.A(net827),
    .B(_2675_),
    .C(\hvsync_gen.vpos[9] ),
    .Y(_2319_));
 sg13g2_a21oi_1 _6660_ (.A1(_0033_),
    .A2(_3051_),
    .Y(_2320_),
    .B1(net900));
 sg13g2_nor2_1 _6661_ (.A(\hvsync_gen.hpos[9] ),
    .B(_2633_),
    .Y(_2321_));
 sg13g2_nor3_2 _6662_ (.A(net897),
    .B(\hvsync_gen.hpos[9] ),
    .C(_2633_),
    .Y(_2322_));
 sg13g2_a22oi_1 _6663_ (.Y(_2323_),
    .B1(_2322_),
    .B2(\hvsync_gen.vpos[6] ),
    .A2(_2318_),
    .A1(_2316_));
 sg13g2_nand4_1 _6664_ (.B(_2319_),
    .C(_2320_),
    .A(_2312_),
    .Y(_2324_),
    .D(_2323_));
 sg13g2_and2_1 _6665_ (.A(net835),
    .B(net837),
    .X(_2325_));
 sg13g2_and2_1 _6666_ (.A(net831),
    .B(net830),
    .X(_2326_));
 sg13g2_nand3_1 _6667_ (.B(_2325_),
    .C(_2326_),
    .A(net833),
    .Y(_2327_));
 sg13g2_nand2b_1 _6668_ (.Y(_2328_),
    .B(_2327_),
    .A_N(net827));
 sg13g2_nor2_1 _6669_ (.A(_2644_),
    .B(_3063_),
    .Y(_2329_));
 sg13g2_nand2b_1 _6670_ (.Y(_2330_),
    .B(_3062_),
    .A_N(net835));
 sg13g2_nand3_1 _6671_ (.B(_3015_),
    .C(_3032_),
    .A(_0033_),
    .Y(_2331_));
 sg13g2_a221oi_1 _6672_ (.B2(_0021_),
    .C1(_2331_),
    .B1(_2328_),
    .A1(net896),
    .Y(_2332_),
    .A2(_3275_));
 sg13g2_o21ai_1 _6673_ (.B1(_2332_),
    .Y(_2333_),
    .A1(_2329_),
    .A2(_2330_));
 sg13g2_and2_1 _6674_ (.A(net914),
    .B(\title_r_pixels_in_scanline[2] ),
    .X(_2334_));
 sg13g2_a21oi_1 _6675_ (.A1(_2301_),
    .A2(_2314_),
    .Y(_2335_),
    .B1(_2302_));
 sg13g2_a21oi_1 _6676_ (.A1(_2313_),
    .A2(_2335_),
    .Y(_2336_),
    .B1(_2334_));
 sg13g2_nand4_1 _6677_ (.B(_2303_),
    .C(_2313_),
    .A(net902),
    .Y(_2337_),
    .D(_2315_));
 sg13g2_o21ai_1 _6678_ (.B1(_2337_),
    .Y(_2338_),
    .A1(net913),
    .A2(\title_r_pixels_in_scanline[3] ));
 sg13g2_a22oi_1 _6679_ (.Y(_2339_),
    .B1(\title_r_pixels_in_scanline[3] ),
    .B2(net912),
    .A2(\title_r_pixels_in_scanline[4] ),
    .A1(net908));
 sg13g2_o21ai_1 _6680_ (.B1(_2339_),
    .Y(_2340_),
    .A1(_2336_),
    .A2(_2338_));
 sg13g2_o21ai_1 _6681_ (.B1(_2340_),
    .Y(_2341_),
    .A1(net908),
    .A2(\title_r_pixels_in_scanline[4] ));
 sg13g2_o21ai_1 _6682_ (.B1(_2297_),
    .Y(_2342_),
    .A1(_2298_),
    .A2(_2341_));
 sg13g2_nand4_1 _6683_ (.B(_2319_),
    .C(_2322_),
    .A(_3015_),
    .Y(_2343_),
    .D(_2342_));
 sg13g2_nand3_1 _6684_ (.B(_2333_),
    .C(_2343_),
    .A(_2324_),
    .Y(_2344_));
 sg13g2_o21ai_1 _6685_ (.B1(net860),
    .Y(_2345_),
    .A1(_2407_),
    .A2(_0322_));
 sg13g2_and3_1 _6686_ (.X(_2346_),
    .A(net858),
    .B(_2344_),
    .C(_2345_));
 sg13g2_nor2_1 _6687_ (.A(_3525_),
    .B(_2346_),
    .Y(_2347_));
 sg13g2_nand4_1 _6688_ (.B(_2272_),
    .C(_2277_),
    .A(_2242_),
    .Y(_2348_),
    .D(_2347_));
 sg13g2_nand2_2 _6689_ (.Y(_2349_),
    .A(net229),
    .B(_3521_));
 sg13g2_nand3_1 _6690_ (.B(_2272_),
    .C(_2349_),
    .A(_2242_),
    .Y(_2350_));
 sg13g2_inv_1 _6691_ (.Y(_2351_),
    .A(_2350_));
 sg13g2_nand3b_1 _6692_ (.B(_2348_),
    .C(_2350_),
    .Y(_2352_),
    .A_N(_1829_));
 sg13g2_a21oi_1 _6693_ (.A1(_2295_),
    .A2(_2352_),
    .Y(_2353_),
    .B1(_3522_));
 sg13g2_o21ai_1 _6694_ (.B1(_3520_),
    .Y(_2354_),
    .A1(_2279_),
    .A2(_2353_));
 sg13g2_xor2_1 _6695_ (.B(_2263_),
    .A(_2252_),
    .X(_2355_));
 sg13g2_xnor2_1 _6696_ (.Y(_2357_),
    .A(_2180_),
    .B(_2184_));
 sg13g2_nand2_1 _6697_ (.Y(_2358_),
    .A(net754),
    .B(_2357_));
 sg13g2_o21ai_1 _6698_ (.B1(_2358_),
    .Y(_2359_),
    .A1(net754),
    .A2(_2355_));
 sg13g2_nor2b_1 _6699_ (.A(_2293_),
    .B_N(_2359_),
    .Y(_2360_));
 sg13g2_o21ai_1 _6700_ (.B1(_3516_),
    .Y(_2361_),
    .A1(_2344_),
    .A2(_2360_));
 sg13g2_inv_1 _6701_ (.Y(_2362_),
    .A(_2361_));
 sg13g2_nand2b_1 _6702_ (.Y(_2363_),
    .B(_2261_),
    .A_N(_2260_));
 sg13g2_nand3_1 _6703_ (.B(_2262_),
    .C(_2363_),
    .A(_2241_),
    .Y(_2364_));
 sg13g2_xnor2_1 _6704_ (.Y(_2365_),
    .A(_2177_),
    .B(_2179_));
 sg13g2_o21ai_1 _6705_ (.B1(_2364_),
    .Y(_2366_),
    .A1(_2241_),
    .A2(_2365_));
 sg13g2_and4_1 _6706_ (.A(_2285_),
    .B(_2291_),
    .C(_2359_),
    .D(_2366_),
    .X(_2368_));
 sg13g2_xnor2_1 _6707_ (.Y(_2369_),
    .A(_2258_),
    .B(_2259_));
 sg13g2_nand3_1 _6708_ (.B(_2175_),
    .C(_2176_),
    .A(_2172_),
    .Y(_2370_));
 sg13g2_nor2_1 _6709_ (.A(_2177_),
    .B(_2241_),
    .Y(_2371_));
 sg13g2_a22oi_1 _6710_ (.Y(_2372_),
    .B1(_2370_),
    .B2(_2371_),
    .A2(_2369_),
    .A1(_2241_));
 sg13g2_nor2_1 _6711_ (.A(_3519_),
    .B(_2372_),
    .Y(_2373_));
 sg13g2_a21oi_1 _6712_ (.A1(_2368_),
    .A2(_2373_),
    .Y(_2374_),
    .B1(_2362_));
 sg13g2_a21oi_1 _6713_ (.A1(_2354_),
    .A2(_2374_),
    .Y(_0084_),
    .B1(_3514_));
 sg13g2_or2_1 _6714_ (.X(_2375_),
    .B(_2274_),
    .A(_3526_));
 sg13g2_nor2_1 _6715_ (.A(_2346_),
    .B(_2349_),
    .Y(_2376_));
 sg13g2_nor2_1 _6716_ (.A(_3525_),
    .B(_2376_),
    .Y(_2378_));
 sg13g2_nand2_1 _6717_ (.Y(_2379_),
    .A(_2350_),
    .B(_2378_));
 sg13g2_a221oi_1 _6718_ (.B2(_2379_),
    .C1(_1829_),
    .B1(_2375_),
    .A1(net852),
    .Y(_2380_),
    .A2(net850));
 sg13g2_o21ai_1 _6719_ (.B1(net716),
    .Y(_2381_),
    .A1(_0057_),
    .A2(_3164_));
 sg13g2_nor2_1 _6720_ (.A(net754),
    .B(_2259_),
    .Y(_2382_));
 sg13g2_xnor2_1 _6721_ (.Y(_2383_),
    .A(_2173_),
    .B(_2174_));
 sg13g2_a22oi_1 _6722_ (.Y(_2384_),
    .B1(_2383_),
    .B2(net754),
    .A2(_2382_),
    .A1(_2381_));
 sg13g2_nand4_1 _6723_ (.B(_2366_),
    .C(_2373_),
    .A(_2359_),
    .Y(_2385_),
    .D(_2384_));
 sg13g2_nor3_2 _6724_ (.A(_2277_),
    .B(_2293_),
    .C(_2385_),
    .Y(_2386_));
 sg13g2_o21ai_1 _6725_ (.B1(_3517_),
    .Y(_2387_),
    .A1(_2380_),
    .A2(_2386_));
 sg13g2_a21oi_1 _6726_ (.A1(_2361_),
    .A2(_2387_),
    .Y(_0085_),
    .B1(_3514_));
 sg13g2_mux2_1 _6727_ (.A0(_2286_),
    .A1(net708),
    .S(_2278_),
    .X(_2389_));
 sg13g2_a221oi_1 _6728_ (.B2(_2389_),
    .C1(_3524_),
    .B1(_2376_),
    .A1(_2047_),
    .Y(_2390_),
    .A2(_2351_));
 sg13g2_nand4_1 _6729_ (.B(_1829_),
    .C(_2294_),
    .A(_1256_),
    .Y(_2391_),
    .D(_2359_));
 sg13g2_nand2_1 _6730_ (.Y(_2392_),
    .A(_3525_),
    .B(_2285_));
 sg13g2_nand3b_1 _6731_ (.B(_2391_),
    .C(_2392_),
    .Y(_2393_),
    .A_N(_3522_));
 sg13g2_a221oi_1 _6732_ (.B2(_2389_),
    .C1(_3516_),
    .B1(_3522_),
    .A1(net850),
    .Y(_2394_),
    .A2(_3518_));
 sg13g2_o21ai_1 _6733_ (.B1(_2394_),
    .Y(_2395_),
    .A1(_2390_),
    .A2(_2393_));
 sg13g2_a21oi_1 _6734_ (.A1(_2361_),
    .A2(_2395_),
    .Y(_0086_),
    .B1(_3514_));
 sg13g2_and2_1 _6735_ (.A(_2277_),
    .B(_2349_),
    .X(_2396_));
 sg13g2_a21oi_1 _6736_ (.A1(_2277_),
    .A2(_2349_),
    .Y(_2398_),
    .B1(_1829_));
 sg13g2_nand2_1 _6737_ (.Y(_2399_),
    .A(_2348_),
    .B(_2398_));
 sg13g2_a22oi_1 _6738_ (.Y(_2400_),
    .B1(_2295_),
    .B2(_2399_),
    .A2(net850),
    .A1(net852));
 sg13g2_nand4_1 _6739_ (.B(_3518_),
    .C(_2368_),
    .A(_0034_),
    .Y(_2401_),
    .D(_2384_));
 sg13g2_nand2b_1 _6740_ (.Y(_2402_),
    .B(_2401_),
    .A_N(_2279_));
 sg13g2_o21ai_1 _6741_ (.B1(_3517_),
    .Y(_2403_),
    .A1(_2400_),
    .A2(_2402_));
 sg13g2_a21oi_1 _6742_ (.A1(_2361_),
    .A2(_2403_),
    .Y(_0087_),
    .B1(_3514_));
 sg13g2_nand2b_1 _6743_ (.Y(_2404_),
    .B(_2378_),
    .A_N(_2396_));
 sg13g2_a221oi_1 _6744_ (.B2(_2404_),
    .C1(_1829_),
    .B1(_2392_),
    .A1(net852),
    .Y(_2405_),
    .A2(net850));
 sg13g2_o21ai_1 _6745_ (.B1(_3517_),
    .Y(_2406_),
    .A1(_2386_),
    .A2(_2405_));
 sg13g2_a21oi_1 _6746_ (.A1(_2361_),
    .A2(_2406_),
    .Y(_0088_),
    .B1(_3514_));
 sg13g2_nor2_1 _6747_ (.A(_3522_),
    .B(_2376_),
    .Y(_2408_));
 sg13g2_a21oi_1 _6748_ (.A1(_1144_),
    .A2(_2278_),
    .Y(_2409_),
    .B1(_2408_));
 sg13g2_o21ai_1 _6749_ (.B1(_2409_),
    .Y(_2410_),
    .A1(_2278_),
    .A2(_2292_));
 sg13g2_nor2b_1 _6750_ (.A(_1985_),
    .B_N(_2396_),
    .Y(_2411_));
 sg13g2_a21oi_1 _6751_ (.A1(_3525_),
    .A2(_2291_),
    .Y(_2412_),
    .B1(_3522_));
 sg13g2_o21ai_1 _6752_ (.B1(_2412_),
    .Y(_2413_),
    .A1(_3524_),
    .A2(_2411_));
 sg13g2_nand3_1 _6753_ (.B(_2410_),
    .C(_2413_),
    .A(_3520_),
    .Y(_2414_));
 sg13g2_a21oi_1 _6754_ (.A1(_2361_),
    .A2(_2414_),
    .Y(_0089_),
    .B1(_3514_));
 sg13g2_nor2_1 _6755_ (.A(net165),
    .B(net199),
    .Y(_2415_));
 sg13g2_xor2_1 _6756_ (.B(\r1[14] ),
    .A(\r1[15] ),
    .X(_2417_));
 sg13g2_xnor2_1 _6757_ (.Y(_2418_),
    .A(_0411_),
    .B(_2417_));
 sg13g2_xnor2_1 _6758_ (.Y(_2419_),
    .A(\r1[16] ),
    .B(\r1[17] ));
 sg13g2_xnor2_1 _6759_ (.Y(_2420_),
    .A(_2418_),
    .B(_2419_));
 sg13g2_xnor2_1 _6760_ (.Y(_2421_),
    .A(net844),
    .B(\r1[10] ));
 sg13g2_xor2_1 _6761_ (.B(\r1[8] ),
    .A(\r1[9] ),
    .X(_2422_));
 sg13g2_xnor2_1 _6762_ (.Y(_2423_),
    .A(_2421_),
    .B(_2422_));
 sg13g2_xnor2_1 _6763_ (.Y(_2424_),
    .A(\r1[5] ),
    .B(net846));
 sg13g2_xor2_1 _6764_ (.B(\r1[0] ),
    .A(\r1[1] ),
    .X(_2425_));
 sg13g2_xor2_1 _6765_ (.B(\r1[6] ),
    .A(\r1[7] ),
    .X(_2426_));
 sg13g2_xnor2_1 _6766_ (.Y(_2428_),
    .A(_2425_),
    .B(_2426_));
 sg13g2_xnor2_1 _6767_ (.Y(_2429_),
    .A(net847),
    .B(net848));
 sg13g2_xnor2_1 _6768_ (.Y(_2430_),
    .A(_2424_),
    .B(_2429_));
 sg13g2_xnor2_1 _6769_ (.Y(_2431_),
    .A(_2428_),
    .B(_2430_));
 sg13g2_xnor2_1 _6770_ (.Y(_2432_),
    .A(_2423_),
    .B(_2431_));
 sg13g2_xnor2_1 _6771_ (.Y(_2433_),
    .A(_2420_),
    .B(_2432_));
 sg13g2_nor3_1 _6772_ (.A(net767),
    .B(_2415_),
    .C(_2433_),
    .Y(_2434_));
 sg13g2_o21ai_1 _6773_ (.B1(net926),
    .Y(_2435_),
    .A1(net211),
    .A2(_2434_));
 sg13g2_a21oi_1 _6774_ (.A1(net211),
    .A2(_2434_),
    .Y(_0090_),
    .B1(_2435_));
 sg13g2_nand2b_1 _6775_ (.Y(_2436_),
    .B(_2415_),
    .A_N(net184));
 sg13g2_o21ai_1 _6776_ (.B1(net925),
    .Y(_2438_),
    .A1(net184),
    .A2(net768));
 sg13g2_a21oi_1 _6777_ (.A1(net768),
    .A2(_2436_),
    .Y(_0091_),
    .B1(_2438_));
 sg13g2_a21oi_1 _6778_ (.A1(net184),
    .A2(_2415_),
    .Y(_2439_),
    .B1(net767));
 sg13g2_o21ai_1 _6779_ (.B1(net925),
    .Y(_2440_),
    .A1(\noise_counter[1] ),
    .A2(net768));
 sg13g2_nor2_1 _6780_ (.A(net185),
    .B(_2440_),
    .Y(_0092_));
 sg13g2_and3_1 _6781_ (.X(_0093_),
    .A(net165),
    .B(net925),
    .C(net767));
 sg13g2_nand2b_1 _6782_ (.Y(_2441_),
    .B(\note2_freq[1] ),
    .A_N(\note2_counter[1] ));
 sg13g2_nand3b_1 _6783_ (.B(_2441_),
    .C(\note2_counter[0] ),
    .Y(_2442_),
    .A_N(\note2_freq[0] ));
 sg13g2_nand2b_1 _6784_ (.Y(_2443_),
    .B(\note2_counter[1] ),
    .A_N(\note2_freq[1] ));
 sg13g2_nand3_1 _6785_ (.B(_2442_),
    .C(_2443_),
    .A(\note2_counter[2] ),
    .Y(_2444_));
 sg13g2_o21ai_1 _6786_ (.B1(_2444_),
    .Y(_2446_),
    .A1(\note2_counter[3] ),
    .A2(_2726_));
 sg13g2_a22oi_1 _6787_ (.Y(_2447_),
    .B1(_2726_),
    .B2(\note2_counter[3] ),
    .A2(_2716_),
    .A1(\note2_counter[4] ));
 sg13g2_o21ai_1 _6788_ (.B1(_2447_),
    .Y(_2448_),
    .A1(_0028_),
    .A2(_2446_));
 sg13g2_a22oi_1 _6789_ (.Y(_2449_),
    .B1(\note2_freq[4] ),
    .B2(_2543_),
    .A2(\note2_freq[5] ),
    .A1(_2536_));
 sg13g2_a22oi_1 _6790_ (.Y(_2450_),
    .B1(_2448_),
    .B2(_2449_),
    .A2(_2705_),
    .A1(\note2_counter[5] ));
 sg13g2_a21oi_1 _6791_ (.A1(_2529_),
    .A2(\note2_freq[6] ),
    .Y(_2451_),
    .B1(_2450_));
 sg13g2_nand2b_1 _6792_ (.Y(_2452_),
    .B(\note2_counter[7] ),
    .A_N(\note2_freq[7] ));
 sg13g2_o21ai_1 _6793_ (.B1(_2452_),
    .Y(_2453_),
    .A1(_2529_),
    .A2(\note2_freq[6] ));
 sg13g2_a22oi_1 _6794_ (.Y(_2454_),
    .B1(\note2_freq[7] ),
    .B2(_2522_),
    .A2(\note2_freq[8] ),
    .A1(_2514_));
 sg13g2_o21ai_1 _6795_ (.B1(_2454_),
    .Y(_2455_),
    .A1(_2451_),
    .A2(_2453_));
 sg13g2_o21ai_1 _6796_ (.B1(_2455_),
    .Y(_2457_),
    .A1(_2514_),
    .A2(\note2_freq[8] ));
 sg13g2_nor2_1 _6797_ (.A(_3061_),
    .B(_2457_),
    .Y(_2458_));
 sg13g2_o21ai_1 _6798_ (.B1(net926),
    .Y(_2459_),
    .A1(net187),
    .A2(_2458_));
 sg13g2_a21oi_1 _6799_ (.A1(net187),
    .A2(net769),
    .Y(_0094_),
    .B1(_2459_));
 sg13g2_nand2_2 _6800_ (.Y(_2460_),
    .A(net769),
    .B(_2457_));
 sg13g2_nand2_2 _6801_ (.Y(_2461_),
    .A(net929),
    .B(_2460_));
 sg13g2_a21oi_1 _6802_ (.A1(\note2_counter[0] ),
    .A2(net769),
    .Y(_2462_),
    .B1(net181));
 sg13g2_nand2_1 _6803_ (.Y(_2463_),
    .A(net181),
    .B(net187));
 sg13g2_nor2_1 _6804_ (.A(_3061_),
    .B(_2463_),
    .Y(_2464_));
 sg13g2_nor3_1 _6805_ (.A(_2461_),
    .B(net182),
    .C(_2464_),
    .Y(_0095_));
 sg13g2_xor2_1 _6806_ (.B(_2463_),
    .A(_0028_),
    .X(_2466_));
 sg13g2_a22oi_1 _6807_ (.Y(_2467_),
    .B1(_2458_),
    .B2(_2466_),
    .A2(_3061_),
    .A1(net192));
 sg13g2_nor2_1 _6808_ (.A(net923),
    .B(net193),
    .Y(_0096_));
 sg13g2_and3_1 _6809_ (.X(_2468_),
    .A(net178),
    .B(net192),
    .C(_2464_));
 sg13g2_a21oi_1 _6810_ (.A1(\note2_counter[2] ),
    .A2(_2464_),
    .Y(_2469_),
    .B1(net178));
 sg13g2_nor3_1 _6811_ (.A(_2461_),
    .B(_2468_),
    .C(net179),
    .Y(_0097_));
 sg13g2_xnor2_1 _6812_ (.Y(_2470_),
    .A(net208),
    .B(_2468_));
 sg13g2_nor2_1 _6813_ (.A(_2461_),
    .B(_2470_),
    .Y(_0098_));
 sg13g2_and3_1 _6814_ (.X(_2471_),
    .A(net175),
    .B(\note2_counter[4] ),
    .C(_2468_));
 sg13g2_a21oi_1 _6815_ (.A1(\note2_counter[4] ),
    .A2(_2468_),
    .Y(_2472_),
    .B1(net175));
 sg13g2_nor3_1 _6816_ (.A(_2461_),
    .B(_2471_),
    .C(net176),
    .Y(_0099_));
 sg13g2_and2_1 _6817_ (.A(net190),
    .B(_2471_),
    .X(_2474_));
 sg13g2_nor2_1 _6818_ (.A(net190),
    .B(_2471_),
    .Y(_2475_));
 sg13g2_nor3_1 _6819_ (.A(_2461_),
    .B(_2474_),
    .C(net191),
    .Y(_0100_));
 sg13g2_nand2_1 _6820_ (.Y(_2476_),
    .A(net201),
    .B(_2474_));
 sg13g2_xnor2_1 _6821_ (.Y(_2477_),
    .A(net201),
    .B(_2474_));
 sg13g2_nor2_1 _6822_ (.A(_2461_),
    .B(_2477_),
    .Y(_0101_));
 sg13g2_xnor2_1 _6823_ (.Y(_2478_),
    .A(_2514_),
    .B(_2476_));
 sg13g2_nor2_1 _6824_ (.A(_2461_),
    .B(_2478_),
    .Y(_0102_));
 sg13g2_o21ai_1 _6825_ (.B1(net929),
    .Y(_2479_),
    .A1(net166),
    .A2(_2460_));
 sg13g2_a21oi_1 _6826_ (.A1(_2507_),
    .A2(_2460_),
    .Y(_0103_),
    .B1(_2479_));
 sg13g2_nor2_1 _6827_ (.A(_2473_),
    .B(\note_freq[7] ),
    .Y(_2481_));
 sg13g2_nor2b_1 _6828_ (.A(\note_freq[0] ),
    .B_N(\note_counter[0] ),
    .Y(_2482_));
 sg13g2_o21ai_1 _6829_ (.B1(_2482_),
    .Y(_2483_),
    .A1(\note_counter[1] ),
    .A2(_2747_));
 sg13g2_a22oi_1 _6830_ (.Y(_2484_),
    .B1(_2757_),
    .B2(\note_counter[2] ),
    .A2(_2747_),
    .A1(\note_counter[1] ));
 sg13g2_a22oi_1 _6831_ (.Y(_2485_),
    .B1(_2483_),
    .B2(_2484_),
    .A2(\note_freq[2] ),
    .A1(_2500_));
 sg13g2_o21ai_1 _6832_ (.B1(_2485_),
    .Y(_2486_),
    .A1(\note_counter[3] ),
    .A2(_2747_));
 sg13g2_a22oi_1 _6833_ (.Y(_2487_),
    .B1(_2747_),
    .B2(\note_counter[3] ),
    .A2(_2737_),
    .A1(\note_counter[4] ));
 sg13g2_nor2b_1 _6834_ (.A(\note_counter[5] ),
    .B_N(\note_freq[5] ),
    .Y(_2488_));
 sg13g2_a221oi_1 _6835_ (.B2(_2487_),
    .C1(_2488_),
    .B1(_2486_),
    .A1(_2490_),
    .Y(_2489_),
    .A2(\note_freq[4] ));
 sg13g2_nand2b_1 _6836_ (.Y(_2491_),
    .B(\note_counter[5] ),
    .A_N(\note_freq[5] ));
 sg13g2_o21ai_1 _6837_ (.B1(_2491_),
    .Y(_2492_),
    .A1(_2480_),
    .A2(\note_freq[6] ));
 sg13g2_nor2_1 _6838_ (.A(_2489_),
    .B(_2492_),
    .Y(_2493_));
 sg13g2_a221oi_1 _6839_ (.B2(_2480_),
    .C1(_2493_),
    .B1(\note_freq[6] ),
    .A1(_2473_),
    .Y(_2494_),
    .A2(\note_freq[7] ));
 sg13g2_o21ai_1 _6840_ (.B1(net768),
    .Y(_2495_),
    .A1(_2481_),
    .A2(_2494_));
 sg13g2_nand2_2 _6841_ (.Y(_2496_),
    .A(net925),
    .B(_2495_));
 sg13g2_xnor2_1 _6842_ (.Y(_2497_),
    .A(net198),
    .B(net768));
 sg13g2_nor2_1 _6843_ (.A(_2496_),
    .B(_2497_),
    .Y(_0104_));
 sg13g2_and3_1 _6844_ (.X(_2498_),
    .A(net172),
    .B(\note_counter[0] ),
    .C(net768));
 sg13g2_a21oi_1 _6845_ (.A1(\note_counter[0] ),
    .A2(net768),
    .Y(_2499_),
    .B1(net172));
 sg13g2_nor3_1 _6846_ (.A(_2496_),
    .B(_2498_),
    .C(net173),
    .Y(_0105_));
 sg13g2_and2_1 _6847_ (.A(net195),
    .B(_2498_),
    .X(_2501_));
 sg13g2_nor2_1 _6848_ (.A(net195),
    .B(_2498_),
    .Y(_2502_));
 sg13g2_nor3_1 _6849_ (.A(_2496_),
    .B(_2501_),
    .C(net196),
    .Y(_0106_));
 sg13g2_and2_1 _6850_ (.A(net188),
    .B(_2501_),
    .X(_2503_));
 sg13g2_nor2_1 _6851_ (.A(net188),
    .B(_2501_),
    .Y(_2504_));
 sg13g2_nor3_1 _6852_ (.A(_2496_),
    .B(_2503_),
    .C(net189),
    .Y(_0107_));
 sg13g2_and2_1 _6853_ (.A(net194),
    .B(_2503_),
    .X(_2505_));
 sg13g2_nor2_1 _6854_ (.A(net194),
    .B(_2503_),
    .Y(_2506_));
 sg13g2_nor3_1 _6855_ (.A(_2496_),
    .B(_2505_),
    .C(_2506_),
    .Y(_0108_));
 sg13g2_and2_1 _6856_ (.A(net197),
    .B(_2505_),
    .X(_2508_));
 sg13g2_nor2_1 _6857_ (.A(net197),
    .B(_2505_),
    .Y(_2509_));
 sg13g2_nor3_1 _6858_ (.A(_2496_),
    .B(_2508_),
    .C(_2509_),
    .Y(_0109_));
 sg13g2_nand2_1 _6859_ (.Y(_2510_),
    .A(net200),
    .B(_2508_));
 sg13g2_xnor2_1 _6860_ (.Y(_2511_),
    .A(net200),
    .B(_2508_));
 sg13g2_nor2_1 _6861_ (.A(_2496_),
    .B(_2511_),
    .Y(_0110_));
 sg13g2_xnor2_1 _6862_ (.Y(_2512_),
    .A(_2473_),
    .B(_2510_));
 sg13g2_nor2_1 _6863_ (.A(_2496_),
    .B(_2512_),
    .Y(_0111_));
 sg13g2_o21ai_1 _6864_ (.B1(net925),
    .Y(_2513_),
    .A1(net168),
    .A2(_2495_));
 sg13g2_a21oi_1 _6865_ (.A1(_2465_),
    .A2(_2495_),
    .Y(_0112_),
    .B1(_2513_));
 sg13g2_nor3_1 _6866_ (.A(_2557_),
    .B(_2568_),
    .C(_2579_),
    .Y(_2515_));
 sg13g2_and3_2 _6867_ (.X(_2516_),
    .A(net913),
    .B(net909),
    .C(_2515_));
 sg13g2_and4_2 _6868_ (.A(_2601_),
    .B(_3054_),
    .C(_3058_),
    .D(_2516_),
    .X(_2517_));
 sg13g2_nor2_1 _6869_ (.A(net924),
    .B(_2517_),
    .Y(_2518_));
 sg13g2_nand2b_2 _6870_ (.Y(_2519_),
    .B(net929),
    .A_N(_2517_));
 sg13g2_and2_1 _6871_ (.A(net159),
    .B(net745),
    .X(_0113_));
 sg13g2_o21ai_1 _6872_ (.B1(net745),
    .Y(_2520_),
    .A1(_2557_),
    .A2(_2568_));
 sg13g2_a21oi_1 _6873_ (.A1(_2557_),
    .A2(_2568_),
    .Y(_0114_),
    .B1(_2520_));
 sg13g2_a21oi_1 _6874_ (.A1(net915),
    .A2(net916),
    .Y(_2521_),
    .B1(net914));
 sg13g2_nor3_1 _6875_ (.A(net924),
    .B(_2515_),
    .C(net231),
    .Y(_0115_));
 sg13g2_nand3b_1 _6876_ (.B(net916),
    .C(net915),
    .Y(_2523_),
    .A_N(net266));
 sg13g2_xor2_1 _6877_ (.B(_2523_),
    .A(net911),
    .X(_2524_));
 sg13g2_nor2_1 _6878_ (.A(_2519_),
    .B(_2524_),
    .Y(_0116_));
 sg13g2_a21oi_1 _6879_ (.A1(net911),
    .A2(_2515_),
    .Y(_2525_),
    .B1(net909));
 sg13g2_nor3_1 _6880_ (.A(net924),
    .B(_2516_),
    .C(_2525_),
    .Y(_0117_));
 sg13g2_nand2_2 _6881_ (.Y(_2526_),
    .A(net906),
    .B(_2516_));
 sg13g2_o21ai_1 _6882_ (.B1(net745),
    .Y(_2527_),
    .A1(net906),
    .A2(_2516_));
 sg13g2_nor2b_1 _6883_ (.A(_2527_),
    .B_N(_2526_),
    .Y(_0118_));
 sg13g2_o21ai_1 _6884_ (.B1(net745),
    .Y(_2528_),
    .A1(net815),
    .A2(_2526_));
 sg13g2_a21oi_1 _6885_ (.A1(net815),
    .A2(_2526_),
    .Y(_0119_),
    .B1(_2528_));
 sg13g2_nor2_1 _6886_ (.A(net212),
    .B(_2526_),
    .Y(_2530_));
 sg13g2_xnor2_1 _6887_ (.Y(_2531_),
    .A(net897),
    .B(_2530_));
 sg13g2_nor2_1 _6888_ (.A(_2519_),
    .B(_2531_),
    .Y(_0120_));
 sg13g2_nand4_1 _6889_ (.B(net897),
    .C(net900),
    .A(net906),
    .Y(_2532_),
    .D(_2516_));
 sg13g2_o21ai_1 _6890_ (.B1(_2518_),
    .Y(_2533_),
    .A1(_2633_),
    .A2(_2532_));
 sg13g2_a21oi_1 _6891_ (.A1(_2633_),
    .A2(_2532_),
    .Y(_0121_),
    .B1(_2533_));
 sg13g2_nor2_1 _6892_ (.A(net206),
    .B(_2532_),
    .Y(_2534_));
 sg13g2_xnor2_1 _6893_ (.Y(_2535_),
    .A(\hvsync_gen.hpos[9] ),
    .B(_2534_));
 sg13g2_nor2_1 _6894_ (.A(_2519_),
    .B(net207),
    .Y(_0122_));
 sg13g2_and2_1 _6895_ (.A(net930),
    .B(net205),
    .X(_0123_));
 sg13g2_and2_1 _6896_ (.A(net930),
    .B(net164),
    .X(_0124_));
 sg13g2_a21oi_1 _6897_ (.A1(net849),
    .A2(_3067_),
    .Y(_2537_),
    .B1(net894));
 sg13g2_nand3_1 _6898_ (.B(net893),
    .C(_3067_),
    .A(net849),
    .Y(_2538_));
 sg13g2_nand2_1 _6899_ (.Y(_2539_),
    .A(net927),
    .B(_2538_));
 sg13g2_nor2_2 _6900_ (.A(_2537_),
    .B(_2539_),
    .Y(_0125_));
 sg13g2_o21ai_1 _6901_ (.B1(net927),
    .Y(_2540_),
    .A1(net816),
    .A2(_2538_));
 sg13g2_a21oi_1 _6902_ (.A1(net816),
    .A2(_2538_),
    .Y(_0126_),
    .B1(_2540_));
 sg13g2_nor2_1 _6903_ (.A(net260),
    .B(_2538_),
    .Y(_2541_));
 sg13g2_o21ai_1 _6904_ (.B1(net927),
    .Y(_2542_),
    .A1(net879),
    .A2(_2541_));
 sg13g2_a21oi_1 _6905_ (.A1(net879),
    .A2(_2541_),
    .Y(_0127_),
    .B1(_2542_));
 sg13g2_a21oi_1 _6906_ (.A1(net874),
    .A2(_3068_),
    .Y(_2544_),
    .B1(_3078_));
 sg13g2_nor2_1 _6907_ (.A(net923),
    .B(_2544_),
    .Y(_0128_));
 sg13g2_nand2_1 _6908_ (.Y(_2545_),
    .A(net867),
    .B(_3068_));
 sg13g2_a21oi_1 _6909_ (.A1(_3083_),
    .A2(_2545_),
    .Y(_0129_),
    .B1(net923));
 sg13g2_nand2_1 _6910_ (.Y(_2546_),
    .A(net264),
    .B(_3068_));
 sg13g2_a21oi_1 _6911_ (.A1(_3073_),
    .A2(_2546_),
    .Y(_0130_),
    .B1(net923));
 sg13g2_nand2_1 _6912_ (.Y(_2547_),
    .A(net289),
    .B(_3068_));
 sg13g2_a21oi_1 _6913_ (.A1(_3090_),
    .A2(_2547_),
    .Y(_0131_),
    .B1(net923));
 sg13g2_nor2_1 _6914_ (.A(net224),
    .B(net753),
    .Y(_2548_));
 sg13g2_o21ai_1 _6915_ (.B1(_0030_),
    .Y(_2549_),
    .A1(_3070_),
    .A2(_3096_));
 sg13g2_nor2_1 _6916_ (.A(_3068_),
    .B(_2549_),
    .Y(_2551_));
 sg13g2_nor3_1 _6917_ (.A(_3099_),
    .B(_2548_),
    .C(_2551_),
    .Y(_0132_));
 sg13g2_o21ai_1 _6918_ (.B1(net930),
    .Y(_2552_),
    .A1(net851),
    .A2(_3098_));
 sg13g2_a21oi_1 _6919_ (.A1(net851),
    .A2(_3098_),
    .Y(_0133_),
    .B1(_2552_));
 sg13g2_nand2b_1 _6920_ (.Y(_2553_),
    .B(_3521_),
    .A_N(_3097_));
 sg13g2_o21ai_1 _6921_ (.B1(net930),
    .Y(_2554_),
    .A1(_3097_),
    .A2(_2349_));
 sg13g2_a21oi_1 _6922_ (.A1(_2388_),
    .A2(_2553_),
    .Y(_0134_),
    .B1(_2554_));
 sg13g2_o21ai_1 _6923_ (.B1(net929),
    .Y(_2555_),
    .A1(net849),
    .A2(_3067_));
 sg13g2_a21oi_1 _6924_ (.A1(_2377_),
    .A2(net753),
    .Y(_0135_),
    .B1(_2555_));
 sg13g2_nor2_1 _6925_ (.A(\center_y[0] ),
    .B(net911),
    .Y(_2556_));
 sg13g2_nor2_1 _6926_ (.A(net849),
    .B(net914),
    .Y(_2558_));
 sg13g2_a22oi_1 _6927_ (.Y(_2559_),
    .B1(net908),
    .B2(net889),
    .A2(net910),
    .A1(net895));
 sg13g2_o21ai_1 _6928_ (.B1(_2559_),
    .Y(_2560_),
    .A1(_2556_),
    .A2(_2558_));
 sg13g2_a22oi_1 _6929_ (.Y(_2561_),
    .B1(_2601_),
    .B2(_2437_),
    .A2(_2590_),
    .A1(_2445_));
 sg13g2_nand2_1 _6930_ (.Y(_2562_),
    .A(net880),
    .B(net904));
 sg13g2_xor2_1 _6931_ (.B(net901),
    .A(\center_x[2] ),
    .X(_2563_));
 sg13g2_nand3_1 _6932_ (.B(_2562_),
    .C(_2563_),
    .A(_0022_),
    .Y(_2564_));
 sg13g2_a21oi_1 _6933_ (.A1(_2560_),
    .A2(_2561_),
    .Y(_2565_),
    .B1(_2564_));
 sg13g2_a21o_1 _6934_ (.A2(_3058_),
    .A1(net817),
    .B1(_2565_),
    .X(_2566_));
 sg13g2_and2_1 _6935_ (.A(net840),
    .B(net838),
    .X(_2567_));
 sg13g2_and2_1 _6936_ (.A(net837),
    .B(_2567_),
    .X(_2569_));
 sg13g2_o21ai_1 _6937_ (.B1(\hvsync_gen.vpos[8] ),
    .Y(_2570_),
    .A1(_2330_),
    .A2(_2569_));
 sg13g2_nor4_1 _6938_ (.A(net840),
    .B(net835),
    .C(_2644_),
    .D(_3040_),
    .Y(_2571_));
 sg13g2_nor4_1 _6939_ (.A(\hvsync_gen.hpos[9] ),
    .B(net896),
    .C(\hvsync_gen.vpos[9] ),
    .D(_2571_),
    .Y(_2572_));
 sg13g2_nand3_1 _6940_ (.B(_2570_),
    .C(_2572_),
    .A(_2566_),
    .Y(_2573_));
 sg13g2_nand2_1 _6941_ (.Y(_2574_),
    .A(net816),
    .B(_2601_));
 sg13g2_nand2b_1 _6942_ (.Y(_2575_),
    .B(_0029_),
    .A_N(net849));
 sg13g2_nor2b_1 _6943_ (.A(_0029_),
    .B_N(net849),
    .Y(_2576_));
 sg13g2_a221oi_1 _6944_ (.B2(net910),
    .C1(_2576_),
    .B1(_2575_),
    .A1(net895),
    .Y(_2577_),
    .A2(net907));
 sg13g2_o21ai_1 _6945_ (.B1(_2574_),
    .Y(_2578_),
    .A1(net895),
    .A2(net907));
 sg13g2_a22oi_1 _6946_ (.Y(_2580_),
    .B1(net900),
    .B2(net880),
    .A2(net903),
    .A1(net889));
 sg13g2_o21ai_1 _6947_ (.B1(_2580_),
    .Y(_2581_),
    .A1(_2577_),
    .A2(_2578_));
 sg13g2_o21ai_1 _6948_ (.B1(_2581_),
    .Y(_2582_),
    .A1(net880),
    .A2(net900));
 sg13g2_nand3_1 _6949_ (.B(net897),
    .C(_3059_),
    .A(noise),
    .Y(_2583_));
 sg13g2_nor3_1 _6950_ (.A(_3516_),
    .B(_3527_),
    .C(_2583_),
    .Y(_2584_));
 sg13g2_a21oi_1 _6951_ (.A1(_3024_),
    .A2(_3527_),
    .Y(_2585_),
    .B1(_0022_));
 sg13g2_nor2_1 _6952_ (.A(_3024_),
    .B(_3527_),
    .Y(_2586_));
 sg13g2_o21ai_1 _6953_ (.B1(_2586_),
    .Y(_2587_),
    .A1(net903),
    .A2(_3015_));
 sg13g2_nand3_1 _6954_ (.B(_3047_),
    .C(_2587_),
    .A(note2),
    .Y(_2588_));
 sg13g2_o21ai_1 _6955_ (.B1(net849),
    .Y(_2589_),
    .A1(net910),
    .A2(net908));
 sg13g2_a22oi_1 _6956_ (.Y(_2591_),
    .B1(net903),
    .B2(net895),
    .A2(net907),
    .A1(net910));
 sg13g2_nor2_1 _6957_ (.A(net895),
    .B(net903),
    .Y(_2592_));
 sg13g2_a221oi_1 _6958_ (.B2(_2591_),
    .C1(_2592_),
    .B1(_2589_),
    .A1(net816),
    .Y(_2593_),
    .A2(net815));
 sg13g2_a22oi_1 _6959_ (.Y(_2594_),
    .B1(net901),
    .B2(net889),
    .A2(net898),
    .A1(net883));
 sg13g2_nand2b_1 _6960_ (.Y(_2595_),
    .B(_2594_),
    .A_N(_2593_));
 sg13g2_o21ai_1 _6961_ (.B1(_2595_),
    .Y(_2596_),
    .A1(net880),
    .A2(net898));
 sg13g2_nand2b_1 _6962_ (.Y(_2597_),
    .B(net850),
    .A_N(_3521_));
 sg13g2_nand4_1 _6963_ (.B(_2321_),
    .C(_2596_),
    .A(note),
    .Y(_2598_),
    .D(_2597_));
 sg13g2_o21ai_1 _6964_ (.B1(_2598_),
    .Y(_2599_),
    .A1(_2585_),
    .A2(_2588_));
 sg13g2_a21oi_1 _6965_ (.A1(_2582_),
    .A2(_2584_),
    .Y(_2600_),
    .B1(_2599_));
 sg13g2_a21oi_2 _6966_ (.B1(net924),
    .Y(_0136_),
    .A2(_2600_),
    .A1(_2573_));
 sg13g2_nor2_1 _6967_ (.A(net767),
    .B(_3143_),
    .Y(_2602_));
 sg13g2_nand2_1 _6968_ (.Y(_2603_),
    .A(net769),
    .B(_3142_));
 sg13g2_nor2b_1 _6969_ (.A(net824),
    .B_N(\r1[0] ),
    .Y(_2604_));
 sg13g2_nor2_1 _6970_ (.A(net255),
    .B(net742),
    .Y(_2605_));
 sg13g2_nor2_1 _6971_ (.A(net778),
    .B(_2605_),
    .Y(_2606_));
 sg13g2_o21ai_1 _6972_ (.B1(_2606_),
    .Y(_2607_),
    .A1(_2602_),
    .A2(_2604_));
 sg13g2_nand2_1 _6973_ (.Y(_2608_),
    .A(_3059_),
    .B(_3584_));
 sg13g2_nor2_1 _6974_ (.A(net903),
    .B(net810),
    .Y(_2609_));
 sg13g2_nand2_1 _6975_ (.Y(_2610_),
    .A(net880),
    .B(_2579_));
 sg13g2_o21ai_1 _6976_ (.B1(_2610_),
    .Y(_2612_),
    .A1(net817),
    .A2(net910));
 sg13g2_nand2_1 _6977_ (.Y(_2613_),
    .A(net817),
    .B(net910));
 sg13g2_o21ai_1 _6978_ (.B1(_2613_),
    .Y(_2614_),
    .A1(net880),
    .A2(_2579_));
 sg13g2_nor2_1 _6979_ (.A(_2612_),
    .B(_2614_),
    .Y(_2615_));
 sg13g2_a22oi_1 _6980_ (.Y(_2616_),
    .B1(net916),
    .B2(_2456_),
    .A2(net915),
    .A1(net816));
 sg13g2_nor2_1 _6981_ (.A(net816),
    .B(net915),
    .Y(_2617_));
 sg13g2_o21ai_1 _6982_ (.B1(_2615_),
    .Y(_2618_),
    .A1(_2616_),
    .A2(_2617_));
 sg13g2_a22oi_1 _6983_ (.Y(_2619_),
    .B1(_2612_),
    .B2(_2613_),
    .A2(_2590_),
    .A1(net818));
 sg13g2_a22oi_1 _6984_ (.Y(_2620_),
    .B1(_2618_),
    .B2(_2619_),
    .A2(net907),
    .A1(net873));
 sg13g2_xnor2_1 _6985_ (.Y(_2621_),
    .A(_3015_),
    .B(net149));
 sg13g2_o21ai_1 _6986_ (.B1(_2621_),
    .Y(_2623_),
    .A1(_2609_),
    .A2(_2620_));
 sg13g2_a21oi_1 _6987_ (.A1(net903),
    .A2(net810),
    .Y(_2624_),
    .B1(_2623_));
 sg13g2_a221oi_1 _6988_ (.B2(net815),
    .C1(_2624_),
    .B1(net150),
    .A1(_0022_),
    .Y(_2625_),
    .A2(net806));
 sg13g2_o21ai_1 _6989_ (.B1(_0033_),
    .Y(_2626_),
    .A1(_3024_),
    .A2(net806));
 sg13g2_a21oi_1 _6990_ (.A1(_3024_),
    .A2(net806),
    .Y(_2627_),
    .B1(_2626_));
 sg13g2_or2_1 _6991_ (.X(_2628_),
    .B(net806),
    .A(_0022_));
 sg13g2_nand2_1 _6992_ (.Y(_2629_),
    .A(_2627_),
    .B(_2628_));
 sg13g2_o21ai_1 _6993_ (.B1(_2608_),
    .Y(_2630_),
    .A1(_2625_),
    .A2(_2629_));
 sg13g2_xor2_1 _6994_ (.B(net907),
    .A(net873),
    .X(_2631_));
 sg13g2_a21oi_1 _6995_ (.A1(_0022_),
    .A2(net806),
    .Y(_2632_),
    .B1(_2609_));
 sg13g2_and2_1 _6996_ (.A(_2616_),
    .B(_2631_),
    .X(_2634_));
 sg13g2_a221oi_1 _6997_ (.B2(net810),
    .C1(_2617_),
    .B1(net904),
    .A1(net895),
    .Y(_2635_),
    .A2(_2568_));
 sg13g2_and4_1 _6998_ (.A(_2621_),
    .B(_2628_),
    .C(_2634_),
    .D(_2635_),
    .X(_2636_));
 sg13g2_nand4_1 _6999_ (.B(_2627_),
    .C(_2632_),
    .A(_2615_),
    .Y(_2637_),
    .D(_2636_));
 sg13g2_and2_2 _7000_ (.A(_2630_),
    .B(_2637_),
    .X(_2638_));
 sg13g2_nand2_1 _7001_ (.Y(_2639_),
    .A(_2630_),
    .B(_2637_));
 sg13g2_nand2_1 _7002_ (.Y(_2640_),
    .A(net893),
    .B(\r1[0] ));
 sg13g2_xnor2_1 _7003_ (.Y(_2641_),
    .A(net894),
    .B(\r1[0] ));
 sg13g2_a21oi_1 _7004_ (.A1(_2638_),
    .A2(_2641_),
    .Y(_2642_),
    .B1(_3106_));
 sg13g2_o21ai_1 _7005_ (.B1(_2642_),
    .Y(_2643_),
    .A1(_2604_),
    .A2(_2638_));
 sg13g2_a21oi_1 _7006_ (.A1(_2607_),
    .A2(_2643_),
    .Y(_0137_),
    .B1(net923));
 sg13g2_nand2b_1 _7007_ (.Y(_2645_),
    .B(\r1[1] ),
    .A_N(net824));
 sg13g2_xor2_1 _7008_ (.B(\r1[1] ),
    .A(net885),
    .X(_2646_));
 sg13g2_nand2b_1 _7009_ (.Y(_2647_),
    .B(_2646_),
    .A_N(_2640_));
 sg13g2_xnor2_1 _7010_ (.Y(_2648_),
    .A(_2640_),
    .B(_2646_));
 sg13g2_a21oi_1 _7011_ (.A1(_2638_),
    .A2(_2648_),
    .Y(_2649_),
    .B1(net775));
 sg13g2_o21ai_1 _7012_ (.B1(_2649_),
    .Y(_2650_),
    .A1(net724),
    .A2(_2645_));
 sg13g2_nand2_1 _7013_ (.Y(_2651_),
    .A(\r1[1] ),
    .B(_1907_));
 sg13g2_nand2_1 _7014_ (.Y(_2652_),
    .A(_2841_),
    .B(_1908_));
 sg13g2_nand2_1 _7015_ (.Y(_2653_),
    .A(_2651_),
    .B(_2652_));
 sg13g2_a21oi_1 _7016_ (.A1(_2605_),
    .A2(_2653_),
    .Y(_2655_),
    .B1(net778));
 sg13g2_nand2b_1 _7017_ (.Y(_2656_),
    .B(net743),
    .A_N(_2645_));
 sg13g2_nand4_1 _7018_ (.B(net744),
    .C(_2651_),
    .A(net255),
    .Y(_2657_),
    .D(_2652_));
 sg13g2_nand3_1 _7019_ (.B(_2656_),
    .C(_2657_),
    .A(_2655_),
    .Y(_2658_));
 sg13g2_and3_1 _7020_ (.X(_0138_),
    .A(net927),
    .B(_2650_),
    .C(_2658_));
 sg13g2_and2_1 _7021_ (.A(net878),
    .B(\r1[2] ),
    .X(_2659_));
 sg13g2_xor2_1 _7022_ (.B(net848),
    .A(net878),
    .X(_2660_));
 sg13g2_o21ai_1 _7023_ (.B1(_2647_),
    .Y(_2661_),
    .A1(net816),
    .A2(_2841_));
 sg13g2_xnor2_1 _7024_ (.Y(_2662_),
    .A(_2660_),
    .B(_2661_));
 sg13g2_nand2b_1 _7025_ (.Y(_2663_),
    .B(net848),
    .A_N(net824));
 sg13g2_nand2_1 _7026_ (.Y(_2665_),
    .A(net723),
    .B(_2663_));
 sg13g2_a21oi_1 _7027_ (.A1(net724),
    .A2(_2662_),
    .Y(_2666_),
    .B1(net775));
 sg13g2_nand2_1 _7028_ (.Y(_2667_),
    .A(net848),
    .B(_1896_));
 sg13g2_xor2_1 _7029_ (.B(_1895_),
    .A(net848),
    .X(_2668_));
 sg13g2_nand2_1 _7030_ (.Y(_2669_),
    .A(\r1[0] ),
    .B(_2652_));
 sg13g2_a21o_1 _7031_ (.A2(_2669_),
    .A1(_2651_),
    .B1(_2668_),
    .X(_2670_));
 sg13g2_nand3_1 _7032_ (.B(_2668_),
    .C(_2669_),
    .A(_2651_),
    .Y(_2671_));
 sg13g2_a21o_1 _7033_ (.A2(_2671_),
    .A1(_2670_),
    .B1(net742),
    .X(_2672_));
 sg13g2_a21oi_1 _7034_ (.A1(net742),
    .A2(_2663_),
    .Y(_2673_),
    .B1(net778));
 sg13g2_a22oi_1 _7035_ (.Y(_2674_),
    .B1(_2672_),
    .B2(_2673_),
    .A2(_2666_),
    .A1(_2665_));
 sg13g2_nor2_1 _7036_ (.A(net923),
    .B(_2674_),
    .Y(_0139_));
 sg13g2_nand2_1 _7037_ (.Y(_2676_),
    .A(net874),
    .B(net847));
 sg13g2_xnor2_1 _7038_ (.Y(_2677_),
    .A(net874),
    .B(\r1[3] ));
 sg13g2_a21oi_1 _7039_ (.A1(_2660_),
    .A2(_2661_),
    .Y(_2678_),
    .B1(_2659_));
 sg13g2_xor2_1 _7040_ (.B(_2678_),
    .A(_2677_),
    .X(_2679_));
 sg13g2_nand2b_1 _7041_ (.Y(_2680_),
    .B(net847),
    .A_N(net824));
 sg13g2_a21oi_1 _7042_ (.A1(net723),
    .A2(_2680_),
    .Y(_2681_),
    .B1(net775));
 sg13g2_o21ai_1 _7043_ (.B1(_2681_),
    .Y(_2682_),
    .A1(net722),
    .A2(_2679_));
 sg13g2_xor2_1 _7044_ (.B(_1893_),
    .A(net847),
    .X(_2683_));
 sg13g2_a21oi_1 _7045_ (.A1(_2667_),
    .A2(_2670_),
    .Y(_2684_),
    .B1(_2683_));
 sg13g2_and3_1 _7046_ (.X(_2686_),
    .A(_2667_),
    .B(_2670_),
    .C(_2683_));
 sg13g2_o21ai_1 _7047_ (.B1(net744),
    .Y(_2687_),
    .A1(_2684_),
    .A2(_2686_));
 sg13g2_a21oi_1 _7048_ (.A1(net742),
    .A2(_2680_),
    .Y(_2688_),
    .B1(net779));
 sg13g2_nand2_1 _7049_ (.Y(_2689_),
    .A(_2687_),
    .B(_2688_));
 sg13g2_a21oi_1 _7050_ (.A1(_2682_),
    .A2(_2689_),
    .Y(_0140_),
    .B1(net923));
 sg13g2_nor2b_1 _7051_ (.A(net867),
    .B_N(\r1[4] ),
    .Y(_2690_));
 sg13g2_xnor2_1 _7052_ (.Y(_2691_),
    .A(net867),
    .B(net846));
 sg13g2_o21ai_1 _7053_ (.B1(_2676_),
    .Y(_2692_),
    .A1(_2677_),
    .A2(_2678_));
 sg13g2_xor2_1 _7054_ (.B(_2692_),
    .A(_2691_),
    .X(_2693_));
 sg13g2_nand2b_1 _7055_ (.Y(_2694_),
    .B(net846),
    .A_N(net823));
 sg13g2_a21oi_1 _7056_ (.A1(net722),
    .A2(_2694_),
    .Y(_2696_),
    .B1(net775));
 sg13g2_o21ai_1 _7057_ (.B1(_2696_),
    .Y(_2697_),
    .A1(net722),
    .A2(_2693_));
 sg13g2_xnor2_1 _7058_ (.Y(_2698_),
    .A(net846),
    .B(_3573_));
 sg13g2_a21oi_1 _7059_ (.A1(net847),
    .A2(_1894_),
    .Y(_2699_),
    .B1(_2684_));
 sg13g2_nor2_1 _7060_ (.A(_2698_),
    .B(_2699_),
    .Y(_2700_));
 sg13g2_xor2_1 _7061_ (.B(_2699_),
    .A(_2698_),
    .X(_2701_));
 sg13g2_a21oi_1 _7062_ (.A1(net742),
    .A2(_2694_),
    .Y(_2702_),
    .B1(net779));
 sg13g2_o21ai_1 _7063_ (.B1(_2702_),
    .Y(_2703_),
    .A1(net742),
    .A2(_2701_));
 sg13g2_a21oi_1 _7064_ (.A1(_2697_),
    .A2(_2703_),
    .Y(_0141_),
    .B1(net920));
 sg13g2_a21oi_1 _7065_ (.A1(net846),
    .A2(_3573_),
    .Y(_2704_),
    .B1(_2700_));
 sg13g2_nor2_1 _7066_ (.A(net845),
    .B(_1862_),
    .Y(_2706_));
 sg13g2_nand2_1 _7067_ (.Y(_2707_),
    .A(net845),
    .B(_1862_));
 sg13g2_nand2b_1 _7068_ (.Y(_2708_),
    .B(_2707_),
    .A_N(_2706_));
 sg13g2_a21oi_1 _7069_ (.A1(_2704_),
    .A2(_2708_),
    .Y(_2709_),
    .B1(net742));
 sg13g2_o21ai_1 _7070_ (.B1(_2709_),
    .Y(_2710_),
    .A1(_2704_),
    .A2(_2708_));
 sg13g2_nor2b_1 _7071_ (.A(net823),
    .B_N(net845),
    .Y(_2711_));
 sg13g2_a21oi_1 _7072_ (.A1(net742),
    .A2(_2711_),
    .Y(_2712_),
    .B1(net779));
 sg13g2_a21oi_1 _7073_ (.A1(_2691_),
    .A2(_2692_),
    .Y(_2713_),
    .B1(_2690_));
 sg13g2_nand2_1 _7074_ (.Y(_2714_),
    .A(net845),
    .B(net807));
 sg13g2_nor2_1 _7075_ (.A(net845),
    .B(net807),
    .Y(_2715_));
 sg13g2_xnor2_1 _7076_ (.Y(_2717_),
    .A(net845),
    .B(net810));
 sg13g2_xnor2_1 _7077_ (.Y(_2718_),
    .A(_2713_),
    .B(_2717_));
 sg13g2_nand2_1 _7078_ (.Y(_2719_),
    .A(net724),
    .B(_2718_));
 sg13g2_a21oi_1 _7079_ (.A1(net722),
    .A2(_2711_),
    .Y(_2720_),
    .B1(net775));
 sg13g2_a221oi_1 _7080_ (.B2(_2720_),
    .C1(net920),
    .B1(_2719_),
    .A1(_2710_),
    .Y(_0142_),
    .A2(_2712_));
 sg13g2_or2_1 _7081_ (.X(_2721_),
    .B(_2715_),
    .A(_2713_));
 sg13g2_nand2_1 _7082_ (.Y(_2722_),
    .A(_2714_),
    .B(_2721_));
 sg13g2_xnor2_1 _7083_ (.Y(_2723_),
    .A(\r1[6] ),
    .B(net146));
 sg13g2_a21oi_1 _7084_ (.A1(_2714_),
    .A2(_2721_),
    .Y(_2724_),
    .B1(_2723_));
 sg13g2_xnor2_1 _7085_ (.Y(_2725_),
    .A(_2722_),
    .B(_2723_));
 sg13g2_nand2b_1 _7086_ (.Y(_2727_),
    .B(\r1[6] ),
    .A_N(net823));
 sg13g2_a21oi_1 _7087_ (.A1(net722),
    .A2(_2727_),
    .Y(_2728_),
    .B1(net775));
 sg13g2_o21ai_1 _7088_ (.B1(_2728_),
    .Y(_2729_),
    .A1(net722),
    .A2(_2725_));
 sg13g2_or2_1 _7089_ (.X(_2730_),
    .B(_2706_),
    .A(_2704_));
 sg13g2_xnor2_1 _7090_ (.Y(_2731_),
    .A(\r1[6] ),
    .B(_1945_));
 sg13g2_a21oi_1 _7091_ (.A1(_2707_),
    .A2(_2730_),
    .Y(_2732_),
    .B1(_2731_));
 sg13g2_and3_1 _7092_ (.X(_2733_),
    .A(_2707_),
    .B(_2730_),
    .C(_2731_));
 sg13g2_o21ai_1 _7093_ (.B1(net744),
    .Y(_2734_),
    .A1(_2732_),
    .A2(_2733_));
 sg13g2_a21oi_1 _7094_ (.A1(net743),
    .A2(_2727_),
    .Y(_2735_),
    .B1(net779));
 sg13g2_nand2_1 _7095_ (.Y(_2736_),
    .A(_2734_),
    .B(_2735_));
 sg13g2_a21oi_1 _7096_ (.A1(_2729_),
    .A2(_2736_),
    .Y(_0143_),
    .B1(net920));
 sg13g2_nand2_1 _7097_ (.Y(_2738_),
    .A(_2820_),
    .B(net805));
 sg13g2_xnor2_1 _7098_ (.Y(_2739_),
    .A(_0040_),
    .B(net805));
 sg13g2_a21oi_1 _7099_ (.A1(_2831_),
    .A2(net147),
    .Y(_2740_),
    .B1(_2724_));
 sg13g2_nand2b_1 _7100_ (.Y(_2741_),
    .B(_2739_),
    .A_N(_2740_));
 sg13g2_xnor2_1 _7101_ (.Y(_2742_),
    .A(_2739_),
    .B(_2740_));
 sg13g2_nand2b_1 _7102_ (.Y(_2743_),
    .B(net285),
    .A_N(net822));
 sg13g2_a21oi_1 _7103_ (.A1(net722),
    .A2(_2743_),
    .Y(_2744_),
    .B1(_3106_));
 sg13g2_o21ai_1 _7104_ (.B1(_2744_),
    .Y(_2745_),
    .A1(net722),
    .A2(_2742_));
 sg13g2_nand2_1 _7105_ (.Y(_2746_),
    .A(\r1[7] ),
    .B(_2008_));
 sg13g2_xor2_1 _7106_ (.B(_2008_),
    .A(\r1[7] ),
    .X(_2748_));
 sg13g2_a21oi_1 _7107_ (.A1(_2831_),
    .A2(_1945_),
    .Y(_2749_),
    .B1(_2732_));
 sg13g2_nand2b_1 _7108_ (.Y(_2750_),
    .B(_2748_),
    .A_N(_2749_));
 sg13g2_xnor2_1 _7109_ (.Y(_2751_),
    .A(_2748_),
    .B(_2749_));
 sg13g2_a21oi_1 _7110_ (.A1(net743),
    .A2(_2743_),
    .Y(_2752_),
    .B1(net779));
 sg13g2_o21ai_1 _7111_ (.B1(_2752_),
    .Y(_2753_),
    .A1(net743),
    .A2(_2751_));
 sg13g2_a21oi_1 _7112_ (.A1(_2745_),
    .A2(_2753_),
    .Y(_0144_),
    .B1(net920));
 sg13g2_a21oi_2 _7113_ (.B1(_3594_),
    .Y(_2754_),
    .A2(_2741_),
    .A1(_2738_));
 sg13g2_nand3_1 _7114_ (.B(_2738_),
    .C(_2741_),
    .A(_3594_),
    .Y(_2755_));
 sg13g2_nor2b_1 _7115_ (.A(_2754_),
    .B_N(_2755_),
    .Y(_2756_));
 sg13g2_nand2b_1 _7116_ (.Y(_2758_),
    .B(net273),
    .A_N(net822));
 sg13g2_a21oi_1 _7117_ (.A1(net723),
    .A2(_2758_),
    .Y(_2759_),
    .B1(net774));
 sg13g2_o21ai_1 _7118_ (.B1(_2759_),
    .Y(_2760_),
    .A1(net723),
    .A2(_2756_));
 sg13g2_xnor2_1 _7119_ (.Y(_2761_),
    .A(\r1[8] ),
    .B(_2213_));
 sg13g2_and3_1 _7120_ (.X(_2762_),
    .A(_2746_),
    .B(_2750_),
    .C(_2761_));
 sg13g2_a21oi_1 _7121_ (.A1(_2746_),
    .A2(_2750_),
    .Y(_2763_),
    .B1(_2761_));
 sg13g2_nor2_1 _7122_ (.A(_2762_),
    .B(_2763_),
    .Y(_2764_));
 sg13g2_a21oi_1 _7123_ (.A1(net741),
    .A2(_2758_),
    .Y(_2765_),
    .B1(net777));
 sg13g2_o21ai_1 _7124_ (.B1(_2765_),
    .Y(_2766_),
    .A1(net741),
    .A2(_2764_));
 sg13g2_a21oi_1 _7125_ (.A1(_2760_),
    .A2(_2766_),
    .Y(_0145_),
    .B1(net919));
 sg13g2_a21oi_1 _7126_ (.A1(_2810_),
    .A2(_2213_),
    .Y(_2768_),
    .B1(_2763_));
 sg13g2_o21ai_1 _7127_ (.B1(_2212_),
    .Y(_2769_),
    .A1(_2204_),
    .A2(_2210_));
 sg13g2_o21ai_1 _7128_ (.B1(_2208_),
    .Y(_2770_),
    .A1(net826),
    .A2(_2205_));
 sg13g2_nand3_1 _7129_ (.B(\hvsync_gen.vpos[8] ),
    .C(_3584_),
    .A(net826),
    .Y(_2771_));
 sg13g2_nand2_1 _7130_ (.Y(_2772_),
    .A(\hvsync_gen.vpos[8] ),
    .B(net805));
 sg13g2_or2_1 _7131_ (.X(_2773_),
    .B(\hvsync_gen.vpos[8] ),
    .A(net826));
 sg13g2_o21ai_1 _7132_ (.B1(_2772_),
    .Y(_2774_),
    .A1(net805),
    .A2(_2773_));
 sg13g2_nor2b_1 _7133_ (.A(_2774_),
    .B_N(_2771_),
    .Y(_2775_));
 sg13g2_xnor2_1 _7134_ (.Y(_2776_),
    .A(net761),
    .B(_2775_));
 sg13g2_inv_1 _7135_ (.Y(_2777_),
    .A(_2776_));
 sg13g2_xnor2_1 _7136_ (.Y(_2779_),
    .A(_2770_),
    .B(_2777_));
 sg13g2_nor2b_1 _7137_ (.A(_2779_),
    .B_N(_2769_),
    .Y(_2780_));
 sg13g2_xnor2_1 _7138_ (.Y(_2781_),
    .A(_2769_),
    .B(_2779_));
 sg13g2_nand2_1 _7139_ (.Y(_2782_),
    .A(\r1[9] ),
    .B(_2781_));
 sg13g2_xnor2_1 _7140_ (.Y(_2783_),
    .A(\r1[9] ),
    .B(_2781_));
 sg13g2_or2_1 _7141_ (.X(_2784_),
    .B(_2783_),
    .A(_2768_));
 sg13g2_a21oi_1 _7142_ (.A1(_2768_),
    .A2(_2783_),
    .Y(_2785_),
    .B1(net741));
 sg13g2_nor2b_1 _7143_ (.A(net822),
    .B_N(net293),
    .Y(_2786_));
 sg13g2_a22oi_1 _7144_ (.Y(_2787_),
    .B1(_2786_),
    .B2(net741),
    .A2(_2785_),
    .A1(_2784_));
 sg13g2_nor2_1 _7145_ (.A(_3588_),
    .B(_2754_),
    .Y(_2788_));
 sg13g2_xnor2_1 _7146_ (.Y(_2790_),
    .A(_2789_),
    .B(_2788_));
 sg13g2_nand2_1 _7147_ (.Y(_2791_),
    .A(net724),
    .B(_2790_));
 sg13g2_a21oi_1 _7148_ (.A1(net723),
    .A2(_2786_),
    .Y(_2792_),
    .B1(net774));
 sg13g2_a221oi_1 _7149_ (.B2(_2792_),
    .C1(net919),
    .B1(_2791_),
    .A1(net774),
    .Y(_0146_),
    .A2(_2787_));
 sg13g2_a22oi_1 _7150_ (.Y(_2793_),
    .B1(_2754_),
    .B2(\r1[9] ),
    .A2(_3588_),
    .A1(_2789_));
 sg13g2_xnor2_1 _7151_ (.Y(_2794_),
    .A(_2799_),
    .B(_2793_));
 sg13g2_nand2b_1 _7152_ (.Y(_2795_),
    .B(net276),
    .A_N(net821));
 sg13g2_a21oi_1 _7153_ (.A1(net721),
    .A2(_2795_),
    .Y(_2796_),
    .B1(net773));
 sg13g2_o21ai_1 _7154_ (.B1(_2796_),
    .Y(_2797_),
    .A1(net721),
    .A2(_2794_));
 sg13g2_nand2_1 _7155_ (.Y(_2798_),
    .A(_2782_),
    .B(_2784_));
 sg13g2_a21oi_1 _7156_ (.A1(_2770_),
    .A2(_2777_),
    .Y(_2800_),
    .B1(_2780_));
 sg13g2_xor2_1 _7157_ (.B(_2772_),
    .A(\hvsync_gen.vpos[9] ),
    .X(_2801_));
 sg13g2_nor2_1 _7158_ (.A(net761),
    .B(_2771_),
    .Y(_2802_));
 sg13g2_a21oi_1 _7159_ (.A1(net761),
    .A2(_2774_),
    .Y(_2803_),
    .B1(_2802_));
 sg13g2_xnor2_1 _7160_ (.Y(_2804_),
    .A(_2801_),
    .B(_2803_));
 sg13g2_xnor2_1 _7161_ (.Y(_2805_),
    .A(_2800_),
    .B(_2804_));
 sg13g2_inv_1 _7162_ (.Y(_2806_),
    .A(net711));
 sg13g2_xnor2_1 _7163_ (.Y(_2807_),
    .A(_2778_),
    .B(net712));
 sg13g2_xnor2_1 _7164_ (.Y(_2808_),
    .A(_2798_),
    .B(_2807_));
 sg13g2_nand2_1 _7165_ (.Y(_2809_),
    .A(net744),
    .B(_2808_));
 sg13g2_a21oi_1 _7166_ (.A1(net740),
    .A2(_2795_),
    .Y(_2811_),
    .B1(net776));
 sg13g2_nand2_1 _7167_ (.Y(_2812_),
    .A(_2809_),
    .B(_2811_));
 sg13g2_a21oi_1 _7168_ (.A1(_2797_),
    .A2(_2812_),
    .Y(_0147_),
    .B1(net919));
 sg13g2_nand2b_1 _7169_ (.Y(_2813_),
    .B(net843),
    .A_N(net821));
 sg13g2_nand2_1 _7170_ (.Y(_2814_),
    .A(net811),
    .B(_2813_));
 sg13g2_nand2_1 _7171_ (.Y(_2815_),
    .A(net740),
    .B(_2814_));
 sg13g2_a22oi_1 _7172_ (.Y(_2816_),
    .B1(_2807_),
    .B2(_2798_),
    .A2(net712),
    .A1(_2799_));
 sg13g2_nor2_1 _7173_ (.A(net843),
    .B(net712),
    .Y(_2817_));
 sg13g2_nand2_1 _7174_ (.Y(_2818_),
    .A(net843),
    .B(net712));
 sg13g2_nand2b_1 _7175_ (.Y(_2819_),
    .B(_2818_),
    .A_N(_2817_));
 sg13g2_o21ai_1 _7176_ (.B1(net744),
    .Y(_2821_),
    .A1(_2816_),
    .A2(_2819_));
 sg13g2_a21o_1 _7177_ (.A2(_2819_),
    .A1(_2816_),
    .B1(_2821_),
    .X(_2822_));
 sg13g2_a221oi_1 _7178_ (.B2(_2822_),
    .C1(net776),
    .B1(_2815_),
    .A1(net798),
    .Y(_2823_),
    .A2(_2813_));
 sg13g2_nand3b_1 _7179_ (.B(\r1[10] ),
    .C(net843),
    .Y(_2824_),
    .A_N(_2793_));
 sg13g2_nor2_1 _7180_ (.A(_2778_),
    .B(_2793_),
    .Y(_2825_));
 sg13g2_nor2_1 _7181_ (.A(net721),
    .B(_2824_),
    .Y(_2826_));
 sg13g2_nand2_2 _7182_ (.Y(_2827_),
    .A(net819),
    .B(net721));
 sg13g2_a22oi_1 _7183_ (.Y(_2828_),
    .B1(_2827_),
    .B2(net843),
    .A2(_2825_),
    .A1(net724));
 sg13g2_nor3_1 _7184_ (.A(net773),
    .B(_2826_),
    .C(_2828_),
    .Y(_2829_));
 sg13g2_o21ai_1 _7185_ (.B1(net925),
    .Y(_2830_),
    .A1(_2823_),
    .A2(_2829_));
 sg13g2_inv_1 _7186_ (.Y(_0148_),
    .A(_2830_));
 sg13g2_xor2_1 _7187_ (.B(net711),
    .A(\r1[12] ),
    .X(_2832_));
 sg13g2_o21ai_1 _7188_ (.B1(_2818_),
    .Y(_2833_),
    .A1(_2816_),
    .A2(_2817_));
 sg13g2_nor2b_1 _7189_ (.A(net819),
    .B_N(net277),
    .Y(_2834_));
 sg13g2_a21oi_1 _7190_ (.A1(net739),
    .A2(_2834_),
    .Y(_2835_),
    .B1(net776));
 sg13g2_xor2_1 _7191_ (.B(_2833_),
    .A(_2832_),
    .X(_2836_));
 sg13g2_nand2_1 _7192_ (.Y(_2837_),
    .A(net744),
    .B(_2836_));
 sg13g2_xnor2_1 _7193_ (.Y(_2838_),
    .A(_2871_),
    .B(_2824_));
 sg13g2_nand2_1 _7194_ (.Y(_2839_),
    .A(net721),
    .B(_2834_));
 sg13g2_a21oi_1 _7195_ (.A1(net724),
    .A2(_2838_),
    .Y(_2840_),
    .B1(net773));
 sg13g2_a221oi_1 _7196_ (.B2(_2840_),
    .C1(net919),
    .B1(_2839_),
    .A1(_2835_),
    .Y(_0149_),
    .A2(_2837_));
 sg13g2_a22oi_1 _7197_ (.Y(_2842_),
    .B1(_2832_),
    .B2(_2833_),
    .A2(net711),
    .A1(_2871_));
 sg13g2_nand2_1 _7198_ (.Y(_2843_),
    .A(net842),
    .B(net711));
 sg13g2_nor2_1 _7199_ (.A(net842),
    .B(net711),
    .Y(_2844_));
 sg13g2_xnor2_1 _7200_ (.Y(_2845_),
    .A(net842),
    .B(net711));
 sg13g2_xnor2_1 _7201_ (.Y(_2846_),
    .A(_2842_),
    .B(_2845_));
 sg13g2_nor2b_1 _7202_ (.A(net819),
    .B_N(net842),
    .Y(_2847_));
 sg13g2_a21oi_1 _7203_ (.A1(net739),
    .A2(_2847_),
    .Y(_2848_),
    .B1(net776));
 sg13g2_o21ai_1 _7204_ (.B1(_2848_),
    .Y(_2849_),
    .A1(net739),
    .A2(_2846_));
 sg13g2_a22oi_1 _7205_ (.Y(_2850_),
    .B1(_2827_),
    .B2(net842),
    .A2(_2826_),
    .A1(net277));
 sg13g2_nor3_2 _7206_ (.A(_0410_),
    .B(net721),
    .C(_2824_),
    .Y(_2852_));
 sg13g2_o21ai_1 _7207_ (.B1(net776),
    .Y(_2853_),
    .A1(_2850_),
    .A2(_2852_));
 sg13g2_and3_1 _7208_ (.X(_0150_),
    .A(net925),
    .B(_2849_),
    .C(_2853_));
 sg13g2_a21oi_1 _7209_ (.A1(net290),
    .A2(_2827_),
    .Y(_2854_),
    .B1(_2852_));
 sg13g2_a21oi_1 _7210_ (.A1(net290),
    .A2(_2852_),
    .Y(_2855_),
    .B1(net773));
 sg13g2_nand2b_1 _7211_ (.Y(_2856_),
    .B(_2855_),
    .A_N(_2854_));
 sg13g2_xor2_1 _7212_ (.B(net711),
    .A(\r1[14] ),
    .X(_2857_));
 sg13g2_o21ai_1 _7213_ (.B1(_2843_),
    .Y(_2858_),
    .A1(_2842_),
    .A2(_2844_));
 sg13g2_nand2_1 _7214_ (.Y(_2859_),
    .A(_2857_),
    .B(_2858_));
 sg13g2_xor2_1 _7215_ (.B(_2858_),
    .A(_2857_),
    .X(_2860_));
 sg13g2_nand2b_1 _7216_ (.Y(_2862_),
    .B(\r1[14] ),
    .A_N(net819));
 sg13g2_a21oi_1 _7217_ (.A1(net739),
    .A2(_2862_),
    .Y(_2863_),
    .B1(net776));
 sg13g2_o21ai_1 _7218_ (.B1(_2863_),
    .Y(_2864_),
    .A1(net739),
    .A2(_2860_));
 sg13g2_a21oi_1 _7219_ (.A1(_2856_),
    .A2(_2864_),
    .Y(_0151_),
    .B1(net919));
 sg13g2_o21ai_1 _7220_ (.B1(_2859_),
    .Y(_2865_),
    .A1(_0042_),
    .A2(_2806_));
 sg13g2_xor2_1 _7221_ (.B(net711),
    .A(\r1[15] ),
    .X(_2866_));
 sg13g2_nand2_1 _7222_ (.Y(_2867_),
    .A(_2865_),
    .B(_2866_));
 sg13g2_o21ai_1 _7223_ (.B1(net744),
    .Y(_2868_),
    .A1(_2865_),
    .A2(_2866_));
 sg13g2_nor2b_1 _7224_ (.A(_2868_),
    .B_N(_2867_),
    .Y(_2869_));
 sg13g2_nand2b_1 _7225_ (.Y(_2870_),
    .B(\r1[15] ),
    .A_N(net821));
 sg13g2_o21ai_1 _7226_ (.B1(net766),
    .Y(_2872_),
    .A1(net744),
    .A2(_2870_));
 sg13g2_a21oi_1 _7227_ (.A1(net752),
    .A2(_2870_),
    .Y(_2873_),
    .B1(net776));
 sg13g2_o21ai_1 _7228_ (.B1(_2873_),
    .Y(_2874_),
    .A1(_2869_),
    .A2(_2872_));
 sg13g2_nor2b_1 _7229_ (.A(net282),
    .B_N(_2852_),
    .Y(_2875_));
 sg13g2_a21oi_1 _7230_ (.A1(\r1[15] ),
    .A2(_2827_),
    .Y(_2876_),
    .B1(_2875_));
 sg13g2_a21oi_1 _7231_ (.A1(\r1[15] ),
    .A2(_2875_),
    .Y(_2877_),
    .B1(net773));
 sg13g2_nand2b_1 _7232_ (.Y(_2878_),
    .B(_2877_),
    .A_N(_2876_));
 sg13g2_a21oi_1 _7233_ (.A1(_2874_),
    .A2(net283),
    .Y(_0152_),
    .B1(net919));
 sg13g2_o21ai_1 _7234_ (.B1(_2867_),
    .Y(_2879_),
    .A1(_0036_),
    .A2(_2806_));
 sg13g2_xnor2_1 _7235_ (.Y(_2880_),
    .A(_2979_),
    .B(net712));
 sg13g2_nor2_1 _7236_ (.A(_2879_),
    .B(_2880_),
    .Y(_2882_));
 sg13g2_a21o_1 _7237_ (.A2(_2880_),
    .A1(_2879_),
    .B1(net739),
    .X(_2883_));
 sg13g2_nor2_1 _7238_ (.A(_2882_),
    .B(_2883_),
    .Y(_2884_));
 sg13g2_nor2_1 _7239_ (.A(_2979_),
    .B(net819),
    .Y(_2885_));
 sg13g2_a21oi_1 _7240_ (.A1(net740),
    .A2(_2885_),
    .Y(_2886_),
    .B1(_2884_));
 sg13g2_nand4_1 _7241_ (.B(\r1[14] ),
    .C(net842),
    .A(\r1[15] ),
    .Y(_2887_),
    .D(\r1[12] ));
 sg13g2_nor2_1 _7242_ (.A(_2824_),
    .B(_2887_),
    .Y(_2888_));
 sg13g2_xnor2_1 _7243_ (.Y(_2889_),
    .A(net250),
    .B(_2888_));
 sg13g2_nand2_1 _7244_ (.Y(_2890_),
    .A(net724),
    .B(_2889_));
 sg13g2_a21oi_1 _7245_ (.A1(net721),
    .A2(_2885_),
    .Y(_2891_),
    .B1(net773));
 sg13g2_a221oi_1 _7246_ (.B2(_2891_),
    .C1(net919),
    .B1(_2890_),
    .A1(net773),
    .Y(_0153_),
    .A2(_2886_));
 sg13g2_nor3_1 _7247_ (.A(_2419_),
    .B(_2824_),
    .C(_2887_),
    .Y(_2893_));
 sg13g2_o21ai_1 _7248_ (.B1(net724),
    .Y(_2894_),
    .A1(_2989_),
    .A2(_2888_));
 sg13g2_nand2b_1 _7249_ (.Y(_2895_),
    .B(net248),
    .A_N(net819));
 sg13g2_a21oi_1 _7250_ (.A1(net721),
    .A2(_2895_),
    .Y(_2896_),
    .B1(net773));
 sg13g2_o21ai_1 _7251_ (.B1(_2896_),
    .Y(_2897_),
    .A1(_2893_),
    .A2(_2894_));
 sg13g2_nand2_1 _7252_ (.Y(_2898_),
    .A(_0014_),
    .B(net712));
 sg13g2_or4_1 _7253_ (.A(_2979_),
    .B(net739),
    .C(net712),
    .D(_2867_),
    .X(_2899_));
 sg13g2_o21ai_1 _7254_ (.B1(_2899_),
    .Y(_2900_),
    .A1(_2883_),
    .A2(_2898_));
 sg13g2_a21oi_1 _7255_ (.A1(net819),
    .A2(net739),
    .Y(_2901_),
    .B1(_2989_));
 sg13g2_a21oi_1 _7256_ (.A1(net248),
    .A2(_2900_),
    .Y(_2903_),
    .B1(net776));
 sg13g2_o21ai_1 _7257_ (.B1(_2903_),
    .Y(_2904_),
    .A1(_2900_),
    .A2(_2901_));
 sg13g2_a21oi_1 _7258_ (.A1(_2897_),
    .A2(_2904_),
    .Y(_0154_),
    .B1(net919));
 sg13g2_and2_1 _7259_ (.A(net929),
    .B(_3512_),
    .X(_2905_));
 sg13g2_nand2_2 _7260_ (.Y(_2906_),
    .A(net929),
    .B(_3512_));
 sg13g2_nor2_1 _7261_ (.A(net170),
    .B(_3125_),
    .Y(_2907_));
 sg13g2_nor2_1 _7262_ (.A(\title_r[0] ),
    .B(net795),
    .Y(_2908_));
 sg13g2_nor3_1 _7263_ (.A(_2906_),
    .B(_2907_),
    .C(_2908_),
    .Y(_0155_));
 sg13g2_xor2_1 _7264_ (.B(net916),
    .A(\title_r[1] ),
    .X(_2909_));
 sg13g2_xnor2_1 _7265_ (.Y(_2910_),
    .A(net170),
    .B(_2909_));
 sg13g2_nand3_1 _7266_ (.B(net752),
    .C(_2910_),
    .A(net841),
    .Y(_2912_));
 sg13g2_a22oi_1 _7267_ (.Y(_2913_),
    .B1(_2910_),
    .B2(net795),
    .A2(net752),
    .A1(net841));
 sg13g2_inv_1 _7268_ (.Y(_2914_),
    .A(_2913_));
 sg13g2_a22oi_1 _7269_ (.Y(_2915_),
    .B1(_2912_),
    .B2(_2914_),
    .A2(_3125_),
    .A1(net215));
 sg13g2_nor2_1 _7270_ (.A(_2906_),
    .B(_2915_),
    .Y(_0156_));
 sg13g2_o21ai_1 _7271_ (.B1(_3470_),
    .Y(_2916_),
    .A1(_3471_),
    .A2(_3472_));
 sg13g2_a21oi_1 _7272_ (.A1(_3473_),
    .A2(_2916_),
    .Y(_2917_),
    .B1(net764));
 sg13g2_o21ai_1 _7273_ (.B1(_3424_),
    .Y(_2918_),
    .A1(_3425_),
    .A2(_3426_));
 sg13g2_nor2b_1 _7274_ (.A(_3427_),
    .B_N(_2918_),
    .Y(_2919_));
 sg13g2_nand2_2 _7275_ (.Y(_2920_),
    .A(net793),
    .B(net764));
 sg13g2_nor2_1 _7276_ (.A(net220),
    .B(net793),
    .Y(_2922_));
 sg13g2_o21ai_1 _7277_ (.B1(net734),
    .Y(_2923_),
    .A1(_2919_),
    .A2(_2920_));
 sg13g2_nor3_1 _7278_ (.A(_2917_),
    .B(_2922_),
    .C(_2923_),
    .Y(_0157_));
 sg13g2_or3_1 _7279_ (.A(_3422_),
    .B(_3423_),
    .C(_3427_),
    .X(_2924_));
 sg13g2_nand3_1 _7280_ (.B(_3428_),
    .C(_2924_),
    .A(net764),
    .Y(_2925_));
 sg13g2_nand2_1 _7281_ (.Y(_2926_),
    .A(_3473_),
    .B(_3474_));
 sg13g2_nor2_1 _7282_ (.A(net764),
    .B(_3475_),
    .Y(_2927_));
 sg13g2_a21oi_1 _7283_ (.A1(_2926_),
    .A2(_2927_),
    .Y(_2928_),
    .B1(_3125_));
 sg13g2_o21ai_1 _7284_ (.B1(net734),
    .Y(_2929_),
    .A1(net240),
    .A2(net794));
 sg13g2_a21oi_1 _7285_ (.A1(_2925_),
    .A2(_2928_),
    .Y(_0158_),
    .B1(_2929_));
 sg13g2_nand3_1 _7286_ (.B(_3428_),
    .C(_3429_),
    .A(_3421_),
    .Y(_2931_));
 sg13g2_a21oi_1 _7287_ (.A1(_3430_),
    .A2(_2931_),
    .Y(_2932_),
    .B1(_2920_));
 sg13g2_o21ai_1 _7288_ (.B1(net734),
    .Y(_2933_),
    .A1(net258),
    .A2(net793));
 sg13g2_or3_1 _7289_ (.A(_3469_),
    .B(_3475_),
    .C(_3477_),
    .X(_2934_));
 sg13g2_a21oi_1 _7290_ (.A1(_3478_),
    .A2(_2934_),
    .Y(_2935_),
    .B1(net764));
 sg13g2_nor3_1 _7291_ (.A(_2932_),
    .B(_2933_),
    .C(_2935_),
    .Y(_0159_));
 sg13g2_nand3_1 _7292_ (.B(_3420_),
    .C(_3430_),
    .A(_3419_),
    .Y(_2936_));
 sg13g2_a21oi_1 _7293_ (.A1(_3431_),
    .A2(_2936_),
    .Y(_2937_),
    .B1(_2920_));
 sg13g2_o21ai_1 _7294_ (.B1(net734),
    .Y(_2938_),
    .A1(net292),
    .A2(net794));
 sg13g2_and3_1 _7295_ (.X(_2939_),
    .A(_3466_),
    .B(_3478_),
    .C(_3479_));
 sg13g2_o21ai_1 _7296_ (.B1(net751),
    .Y(_2941_),
    .A1(_3480_),
    .A2(_2939_));
 sg13g2_nor2_1 _7297_ (.A(_2937_),
    .B(_2938_),
    .Y(_2942_));
 sg13g2_and2_1 _7298_ (.A(_2941_),
    .B(_2942_),
    .X(_0160_));
 sg13g2_nand3_1 _7299_ (.B(_3418_),
    .C(_3431_),
    .A(_3417_),
    .Y(_2943_));
 sg13g2_a21oi_1 _7300_ (.A1(_3432_),
    .A2(_2943_),
    .Y(_2944_),
    .B1(_2920_));
 sg13g2_o21ai_1 _7301_ (.B1(net735),
    .Y(_2945_),
    .A1(net253),
    .A2(net794));
 sg13g2_or3_1 _7302_ (.A(_3464_),
    .B(_3480_),
    .C(_3482_),
    .X(_2946_));
 sg13g2_a21oi_1 _7303_ (.A1(_3483_),
    .A2(_2946_),
    .Y(_2947_),
    .B1(net765));
 sg13g2_nor3_1 _7304_ (.A(_2944_),
    .B(_2945_),
    .C(_2947_),
    .Y(_0161_));
 sg13g2_nand3_1 _7305_ (.B(_3416_),
    .C(_3432_),
    .A(_3415_),
    .Y(_2948_));
 sg13g2_nor2b_1 _7306_ (.A(_3433_),
    .B_N(_2948_),
    .Y(_2950_));
 sg13g2_o21ai_1 _7307_ (.B1(net735),
    .Y(_2951_),
    .A1(net244),
    .A2(net794));
 sg13g2_and3_1 _7308_ (.X(_2952_),
    .A(_3461_),
    .B(_3483_),
    .C(_3484_));
 sg13g2_o21ai_1 _7309_ (.B1(net751),
    .Y(_2953_),
    .A1(_3485_),
    .A2(_2952_));
 sg13g2_o21ai_1 _7310_ (.B1(_2953_),
    .Y(_2954_),
    .A1(_2920_),
    .A2(_2950_));
 sg13g2_nor2_1 _7311_ (.A(_2951_),
    .B(_2954_),
    .Y(_0162_));
 sg13g2_or3_1 _7312_ (.A(_3414_),
    .B(_3433_),
    .C(_3435_),
    .X(_2955_));
 sg13g2_a21oi_1 _7313_ (.A1(_3436_),
    .A2(_2955_),
    .Y(_2956_),
    .B1(_2920_));
 sg13g2_o21ai_1 _7314_ (.B1(net735),
    .Y(_2957_),
    .A1(net247),
    .A2(net794));
 sg13g2_a21oi_1 _7315_ (.A1(\title_r[8] ),
    .A2(_3457_),
    .Y(_2958_),
    .B1(_3499_));
 sg13g2_nor2b_1 _7316_ (.A(_3486_),
    .B_N(_2958_),
    .Y(_2960_));
 sg13g2_xnor2_1 _7317_ (.Y(_2961_),
    .A(_3486_),
    .B(_2958_));
 sg13g2_nor2_1 _7318_ (.A(net764),
    .B(_2961_),
    .Y(_2962_));
 sg13g2_nor3_1 _7319_ (.A(_2956_),
    .B(_2957_),
    .C(_2962_),
    .Y(_0163_));
 sg13g2_nand2_1 _7320_ (.Y(_2963_),
    .A(_3434_),
    .B(_3436_));
 sg13g2_xnor2_1 _7321_ (.Y(_2964_),
    .A(_3413_),
    .B(_2963_));
 sg13g2_or3_1 _7322_ (.A(_3497_),
    .B(_3499_),
    .C(_2960_),
    .X(_2965_));
 sg13g2_and2_1 _7323_ (.A(_3497_),
    .B(_2960_),
    .X(_2966_));
 sg13g2_nand3_1 _7324_ (.B(_3500_),
    .C(_2965_),
    .A(net751),
    .Y(_2967_));
 sg13g2_o21ai_1 _7325_ (.B1(net793),
    .Y(_2968_),
    .A1(_2966_),
    .A2(_2967_));
 sg13g2_a21oi_1 _7326_ (.A1(net764),
    .A2(_2964_),
    .Y(_2970_),
    .B1(_2968_));
 sg13g2_o21ai_1 _7327_ (.B1(net735),
    .Y(_2971_),
    .A1(net242),
    .A2(net794));
 sg13g2_nor2_1 _7328_ (.A(_2970_),
    .B(_2971_),
    .Y(_0164_));
 sg13g2_o21ai_1 _7329_ (.B1(_3438_),
    .Y(_2972_),
    .A1(_3437_),
    .A2(_3442_));
 sg13g2_or3_1 _7330_ (.A(_3437_),
    .B(_3438_),
    .C(_3442_),
    .X(_2973_));
 sg13g2_a21oi_1 _7331_ (.A1(_2972_),
    .A2(_2973_),
    .Y(_2974_),
    .B1(_2920_));
 sg13g2_nand2_2 _7332_ (.Y(_2975_),
    .A(net793),
    .B(net734));
 sg13g2_nand2_1 _7333_ (.Y(_2976_),
    .A(net245),
    .B(net734));
 sg13g2_nor3_1 _7334_ (.A(_3501_),
    .B(_3502_),
    .C(_2966_),
    .Y(_2977_));
 sg13g2_o21ai_1 _7335_ (.B1(_3502_),
    .Y(_2978_),
    .A1(_3501_),
    .A2(_2966_));
 sg13g2_nand2b_1 _7336_ (.Y(_2980_),
    .B(_2978_),
    .A_N(_2977_));
 sg13g2_a221oi_1 _7337_ (.B2(net751),
    .C1(_2974_),
    .B1(_2980_),
    .A1(_2975_),
    .Y(_0165_),
    .A2(_2976_));
 sg13g2_o21ai_1 _7338_ (.B1(_2972_),
    .Y(_2981_),
    .A1(_2356_),
    .A2(net899));
 sg13g2_o21ai_1 _7339_ (.B1(net793),
    .Y(_2982_),
    .A1(_3439_),
    .A2(_2981_));
 sg13g2_a21oi_1 _7340_ (.A1(_3439_),
    .A2(_2981_),
    .Y(_2983_),
    .B1(_2982_));
 sg13g2_nor2_1 _7341_ (.A(net751),
    .B(_2983_),
    .Y(_2984_));
 sg13g2_nand2b_1 _7342_ (.Y(_2985_),
    .B(_2978_),
    .A_N(_3493_));
 sg13g2_xnor2_1 _7343_ (.Y(_2986_),
    .A(_3490_),
    .B(_2985_));
 sg13g2_a21oi_1 _7344_ (.A1(net751),
    .A2(_2986_),
    .Y(_2987_),
    .B1(_2984_));
 sg13g2_o21ai_1 _7345_ (.B1(net734),
    .Y(_2988_),
    .A1(net254),
    .A2(net793));
 sg13g2_nor2_1 _7346_ (.A(_2987_),
    .B(_2988_),
    .Y(_0166_));
 sg13g2_xnor2_1 _7347_ (.Y(_2990_),
    .A(_3412_),
    .B(_3445_));
 sg13g2_nor2_1 _7348_ (.A(_2920_),
    .B(_2990_),
    .Y(_2991_));
 sg13g2_nand2_1 _7349_ (.Y(_2992_),
    .A(net236),
    .B(net734));
 sg13g2_xnor2_1 _7350_ (.Y(_2993_),
    .A(_3455_),
    .B(_3506_));
 sg13g2_a221oi_1 _7351_ (.B2(net751),
    .C1(_2991_),
    .B1(_2993_),
    .A1(_2975_),
    .Y(_0167_),
    .A2(_2992_));
 sg13g2_nor2_1 _7352_ (.A(\title_r[8] ),
    .B(\title_r[7] ),
    .Y(_2994_));
 sg13g2_nor3_2 _7353_ (.A(\title_r[6] ),
    .B(\title_r[5] ),
    .C(\title_r[4] ),
    .Y(_2995_));
 sg13g2_nand3_1 _7354_ (.B(\title_r[10] ),
    .C(\title_r[9] ),
    .A(\title_r[11] ),
    .Y(_2996_));
 sg13g2_a21oi_1 _7355_ (.A1(_2994_),
    .A2(_2995_),
    .Y(_2997_),
    .B1(_2996_));
 sg13g2_o21ai_1 _7356_ (.B1(_2550_),
    .Y(_2999_),
    .A1(\title_r[12] ),
    .A2(_2997_));
 sg13g2_o21ai_1 _7357_ (.B1(_2633_),
    .Y(_3000_),
    .A1(_3048_),
    .A2(_3057_));
 sg13g2_nand3_1 _7358_ (.B(_2999_),
    .C(_3000_),
    .A(\hvsync_gen.hpos[9] ),
    .Y(_3001_));
 sg13g2_a21oi_2 _7359_ (.B1(_2975_),
    .Y(_3002_),
    .A2(_3001_),
    .A1(_3133_));
 sg13g2_nand3_1 _7360_ (.B(net765),
    .C(_3002_),
    .A(net160),
    .Y(_3003_));
 sg13g2_o21ai_1 _7361_ (.B1(_3003_),
    .Y(_0168_),
    .A1(_3007_),
    .A2(_3002_));
 sg13g2_and3_1 _7362_ (.X(_3004_),
    .A(net202),
    .B(\title_r_pixels_in_scanline[0] ),
    .C(_3002_));
 sg13g2_nor2_2 _7363_ (.A(net765),
    .B(_2906_),
    .Y(_3005_));
 sg13g2_a21oi_1 _7364_ (.A1(\title_r_pixels_in_scanline[0] ),
    .A2(_3002_),
    .Y(_3006_),
    .B1(net202));
 sg13g2_nor3_1 _7365_ (.A(_3004_),
    .B(_3005_),
    .C(net203),
    .Y(_0169_));
 sg13g2_and2_1 _7366_ (.A(net217),
    .B(_3004_),
    .X(_3008_));
 sg13g2_nor2_1 _7367_ (.A(net217),
    .B(_3004_),
    .Y(_3009_));
 sg13g2_nor3_1 _7368_ (.A(_3005_),
    .B(_3008_),
    .C(net218),
    .Y(_0170_));
 sg13g2_and2_1 _7369_ (.A(net232),
    .B(_3008_),
    .X(_3010_));
 sg13g2_nor2_1 _7370_ (.A(net232),
    .B(_3008_),
    .Y(_3011_));
 sg13g2_nor3_1 _7371_ (.A(_3005_),
    .B(_3010_),
    .C(_3011_),
    .Y(_0171_));
 sg13g2_nand2_1 _7372_ (.Y(_3012_),
    .A(\title_r_pixels_in_scanline[4] ),
    .B(_3010_));
 sg13g2_xnor2_1 _7373_ (.Y(_3013_),
    .A(net239),
    .B(_3010_));
 sg13g2_nor2_1 _7374_ (.A(_3005_),
    .B(_3013_),
    .Y(_0172_));
 sg13g2_xor2_1 _7375_ (.B(_3012_),
    .A(net227),
    .X(_3014_));
 sg13g2_nor2_1 _7376_ (.A(_3005_),
    .B(net228),
    .Y(_0173_));
 sg13g2_nor3_1 _7377_ (.A(net840),
    .B(net838),
    .C(\hvsync_gen.vpos[8] ),
    .Y(_3016_));
 sg13g2_nand4_1 _7378_ (.B(_3062_),
    .C(_2325_),
    .A(\hvsync_gen.vpos[9] ),
    .Y(_3017_),
    .D(_3016_));
 sg13g2_and2_1 _7379_ (.A(net929),
    .B(_3017_),
    .X(_3018_));
 sg13g2_inv_1 _7380_ (.Y(_3019_),
    .A(_3018_));
 sg13g2_nand2_2 _7381_ (.Y(_3020_),
    .A(_2517_),
    .B(_3018_));
 sg13g2_inv_1 _7382_ (.Y(_3021_),
    .A(_3020_));
 sg13g2_a22oi_1 _7383_ (.Y(_3022_),
    .B1(_3021_),
    .B2(net209),
    .A2(net745),
    .A1(net840));
 sg13g2_inv_1 _7384_ (.Y(_0174_),
    .A(net210));
 sg13g2_nor3_1 _7385_ (.A(_3063_),
    .B(_2567_),
    .C(_3020_),
    .Y(_3023_));
 sg13g2_a21o_1 _7386_ (.A2(net745),
    .A1(net838),
    .B1(_3023_),
    .X(_0175_));
 sg13g2_and3_1 _7387_ (.X(_3025_),
    .A(net840),
    .B(net838),
    .C(_2519_));
 sg13g2_o21ai_1 _7388_ (.B1(_2519_),
    .Y(_3026_),
    .A1(_2569_),
    .A2(_3019_));
 sg13g2_o21ai_1 _7389_ (.B1(_3026_),
    .Y(_3027_),
    .A1(net837),
    .A2(_3025_));
 sg13g2_inv_1 _7390_ (.Y(_0176_),
    .A(_3027_));
 sg13g2_and2_1 _7391_ (.A(net835),
    .B(_3026_),
    .X(_3028_));
 sg13g2_nor3_1 _7392_ (.A(net835),
    .B(_2644_),
    .C(net924),
    .Y(_3029_));
 sg13g2_a21o_1 _7393_ (.A2(_3029_),
    .A1(_3025_),
    .B1(_3028_),
    .X(_0177_));
 sg13g2_a21oi_1 _7394_ (.A1(_2325_),
    .A2(_3025_),
    .Y(_3030_),
    .B1(net833));
 sg13g2_nand3_1 _7395_ (.B(net833),
    .C(_2569_),
    .A(net835),
    .Y(_3031_));
 sg13g2_nor2_1 _7396_ (.A(net745),
    .B(_3031_),
    .Y(_3033_));
 sg13g2_a21oi_1 _7397_ (.A1(_2519_),
    .A2(_3019_),
    .Y(_3034_),
    .B1(_3033_));
 sg13g2_nor2b_1 _7398_ (.A(_3030_),
    .B_N(_3034_),
    .Y(_0178_));
 sg13g2_nor3_1 _7399_ (.A(net831),
    .B(_3020_),
    .C(_3031_),
    .Y(_3035_));
 sg13g2_a21o_1 _7400_ (.A2(_3034_),
    .A1(net831),
    .B1(_3035_),
    .X(_0179_));
 sg13g2_a21oi_1 _7401_ (.A1(net831),
    .A2(_3033_),
    .Y(_3036_),
    .B1(net830));
 sg13g2_a221oi_1 _7402_ (.B2(_2326_),
    .C1(_3036_),
    .B1(_3033_),
    .A1(_2519_),
    .Y(_0180_),
    .A2(_3019_));
 sg13g2_nand2_1 _7403_ (.Y(_3037_),
    .A(net827),
    .B(net745));
 sg13g2_nor3_1 _7404_ (.A(_2654_),
    .B(net237),
    .C(_3031_),
    .Y(_3038_));
 sg13g2_xnor2_1 _7405_ (.Y(_3039_),
    .A(net826),
    .B(_3038_));
 sg13g2_o21ai_1 _7406_ (.B1(_3037_),
    .Y(_0181_),
    .A1(_3020_),
    .A2(_3039_));
 sg13g2_a21oi_1 _7407_ (.A1(_3140_),
    .A2(_3018_),
    .Y(_3041_),
    .B1(_3034_));
 sg13g2_nand3_1 _7408_ (.B(_2326_),
    .C(_3033_),
    .A(net826),
    .Y(_3042_));
 sg13g2_a21oi_1 _7409_ (.A1(_2675_),
    .A2(_3042_),
    .Y(_0182_),
    .B1(_3041_));
 sg13g2_nand2b_1 _7410_ (.Y(_3043_),
    .B(net241),
    .A_N(_3041_));
 sg13g2_nand2_1 _7411_ (.Y(_3044_),
    .A(net929),
    .B(_3032_));
 sg13g2_o21ai_1 _7412_ (.B1(_3043_),
    .Y(_0183_),
    .A1(_3042_),
    .A2(_3044_));
 sg13g2_dfrbp_1 _7413_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net30),
    .D(_0061_),
    .Q_N(_3693_),
    .Q(\note2_freq[1] ));
 sg13g2_dfrbp_1 _7414_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net102),
    .D(_0062_),
    .Q_N(_3692_),
    .Q(\note_freq[1] ));
 sg13g2_dfrbp_1 _7415_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net101),
    .D(_0063_),
    .Q_N(_3691_),
    .Q(\r2[0] ));
 sg13g2_dfrbp_1 _7416_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net100),
    .D(_0064_),
    .Q_N(_0023_),
    .Q(\r2[1] ));
 sg13g2_dfrbp_1 _7417_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net99),
    .D(_0065_),
    .Q_N(_0054_),
    .Q(\r2[2] ));
 sg13g2_dfrbp_1 _7418_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net98),
    .D(_0066_),
    .Q_N(_3690_),
    .Q(\r2[3] ));
 sg13g2_dfrbp_1 _7419_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net97),
    .D(_0067_),
    .Q_N(_0052_),
    .Q(\r2[4] ));
 sg13g2_dfrbp_1 _7420_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net96),
    .D(_0068_),
    .Q_N(_3689_),
    .Q(\r2[5] ));
 sg13g2_dfrbp_1 _7421_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net95),
    .D(net272),
    .Q_N(_0051_),
    .Q(\r2[6] ));
 sg13g2_dfrbp_1 _7422_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net94),
    .D(_0070_),
    .Q_N(_3688_),
    .Q(\r2[7] ));
 sg13g2_dfrbp_1 _7423_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net93),
    .D(_0071_),
    .Q_N(_0050_),
    .Q(\r2[8] ));
 sg13g2_dfrbp_1 _7424_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net92),
    .D(_0072_),
    .Q_N(_0025_),
    .Q(\r2[9] ));
 sg13g2_dfrbp_1 _7425_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net91),
    .D(_0073_),
    .Q_N(_0049_),
    .Q(\r2[10] ));
 sg13g2_dfrbp_1 _7426_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net90),
    .D(_0074_),
    .Q_N(_0048_),
    .Q(\r2[11] ));
 sg13g2_dfrbp_1 _7427_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net89),
    .D(_0075_),
    .Q_N(_0047_),
    .Q(\r2[12] ));
 sg13g2_dfrbp_1 _7428_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net88),
    .D(_0076_),
    .Q_N(_0046_),
    .Q(\r2[13] ));
 sg13g2_dfrbp_1 _7429_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net87),
    .D(_0077_),
    .Q_N(_0044_),
    .Q(\r2[14] ));
 sg13g2_dfrbp_1 _7430_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net86),
    .D(_0078_),
    .Q_N(_0043_),
    .Q(\r2[15] ));
 sg13g2_dfrbp_1 _7431_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net85),
    .D(_0079_),
    .Q_N(_0026_),
    .Q(\r2[16] ));
 sg13g2_dfrbp_1 _7432_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net84),
    .D(_0080_),
    .Q_N(_0013_),
    .Q(\r2[17] ));
 sg13g2_dfrbp_1 _7433_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net83),
    .D(_0081_),
    .Q_N(_0015_),
    .Q(\r2[18] ));
 sg13g2_dfrbp_1 _7434_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net82),
    .D(_0082_),
    .Q_N(_3687_),
    .Q(\note_freq[0] ));
 sg13g2_dfrbp_1 _7435_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net81),
    .D(_0083_),
    .Q_N(_3686_),
    .Q(\title_r[13] ));
 sg13g2_dfrbp_1 _7436_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net79),
    .D(_0084_),
    .Q_N(_3685_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _7437_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net78),
    .D(_0085_),
    .Q_N(_3684_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _7438_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net77),
    .D(_0086_),
    .Q_N(_3683_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _7439_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net76),
    .D(_0087_),
    .Q_N(_3682_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _7440_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net75),
    .D(_0088_),
    .Q_N(_3681_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _7441_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net31),
    .D(_0089_),
    .Q_N(_3694_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _7442_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net32),
    .D(_0000_),
    .Q_N(_3695_),
    .Q(\note2_freq[0] ));
 sg13g2_dfrbp_1 _7443_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net33),
    .D(_0001_),
    .Q_N(_3696_),
    .Q(\note2_freq[4] ));
 sg13g2_dfrbp_1 _7444_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net34),
    .D(_0002_),
    .Q_N(_3697_),
    .Q(\note2_freq[5] ));
 sg13g2_dfrbp_1 _7445_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net119),
    .D(_0003_),
    .Q_N(_3698_),
    .Q(\note2_freq[6] ));
 sg13g2_dfrbp_1 _7446_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net74),
    .D(_0004_),
    .Q_N(_3680_),
    .Q(\note2_freq[8] ));
 sg13g2_dfrbp_1 _7447_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net73),
    .D(_0090_),
    .Q_N(_3679_),
    .Q(noise));
 sg13g2_dfrbp_1 _7448_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net71),
    .D(_0091_),
    .Q_N(_3678_),
    .Q(\noise_counter[0] ));
 sg13g2_dfrbp_1 _7449_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net69),
    .D(net186),
    .Q_N(_3677_),
    .Q(\noise_counter[1] ));
 sg13g2_dfrbp_1 _7450_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net67),
    .D(_0093_),
    .Q_N(_3676_),
    .Q(\noise_counter[2] ));
 sg13g2_dfrbp_1 _7451_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net65),
    .D(_0094_),
    .Q_N(_3675_),
    .Q(\note2_counter[0] ));
 sg13g2_dfrbp_1 _7452_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net63),
    .D(net183),
    .Q_N(_3674_),
    .Q(\note2_counter[1] ));
 sg13g2_dfrbp_1 _7453_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net61),
    .D(_0096_),
    .Q_N(_0028_),
    .Q(\note2_counter[2] ));
 sg13g2_dfrbp_1 _7454_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net59),
    .D(net180),
    .Q_N(_3673_),
    .Q(\note2_counter[3] ));
 sg13g2_dfrbp_1 _7455_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net57),
    .D(_0098_),
    .Q_N(_3672_),
    .Q(\note2_counter[4] ));
 sg13g2_dfrbp_1 _7456_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net55),
    .D(net177),
    .Q_N(_3671_),
    .Q(\note2_counter[5] ));
 sg13g2_dfrbp_1 _7457_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net53),
    .D(_0100_),
    .Q_N(_3670_),
    .Q(\note2_counter[6] ));
 sg13g2_dfrbp_1 _7458_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net51),
    .D(_0101_),
    .Q_N(_3669_),
    .Q(\note2_counter[7] ));
 sg13g2_dfrbp_1 _7459_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net49),
    .D(_0102_),
    .Q_N(_3668_),
    .Q(\note2_counter[8] ));
 sg13g2_dfrbp_1 _7460_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net47),
    .D(net167),
    .Q_N(_0056_),
    .Q(note2));
 sg13g2_dfrbp_1 _7461_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net45),
    .D(_0104_),
    .Q_N(_3667_),
    .Q(\note_counter[0] ));
 sg13g2_dfrbp_1 _7462_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net43),
    .D(net174),
    .Q_N(_3666_),
    .Q(\note_counter[1] ));
 sg13g2_dfrbp_1 _7463_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net41),
    .D(_0106_),
    .Q_N(_3665_),
    .Q(\note_counter[2] ));
 sg13g2_dfrbp_1 _7464_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net39),
    .D(_0107_),
    .Q_N(_3664_),
    .Q(\note_counter[3] ));
 sg13g2_dfrbp_1 _7465_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net37),
    .D(_0108_),
    .Q_N(_3663_),
    .Q(\note_counter[4] ));
 sg13g2_dfrbp_1 _7466_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net35),
    .D(_0109_),
    .Q_N(_3662_),
    .Q(\note_counter[5] ));
 sg13g2_dfrbp_1 _7467_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net28),
    .D(_0110_),
    .Q_N(_3661_),
    .Q(\note_counter[6] ));
 sg13g2_dfrbp_1 _7468_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net26),
    .D(_0111_),
    .Q_N(_3660_),
    .Q(\note_counter[7] ));
 sg13g2_dfrbp_1 _7469_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net24),
    .D(net169),
    .Q_N(_0055_),
    .Q(note));
 sg13g2_dfrbp_1 _7470_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net22),
    .D(_0113_),
    .Q_N(_0060_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _7471_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net21),
    .D(net222),
    .Q_N(_3659_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _7472_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net20),
    .D(_0115_),
    .Q_N(_0029_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _7473_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net19),
    .D(_0116_),
    .Q_N(_3658_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _7474_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net18),
    .D(_0117_),
    .Q_N(_3657_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _7475_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net17),
    .D(_0118_),
    .Q_N(_3656_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _7476_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net16),
    .D(_0119_),
    .Q_N(_0019_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _7477_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net15),
    .D(_0120_),
    .Q_N(_0022_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _7478_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net14),
    .D(_0121_),
    .Q_N(_0021_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _7479_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net13),
    .D(_0122_),
    .Q_N(_0033_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _7480_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net12),
    .D(_0123_),
    .Q_N(_3655_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _7481_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net11),
    .D(_0124_),
    .Q_N(_3654_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _7482_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net10),
    .D(_0125_),
    .Q_N(_0035_),
    .Q(\center_y[0] ));
 sg13g2_dfrbp_1 _7483_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net8),
    .D(_0126_),
    .Q_N(_0012_),
    .Q(\center_x[0] ));
 sg13g2_dfrbp_1 _7484_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net6),
    .D(net261),
    .Q_N(_0053_),
    .Q(\center_x[1] ));
 sg13g2_dfrbp_1 _7485_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net4),
    .D(_0128_),
    .Q_N(_0032_),
    .Q(\center_x[2] ));
 sg13g2_dfrbp_1 _7486_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net2),
    .D(_0129_),
    .Q_N(_0031_),
    .Q(\center_x[3] ));
 sg13g2_dfrbp_1 _7487_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net137),
    .D(net265),
    .Q_N(_0018_),
    .Q(\center_x[4] ));
 sg13g2_dfrbp_1 _7488_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net129),
    .D(_0131_),
    .Q_N(_0020_),
    .Q(\center_x[5] ));
 sg13g2_dfrbp_1 _7489_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net127),
    .D(net225),
    .Q_N(_0030_),
    .Q(\frame_counter[7] ));
 sg13g2_dfrbp_1 _7490_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net125),
    .D(net257),
    .Q_N(_0017_),
    .Q(\frame_counter[8] ));
 sg13g2_dfrbp_1 _7491_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net123),
    .D(_0134_),
    .Q_N(_0034_),
    .Q(\frame_counter[9] ));
 sg13g2_dfrbp_1 _7492_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net121),
    .D(net163),
    .Q_N(\envelopeA[0] ),
    .Q(frame_counter_frac));
 sg13g2_dfrbp_1 _7493_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net118),
    .D(_0136_),
    .Q_N(_3653_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _7494_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net117),
    .D(_0137_),
    .Q_N(_0027_),
    .Q(\r1[0] ));
 sg13g2_dfrbp_1 _7495_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net116),
    .D(_0138_),
    .Q_N(_3652_),
    .Q(\r1[1] ));
 sg13g2_dfrbp_1 _7496_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net115),
    .D(_0139_),
    .Q_N(_3651_),
    .Q(\r1[2] ));
 sg13g2_dfrbp_1 _7497_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net114),
    .D(_0140_),
    .Q_N(_3650_),
    .Q(\r1[3] ));
 sg13g2_dfrbp_1 _7498_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net113),
    .D(_0141_),
    .Q_N(_3649_),
    .Q(\r1[4] ));
 sg13g2_dfrbp_1 _7499_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net112),
    .D(_0142_),
    .Q_N(_3648_),
    .Q(\r1[5] ));
 sg13g2_dfrbp_1 _7500_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net111),
    .D(_0143_),
    .Q_N(_0041_),
    .Q(\r1[6] ));
 sg13g2_dfrbp_1 _7501_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net110),
    .D(_0144_),
    .Q_N(_0040_),
    .Q(\r1[7] ));
 sg13g2_dfrbp_1 _7502_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net109),
    .D(_0145_),
    .Q_N(_0039_),
    .Q(\r1[8] ));
 sg13g2_dfrbp_1 _7503_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net108),
    .D(_0146_),
    .Q_N(_0038_),
    .Q(\r1[9] ));
 sg13g2_dfrbp_1 _7504_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net107),
    .D(_0147_),
    .Q_N(_0037_),
    .Q(\r1[10] ));
 sg13g2_dfrbp_1 _7505_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net106),
    .D(_0148_),
    .Q_N(_3647_),
    .Q(\r1[11] ));
 sg13g2_dfrbp_1 _7506_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net105),
    .D(net278),
    .Q_N(_0045_),
    .Q(\r1[12] ));
 sg13g2_dfrbp_1 _7507_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net104),
    .D(_0150_),
    .Q_N(_3646_),
    .Q(\r1[13] ));
 sg13g2_dfrbp_1 _7508_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net103),
    .D(net291),
    .Q_N(_0042_),
    .Q(\r1[14] ));
 sg13g2_dfrbp_1 _7509_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net80),
    .D(_0152_),
    .Q_N(_0036_),
    .Q(\r1[15] ));
 sg13g2_dfrbp_1 _7510_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net72),
    .D(_0153_),
    .Q_N(_0014_),
    .Q(\r1[16] ));
 sg13g2_dfrbp_1 _7511_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net70),
    .D(_0154_),
    .Q_N(_0016_),
    .Q(\r1[17] ));
 sg13g2_dfrbp_1 _7512_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net68),
    .D(net171),
    .Q_N(_0059_),
    .Q(\title_r[0] ));
 sg13g2_dfrbp_1 _7513_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net64),
    .D(_0156_),
    .Q_N(_3645_),
    .Q(\title_r[1] ));
 sg13g2_dfrbp_1 _7514_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net60),
    .D(_0157_),
    .Q_N(_3644_),
    .Q(\title_r[2] ));
 sg13g2_dfrbp_1 _7515_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net56),
    .D(_0158_),
    .Q_N(_3643_),
    .Q(\title_r[3] ));
 sg13g2_dfrbp_1 _7516_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net52),
    .D(_0159_),
    .Q_N(_3642_),
    .Q(\title_r[4] ));
 sg13g2_dfrbp_1 _7517_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net48),
    .D(_0160_),
    .Q_N(_3641_),
    .Q(\title_r[5] ));
 sg13g2_dfrbp_1 _7518_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net44),
    .D(_0161_),
    .Q_N(_3640_),
    .Q(\title_r[6] ));
 sg13g2_dfrbp_1 _7519_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net40),
    .D(_0162_),
    .Q_N(_3639_),
    .Q(\title_r[7] ));
 sg13g2_dfrbp_1 _7520_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net36),
    .D(_0163_),
    .Q_N(_3638_),
    .Q(\title_r[8] ));
 sg13g2_dfrbp_1 _7521_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net27),
    .D(_0164_),
    .Q_N(_3637_),
    .Q(\title_r[9] ));
 sg13g2_dfrbp_1 _7522_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net23),
    .D(_0165_),
    .Q_N(_3636_),
    .Q(\title_r[10] ));
 sg13g2_dfrbp_1 _7523_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net7),
    .D(_0166_),
    .Q_N(_3635_),
    .Q(\title_r[11] ));
 sg13g2_dfrbp_1 _7524_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net3),
    .D(_0167_),
    .Q_N(_3634_),
    .Q(\title_r[12] ));
 sg13g2_dfrbp_1 _7525_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net136),
    .D(net161),
    .Q_N(_0058_),
    .Q(\title_r_pixels_in_scanline[0] ));
 sg13g2_dfrbp_1 _7526_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net126),
    .D(net204),
    .Q_N(_3633_),
    .Q(\title_r_pixels_in_scanline[1] ));
 sg13g2_dfrbp_1 _7527_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net122),
    .D(_0170_),
    .Q_N(_3632_),
    .Q(\title_r_pixels_in_scanline[2] ));
 sg13g2_dfrbp_1 _7528_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net66),
    .D(_0171_),
    .Q_N(_3631_),
    .Q(\title_r_pixels_in_scanline[3] ));
 sg13g2_dfrbp_1 _7529_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net58),
    .D(_0172_),
    .Q_N(_3630_),
    .Q(\title_r_pixels_in_scanline[4] ));
 sg13g2_dfrbp_1 _7530_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net130),
    .D(_0173_),
    .Q_N(_3699_),
    .Q(\title_r_pixels_in_scanline[5] ));
 sg13g2_dfrbp_1 _7531_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net50),
    .D(_0010_),
    .Q_N(_3629_),
    .Q(hsync));
 sg13g2_dfrbp_1 _7532_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net42),
    .D(_0174_),
    .Q_N(_0057_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _7533_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net29),
    .D(_0175_),
    .Q_N(_3628_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _7534_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net9),
    .D(_0176_),
    .Q_N(_3627_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _7535_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net1),
    .D(_0177_),
    .Q_N(_3626_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _7536_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net124),
    .D(_0178_),
    .Q_N(_3625_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _7537_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net62),
    .D(_0179_),
    .Q_N(_3624_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _7538_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net46),
    .D(_0180_),
    .Q_N(_0024_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _7539_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net25),
    .D(_0181_),
    .Q_N(_3623_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _7540_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net128),
    .D(_0182_),
    .Q_N(_3622_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _7541_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net131),
    .D(_0183_),
    .Q_N(_3700_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _7542_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net132),
    .D(net235),
    .Q_N(_3701_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _7543_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net133),
    .D(_0005_),
    .Q_N(_3702_),
    .Q(\note_freq[2] ));
 sg13g2_dfrbp_1 _7544_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net134),
    .D(_0006_),
    .Q_N(_3703_),
    .Q(\note_freq[4] ));
 sg13g2_dfrbp_1 _7545_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net135),
    .D(_0007_),
    .Q_N(_3704_),
    .Q(\note_freq[5] ));
 sg13g2_dfrbp_1 _7546_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net38),
    .D(_0008_),
    .Q_N(_3705_),
    .Q(\note_freq[6] ));
 sg13g2_dfrbp_1 _7547_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net54),
    .D(_0009_),
    .Q_N(_3621_),
    .Q(\note_freq[7] ));
 sg13g2_dfrbp_1 _7548_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net5),
    .D(_0184_),
    .Q_N(_3620_),
    .Q(\note2_freq[7] ));
 sg13g2_dfrbp_1 _7549_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net120),
    .D(_0185_),
    .Q_N(_3619_),
    .Q(\note2_freq[3] ));
 sg13g2_tiehi _7486__2 (.L_HI(net2));
 sg13g2_tiehi _7524__3 (.L_HI(net3));
 sg13g2_tiehi _7485__4 (.L_HI(net4));
 sg13g2_tiehi _7548__5 (.L_HI(net5));
 sg13g2_tiehi _7484__6 (.L_HI(net6));
 sg13g2_tiehi _7523__7 (.L_HI(net7));
 sg13g2_tiehi _7483__8 (.L_HI(net8));
 sg13g2_tiehi _7534__9 (.L_HI(net9));
 sg13g2_tiehi _7482__10 (.L_HI(net10));
 sg13g2_tiehi _7481__11 (.L_HI(net11));
 sg13g2_tiehi _7480__12 (.L_HI(net12));
 sg13g2_tiehi _7479__13 (.L_HI(net13));
 sg13g2_tiehi _7478__14 (.L_HI(net14));
 sg13g2_tiehi _7477__15 (.L_HI(net15));
 sg13g2_tiehi _7476__16 (.L_HI(net16));
 sg13g2_tiehi _7475__17 (.L_HI(net17));
 sg13g2_tiehi _7474__18 (.L_HI(net18));
 sg13g2_tiehi _7473__19 (.L_HI(net19));
 sg13g2_tiehi _7472__20 (.L_HI(net20));
 sg13g2_tiehi _7471__21 (.L_HI(net21));
 sg13g2_tiehi _7470__22 (.L_HI(net22));
 sg13g2_tiehi _7522__23 (.L_HI(net23));
 sg13g2_tiehi _7469__24 (.L_HI(net24));
 sg13g2_tiehi _7539__25 (.L_HI(net25));
 sg13g2_tiehi _7468__26 (.L_HI(net26));
 sg13g2_tiehi _7521__27 (.L_HI(net27));
 sg13g2_tiehi _7467__28 (.L_HI(net28));
 sg13g2_tiehi _7533__29 (.L_HI(net29));
 sg13g2_tiehi _7413__30 (.L_HI(net30));
 sg13g2_tiehi _7441__31 (.L_HI(net31));
 sg13g2_tiehi _7442__32 (.L_HI(net32));
 sg13g2_tiehi _7443__33 (.L_HI(net33));
 sg13g2_tiehi _7444__34 (.L_HI(net34));
 sg13g2_tiehi _7466__35 (.L_HI(net35));
 sg13g2_tiehi _7520__36 (.L_HI(net36));
 sg13g2_tiehi _7465__37 (.L_HI(net37));
 sg13g2_tiehi _7546__38 (.L_HI(net38));
 sg13g2_tiehi _7464__39 (.L_HI(net39));
 sg13g2_tiehi _7519__40 (.L_HI(net40));
 sg13g2_tiehi _7463__41 (.L_HI(net41));
 sg13g2_tiehi _7532__42 (.L_HI(net42));
 sg13g2_tiehi _7462__43 (.L_HI(net43));
 sg13g2_tiehi _7518__44 (.L_HI(net44));
 sg13g2_tiehi _7461__45 (.L_HI(net45));
 sg13g2_tiehi _7538__46 (.L_HI(net46));
 sg13g2_tiehi _7460__47 (.L_HI(net47));
 sg13g2_tiehi _7517__48 (.L_HI(net48));
 sg13g2_tiehi _7459__49 (.L_HI(net49));
 sg13g2_tiehi _7531__50 (.L_HI(net50));
 sg13g2_tiehi _7458__51 (.L_HI(net51));
 sg13g2_tiehi _7516__52 (.L_HI(net52));
 sg13g2_tiehi _7457__53 (.L_HI(net53));
 sg13g2_tiehi _7547__54 (.L_HI(net54));
 sg13g2_tiehi _7456__55 (.L_HI(net55));
 sg13g2_tiehi _7515__56 (.L_HI(net56));
 sg13g2_tiehi _7455__57 (.L_HI(net57));
 sg13g2_tiehi _7529__58 (.L_HI(net58));
 sg13g2_tiehi _7454__59 (.L_HI(net59));
 sg13g2_tiehi _7514__60 (.L_HI(net60));
 sg13g2_tiehi _7453__61 (.L_HI(net61));
 sg13g2_tiehi _7537__62 (.L_HI(net62));
 sg13g2_tiehi _7452__63 (.L_HI(net63));
 sg13g2_tiehi _7513__64 (.L_HI(net64));
 sg13g2_tiehi _7451__65 (.L_HI(net65));
 sg13g2_tiehi _7528__66 (.L_HI(net66));
 sg13g2_tiehi _7450__67 (.L_HI(net67));
 sg13g2_tiehi _7512__68 (.L_HI(net68));
 sg13g2_tiehi _7449__69 (.L_HI(net69));
 sg13g2_tiehi _7511__70 (.L_HI(net70));
 sg13g2_tiehi _7448__71 (.L_HI(net71));
 sg13g2_tiehi _7510__72 (.L_HI(net72));
 sg13g2_tiehi _7447__73 (.L_HI(net73));
 sg13g2_tiehi _7446__74 (.L_HI(net74));
 sg13g2_tiehi _7440__75 (.L_HI(net75));
 sg13g2_tiehi _7439__76 (.L_HI(net76));
 sg13g2_tiehi _7438__77 (.L_HI(net77));
 sg13g2_tiehi _7437__78 (.L_HI(net78));
 sg13g2_tiehi _7436__79 (.L_HI(net79));
 sg13g2_tiehi _7509__80 (.L_HI(net80));
 sg13g2_tiehi _7435__81 (.L_HI(net81));
 sg13g2_tiehi _7434__82 (.L_HI(net82));
 sg13g2_tiehi _7433__83 (.L_HI(net83));
 sg13g2_tiehi _7432__84 (.L_HI(net84));
 sg13g2_tiehi _7431__85 (.L_HI(net85));
 sg13g2_tiehi _7430__86 (.L_HI(net86));
 sg13g2_tiehi _7429__87 (.L_HI(net87));
 sg13g2_tiehi _7428__88 (.L_HI(net88));
 sg13g2_tiehi _7427__89 (.L_HI(net89));
 sg13g2_tiehi _7426__90 (.L_HI(net90));
 sg13g2_tiehi _7425__91 (.L_HI(net91));
 sg13g2_tiehi _7424__92 (.L_HI(net92));
 sg13g2_tiehi _7423__93 (.L_HI(net93));
 sg13g2_tiehi _7422__94 (.L_HI(net94));
 sg13g2_tiehi _7421__95 (.L_HI(net95));
 sg13g2_tiehi _7420__96 (.L_HI(net96));
 sg13g2_tiehi _7419__97 (.L_HI(net97));
 sg13g2_tiehi _7418__98 (.L_HI(net98));
 sg13g2_tiehi _7417__99 (.L_HI(net99));
 sg13g2_tiehi _7416__100 (.L_HI(net100));
 sg13g2_tiehi _7415__101 (.L_HI(net101));
 sg13g2_tiehi _7414__102 (.L_HI(net102));
 sg13g2_tiehi _7508__103 (.L_HI(net103));
 sg13g2_tiehi _7507__104 (.L_HI(net104));
 sg13g2_tiehi _7506__105 (.L_HI(net105));
 sg13g2_tiehi _7505__106 (.L_HI(net106));
 sg13g2_tiehi _7504__107 (.L_HI(net107));
 sg13g2_tiehi _7503__108 (.L_HI(net108));
 sg13g2_tiehi _7502__109 (.L_HI(net109));
 sg13g2_tiehi _7501__110 (.L_HI(net110));
 sg13g2_tiehi _7500__111 (.L_HI(net111));
 sg13g2_tiehi _7499__112 (.L_HI(net112));
 sg13g2_tiehi _7498__113 (.L_HI(net113));
 sg13g2_tiehi _7497__114 (.L_HI(net114));
 sg13g2_tiehi _7496__115 (.L_HI(net115));
 sg13g2_tiehi _7495__116 (.L_HI(net116));
 sg13g2_tiehi _7494__117 (.L_HI(net117));
 sg13g2_tiehi _7493__118 (.L_HI(net118));
 sg13g2_tiehi _7445__119 (.L_HI(net119));
 sg13g2_tiehi _7549__120 (.L_HI(net120));
 sg13g2_tiehi _7492__121 (.L_HI(net121));
 sg13g2_tiehi _7527__122 (.L_HI(net122));
 sg13g2_tiehi _7491__123 (.L_HI(net123));
 sg13g2_tiehi _7536__124 (.L_HI(net124));
 sg13g2_tiehi _7490__125 (.L_HI(net125));
 sg13g2_tiehi _7526__126 (.L_HI(net126));
 sg13g2_tiehi _7489__127 (.L_HI(net127));
 sg13g2_tiehi _7540__128 (.L_HI(net128));
 sg13g2_tiehi _7488__129 (.L_HI(net129));
 sg13g2_tiehi _7530__130 (.L_HI(net130));
 sg13g2_tiehi _7541__131 (.L_HI(net131));
 sg13g2_tiehi _7542__132 (.L_HI(net132));
 sg13g2_tiehi _7543__133 (.L_HI(net133));
 sg13g2_tiehi _7544__134 (.L_HI(net134));
 sg13g2_tiehi _7545__135 (.L_HI(net135));
 sg13g2_tiehi _7525__136 (.L_HI(net136));
 sg13g2_tiehi _7487__137 (.L_HI(net137));
 sg13g2_tiehi tt_um_rejunity_vga_test01_138 (.L_HI(net138));
 sg13g2_tiehi tt_um_rejunity_vga_test01_139 (.L_HI(net139));
 sg13g2_tiehi tt_um_rejunity_vga_test01_140 (.L_HI(net140));
 sg13g2_tiehi tt_um_rejunity_vga_test01_141 (.L_HI(net141));
 sg13g2_tiehi tt_um_rejunity_vga_test01_142 (.L_HI(net142));
 sg13g2_tiehi tt_um_rejunity_vga_test01_143 (.L_HI(net143));
 sg13g2_tiehi tt_um_rejunity_vga_test01_144 (.L_HI(net144));
 sg13g2_tiehi tt_um_rejunity_vga_test01_145 (.L_HI(net145));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _7695_ (.A(uio_out[7]),
    .X(uio_out[0]));
 sg13g2_buf_1 _7696_ (.A(uio_out[7]),
    .X(uio_out[1]));
 sg13g2_buf_1 _7697_ (.A(uio_out[7]),
    .X(uio_out[2]));
 sg13g2_buf_1 _7698_ (.A(uio_out[7]),
    .X(uio_out[3]));
 sg13g2_buf_1 _7699_ (.A(uio_out[7]),
    .X(uio_out[4]));
 sg13g2_buf_1 _7700_ (.A(uio_out[7]),
    .X(uio_out[5]));
 sg13g2_buf_1 _7701_ (.A(uio_out[7]),
    .X(uio_out[6]));
 sg13g2_buf_8 fanout704 (.A(_1662_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_1515_),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(_1256_));
 sg13g2_buf_2 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(_1212_));
 sg13g2_buf_2 fanout709 (.A(_1157_),
    .X(net709));
 sg13g2_buf_1 fanout710 (.A(_1157_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(net712),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_2805_),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(_0477_));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(_0427_));
 sg13g2_buf_4 fanout715 (.X(net715),
    .A(_0362_));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(_0276_));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(net718));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(_3302_));
 sg13g2_buf_2 fanout719 (.A(_0312_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_0312_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(net723),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net723),
    .X(net722));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(_2639_));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(_2638_));
 sg13g2_buf_2 fanout725 (.A(_0336_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_0327_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_0373_),
    .X(net727));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(_3131_));
 sg13g2_buf_2 fanout729 (.A(_0564_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(net731),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(net733),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_3130_),
    .X(net733));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(_2905_));
 sg13g2_buf_1 fanout735 (.A(_2905_),
    .X(net735));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(_3152_));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(_3147_));
 sg13g2_buf_1 fanout738 (.A(_3147_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(net740),
    .X(net739));
 sg13g2_buf_1 fanout740 (.A(net741),
    .X(net740));
 sg13g2_buf_1 fanout741 (.A(_2603_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_2603_),
    .X(net743));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(_2602_));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(_2518_));
 sg13g2_buf_2 fanout746 (.A(_0379_),
    .X(net746));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(_0379_));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(_3146_));
 sg13g2_buf_4 fanout749 (.X(net749),
    .A(_3145_));
 sg13g2_buf_2 fanout750 (.A(_3145_),
    .X(net750));
 sg13g2_buf_4 fanout751 (.X(net751),
    .A(net752));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(_3134_));
 sg13g2_buf_2 fanout753 (.A(_3067_),
    .X(net753));
 sg13g2_buf_4 fanout754 (.X(net754),
    .A(_2240_));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(_0374_));
 sg13g2_buf_2 fanout756 (.A(_0374_),
    .X(net756));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(_0324_));
 sg13g2_buf_2 fanout758 (.A(_0324_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_3576_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_3575_),
    .X(net760));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(_3560_));
 sg13g2_buf_2 fanout762 (.A(_3560_),
    .X(net762));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(_3178_));
 sg13g2_buf_4 fanout764 (.X(net764),
    .A(net765));
 sg13g2_buf_2 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_4 fanout766 (.X(net766),
    .A(_3135_));
 sg13g2_buf_4 fanout767 (.X(net767),
    .A(_3061_));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(_3060_));
 sg13g2_buf_2 fanout769 (.A(_3060_),
    .X(net769));
 sg13g2_buf_4 fanout770 (.X(net770),
    .A(_1830_));
 sg13g2_buf_2 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_4 fanout772 (.X(net772),
    .A(_0330_));
 sg13g2_buf_2 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(net775));
 sg13g2_buf_2 fanout775 (.A(_3106_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_4 fanout777 (.X(net777),
    .A(net780));
 sg13g2_buf_4 fanout778 (.X(net778),
    .A(net779));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(net780));
 sg13g2_buf_2 fanout780 (.A(_3105_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_0815_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_0679_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_0644_),
    .X(net783));
 sg13g2_buf_4 fanout784 (.X(net784),
    .A(_0334_));
 sg13g2_buf_4 fanout785 (.X(net785),
    .A(_0333_));
 sg13g2_buf_2 fanout786 (.A(_0333_),
    .X(net786));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(_0291_));
 sg13g2_buf_2 fanout788 (.A(_0291_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(net790),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_3579_),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_3523_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_3523_),
    .X(net792));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(net795));
 sg13g2_buf_2 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_3124_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(_3095_),
    .X(net797));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(net799));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(_3052_));
 sg13g2_buf_2 fanout800 (.A(net801),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_0377_),
    .X(net801));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_0279_));
 sg13g2_buf_1 fanout803 (.A(_0279_),
    .X(net803));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(_0278_));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(_3583_));
 sg13g2_buf_2 fanout806 (.A(_3583_),
    .X(net806));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(_3582_));
 sg13g2_buf_2 fanout808 (.A(net809),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(net810),
    .X(net809));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(_3581_));
 sg13g2_buf_4 fanout811 (.X(net811),
    .A(_3053_));
 sg13g2_buf_2 fanout812 (.A(net813),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_2969_),
    .X(net813));
 sg13g2_buf_4 fanout814 (.X(net814),
    .A(_2969_));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(_2611_));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(_2445_));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(_2427_));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(_2416_));
 sg13g2_buf_2 fanout819 (.A(net821),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(net822),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(net825),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net825),
    .X(net823));
 sg13g2_buf_1 fanout824 (.A(net825),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(\hvsync_gen.vsync ),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(net233),
    .X(net826));
 sg13g2_buf_1 fanout827 (.A(net233),
    .X(net827));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(\hvsync_gen.vpos[6] ));
 sg13g2_buf_1 fanout829 (.A(\hvsync_gen.vpos[6] ),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(\hvsync_gen.vpos[6] ),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(\hvsync_gen.vpos[5] ),
    .X(net832));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(net834));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(\hvsync_gen.vpos[4] ));
 sg13g2_buf_2 fanout835 (.A(net836),
    .X(net835));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(\hvsync_gen.vpos[3] ));
 sg13g2_buf_2 fanout837 (.A(\hvsync_gen.vpos[2] ),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(net839),
    .X(net838));
 sg13g2_buf_4 fanout839 (.X(net839),
    .A(\hvsync_gen.vpos[1] ));
 sg13g2_buf_2 fanout840 (.A(\hvsync_gen.vpos[0] ),
    .X(net840));
 sg13g2_buf_1 fanout841 (.A(\hvsync_gen.vpos[0] ),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(\r1[13] ),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(\r1[11] ),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(\r1[11] ),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(\r1[5] ),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(\r1[4] ),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(\r1[3] ),
    .X(net847));
 sg13g2_buf_4 fanout848 (.X(net848),
    .A(\r1[2] ));
 sg13g2_buf_4 fanout849 (.X(net849),
    .A(net286));
 sg13g2_buf_2 fanout850 (.A(_0034_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(net256),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(\frame_counter[7] ),
    .X(net852));
 sg13g2_buf_4 fanout853 (.X(net853),
    .A(_0020_));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(\center_x[5] ));
 sg13g2_buf_2 fanout855 (.A(net857),
    .X(net855));
 sg13g2_buf_1 fanout856 (.A(net857),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(net858),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(\center_x[5] ),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_0018_),
    .X(net861));
 sg13g2_buf_4 fanout862 (.X(net862),
    .A(\center_x[4] ));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(\center_x[4] ));
 sg13g2_buf_2 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(net866),
    .X(net865));
 sg13g2_buf_4 fanout866 (.X(net866),
    .A(\center_x[4] ));
 sg13g2_buf_4 fanout867 (.X(net867),
    .A(net868));
 sg13g2_buf_2 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_4 fanout869 (.X(net869),
    .A(\center_x[3] ));
 sg13g2_buf_2 fanout870 (.A(net871),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(net872),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_4 fanout873 (.X(net873),
    .A(\center_x[3] ));
 sg13g2_buf_4 fanout874 (.X(net874),
    .A(net875));
 sg13g2_buf_2 fanout875 (.A(\center_x[2] ),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net877),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(\center_x[2] ),
    .X(net877));
 sg13g2_buf_4 fanout878 (.X(net878),
    .A(net879));
 sg13g2_buf_4 fanout879 (.X(net879),
    .A(\center_x[1] ));
 sg13g2_buf_2 fanout880 (.A(net883),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net882),
    .X(net881));
 sg13g2_buf_1 fanout882 (.A(net883),
    .X(net882));
 sg13g2_buf_4 fanout883 (.X(net883),
    .A(\center_x[1] ));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(net885));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(\center_x[0] ));
 sg13g2_buf_2 fanout886 (.A(net887),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net889),
    .X(net888));
 sg13g2_buf_4 fanout889 (.X(net889),
    .A(\center_x[0] ));
 sg13g2_buf_4 fanout890 (.X(net890),
    .A(net891));
 sg13g2_buf_4 fanout891 (.X(net891),
    .A(net892));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(_0035_));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(net895));
 sg13g2_buf_2 fanout894 (.A(net895),
    .X(net894));
 sg13g2_buf_4 fanout895 (.X(net895),
    .A(\center_y[0] ));
 sg13g2_buf_2 fanout896 (.A(\hvsync_gen.hpos[8] ),
    .X(net896));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(net898));
 sg13g2_buf_2 fanout898 (.A(\hvsync_gen.hpos[7] ),
    .X(net898));
 sg13g2_buf_4 fanout899 (.X(net899),
    .A(net902));
 sg13g2_buf_2 fanout900 (.A(net902),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(net902),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(\hvsync_gen.hpos[6] ),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(net905),
    .X(net903));
 sg13g2_buf_1 fanout904 (.A(net905),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(net906),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(net246),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net908),
    .X(net907));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(net909));
 sg13g2_buf_2 fanout909 (.A(net223),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(net911),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(net913),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(\hvsync_gen.hpos[3] ),
    .X(net913));
 sg13g2_buf_4 fanout914 (.X(net914),
    .A(net230));
 sg13g2_buf_2 fanout915 (.A(net221),
    .X(net915));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(\hvsync_gen.hpos[0] ));
 sg13g2_buf_2 fanout917 (.A(\r2[9] ),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(net922),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(net922),
    .X(net919));
 sg13g2_buf_4 fanout920 (.X(net920),
    .A(net922));
 sg13g2_buf_2 fanout921 (.A(net922),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_2685_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_2685_),
    .X(net923));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(_2685_));
 sg13g2_buf_4 fanout925 (.X(net925),
    .A(net928));
 sg13g2_buf_4 fanout926 (.X(net926),
    .A(net928));
 sg13g2_buf_1 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_4 fanout928 (.X(net928),
    .A(rst_n));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(rst_n));
 sg13g2_buf_2 fanout930 (.A(rst_n),
    .X(net930));
 sg13g2_tiehi _7535__1 (.L_HI(net1));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_29__leaf_clk));
 sg13g2_dlygate4sd1_1 rebuffer1 (.A(_3591_),
    .X(net146));
 sg13g2_buf_1 rebuffer2 (.A(net146),
    .X(net147));
 sg13g2_dlygate4sd1_1 rebuffer3 (.A(_3591_),
    .X(net148));
 sg13g2_dlygate4sd1_1 rebuffer4 (.A(net148),
    .X(net149));
 sg13g2_dlygate4sd1_1 rebuffer5 (.A(net149),
    .X(net150));
 sg13g2_buf_2 rebuffer6 (.A(_0965_),
    .X(net151));
 sg13g2_buf_2 rebuffer7 (.A(_3608_),
    .X(net152));
 sg13g2_buf_1 rebuffer8 (.A(net152),
    .X(net153));
 sg13g2_dlygate4sd1_1 rebuffer9 (.A(_3589_),
    .X(net154));
 sg13g2_dlygate4sd1_1 rebuffer10 (.A(net154),
    .X(net155));
 sg13g2_dlygate4sd1_1 rebuffer11 (.A(_1211_),
    .X(net156));
 sg13g2_dlygate4sd1_1 rebuffer12 (.A(_0264_),
    .X(net157));
 sg13g2_dlygate4sd1_1 rebuffer13 (.A(_1375_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0060_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0058_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0168_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold17 (.A(\envelopeA[0] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0135_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold19 (.A(hsync),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold20 (.A(\noise_counter[2] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0056_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0103_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0055_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0112_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0059_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0155_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold27 (.A(\note_counter[1] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold28 (.A(_2499_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0105_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold30 (.A(\note2_counter[5] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold31 (.A(_2472_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0099_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold33 (.A(\note2_counter[3] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold34 (.A(_2469_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0097_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold36 (.A(\note2_counter[1] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold37 (.A(_2462_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0095_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold39 (.A(\noise_counter[0] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold40 (.A(_2439_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0092_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold42 (.A(\note2_counter[0] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold43 (.A(\note_counter[3] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold44 (.A(_2504_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold45 (.A(\note2_counter[6] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold46 (.A(_2475_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold47 (.A(\note2_counter[2] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold48 (.A(_2467_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold49 (.A(\note_counter[4] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold50 (.A(\note_counter[2] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold51 (.A(_2502_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold52 (.A(\note_counter[5] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold53 (.A(\note_counter[0] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold54 (.A(\noise_counter[1] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold55 (.A(\note_counter[6] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold56 (.A(\note2_counter[7] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold57 (.A(\title_r_pixels_in_scanline[1] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold58 (.A(_3006_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0169_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold60 (.A(\hvsync_gen.vsync ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0021_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold62 (.A(_2535_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold63 (.A(\note2_counter[4] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0057_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold65 (.A(_3022_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold66 (.A(noise),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0019_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0033_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold69 (.A(_3050_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold70 (.A(\title_r[1] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold71 (.A(\note2_counter[8] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold72 (.A(\title_r_pixels_in_scanline[2] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold73 (.A(_3009_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold74 (.A(\note_counter[7] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold75 (.A(\title_r[2] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold76 (.A(\hvsync_gen.hpos[1] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0114_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold78 (.A(\hvsync_gen.hpos[4] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold79 (.A(\frame_counter[7] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0132_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold81 (.A(\r2[12] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold82 (.A(\title_r_pixels_in_scanline[5] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold83 (.A(_3014_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold84 (.A(\frame_counter[9] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold85 (.A(\hvsync_gen.hpos[2] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold86 (.A(_2521_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold87 (.A(\title_r_pixels_in_scanline[3] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold88 (.A(\hvsync_gen.vpos[7] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold89 (.A(_3045_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0011_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold91 (.A(\title_r[12] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0024_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold93 (.A(\r2[15] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold94 (.A(\title_r_pixels_in_scanline[4] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold95 (.A(\title_r[3] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold96 (.A(\hvsync_gen.vpos[9] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold97 (.A(\title_r[9] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold98 (.A(\title_r[13] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold99 (.A(\title_r[7] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold100 (.A(\title_r[10] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold101 (.A(\hvsync_gen.hpos[5] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold102 (.A(\title_r[8] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold103 (.A(\r1[17] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold104 (.A(\r2[13] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0014_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0015_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold107 (.A(_3411_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold108 (.A(\title_r[6] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold109 (.A(\title_r[11] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0027_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold111 (.A(\frame_counter[8] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0133_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold113 (.A(\title_r[4] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold114 (.A(\hvsync_gen.vpos[8] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0012_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0127_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0031_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold119 (.A(net862),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0130_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0029_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold122 (.A(\r2[2] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0048_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold124 (.A(_3326_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold125 (.A(\r2[16] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold126 (.A(\r2[6] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0069_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold128 (.A(\r1[8] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold129 (.A(\r2[14] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold130 (.A(_3362_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold131 (.A(\r1[10] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold132 (.A(\r1[12] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0149_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold134 (.A(\r2[4] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold135 (.A(\r2[8] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold136 (.A(_3285_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0042_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold138 (.A(_2878_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold139 (.A(\r2[10] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold140 (.A(\r1[7] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold141 (.A(frame_counter_frac),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold142 (.A(\r2[0] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold144 (.A(net854),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold145 (.A(\r1[14] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0151_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold147 (.A(\title_r[5] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold148 (.A(\r1[9] ),
    .X(net293));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_fill_2 FILLER_0_101 ();
 sg13g2_decap_8 FILLER_0_115 ();
 sg13g2_decap_8 FILLER_0_122 ();
 sg13g2_fill_1 FILLER_0_129 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_fill_1 FILLER_0_141 ();
 sg13g2_decap_8 FILLER_0_146 ();
 sg13g2_decap_8 FILLER_0_153 ();
 sg13g2_decap_4 FILLER_0_160 ();
 sg13g2_fill_2 FILLER_0_173 ();
 sg13g2_fill_2 FILLER_0_180 ();
 sg13g2_fill_1 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_fill_2 FILLER_0_219 ();
 sg13g2_decap_4 FILLER_0_226 ();
 sg13g2_fill_2 FILLER_0_230 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_fill_2 FILLER_0_253 ();
 sg13g2_fill_1 FILLER_0_255 ();
 sg13g2_decap_4 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_4 FILLER_0_283 ();
 sg13g2_fill_1 FILLER_0_295 ();
 sg13g2_fill_2 FILLER_0_300 ();
 sg13g2_fill_1 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_decap_4 FILLER_0_314 ();
 sg13g2_fill_2 FILLER_0_318 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_4 FILLER_1_63 ();
 sg13g2_fill_2 FILLER_1_67 ();
 sg13g2_fill_1 FILLER_1_145 ();
 sg13g2_fill_1 FILLER_1_192 ();
 sg13g2_decap_4 FILLER_1_198 ();
 sg13g2_fill_1 FILLER_1_202 ();
 sg13g2_fill_1 FILLER_1_208 ();
 sg13g2_fill_2 FILLER_1_247 ();
 sg13g2_fill_1 FILLER_1_249 ();
 sg13g2_fill_2 FILLER_1_258 ();
 sg13g2_fill_1 FILLER_1_265 ();
 sg13g2_fill_1 FILLER_1_289 ();
 sg13g2_fill_2 FILLER_1_300 ();
 sg13g2_fill_1 FILLER_1_302 ();
 sg13g2_fill_1 FILLER_1_320 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_4 FILLER_2_63 ();
 sg13g2_fill_1 FILLER_2_67 ();
 sg13g2_fill_1 FILLER_2_94 ();
 sg13g2_fill_2 FILLER_2_100 ();
 sg13g2_fill_2 FILLER_2_201 ();
 sg13g2_fill_2 FILLER_2_224 ();
 sg13g2_fill_2 FILLER_2_281 ();
 sg13g2_fill_1 FILLER_2_300 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_56 ();
 sg13g2_fill_1 FILLER_3_58 ();
 sg13g2_fill_1 FILLER_3_85 ();
 sg13g2_fill_2 FILLER_3_94 ();
 sg13g2_fill_2 FILLER_3_109 ();
 sg13g2_fill_1 FILLER_3_242 ();
 sg13g2_fill_1 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_fill_2 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_4 FILLER_4_49 ();
 sg13g2_fill_1 FILLER_4_53 ();
 sg13g2_fill_2 FILLER_4_122 ();
 sg13g2_fill_2 FILLER_4_160 ();
 sg13g2_fill_1 FILLER_4_162 ();
 sg13g2_fill_1 FILLER_4_215 ();
 sg13g2_fill_2 FILLER_4_253 ();
 sg13g2_fill_1 FILLER_4_255 ();
 sg13g2_fill_1 FILLER_4_281 ();
 sg13g2_fill_2 FILLER_4_293 ();
 sg13g2_fill_1 FILLER_4_295 ();
 sg13g2_fill_1 FILLER_4_336 ();
 sg13g2_fill_2 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_4 FILLER_5_56 ();
 sg13g2_decap_4 FILLER_5_73 ();
 sg13g2_fill_2 FILLER_5_91 ();
 sg13g2_fill_2 FILLER_5_98 ();
 sg13g2_fill_2 FILLER_5_127 ();
 sg13g2_fill_2 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_151 ();
 sg13g2_decap_4 FILLER_5_158 ();
 sg13g2_fill_1 FILLER_5_167 ();
 sg13g2_fill_1 FILLER_5_173 ();
 sg13g2_fill_2 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_241 ();
 sg13g2_fill_1 FILLER_5_243 ();
 sg13g2_fill_2 FILLER_5_288 ();
 sg13g2_fill_2 FILLER_5_303 ();
 sg13g2_fill_2 FILLER_5_317 ();
 sg13g2_fill_1 FILLER_5_319 ();
 sg13g2_fill_1 FILLER_5_328 ();
 sg13g2_fill_2 FILLER_5_351 ();
 sg13g2_fill_1 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_4 FILLER_6_42 ();
 sg13g2_fill_2 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_fill_1 FILLER_6_82 ();
 sg13g2_fill_2 FILLER_6_114 ();
 sg13g2_fill_1 FILLER_6_116 ();
 sg13g2_fill_1 FILLER_6_122 ();
 sg13g2_fill_2 FILLER_6_143 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_fill_2 FILLER_6_162 ();
 sg13g2_fill_1 FILLER_6_164 ();
 sg13g2_decap_8 FILLER_6_197 ();
 sg13g2_decap_4 FILLER_6_204 ();
 sg13g2_fill_2 FILLER_6_208 ();
 sg13g2_fill_2 FILLER_6_218 ();
 sg13g2_decap_4 FILLER_6_228 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_fill_2 FILLER_6_259 ();
 sg13g2_fill_2 FILLER_6_265 ();
 sg13g2_decap_8 FILLER_6_271 ();
 sg13g2_fill_2 FILLER_6_278 ();
 sg13g2_fill_1 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_fill_2 FILLER_6_330 ();
 sg13g2_decap_4 FILLER_6_349 ();
 sg13g2_fill_1 FILLER_6_353 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_2 FILLER_7_82 ();
 sg13g2_fill_1 FILLER_7_89 ();
 sg13g2_fill_1 FILLER_7_117 ();
 sg13g2_fill_1 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_185 ();
 sg13g2_fill_2 FILLER_7_234 ();
 sg13g2_fill_1 FILLER_7_236 ();
 sg13g2_decap_8 FILLER_7_251 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_decap_8 FILLER_7_293 ();
 sg13g2_fill_1 FILLER_7_304 ();
 sg13g2_fill_1 FILLER_7_328 ();
 sg13g2_fill_2 FILLER_7_341 ();
 sg13g2_fill_1 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_fill_1 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_77 ();
 sg13g2_fill_1 FILLER_8_79 ();
 sg13g2_fill_1 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_110 ();
 sg13g2_fill_2 FILLER_8_121 ();
 sg13g2_fill_1 FILLER_8_123 ();
 sg13g2_fill_1 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_156 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_fill_2 FILLER_8_237 ();
 sg13g2_fill_1 FILLER_8_239 ();
 sg13g2_fill_2 FILLER_8_245 ();
 sg13g2_fill_1 FILLER_8_247 ();
 sg13g2_fill_1 FILLER_8_253 ();
 sg13g2_fill_2 FILLER_8_276 ();
 sg13g2_fill_1 FILLER_8_278 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_4 FILLER_8_368 ();
 sg13g2_fill_1 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_4 ();
 sg13g2_fill_1 FILLER_9_61 ();
 sg13g2_fill_1 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_123 ();
 sg13g2_fill_2 FILLER_9_133 ();
 sg13g2_fill_1 FILLER_9_135 ();
 sg13g2_decap_4 FILLER_9_141 ();
 sg13g2_fill_2 FILLER_9_145 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_fill_2 FILLER_9_157 ();
 sg13g2_fill_1 FILLER_9_197 ();
 sg13g2_fill_2 FILLER_9_216 ();
 sg13g2_fill_2 FILLER_9_236 ();
 sg13g2_fill_1 FILLER_9_238 ();
 sg13g2_fill_2 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_fill_1 FILLER_9_324 ();
 sg13g2_fill_2 FILLER_9_335 ();
 sg13g2_fill_2 FILLER_9_347 ();
 sg13g2_fill_1 FILLER_9_357 ();
 sg13g2_fill_2 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_fill_2 FILLER_9_377 ();
 sg13g2_fill_1 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_11 ();
 sg13g2_fill_2 FILLER_10_16 ();
 sg13g2_fill_1 FILLER_10_18 ();
 sg13g2_fill_1 FILLER_10_31 ();
 sg13g2_fill_1 FILLER_10_53 ();
 sg13g2_fill_2 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_fill_2 FILLER_10_175 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_fill_2 FILLER_10_271 ();
 sg13g2_fill_1 FILLER_10_327 ();
 sg13g2_fill_2 FILLER_10_335 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_fill_2 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_15 ();
 sg13g2_fill_1 FILLER_11_25 ();
 sg13g2_fill_2 FILLER_11_40 ();
 sg13g2_fill_1 FILLER_11_54 ();
 sg13g2_fill_2 FILLER_11_81 ();
 sg13g2_fill_2 FILLER_11_99 ();
 sg13g2_fill_1 FILLER_11_101 ();
 sg13g2_fill_2 FILLER_11_125 ();
 sg13g2_fill_1 FILLER_11_127 ();
 sg13g2_decap_8 FILLER_11_150 ();
 sg13g2_fill_1 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_193 ();
 sg13g2_fill_2 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_201 ();
 sg13g2_fill_1 FILLER_11_259 ();
 sg13g2_decap_4 FILLER_11_272 ();
 sg13g2_fill_1 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_fill_2 FILLER_11_315 ();
 sg13g2_fill_1 FILLER_11_338 ();
 sg13g2_fill_1 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_60 ();
 sg13g2_fill_1 FILLER_12_65 ();
 sg13g2_fill_2 FILLER_12_70 ();
 sg13g2_fill_2 FILLER_12_81 ();
 sg13g2_fill_2 FILLER_12_96 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_fill_2 FILLER_12_224 ();
 sg13g2_fill_2 FILLER_12_241 ();
 sg13g2_fill_1 FILLER_12_243 ();
 sg13g2_fill_2 FILLER_12_254 ();
 sg13g2_fill_1 FILLER_12_256 ();
 sg13g2_fill_1 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_303 ();
 sg13g2_decap_4 FILLER_12_312 ();
 sg13g2_decap_4 FILLER_12_321 ();
 sg13g2_fill_2 FILLER_12_334 ();
 sg13g2_fill_1 FILLER_12_345 ();
 sg13g2_decap_4 FILLER_12_369 ();
 sg13g2_fill_2 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_69 ();
 sg13g2_fill_1 FILLER_13_76 ();
 sg13g2_fill_1 FILLER_13_83 ();
 sg13g2_decap_8 FILLER_13_92 ();
 sg13g2_decap_4 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_125 ();
 sg13g2_fill_2 FILLER_13_139 ();
 sg13g2_fill_1 FILLER_13_233 ();
 sg13g2_fill_1 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_250 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_283 ();
 sg13g2_fill_1 FILLER_13_285 ();
 sg13g2_fill_2 FILLER_13_311 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_decap_4 FILLER_13_347 ();
 sg13g2_fill_2 FILLER_13_351 ();
 sg13g2_fill_2 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_11 ();
 sg13g2_fill_1 FILLER_14_26 ();
 sg13g2_fill_1 FILLER_14_36 ();
 sg13g2_fill_1 FILLER_14_101 ();
 sg13g2_fill_2 FILLER_14_112 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_fill_1 FILLER_14_197 ();
 sg13g2_fill_2 FILLER_14_216 ();
 sg13g2_fill_1 FILLER_14_223 ();
 sg13g2_decap_4 FILLER_14_234 ();
 sg13g2_fill_2 FILLER_14_238 ();
 sg13g2_fill_2 FILLER_14_255 ();
 sg13g2_decap_8 FILLER_14_267 ();
 sg13g2_decap_8 FILLER_14_274 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_decap_4 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_302 ();
 sg13g2_decap_4 FILLER_14_335 ();
 sg13g2_decap_4 FILLER_14_342 ();
 sg13g2_fill_1 FILLER_14_346 ();
 sg13g2_decap_4 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_15_60 ();
 sg13g2_fill_2 FILLER_15_86 ();
 sg13g2_fill_1 FILLER_15_121 ();
 sg13g2_fill_2 FILLER_15_126 ();
 sg13g2_decap_4 FILLER_15_146 ();
 sg13g2_fill_1 FILLER_15_150 ();
 sg13g2_decap_8 FILLER_15_156 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_2 FILLER_15_186 ();
 sg13g2_fill_1 FILLER_15_188 ();
 sg13g2_fill_2 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_242 ();
 sg13g2_fill_2 FILLER_15_256 ();
 sg13g2_fill_2 FILLER_15_266 ();
 sg13g2_fill_1 FILLER_15_268 ();
 sg13g2_fill_1 FILLER_15_277 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_decap_4 FILLER_15_306 ();
 sg13g2_fill_2 FILLER_15_322 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_fill_2 FILLER_16_104 ();
 sg13g2_fill_1 FILLER_16_106 ();
 sg13g2_fill_2 FILLER_16_143 ();
 sg13g2_fill_1 FILLER_16_145 ();
 sg13g2_fill_2 FILLER_16_151 ();
 sg13g2_fill_2 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_194 ();
 sg13g2_decap_4 FILLER_16_207 ();
 sg13g2_fill_1 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_fill_1 FILLER_16_362 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_1 FILLER_17_17 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_fill_1 FILLER_17_74 ();
 sg13g2_fill_2 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_decap_4 FILLER_17_201 ();
 sg13g2_fill_2 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_291 ();
 sg13g2_fill_1 FILLER_17_301 ();
 sg13g2_fill_2 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_313 ();
 sg13g2_fill_2 FILLER_17_320 ();
 sg13g2_fill_1 FILLER_17_322 ();
 sg13g2_fill_2 FILLER_17_334 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_fill_1 FILLER_17_346 ();
 sg13g2_fill_2 FILLER_17_360 ();
 sg13g2_fill_2 FILLER_17_371 ();
 sg13g2_fill_1 FILLER_17_373 ();
 sg13g2_fill_2 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_fill_2 FILLER_18_26 ();
 sg13g2_decap_4 FILLER_18_57 ();
 sg13g2_fill_2 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_67 ();
 sg13g2_fill_1 FILLER_18_83 ();
 sg13g2_fill_2 FILLER_18_94 ();
 sg13g2_fill_1 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_120 ();
 sg13g2_fill_1 FILLER_18_122 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_269 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_321 ();
 sg13g2_decap_4 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_decap_4 FILLER_18_364 ();
 sg13g2_fill_2 FILLER_18_368 ();
 sg13g2_fill_1 FILLER_18_383 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_fill_2 FILLER_19_127 ();
 sg13g2_fill_2 FILLER_19_151 ();
 sg13g2_fill_1 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_178 ();
 sg13g2_decap_8 FILLER_19_205 ();
 sg13g2_decap_8 FILLER_19_212 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_263 ();
 sg13g2_fill_1 FILLER_19_265 ();
 sg13g2_fill_2 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_294 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_fill_2 FILLER_19_308 ();
 sg13g2_fill_2 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_fill_1 FILLER_19_344 ();
 sg13g2_fill_2 FILLER_19_353 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_fill_1 FILLER_20_95 ();
 sg13g2_decap_4 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_decap_4 FILLER_20_215 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_4 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_decap_4 FILLER_20_241 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_296 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_313 ();
 sg13g2_fill_1 FILLER_20_315 ();
 sg13g2_fill_2 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_344 ();
 sg13g2_fill_1 FILLER_20_351 ();
 sg13g2_fill_2 FILLER_20_360 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_6 ();
 sg13g2_decap_4 FILLER_21_13 ();
 sg13g2_fill_1 FILLER_21_30 ();
 sg13g2_fill_1 FILLER_21_38 ();
 sg13g2_decap_8 FILLER_21_43 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_fill_1 FILLER_21_52 ();
 sg13g2_fill_1 FILLER_21_79 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_122 ();
 sg13g2_fill_2 FILLER_21_137 ();
 sg13g2_fill_1 FILLER_21_139 ();
 sg13g2_decap_4 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_4 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_283 ();
 sg13g2_fill_2 FILLER_21_298 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_fill_2 FILLER_21_357 ();
 sg13g2_decap_4 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_44 ();
 sg13g2_decap_4 FILLER_22_50 ();
 sg13g2_fill_1 FILLER_22_110 ();
 sg13g2_fill_1 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_129 ();
 sg13g2_decap_8 FILLER_22_136 ();
 sg13g2_fill_2 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_150 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_237 ();
 sg13g2_fill_1 FILLER_22_239 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_fill_1 FILLER_22_334 ();
 sg13g2_decap_4 FILLER_22_339 ();
 sg13g2_fill_2 FILLER_22_371 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_6 ();
 sg13g2_fill_1 FILLER_23_10 ();
 sg13g2_fill_2 FILLER_23_15 ();
 sg13g2_fill_1 FILLER_23_17 ();
 sg13g2_fill_2 FILLER_23_22 ();
 sg13g2_fill_1 FILLER_23_24 ();
 sg13g2_fill_2 FILLER_23_61 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_fill_2 FILLER_23_186 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_326 ();
 sg13g2_fill_1 FILLER_23_328 ();
 sg13g2_decap_4 FILLER_23_333 ();
 sg13g2_decap_4 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_350 ();
 sg13g2_fill_1 FILLER_23_362 ();
 sg13g2_fill_2 FILLER_23_368 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_fill_2 FILLER_24_56 ();
 sg13g2_decap_4 FILLER_24_137 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_2 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_decap_4 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_361 ();
 sg13g2_decap_4 FILLER_24_377 ();
 sg13g2_fill_2 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_53 ();
 sg13g2_fill_2 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_fill_2 FILLER_25_139 ();
 sg13g2_fill_1 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_decap_8 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_245 ();
 sg13g2_fill_1 FILLER_25_247 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_fill_2 FILLER_25_299 ();
 sg13g2_fill_2 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_4 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_fill_2 FILLER_26_62 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_fill_2 FILLER_26_101 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_decap_8 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_155 ();
 sg13g2_decap_4 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_199 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_231 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_fill_2 FILLER_26_261 ();
 sg13g2_fill_1 FILLER_26_263 ();
 sg13g2_fill_2 FILLER_26_283 ();
 sg13g2_fill_1 FILLER_26_293 ();
 sg13g2_decap_4 FILLER_26_347 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_fill_1 FILLER_27_62 ();
 sg13g2_fill_1 FILLER_27_71 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_fill_2 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_fill_2 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_59 ();
 sg13g2_fill_1 FILLER_28_90 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_207 ();
 sg13g2_decap_4 FILLER_28_225 ();
 sg13g2_decap_4 FILLER_28_234 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_decap_4 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_fill_2 FILLER_28_329 ();
 sg13g2_decap_4 FILLER_28_335 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_decap_4 FILLER_28_350 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_93 ();
 sg13g2_fill_1 FILLER_29_95 ();
 sg13g2_fill_2 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_decap_8 FILLER_29_204 ();
 sg13g2_decap_8 FILLER_29_211 ();
 sg13g2_decap_4 FILLER_29_218 ();
 sg13g2_fill_1 FILLER_29_222 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_278 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_decap_4 FILLER_29_295 ();
 sg13g2_fill_2 FILLER_29_299 ();
 sg13g2_fill_2 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_fill_1 FILLER_29_374 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_fill_1 FILLER_30_34 ();
 sg13g2_fill_2 FILLER_30_107 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_fill_2 FILLER_30_164 ();
 sg13g2_fill_2 FILLER_30_191 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_decap_4 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_214 ();
 sg13g2_decap_8 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_decap_4 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_31_74 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_115 ();
 sg13g2_fill_2 FILLER_31_137 ();
 sg13g2_decap_4 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_fill_1 FILLER_32_13 ();
 sg13g2_fill_2 FILLER_32_19 ();
 sg13g2_fill_2 FILLER_32_34 ();
 sg13g2_fill_1 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_131 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_4 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_decap_4 FILLER_32_267 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_fill_2 FILLER_32_302 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_361 ();
 sg13g2_decap_4 FILLER_32_378 ();
 sg13g2_fill_2 FILLER_32_382 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_1 FILLER_33_26 ();
 sg13g2_fill_2 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_decap_8 FILLER_33_167 ();
 sg13g2_fill_2 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_197 ();
 sg13g2_decap_4 FILLER_33_215 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_239 ();
 sg13g2_decap_8 FILLER_33_246 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_decap_4 FILLER_33_289 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_fill_2 FILLER_33_317 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_fill_1 FILLER_34_71 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_118 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_133 ();
 sg13g2_fill_1 FILLER_34_135 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_decap_4 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_fill_2 FILLER_34_329 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_81 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_104 ();
 sg13g2_fill_1 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_163 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_2 FILLER_35_209 ();
 sg13g2_fill_1 FILLER_35_241 ();
 sg13g2_fill_1 FILLER_35_247 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_315 ();
 sg13g2_decap_4 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_361 ();
 sg13g2_fill_2 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_372 ();
 sg13g2_fill_2 FILLER_35_378 ();
 sg13g2_fill_1 FILLER_35_380 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_1 FILLER_36_69 ();
 sg13g2_decap_8 FILLER_36_82 ();
 sg13g2_decap_8 FILLER_36_89 ();
 sg13g2_decap_4 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_100 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_fill_2 FILLER_36_146 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_2 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_2 FILLER_37_26 ();
 sg13g2_decap_8 FILLER_37_80 ();
 sg13g2_fill_2 FILLER_37_87 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_fill_2 FILLER_37_153 ();
 sg13g2_decap_4 FILLER_37_164 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_173 ();
 sg13g2_fill_2 FILLER_37_180 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_decap_8 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_300 ();
 sg13g2_fill_1 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_368 ();
 sg13g2_fill_1 FILLER_37_384 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_2 FILLER_38_17 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_145 ();
 sg13g2_decap_8 FILLER_38_166 ();
 sg13g2_fill_2 FILLER_38_173 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_202 ();
 sg13g2_fill_1 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_209 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_decap_4 FILLER_38_269 ();
 sg13g2_decap_8 FILLER_38_281 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_fill_1 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_fill_2 FILLER_38_348 ();
 sg13g2_fill_2 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_fill_1 FILLER_39_31 ();
 sg13g2_fill_2 FILLER_39_47 ();
 sg13g2_fill_1 FILLER_39_49 ();
 sg13g2_fill_1 FILLER_39_63 ();
 sg13g2_decap_4 FILLER_39_108 ();
 sg13g2_fill_2 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_118 ();
 sg13g2_decap_8 FILLER_39_131 ();
 sg13g2_decap_8 FILLER_39_141 ();
 sg13g2_fill_2 FILLER_39_166 ();
 sg13g2_decap_8 FILLER_39_213 ();
 sg13g2_fill_2 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_256 ();
 sg13g2_decap_8 FILLER_39_263 ();
 sg13g2_fill_2 FILLER_39_270 ();
 sg13g2_fill_1 FILLER_39_272 ();
 sg13g2_fill_1 FILLER_39_281 ();
 sg13g2_decap_8 FILLER_39_302 ();
 sg13g2_fill_2 FILLER_39_338 ();
 sg13g2_fill_2 FILLER_39_345 ();
 sg13g2_fill_1 FILLER_39_347 ();
 sg13g2_fill_2 FILLER_39_361 ();
 sg13g2_fill_1 FILLER_39_363 ();
 sg13g2_decap_8 FILLER_39_396 ();
 sg13g2_decap_4 FILLER_39_403 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_2 FILLER_40_114 ();
 sg13g2_fill_1 FILLER_40_116 ();
 sg13g2_fill_1 FILLER_40_143 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_207 ();
 sg13g2_fill_2 FILLER_40_267 ();
 sg13g2_fill_1 FILLER_40_269 ();
 sg13g2_decap_4 FILLER_40_299 ();
 sg13g2_fill_1 FILLER_40_303 ();
 sg13g2_fill_1 FILLER_40_327 ();
 sg13g2_fill_1 FILLER_40_333 ();
 sg13g2_decap_4 FILLER_40_339 ();
 sg13g2_fill_1 FILLER_40_348 ();
 sg13g2_fill_1 FILLER_40_369 ();
 sg13g2_fill_2 FILLER_40_378 ();
 sg13g2_fill_1 FILLER_40_380 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_22 ();
 sg13g2_fill_1 FILLER_41_54 ();
 sg13g2_fill_2 FILLER_41_64 ();
 sg13g2_fill_1 FILLER_41_66 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_fill_1 FILLER_41_163 ();
 sg13g2_fill_2 FILLER_41_200 ();
 sg13g2_fill_1 FILLER_41_202 ();
 sg13g2_fill_2 FILLER_41_242 ();
 sg13g2_fill_1 FILLER_41_252 ();
 sg13g2_decap_4 FILLER_41_293 ();
 sg13g2_fill_1 FILLER_41_313 ();
 sg13g2_fill_1 FILLER_41_335 ();
 sg13g2_fill_1 FILLER_41_352 ();
 sg13g2_fill_1 FILLER_41_371 ();
 sg13g2_fill_2 FILLER_41_385 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_5 ();
 sg13g2_decap_8 FILLER_42_12 ();
 sg13g2_fill_2 FILLER_42_19 ();
 sg13g2_fill_2 FILLER_42_30 ();
 sg13g2_fill_1 FILLER_42_41 ();
 sg13g2_fill_1 FILLER_42_56 ();
 sg13g2_fill_2 FILLER_42_65 ();
 sg13g2_fill_2 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_91 ();
 sg13g2_decap_4 FILLER_42_96 ();
 sg13g2_fill_1 FILLER_42_100 ();
 sg13g2_fill_2 FILLER_42_109 ();
 sg13g2_decap_4 FILLER_42_116 ();
 sg13g2_fill_1 FILLER_42_139 ();
 sg13g2_fill_1 FILLER_42_151 ();
 sg13g2_fill_2 FILLER_42_158 ();
 sg13g2_fill_1 FILLER_42_170 ();
 sg13g2_decap_4 FILLER_42_179 ();
 sg13g2_fill_2 FILLER_42_183 ();
 sg13g2_fill_2 FILLER_42_189 ();
 sg13g2_fill_1 FILLER_42_191 ();
 sg13g2_decap_4 FILLER_42_264 ();
 sg13g2_fill_2 FILLER_42_268 ();
 sg13g2_fill_2 FILLER_42_298 ();
 sg13g2_fill_2 FILLER_42_306 ();
 sg13g2_decap_8 FILLER_42_334 ();
 sg13g2_decap_8 FILLER_42_341 ();
 sg13g2_fill_2 FILLER_42_348 ();
 sg13g2_decap_8 FILLER_42_353 ();
 sg13g2_decap_4 FILLER_42_360 ();
 sg13g2_fill_2 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_4 FILLER_42_403 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_4 FILLER_43_26 ();
 sg13g2_fill_2 FILLER_43_43 ();
 sg13g2_fill_1 FILLER_43_68 ();
 sg13g2_fill_1 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_90 ();
 sg13g2_decap_4 FILLER_43_96 ();
 sg13g2_fill_1 FILLER_43_100 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_4 FILLER_43_119 ();
 sg13g2_decap_4 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_165 ();
 sg13g2_decap_4 FILLER_43_170 ();
 sg13g2_fill_1 FILLER_43_203 ();
 sg13g2_fill_1 FILLER_43_219 ();
 sg13g2_decap_4 FILLER_43_229 ();
 sg13g2_fill_2 FILLER_43_238 ();
 sg13g2_fill_1 FILLER_43_240 ();
 sg13g2_decap_4 FILLER_43_246 ();
 sg13g2_fill_1 FILLER_43_250 ();
 sg13g2_decap_4 FILLER_43_259 ();
 sg13g2_fill_1 FILLER_43_263 ();
 sg13g2_fill_1 FILLER_43_276 ();
 sg13g2_decap_8 FILLER_43_326 ();
 sg13g2_decap_8 FILLER_43_333 ();
 sg13g2_decap_8 FILLER_43_340 ();
 sg13g2_decap_8 FILLER_43_347 ();
 sg13g2_decap_8 FILLER_43_354 ();
 sg13g2_decap_8 FILLER_43_361 ();
 sg13g2_decap_8 FILLER_43_368 ();
 sg13g2_decap_4 FILLER_43_375 ();
 sg13g2_decap_8 FILLER_43_393 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_4 FILLER_44_26 ();
 sg13g2_fill_1 FILLER_44_30 ();
 sg13g2_fill_2 FILLER_44_57 ();
 sg13g2_fill_2 FILLER_44_73 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_fill_2 FILLER_44_101 ();
 sg13g2_fill_2 FILLER_44_130 ();
 sg13g2_decap_4 FILLER_44_142 ();
 sg13g2_decap_8 FILLER_44_188 ();
 sg13g2_fill_2 FILLER_44_195 ();
 sg13g2_fill_1 FILLER_44_197 ();
 sg13g2_fill_2 FILLER_44_203 ();
 sg13g2_fill_1 FILLER_44_205 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_fill_1 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_222 ();
 sg13g2_fill_1 FILLER_44_237 ();
 sg13g2_fill_2 FILLER_44_245 ();
 sg13g2_decap_4 FILLER_44_259 ();
 sg13g2_fill_1 FILLER_44_263 ();
 sg13g2_decap_4 FILLER_44_270 ();
 sg13g2_fill_2 FILLER_44_306 ();
 sg13g2_fill_1 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_330 ();
 sg13g2_decap_4 FILLER_44_349 ();
 sg13g2_fill_1 FILLER_44_373 ();
 sg13g2_fill_2 FILLER_44_378 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_19 ();
 sg13g2_fill_1 FILLER_45_38 ();
 sg13g2_fill_2 FILLER_45_73 ();
 sg13g2_fill_2 FILLER_45_90 ();
 sg13g2_fill_2 FILLER_45_129 ();
 sg13g2_decap_4 FILLER_45_136 ();
 sg13g2_fill_2 FILLER_45_140 ();
 sg13g2_fill_1 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_173 ();
 sg13g2_fill_1 FILLER_45_180 ();
 sg13g2_fill_1 FILLER_45_189 ();
 sg13g2_fill_1 FILLER_45_194 ();
 sg13g2_fill_2 FILLER_45_220 ();
 sg13g2_fill_2 FILLER_45_239 ();
 sg13g2_fill_2 FILLER_45_247 ();
 sg13g2_fill_1 FILLER_45_263 ();
 sg13g2_fill_2 FILLER_45_282 ();
 sg13g2_fill_1 FILLER_45_284 ();
 sg13g2_fill_2 FILLER_45_290 ();
 sg13g2_decap_8 FILLER_45_305 ();
 sg13g2_decap_8 FILLER_45_312 ();
 sg13g2_decap_8 FILLER_45_319 ();
 sg13g2_fill_1 FILLER_45_351 ();
 sg13g2_fill_2 FILLER_45_373 ();
 sg13g2_fill_2 FILLER_45_383 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_4 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_18 ();
 sg13g2_decap_4 FILLER_46_141 ();
 sg13g2_fill_2 FILLER_46_150 ();
 sg13g2_fill_2 FILLER_46_156 ();
 sg13g2_decap_8 FILLER_46_163 ();
 sg13g2_fill_2 FILLER_46_170 ();
 sg13g2_fill_2 FILLER_46_177 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_decap_4 FILLER_46_226 ();
 sg13g2_fill_1 FILLER_46_230 ();
 sg13g2_decap_8 FILLER_46_251 ();
 sg13g2_decap_8 FILLER_46_258 ();
 sg13g2_decap_8 FILLER_46_265 ();
 sg13g2_fill_2 FILLER_46_301 ();
 sg13g2_fill_2 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_fill_1 FILLER_46_322 ();
 sg13g2_fill_1 FILLER_46_365 ();
 sg13g2_fill_2 FILLER_46_386 ();
 sg13g2_fill_1 FILLER_47_60 ();
 sg13g2_fill_2 FILLER_47_68 ();
 sg13g2_fill_2 FILLER_47_91 ();
 sg13g2_fill_1 FILLER_47_124 ();
 sg13g2_fill_2 FILLER_47_133 ();
 sg13g2_decap_4 FILLER_47_148 ();
 sg13g2_fill_2 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_fill_1 FILLER_47_201 ();
 sg13g2_fill_2 FILLER_47_250 ();
 sg13g2_fill_1 FILLER_47_252 ();
 sg13g2_fill_2 FILLER_47_265 ();
 sg13g2_fill_2 FILLER_47_272 ();
 sg13g2_fill_1 FILLER_47_324 ();
 sg13g2_fill_2 FILLER_47_337 ();
 sg13g2_fill_2 FILLER_47_385 ();
 sg13g2_fill_1 FILLER_47_395 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_fill_2 FILLER_48_36 ();
 sg13g2_fill_2 FILLER_48_78 ();
 sg13g2_fill_1 FILLER_48_80 ();
 sg13g2_fill_2 FILLER_48_101 ();
 sg13g2_fill_1 FILLER_48_103 ();
 sg13g2_decap_4 FILLER_48_108 ();
 sg13g2_fill_1 FILLER_48_112 ();
 sg13g2_fill_2 FILLER_48_121 ();
 sg13g2_fill_1 FILLER_48_123 ();
 sg13g2_fill_1 FILLER_48_169 ();
 sg13g2_decap_8 FILLER_48_195 ();
 sg13g2_decap_8 FILLER_48_207 ();
 sg13g2_decap_8 FILLER_48_214 ();
 sg13g2_decap_4 FILLER_48_221 ();
 sg13g2_fill_1 FILLER_48_225 ();
 sg13g2_decap_4 FILLER_48_231 ();
 sg13g2_fill_2 FILLER_48_240 ();
 sg13g2_fill_2 FILLER_48_250 ();
 sg13g2_fill_2 FILLER_48_257 ();
 sg13g2_fill_1 FILLER_48_259 ();
 sg13g2_fill_2 FILLER_48_309 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_fill_2 FILLER_48_330 ();
 sg13g2_fill_1 FILLER_48_332 ();
 sg13g2_fill_1 FILLER_48_345 ();
 sg13g2_decap_4 FILLER_48_349 ();
 sg13g2_fill_2 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_359 ();
 sg13g2_fill_1 FILLER_48_361 ();
 sg13g2_fill_1 FILLER_48_377 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_4 FILLER_49_3 ();
 sg13g2_fill_1 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_28 ();
 sg13g2_fill_2 FILLER_49_52 ();
 sg13g2_fill_2 FILLER_49_85 ();
 sg13g2_fill_1 FILLER_49_103 ();
 sg13g2_decap_4 FILLER_49_108 ();
 sg13g2_fill_2 FILLER_49_112 ();
 sg13g2_fill_2 FILLER_49_161 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_4 FILLER_49_196 ();
 sg13g2_fill_2 FILLER_49_209 ();
 sg13g2_fill_1 FILLER_49_211 ();
 sg13g2_fill_2 FILLER_49_237 ();
 sg13g2_fill_2 FILLER_49_243 ();
 sg13g2_fill_2 FILLER_49_262 ();
 sg13g2_fill_1 FILLER_49_264 ();
 sg13g2_fill_1 FILLER_49_339 ();
 sg13g2_fill_2 FILLER_49_356 ();
 sg13g2_decap_4 FILLER_49_375 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_22 ();
 sg13g2_fill_2 FILLER_50_56 ();
 sg13g2_fill_1 FILLER_50_69 ();
 sg13g2_fill_1 FILLER_50_84 ();
 sg13g2_fill_1 FILLER_50_106 ();
 sg13g2_fill_1 FILLER_50_114 ();
 sg13g2_fill_2 FILLER_50_124 ();
 sg13g2_decap_8 FILLER_50_185 ();
 sg13g2_fill_2 FILLER_50_192 ();
 sg13g2_fill_1 FILLER_50_223 ();
 sg13g2_fill_2 FILLER_50_240 ();
 sg13g2_fill_2 FILLER_50_268 ();
 sg13g2_fill_2 FILLER_50_282 ();
 sg13g2_fill_1 FILLER_50_284 ();
 sg13g2_decap_4 FILLER_50_303 ();
 sg13g2_fill_1 FILLER_50_307 ();
 sg13g2_decap_8 FILLER_50_312 ();
 sg13g2_fill_2 FILLER_50_348 ();
 sg13g2_fill_1 FILLER_50_366 ();
 sg13g2_fill_2 FILLER_50_389 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_26 ();
 sg13g2_fill_2 FILLER_51_75 ();
 sg13g2_fill_1 FILLER_51_93 ();
 sg13g2_fill_1 FILLER_51_169 ();
 sg13g2_fill_1 FILLER_51_193 ();
 sg13g2_fill_1 FILLER_51_240 ();
 sg13g2_fill_1 FILLER_51_250 ();
 sg13g2_decap_8 FILLER_51_260 ();
 sg13g2_decap_8 FILLER_51_267 ();
 sg13g2_decap_8 FILLER_51_274 ();
 sg13g2_decap_8 FILLER_51_281 ();
 sg13g2_decap_4 FILLER_51_293 ();
 sg13g2_fill_2 FILLER_51_297 ();
 sg13g2_decap_8 FILLER_51_308 ();
 sg13g2_fill_2 FILLER_51_315 ();
 sg13g2_fill_1 FILLER_51_317 ();
 sg13g2_fill_1 FILLER_51_337 ();
 sg13g2_fill_1 FILLER_51_361 ();
 sg13g2_fill_2 FILLER_51_378 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_fill_2 FILLER_52_31 ();
 sg13g2_fill_2 FILLER_52_56 ();
 sg13g2_fill_1 FILLER_52_76 ();
 sg13g2_fill_1 FILLER_52_86 ();
 sg13g2_fill_2 FILLER_52_96 ();
 sg13g2_fill_1 FILLER_52_98 ();
 sg13g2_fill_2 FILLER_52_106 ();
 sg13g2_fill_1 FILLER_52_108 ();
 sg13g2_fill_1 FILLER_52_133 ();
 sg13g2_fill_2 FILLER_52_155 ();
 sg13g2_fill_2 FILLER_52_162 ();
 sg13g2_fill_1 FILLER_52_164 ();
 sg13g2_fill_2 FILLER_52_190 ();
 sg13g2_fill_1 FILLER_52_192 ();
 sg13g2_fill_1 FILLER_52_203 ();
 sg13g2_fill_1 FILLER_52_225 ();
 sg13g2_decap_8 FILLER_52_231 ();
 sg13g2_decap_4 FILLER_52_238 ();
 sg13g2_decap_8 FILLER_52_256 ();
 sg13g2_decap_8 FILLER_52_263 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_decap_8 FILLER_52_279 ();
 sg13g2_decap_4 FILLER_52_286 ();
 sg13g2_decap_8 FILLER_52_299 ();
 sg13g2_decap_8 FILLER_52_306 ();
 sg13g2_fill_1 FILLER_52_313 ();
 sg13g2_fill_2 FILLER_52_343 ();
 sg13g2_fill_1 FILLER_52_345 ();
 sg13g2_fill_1 FILLER_52_354 ();
 sg13g2_fill_1 FILLER_52_363 ();
 sg13g2_decap_4 FILLER_52_381 ();
 sg13g2_fill_1 FILLER_52_397 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_18 ();
 sg13g2_fill_1 FILLER_53_20 ();
 sg13g2_fill_2 FILLER_53_73 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_fill_2 FILLER_53_112 ();
 sg13g2_fill_2 FILLER_53_129 ();
 sg13g2_fill_1 FILLER_53_131 ();
 sg13g2_decap_8 FILLER_53_193 ();
 sg13g2_decap_4 FILLER_53_200 ();
 sg13g2_fill_2 FILLER_53_208 ();
 sg13g2_fill_2 FILLER_53_218 ();
 sg13g2_fill_2 FILLER_53_241 ();
 sg13g2_fill_1 FILLER_53_243 ();
 sg13g2_decap_4 FILLER_53_264 ();
 sg13g2_decap_4 FILLER_53_277 ();
 sg13g2_fill_2 FILLER_53_299 ();
 sg13g2_decap_4 FILLER_53_317 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_fill_1 FILLER_53_332 ();
 sg13g2_fill_2 FILLER_53_346 ();
 sg13g2_fill_1 FILLER_53_348 ();
 sg13g2_fill_1 FILLER_53_362 ();
 sg13g2_decap_4 FILLER_53_380 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_fill_2 FILLER_54_30 ();
 sg13g2_fill_1 FILLER_54_32 ();
 sg13g2_fill_1 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_88 ();
 sg13g2_fill_2 FILLER_54_99 ();
 sg13g2_fill_2 FILLER_54_111 ();
 sg13g2_fill_2 FILLER_54_127 ();
 sg13g2_fill_1 FILLER_54_129 ();
 sg13g2_fill_2 FILLER_54_149 ();
 sg13g2_fill_1 FILLER_54_178 ();
 sg13g2_fill_1 FILLER_54_196 ();
 sg13g2_fill_2 FILLER_54_241 ();
 sg13g2_fill_1 FILLER_54_243 ();
 sg13g2_fill_2 FILLER_54_271 ();
 sg13g2_decap_4 FILLER_54_316 ();
 sg13g2_decap_4 FILLER_54_323 ();
 sg13g2_decap_4 FILLER_54_330 ();
 sg13g2_decap_4 FILLER_54_357 ();
 sg13g2_decap_4 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_380 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_18 ();
 sg13g2_fill_1 FILLER_55_93 ();
 sg13g2_fill_1 FILLER_55_102 ();
 sg13g2_fill_2 FILLER_55_111 ();
 sg13g2_decap_4 FILLER_55_135 ();
 sg13g2_fill_1 FILLER_55_185 ();
 sg13g2_fill_2 FILLER_55_216 ();
 sg13g2_fill_1 FILLER_55_218 ();
 sg13g2_fill_1 FILLER_55_232 ();
 sg13g2_fill_1 FILLER_55_278 ();
 sg13g2_decap_4 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_318 ();
 sg13g2_fill_1 FILLER_55_328 ();
 sg13g2_fill_2 FILLER_55_337 ();
 sg13g2_fill_1 FILLER_55_339 ();
 sg13g2_fill_1 FILLER_55_350 ();
 sg13g2_fill_2 FILLER_55_377 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_5 ();
 sg13g2_fill_1 FILLER_56_22 ();
 sg13g2_fill_2 FILLER_56_28 ();
 sg13g2_fill_1 FILLER_56_30 ();
 sg13g2_decap_4 FILLER_56_128 ();
 sg13g2_decap_4 FILLER_56_164 ();
 sg13g2_decap_8 FILLER_56_180 ();
 sg13g2_fill_1 FILLER_56_187 ();
 sg13g2_decap_8 FILLER_56_212 ();
 sg13g2_fill_1 FILLER_56_219 ();
 sg13g2_decap_4 FILLER_56_224 ();
 sg13g2_fill_1 FILLER_56_228 ();
 sg13g2_decap_8 FILLER_56_233 ();
 sg13g2_decap_4 FILLER_56_240 ();
 sg13g2_fill_2 FILLER_56_244 ();
 sg13g2_fill_2 FILLER_56_271 ();
 sg13g2_fill_1 FILLER_56_273 ();
 sg13g2_fill_1 FILLER_56_312 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_2 FILLER_57_20 ();
 sg13g2_decap_8 FILLER_57_26 ();
 sg13g2_decap_4 FILLER_57_33 ();
 sg13g2_fill_1 FILLER_57_37 ();
 sg13g2_fill_2 FILLER_57_104 ();
 sg13g2_fill_2 FILLER_57_134 ();
 sg13g2_decap_8 FILLER_57_170 ();
 sg13g2_fill_2 FILLER_57_177 ();
 sg13g2_fill_1 FILLER_57_179 ();
 sg13g2_decap_8 FILLER_57_206 ();
 sg13g2_decap_8 FILLER_57_213 ();
 sg13g2_decap_8 FILLER_57_243 ();
 sg13g2_decap_4 FILLER_57_250 ();
 sg13g2_fill_1 FILLER_57_254 ();
 sg13g2_decap_4 FILLER_57_264 ();
 sg13g2_fill_2 FILLER_57_268 ();
 sg13g2_fill_2 FILLER_57_300 ();
 sg13g2_fill_1 FILLER_57_302 ();
 sg13g2_fill_2 FILLER_57_331 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_fill_1 FILLER_58_42 ();
 sg13g2_fill_1 FILLER_58_60 ();
 sg13g2_fill_1 FILLER_58_83 ();
 sg13g2_fill_2 FILLER_58_119 ();
 sg13g2_fill_1 FILLER_58_121 ();
 sg13g2_fill_2 FILLER_58_130 ();
 sg13g2_fill_1 FILLER_58_140 ();
 sg13g2_fill_2 FILLER_58_147 ();
 sg13g2_fill_1 FILLER_58_149 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_182 ();
 sg13g2_fill_1 FILLER_58_184 ();
 sg13g2_fill_1 FILLER_58_201 ();
 sg13g2_decap_8 FILLER_58_211 ();
 sg13g2_fill_1 FILLER_58_222 ();
 sg13g2_decap_4 FILLER_58_253 ();
 sg13g2_fill_1 FILLER_58_257 ();
 sg13g2_fill_2 FILLER_58_267 ();
 sg13g2_fill_1 FILLER_58_269 ();
 sg13g2_decap_4 FILLER_58_294 ();
 sg13g2_decap_4 FILLER_58_308 ();
 sg13g2_fill_2 FILLER_58_312 ();
 sg13g2_fill_2 FILLER_58_332 ();
 sg13g2_fill_1 FILLER_58_334 ();
 sg13g2_decap_8 FILLER_58_346 ();
 sg13g2_fill_2 FILLER_58_353 ();
 sg13g2_decap_8 FILLER_58_359 ();
 sg13g2_decap_4 FILLER_58_366 ();
 sg13g2_decap_8 FILLER_58_380 ();
 sg13g2_decap_8 FILLER_58_387 ();
 sg13g2_fill_1 FILLER_58_394 ();
 sg13g2_decap_4 FILLER_58_405 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_2 ();
 sg13g2_fill_2 FILLER_59_18 ();
 sg13g2_fill_1 FILLER_59_20 ();
 sg13g2_fill_2 FILLER_59_39 ();
 sg13g2_fill_2 FILLER_59_69 ();
 sg13g2_fill_1 FILLER_59_88 ();
 sg13g2_fill_2 FILLER_59_104 ();
 sg13g2_fill_1 FILLER_59_133 ();
 sg13g2_fill_2 FILLER_59_148 ();
 sg13g2_fill_1 FILLER_59_171 ();
 sg13g2_fill_2 FILLER_59_213 ();
 sg13g2_fill_1 FILLER_59_215 ();
 sg13g2_fill_2 FILLER_59_251 ();
 sg13g2_fill_1 FILLER_59_266 ();
 sg13g2_decap_4 FILLER_59_288 ();
 sg13g2_decap_8 FILLER_59_296 ();
 sg13g2_fill_2 FILLER_59_303 ();
 sg13g2_fill_1 FILLER_59_328 ();
 sg13g2_decap_4 FILLER_59_333 ();
 sg13g2_fill_1 FILLER_59_337 ();
 sg13g2_decap_8 FILLER_59_353 ();
 sg13g2_decap_8 FILLER_59_360 ();
 sg13g2_fill_2 FILLER_59_367 ();
 sg13g2_fill_1 FILLER_59_369 ();
 sg13g2_decap_4 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_22 ();
 sg13g2_decap_4 FILLER_60_39 ();
 sg13g2_fill_1 FILLER_60_43 ();
 sg13g2_fill_1 FILLER_60_49 ();
 sg13g2_fill_2 FILLER_60_64 ();
 sg13g2_fill_1 FILLER_60_66 ();
 sg13g2_fill_1 FILLER_60_89 ();
 sg13g2_fill_2 FILLER_60_95 ();
 sg13g2_fill_1 FILLER_60_97 ();
 sg13g2_fill_1 FILLER_60_111 ();
 sg13g2_fill_1 FILLER_60_117 ();
 sg13g2_fill_1 FILLER_60_138 ();
 sg13g2_fill_2 FILLER_60_143 ();
 sg13g2_fill_2 FILLER_60_187 ();
 sg13g2_fill_1 FILLER_60_189 ();
 sg13g2_fill_2 FILLER_60_203 ();
 sg13g2_fill_1 FILLER_60_205 ();
 sg13g2_fill_1 FILLER_60_211 ();
 sg13g2_fill_1 FILLER_60_253 ();
 sg13g2_fill_2 FILLER_60_304 ();
 sg13g2_fill_2 FILLER_60_337 ();
 sg13g2_fill_2 FILLER_60_355 ();
 sg13g2_fill_1 FILLER_60_384 ();
 sg13g2_fill_1 FILLER_60_395 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_decap_4 FILLER_61_25 ();
 sg13g2_fill_1 FILLER_61_29 ();
 sg13g2_fill_2 FILLER_61_39 ();
 sg13g2_fill_1 FILLER_61_76 ();
 sg13g2_fill_1 FILLER_61_85 ();
 sg13g2_fill_2 FILLER_61_117 ();
 sg13g2_fill_1 FILLER_61_142 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_decap_8 FILLER_61_202 ();
 sg13g2_fill_2 FILLER_61_209 ();
 sg13g2_fill_1 FILLER_61_254 ();
 sg13g2_fill_2 FILLER_61_273 ();
 sg13g2_decap_8 FILLER_61_283 ();
 sg13g2_fill_2 FILLER_61_290 ();
 sg13g2_fill_1 FILLER_61_292 ();
 sg13g2_decap_4 FILLER_61_305 ();
 sg13g2_fill_2 FILLER_61_309 ();
 sg13g2_fill_2 FILLER_61_320 ();
 sg13g2_fill_2 FILLER_61_373 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_18 ();
 sg13g2_fill_1 FILLER_62_44 ();
 sg13g2_fill_2 FILLER_62_76 ();
 sg13g2_fill_2 FILLER_62_86 ();
 sg13g2_decap_4 FILLER_62_135 ();
 sg13g2_fill_1 FILLER_62_150 ();
 sg13g2_decap_8 FILLER_62_181 ();
 sg13g2_decap_4 FILLER_62_206 ();
 sg13g2_fill_1 FILLER_62_210 ();
 sg13g2_decap_4 FILLER_62_220 ();
 sg13g2_fill_1 FILLER_62_224 ();
 sg13g2_fill_2 FILLER_62_246 ();
 sg13g2_decap_8 FILLER_62_253 ();
 sg13g2_decap_8 FILLER_62_260 ();
 sg13g2_decap_8 FILLER_62_267 ();
 sg13g2_fill_2 FILLER_62_290 ();
 sg13g2_fill_1 FILLER_62_292 ();
 sg13g2_decap_8 FILLER_62_324 ();
 sg13g2_fill_2 FILLER_62_331 ();
 sg13g2_fill_1 FILLER_62_338 ();
 sg13g2_decap_4 FILLER_62_349 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_fill_2 FILLER_63_52 ();
 sg13g2_fill_1 FILLER_63_97 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_fill_2 FILLER_63_135 ();
 sg13g2_fill_1 FILLER_63_137 ();
 sg13g2_fill_1 FILLER_63_159 ();
 sg13g2_fill_1 FILLER_63_165 ();
 sg13g2_decap_8 FILLER_63_171 ();
 sg13g2_fill_2 FILLER_63_185 ();
 sg13g2_fill_1 FILLER_63_187 ();
 sg13g2_fill_1 FILLER_63_214 ();
 sg13g2_fill_1 FILLER_63_228 ();
 sg13g2_fill_1 FILLER_63_246 ();
 sg13g2_fill_1 FILLER_63_270 ();
 sg13g2_fill_1 FILLER_63_295 ();
 sg13g2_decap_8 FILLER_63_338 ();
 sg13g2_fill_2 FILLER_63_345 ();
 sg13g2_decap_4 FILLER_63_352 ();
 sg13g2_fill_1 FILLER_63_356 ();
 sg13g2_fill_2 FILLER_63_382 ();
 sg13g2_fill_1 FILLER_63_384 ();
 sg13g2_fill_2 FILLER_63_390 ();
 sg13g2_fill_1 FILLER_63_396 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_fill_1 FILLER_64_26 ();
 sg13g2_fill_2 FILLER_64_35 ();
 sg13g2_fill_1 FILLER_64_37 ();
 sg13g2_fill_2 FILLER_64_64 ();
 sg13g2_fill_2 FILLER_64_71 ();
 sg13g2_fill_2 FILLER_64_93 ();
 sg13g2_fill_2 FILLER_64_100 ();
 sg13g2_fill_2 FILLER_64_133 ();
 sg13g2_decap_4 FILLER_64_169 ();
 sg13g2_fill_2 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_184 ();
 sg13g2_decap_4 FILLER_64_219 ();
 sg13g2_fill_2 FILLER_64_239 ();
 sg13g2_fill_2 FILLER_64_246 ();
 sg13g2_fill_2 FILLER_64_273 ();
 sg13g2_fill_2 FILLER_64_284 ();
 sg13g2_fill_1 FILLER_64_286 ();
 sg13g2_fill_2 FILLER_64_296 ();
 sg13g2_fill_2 FILLER_64_308 ();
 sg13g2_decap_4 FILLER_64_340 ();
 sg13g2_decap_4 FILLER_64_349 ();
 sg13g2_fill_2 FILLER_64_361 ();
 sg13g2_fill_1 FILLER_64_363 ();
 sg13g2_fill_2 FILLER_64_382 ();
 sg13g2_fill_1 FILLER_64_384 ();
 sg13g2_fill_1 FILLER_64_394 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_34 ();
 sg13g2_fill_1 FILLER_65_46 ();
 sg13g2_fill_1 FILLER_65_61 ();
 sg13g2_fill_2 FILLER_65_80 ();
 sg13g2_fill_1 FILLER_65_82 ();
 sg13g2_fill_1 FILLER_65_88 ();
 sg13g2_fill_2 FILLER_65_107 ();
 sg13g2_fill_1 FILLER_65_109 ();
 sg13g2_fill_1 FILLER_65_144 ();
 sg13g2_fill_2 FILLER_65_149 ();
 sg13g2_decap_8 FILLER_65_162 ();
 sg13g2_fill_1 FILLER_65_169 ();
 sg13g2_fill_1 FILLER_65_195 ();
 sg13g2_decap_8 FILLER_65_212 ();
 sg13g2_fill_1 FILLER_65_219 ();
 sg13g2_decap_8 FILLER_65_225 ();
 sg13g2_decap_8 FILLER_65_232 ();
 sg13g2_decap_4 FILLER_65_239 ();
 sg13g2_fill_2 FILLER_65_247 ();
 sg13g2_decap_8 FILLER_65_275 ();
 sg13g2_fill_2 FILLER_65_282 ();
 sg13g2_fill_1 FILLER_65_284 ();
 sg13g2_fill_1 FILLER_65_305 ();
 sg13g2_fill_2 FILLER_65_322 ();
 sg13g2_fill_2 FILLER_65_351 ();
 sg13g2_decap_4 FILLER_65_361 ();
 sg13g2_fill_1 FILLER_65_365 ();
 sg13g2_fill_2 FILLER_65_374 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_24 ();
 sg13g2_fill_2 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_37 ();
 sg13g2_fill_1 FILLER_66_74 ();
 sg13g2_fill_2 FILLER_66_90 ();
 sg13g2_fill_1 FILLER_66_92 ();
 sg13g2_fill_2 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_111 ();
 sg13g2_fill_2 FILLER_66_118 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_decap_8 FILLER_66_125 ();
 sg13g2_decap_4 FILLER_66_132 ();
 sg13g2_fill_1 FILLER_66_136 ();
 sg13g2_fill_2 FILLER_66_149 ();
 sg13g2_decap_4 FILLER_66_156 ();
 sg13g2_fill_2 FILLER_66_160 ();
 sg13g2_decap_8 FILLER_66_190 ();
 sg13g2_decap_8 FILLER_66_197 ();
 sg13g2_decap_8 FILLER_66_204 ();
 sg13g2_decap_4 FILLER_66_211 ();
 sg13g2_decap_8 FILLER_66_223 ();
 sg13g2_fill_2 FILLER_66_230 ();
 sg13g2_decap_8 FILLER_66_248 ();
 sg13g2_decap_8 FILLER_66_272 ();
 sg13g2_decap_4 FILLER_66_279 ();
 sg13g2_decap_4 FILLER_66_293 ();
 sg13g2_fill_2 FILLER_66_297 ();
 sg13g2_decap_8 FILLER_66_321 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_fill_1 FILLER_66_344 ();
 sg13g2_fill_1 FILLER_66_357 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_fill_2 FILLER_67_26 ();
 sg13g2_fill_2 FILLER_67_93 ();
 sg13g2_fill_1 FILLER_67_95 ();
 sg13g2_decap_4 FILLER_67_114 ();
 sg13g2_fill_1 FILLER_67_118 ();
 sg13g2_fill_1 FILLER_67_134 ();
 sg13g2_fill_1 FILLER_67_143 ();
 sg13g2_fill_1 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_205 ();
 sg13g2_decap_8 FILLER_67_212 ();
 sg13g2_decap_8 FILLER_67_219 ();
 sg13g2_fill_1 FILLER_67_254 ();
 sg13g2_fill_2 FILLER_67_290 ();
 sg13g2_fill_2 FILLER_67_313 ();
 sg13g2_fill_1 FILLER_67_315 ();
 sg13g2_fill_2 FILLER_67_321 ();
 sg13g2_fill_1 FILLER_67_323 ();
 sg13g2_fill_2 FILLER_67_337 ();
 sg13g2_fill_2 FILLER_67_347 ();
 sg13g2_fill_2 FILLER_67_354 ();
 sg13g2_fill_1 FILLER_67_383 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_20 ();
 sg13g2_fill_1 FILLER_68_26 ();
 sg13g2_fill_1 FILLER_68_63 ();
 sg13g2_fill_1 FILLER_68_72 ();
 sg13g2_fill_1 FILLER_68_77 ();
 sg13g2_fill_2 FILLER_68_97 ();
 sg13g2_fill_1 FILLER_68_99 ();
 sg13g2_fill_2 FILLER_68_105 ();
 sg13g2_fill_2 FILLER_68_117 ();
 sg13g2_fill_1 FILLER_68_127 ();
 sg13g2_fill_1 FILLER_68_167 ();
 sg13g2_fill_1 FILLER_68_181 ();
 sg13g2_fill_1 FILLER_68_186 ();
 sg13g2_decap_4 FILLER_68_211 ();
 sg13g2_fill_1 FILLER_68_215 ();
 sg13g2_decap_4 FILLER_68_271 ();
 sg13g2_fill_1 FILLER_68_280 ();
 sg13g2_decap_8 FILLER_68_294 ();
 sg13g2_decap_8 FILLER_68_301 ();
 sg13g2_fill_1 FILLER_68_308 ();
 sg13g2_fill_2 FILLER_68_331 ();
 sg13g2_fill_1 FILLER_68_333 ();
 sg13g2_fill_1 FILLER_68_344 ();
 sg13g2_fill_2 FILLER_68_380 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_17 ();
 sg13g2_fill_1 FILLER_69_19 ();
 sg13g2_fill_2 FILLER_69_25 ();
 sg13g2_fill_1 FILLER_69_27 ();
 sg13g2_fill_1 FILLER_69_44 ();
 sg13g2_fill_1 FILLER_69_57 ();
 sg13g2_fill_2 FILLER_69_86 ();
 sg13g2_fill_1 FILLER_69_102 ();
 sg13g2_fill_2 FILLER_69_144 ();
 sg13g2_fill_2 FILLER_69_160 ();
 sg13g2_fill_1 FILLER_69_162 ();
 sg13g2_fill_2 FILLER_69_183 ();
 sg13g2_fill_2 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_193 ();
 sg13g2_fill_2 FILLER_69_212 ();
 sg13g2_fill_1 FILLER_69_214 ();
 sg13g2_fill_1 FILLER_69_263 ();
 sg13g2_decap_8 FILLER_69_276 ();
 sg13g2_fill_2 FILLER_69_283 ();
 sg13g2_fill_1 FILLER_69_302 ();
 sg13g2_decap_8 FILLER_69_339 ();
 sg13g2_fill_1 FILLER_69_355 ();
 sg13g2_fill_2 FILLER_69_360 ();
 sg13g2_fill_1 FILLER_69_380 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_25 ();
 sg13g2_fill_1 FILLER_70_27 ();
 sg13g2_fill_2 FILLER_70_33 ();
 sg13g2_fill_2 FILLER_70_102 ();
 sg13g2_fill_1 FILLER_70_104 ();
 sg13g2_fill_1 FILLER_70_128 ();
 sg13g2_fill_1 FILLER_70_143 ();
 sg13g2_fill_2 FILLER_70_174 ();
 sg13g2_fill_1 FILLER_70_176 ();
 sg13g2_fill_2 FILLER_70_184 ();
 sg13g2_fill_2 FILLER_70_191 ();
 sg13g2_fill_1 FILLER_70_268 ();
 sg13g2_decap_8 FILLER_70_276 ();
 sg13g2_fill_1 FILLER_70_283 ();
 sg13g2_fill_2 FILLER_70_297 ();
 sg13g2_fill_2 FILLER_70_325 ();
 sg13g2_fill_1 FILLER_70_327 ();
 sg13g2_decap_8 FILLER_70_345 ();
 sg13g2_decap_8 FILLER_70_352 ();
 sg13g2_fill_1 FILLER_70_359 ();
 sg13g2_fill_2 FILLER_70_386 ();
 sg13g2_fill_1 FILLER_70_388 ();
 sg13g2_decap_8 FILLER_70_401 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_fill_1 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_22 ();
 sg13g2_fill_2 FILLER_71_29 ();
 sg13g2_fill_1 FILLER_71_60 ();
 sg13g2_fill_1 FILLER_71_108 ();
 sg13g2_fill_2 FILLER_71_124 ();
 sg13g2_fill_2 FILLER_71_146 ();
 sg13g2_fill_1 FILLER_71_158 ();
 sg13g2_fill_1 FILLER_71_198 ();
 sg13g2_fill_2 FILLER_71_211 ();
 sg13g2_fill_1 FILLER_71_213 ();
 sg13g2_fill_1 FILLER_71_239 ();
 sg13g2_fill_2 FILLER_71_265 ();
 sg13g2_fill_1 FILLER_71_267 ();
 sg13g2_decap_4 FILLER_71_275 ();
 sg13g2_fill_2 FILLER_71_299 ();
 sg13g2_fill_1 FILLER_71_301 ();
 sg13g2_fill_2 FILLER_71_323 ();
 sg13g2_decap_4 FILLER_71_342 ();
 sg13g2_fill_1 FILLER_71_346 ();
 sg13g2_decap_4 FILLER_71_367 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_71_382 ();
 sg13g2_decap_8 FILLER_71_401 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_fill_2 FILLER_72_26 ();
 sg13g2_fill_1 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_59 ();
 sg13g2_fill_2 FILLER_72_87 ();
 sg13g2_fill_1 FILLER_72_104 ();
 sg13g2_fill_2 FILLER_72_148 ();
 sg13g2_fill_2 FILLER_72_157 ();
 sg13g2_fill_2 FILLER_72_199 ();
 sg13g2_fill_1 FILLER_72_210 ();
 sg13g2_fill_2 FILLER_72_226 ();
 sg13g2_decap_8 FILLER_72_233 ();
 sg13g2_fill_2 FILLER_72_240 ();
 sg13g2_decap_8 FILLER_72_275 ();
 sg13g2_fill_1 FILLER_72_282 ();
 sg13g2_fill_2 FILLER_72_308 ();
 sg13g2_fill_1 FILLER_72_351 ();
 sg13g2_fill_1 FILLER_72_360 ();
 sg13g2_fill_1 FILLER_72_374 ();
 sg13g2_fill_1 FILLER_72_387 ();
 sg13g2_decap_4 FILLER_72_405 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_9 ();
 sg13g2_fill_1 FILLER_73_11 ();
 sg13g2_fill_2 FILLER_73_28 ();
 sg13g2_fill_2 FILLER_73_55 ();
 sg13g2_fill_1 FILLER_73_57 ();
 sg13g2_fill_2 FILLER_73_82 ();
 sg13g2_fill_1 FILLER_73_84 ();
 sg13g2_fill_2 FILLER_73_99 ();
 sg13g2_fill_2 FILLER_73_132 ();
 sg13g2_fill_1 FILLER_73_134 ();
 sg13g2_decap_4 FILLER_73_211 ();
 sg13g2_decap_4 FILLER_73_240 ();
 sg13g2_fill_1 FILLER_73_244 ();
 sg13g2_decap_8 FILLER_73_264 ();
 sg13g2_decap_4 FILLER_73_271 ();
 sg13g2_fill_1 FILLER_73_275 ();
 sg13g2_fill_2 FILLER_73_281 ();
 sg13g2_decap_4 FILLER_73_296 ();
 sg13g2_fill_1 FILLER_73_300 ();
 sg13g2_fill_2 FILLER_73_310 ();
 sg13g2_fill_1 FILLER_73_312 ();
 sg13g2_fill_2 FILLER_73_326 ();
 sg13g2_fill_1 FILLER_73_346 ();
 sg13g2_fill_2 FILLER_73_386 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_118 ();
 sg13g2_fill_1 FILLER_74_189 ();
 sg13g2_decap_4 FILLER_74_209 ();
 sg13g2_fill_2 FILLER_74_213 ();
 sg13g2_fill_2 FILLER_74_223 ();
 sg13g2_fill_1 FILLER_74_225 ();
 sg13g2_decap_4 FILLER_74_252 ();
 sg13g2_fill_2 FILLER_74_273 ();
 sg13g2_fill_1 FILLER_74_275 ();
 sg13g2_decap_8 FILLER_74_291 ();
 sg13g2_decap_4 FILLER_74_298 ();
 sg13g2_fill_2 FILLER_74_328 ();
 sg13g2_fill_1 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_374 ();
 sg13g2_fill_1 FILLER_75_50 ();
 sg13g2_fill_1 FILLER_75_67 ();
 sg13g2_fill_2 FILLER_75_104 ();
 sg13g2_fill_2 FILLER_75_141 ();
 sg13g2_fill_2 FILLER_75_158 ();
 sg13g2_decap_4 FILLER_75_169 ();
 sg13g2_decap_8 FILLER_75_195 ();
 sg13g2_decap_4 FILLER_75_202 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_fill_2 FILLER_75_256 ();
 sg13g2_fill_2 FILLER_75_279 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_fill_2 FILLER_75_307 ();
 sg13g2_fill_1 FILLER_75_309 ();
 sg13g2_decap_8 FILLER_75_323 ();
 sg13g2_fill_1 FILLER_75_334 ();
 sg13g2_fill_2 FILLER_75_357 ();
 sg13g2_decap_4 FILLER_75_363 ();
 sg13g2_fill_2 FILLER_75_367 ();
 sg13g2_fill_1 FILLER_75_373 ();
 sg13g2_fill_2 FILLER_75_386 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_fill_1 FILLER_76_42 ();
 sg13g2_fill_2 FILLER_76_102 ();
 sg13g2_fill_2 FILLER_76_118 ();
 sg13g2_fill_1 FILLER_76_120 ();
 sg13g2_decap_4 FILLER_76_151 ();
 sg13g2_fill_1 FILLER_76_170 ();
 sg13g2_decap_8 FILLER_76_181 ();
 sg13g2_decap_4 FILLER_76_188 ();
 sg13g2_fill_1 FILLER_76_192 ();
 sg13g2_fill_2 FILLER_76_212 ();
 sg13g2_fill_1 FILLER_76_240 ();
 sg13g2_fill_2 FILLER_76_246 ();
 sg13g2_fill_2 FILLER_76_297 ();
 sg13g2_decap_8 FILLER_76_307 ();
 sg13g2_decap_8 FILLER_76_314 ();
 sg13g2_fill_1 FILLER_76_338 ();
 sg13g2_decap_4 FILLER_76_351 ();
 sg13g2_fill_1 FILLER_76_355 ();
 sg13g2_fill_2 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_7 ();
 sg13g2_fill_1 FILLER_77_117 ();
 sg13g2_fill_1 FILLER_77_171 ();
 sg13g2_fill_2 FILLER_77_177 ();
 sg13g2_fill_1 FILLER_77_179 ();
 sg13g2_fill_1 FILLER_77_184 ();
 sg13g2_fill_1 FILLER_77_189 ();
 sg13g2_fill_2 FILLER_77_212 ();
 sg13g2_fill_1 FILLER_77_214 ();
 sg13g2_fill_2 FILLER_77_246 ();
 sg13g2_fill_1 FILLER_77_256 ();
 sg13g2_fill_1 FILLER_77_264 ();
 sg13g2_fill_2 FILLER_77_356 ();
 sg13g2_fill_1 FILLER_77_358 ();
 sg13g2_decap_4 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_fill_2 FILLER_78_21 ();
 sg13g2_fill_2 FILLER_78_58 ();
 sg13g2_fill_1 FILLER_78_60 ();
 sg13g2_fill_2 FILLER_78_87 ();
 sg13g2_fill_2 FILLER_78_115 ();
 sg13g2_fill_1 FILLER_78_117 ();
 sg13g2_decap_4 FILLER_78_170 ();
 sg13g2_fill_2 FILLER_78_200 ();
 sg13g2_fill_1 FILLER_78_202 ();
 sg13g2_fill_1 FILLER_78_266 ();
 sg13g2_fill_1 FILLER_78_275 ();
 sg13g2_fill_2 FILLER_78_288 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_45 ();
 sg13g2_fill_2 FILLER_79_72 ();
 sg13g2_decap_4 FILLER_79_202 ();
 sg13g2_fill_2 FILLER_79_206 ();
 sg13g2_fill_2 FILLER_79_225 ();
 sg13g2_fill_1 FILLER_79_227 ();
 sg13g2_fill_1 FILLER_79_245 ();
 sg13g2_fill_2 FILLER_79_250 ();
 sg13g2_fill_2 FILLER_79_262 ();
 sg13g2_fill_2 FILLER_79_292 ();
 sg13g2_fill_1 FILLER_79_312 ();
 sg13g2_fill_2 FILLER_79_323 ();
 sg13g2_fill_1 FILLER_79_325 ();
 sg13g2_fill_2 FILLER_79_331 ();
 sg13g2_fill_1 FILLER_79_333 ();
 sg13g2_fill_2 FILLER_79_338 ();
 sg13g2_fill_2 FILLER_79_360 ();
 sg13g2_fill_1 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_decap_4 FILLER_79_405 ();
 sg13g2_decap_4 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_4 ();
 sg13g2_fill_1 FILLER_80_113 ();
 sg13g2_decap_8 FILLER_80_146 ();
 sg13g2_decap_4 FILLER_80_153 ();
 sg13g2_fill_1 FILLER_80_157 ();
 sg13g2_fill_2 FILLER_80_166 ();
 sg13g2_fill_1 FILLER_80_168 ();
 sg13g2_decap_8 FILLER_80_195 ();
 sg13g2_decap_8 FILLER_80_202 ();
 sg13g2_decap_8 FILLER_80_209 ();
 sg13g2_decap_8 FILLER_80_216 ();
 sg13g2_fill_2 FILLER_80_223 ();
 sg13g2_fill_1 FILLER_80_230 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_decap_8 FILLER_80_249 ();
 sg13g2_fill_2 FILLER_80_256 ();
 sg13g2_fill_1 FILLER_80_258 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_fill_2 FILLER_80_278 ();
 sg13g2_fill_1 FILLER_80_280 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_305 ();
 sg13g2_decap_4 FILLER_80_312 ();
 sg13g2_fill_2 FILLER_80_316 ();
 sg13g2_decap_8 FILLER_80_322 ();
 sg13g2_fill_1 FILLER_80_329 ();
 sg13g2_decap_8 FILLER_80_334 ();
 sg13g2_fill_1 FILLER_80_341 ();
 sg13g2_fill_2 FILLER_80_346 ();
 sg13g2_fill_1 FILLER_80_348 ();
 sg13g2_decap_8 FILLER_80_354 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_decap_8 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_389 ();
 sg13g2_decap_8 FILLER_80_396 ();
 sg13g2_decap_4 FILLER_80_403 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net138;
 assign uio_oe[1] = net139;
 assign uio_oe[2] = net140;
 assign uio_oe[3] = net141;
 assign uio_oe[4] = net142;
 assign uio_oe[5] = net143;
 assign uio_oe[6] = net144;
 assign uio_oe[7] = net145;
endmodule

module tt_um_resfuzzy (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire clknet_0_clk;
 wire \top.controller.count[0] ;
 wire \top.controller.count[1] ;
 wire \top.controller.ef1 ;
 wire \top.controller.r1[0] ;
 wire \top.controller.r1[1] ;
 wire \top.controller.r1[2] ;
 wire \top.controller.r1[3] ;
 wire \top.controller.r1[4] ;
 wire \top.controller.r1[5] ;
 wire \top.controller.r1[6] ;
 wire \top.controller.r1[7] ;
 wire \top.controller.r2[0] ;
 wire \top.controller.r2[1] ;
 wire \top.controller.r2[2] ;
 wire \top.controller.r2[3] ;
 wire \top.controller.r2[4] ;
 wire \top.controller.r2[5] ;
 wire \top.controller.r2[6] ;
 wire \top.controller.r2[7] ;
 wire \top.controller.s1[0] ;
 wire \top.controller.s1[1] ;
 wire \top.controller.s1[2] ;
 wire \top.controller.s1[3] ;
 wire \top.controller.s1[4] ;
 wire \top.controller.s1[5] ;
 wire \top.controller.s1[6] ;
 wire \top.controller.s1[7] ;
 wire \top.controller.s2[0] ;
 wire \top.controller.s2[1] ;
 wire \top.controller.s2[2] ;
 wire \top.controller.s2[3] ;
 wire \top.controller.s2[4] ;
 wire \top.controller.s2[5] ;
 wire \top.controller.s2[6] ;
 wire \top.controller.s2[7] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;

 sg13g2_inv_1 _1001_ (.Y(_0063_),
    .A(net8));
 sg13g2_inv_1 _1002_ (.Y(_0064_),
    .A(net7));
 sg13g2_inv_1 _1003_ (.Y(_0065_),
    .A(net6));
 sg13g2_inv_1 _1004_ (.Y(_0066_),
    .A(net5));
 sg13g2_inv_1 _1005_ (.Y(_0067_),
    .A(net4));
 sg13g2_inv_1 _1006_ (.Y(_0068_),
    .A(net3));
 sg13g2_inv_1 _1007_ (.Y(_0069_),
    .A(net2));
 sg13g2_inv_1 _1008_ (.Y(_0070_),
    .A(net1));
 sg13g2_inv_1 _1009_ (.Y(_0071_),
    .A(net76));
 sg13g2_inv_1 _1010_ (.Y(_0072_),
    .A(net79));
 sg13g2_inv_1 _1011_ (.Y(_0073_),
    .A(net72));
 sg13g2_inv_1 _1012_ (.Y(_0074_),
    .A(net73));
 sg13g2_inv_1 _1013_ (.Y(_0075_),
    .A(net85));
 sg13g2_inv_1 _1014_ (.Y(_0076_),
    .A(net88));
 sg13g2_inv_1 _1015_ (.Y(_0077_),
    .A(net107));
 sg13g2_inv_1 _1016_ (.Y(_0078_),
    .A(net92));
 sg13g2_inv_1 _1017_ (.Y(_0079_),
    .A(\top.controller.ef1 ));
 sg13g2_inv_1 _1018_ (.Y(_0080_),
    .A(net98));
 sg13g2_inv_1 _1019_ (.Y(_0081_),
    .A(net166));
 sg13g2_inv_2 _1020_ (.Y(_0082_),
    .A(net91));
 sg13g2_inv_1 _1021_ (.Y(_0083_),
    .A(net74));
 sg13g2_inv_1 _1022_ (.Y(_0084_),
    .A(_0000_));
 sg13g2_inv_1 _1023_ (.Y(_0085_),
    .A(net150));
 sg13g2_inv_1 _1024_ (.Y(_0086_),
    .A(net147));
 sg13g2_nand2_1 _1025_ (.Y(_0087_),
    .A(net70),
    .B(_0080_));
 sg13g2_and3_1 _1026_ (.X(_0012_),
    .A(net166),
    .B(net68),
    .C(_0087_));
 sg13g2_nor3_1 _1027_ (.A(net70),
    .B(_0080_),
    .C(net158),
    .Y(_0013_));
 sg13g2_nand2_1 _1028_ (.Y(_0088_),
    .A(net144),
    .B(net80));
 sg13g2_nor2_2 _1029_ (.A(\top.controller.s2[0] ),
    .B(\top.controller.s2[1] ),
    .Y(_0089_));
 sg13g2_or2_1 _1030_ (.X(_0090_),
    .B(\top.controller.s2[1] ),
    .A(\top.controller.s2[0] ));
 sg13g2_nor2_1 _1031_ (.A(net150),
    .B(net148),
    .Y(_0091_));
 sg13g2_or2_2 _1032_ (.X(_0092_),
    .B(net148),
    .A(\top.controller.s2[2] ));
 sg13g2_a21oi_1 _1033_ (.A1(_0089_),
    .A2(_0091_),
    .Y(_0093_),
    .B1(_0086_));
 sg13g2_o21ai_1 _1034_ (.B1(net145),
    .Y(_0094_),
    .A1(\top.controller.s2[5] ),
    .A2(_0093_));
 sg13g2_nand2b_2 _1035_ (.Y(_0095_),
    .B(_0094_),
    .A_N(\top.controller.s2[7] ));
 sg13g2_inv_1 _1036_ (.Y(_0096_),
    .A(_0095_));
 sg13g2_o21ai_1 _1037_ (.B1(net150),
    .Y(_0097_),
    .A1(\top.controller.s2[0] ),
    .A2(\top.controller.s2[1] ));
 sg13g2_inv_1 _1038_ (.Y(_0098_),
    .A(_0097_));
 sg13g2_nor2b_1 _1039_ (.A(net149),
    .B_N(_0097_),
    .Y(_0099_));
 sg13g2_nor2b_2 _1040_ (.A(\top.controller.s2[4] ),
    .B_N(net146),
    .Y(_0100_));
 sg13g2_nand3b_1 _1041_ (.B(_0097_),
    .C(_0100_),
    .Y(_0101_),
    .A_N(\top.controller.s2[3] ));
 sg13g2_nor2b_1 _1042_ (.A(_0006_),
    .B_N(net145),
    .Y(_0102_));
 sg13g2_a21o_2 _1043_ (.A2(_0102_),
    .A1(_0101_),
    .B1(\top.controller.s2[7] ),
    .X(_0103_));
 sg13g2_nor2_1 _1044_ (.A(\top.controller.s2[7] ),
    .B(net145),
    .Y(_0104_));
 sg13g2_and2_1 _1045_ (.A(\top.controller.s2[5] ),
    .B(net147),
    .X(_0105_));
 sg13g2_and2_1 _1046_ (.A(\top.controller.s2[0] ),
    .B(\top.controller.s2[1] ),
    .X(_0106_));
 sg13g2_o21ai_1 _1047_ (.B1(_0105_),
    .Y(_0107_),
    .A1(_0092_),
    .A2(_0106_));
 sg13g2_and2_1 _1048_ (.A(net143),
    .B(_0107_),
    .X(_0108_));
 sg13g2_nand2_2 _1049_ (.Y(_0109_),
    .A(net143),
    .B(_0107_));
 sg13g2_or3_1 _1050_ (.A(net149),
    .B(\top.controller.s2[5] ),
    .C(\top.controller.s2[4] ),
    .X(_0110_));
 sg13g2_and2_2 _1051_ (.A(net150),
    .B(\top.controller.s2[1] ),
    .X(_0111_));
 sg13g2_nand3_1 _1052_ (.B(\top.controller.s2[0] ),
    .C(\top.controller.s2[1] ),
    .A(net150),
    .Y(_0112_));
 sg13g2_nor4_1 _1053_ (.A(net149),
    .B(net146),
    .C(net147),
    .D(\top.controller.s2[7] ),
    .Y(_0113_));
 sg13g2_a21oi_2 _1054_ (.B1(net143),
    .Y(_0114_),
    .A2(_0113_),
    .A1(_0112_));
 sg13g2_a21oi_2 _1055_ (.B1(_0114_),
    .Y(_0115_),
    .A2(_0107_),
    .A1(net143));
 sg13g2_nand2_1 _1056_ (.Y(_0116_),
    .A(net149),
    .B(net147));
 sg13g2_xnor2_1 _1057_ (.Y(_0117_),
    .A(net148),
    .B(net147));
 sg13g2_or2_2 _1058_ (.X(_0118_),
    .B(_0103_),
    .A(_0094_));
 sg13g2_nor2_1 _1059_ (.A(net148),
    .B(_0111_),
    .Y(_0119_));
 sg13g2_xnor2_1 _1060_ (.Y(_0120_),
    .A(_0008_),
    .B(_0119_));
 sg13g2_mux2_1 _1061_ (.A0(_0117_),
    .A1(_0120_),
    .S(_0115_),
    .X(_0121_));
 sg13g2_nor3_2 _1062_ (.A(net147),
    .B(_0090_),
    .C(_0092_),
    .Y(_0122_));
 sg13g2_nor3_2 _1063_ (.A(net146),
    .B(\top.controller.s2[7] ),
    .C(\top.controller.s2[6] ),
    .Y(_0123_));
 sg13g2_o21ai_1 _1064_ (.B1(_0123_),
    .Y(_0124_),
    .A1(_0086_),
    .A2(_0099_));
 sg13g2_nor2_1 _1065_ (.A(_0122_),
    .B(_0124_),
    .Y(_0125_));
 sg13g2_inv_1 _1066_ (.Y(_0126_),
    .A(_0125_));
 sg13g2_xnor2_1 _1067_ (.Y(_0127_),
    .A(_0008_),
    .B(_0092_));
 sg13g2_nor3_1 _1068_ (.A(_0094_),
    .B(_0103_),
    .C(_0127_),
    .Y(_0128_));
 sg13g2_a21oi_1 _1069_ (.A1(_0118_),
    .A2(_0121_),
    .Y(_0129_),
    .B1(_0128_));
 sg13g2_o21ai_1 _1070_ (.B1(_0129_),
    .Y(_0130_),
    .A1(_0093_),
    .A2(_0126_));
 sg13g2_nor3_1 _1071_ (.A(net149),
    .B(net147),
    .C(_0111_),
    .Y(_0131_));
 sg13g2_nor2_1 _1072_ (.A(_0110_),
    .B(_0111_),
    .Y(_0132_));
 sg13g2_xor2_1 _1073_ (.B(_0132_),
    .A(_0007_),
    .X(_0133_));
 sg13g2_o21ai_1 _1074_ (.B1(net146),
    .Y(_0134_),
    .A1(net148),
    .A2(\top.controller.s2[4] ));
 sg13g2_nand2b_1 _1075_ (.Y(_0135_),
    .B(_0134_),
    .A_N(net145));
 sg13g2_xor2_1 _1076_ (.B(_0134_),
    .A(net145),
    .X(_0136_));
 sg13g2_a21oi_1 _1077_ (.A1(_0115_),
    .A2(_0133_),
    .Y(_0137_),
    .B1(_0136_));
 sg13g2_and2_1 _1078_ (.A(_0092_),
    .B(_0100_),
    .X(_0138_));
 sg13g2_nand2_1 _1079_ (.Y(_0139_),
    .A(_0092_),
    .B(_0100_));
 sg13g2_nor3_1 _1080_ (.A(_0094_),
    .B(_0103_),
    .C(_0138_),
    .Y(_0140_));
 sg13g2_mux2_2 _1081_ (.A0(_0118_),
    .A1(_0140_),
    .S(_0137_),
    .X(_0141_));
 sg13g2_and2_1 _1082_ (.A(\top.controller.s2[7] ),
    .B(_0135_),
    .X(_0142_));
 sg13g2_nand2_1 _1083_ (.Y(_0143_),
    .A(_0104_),
    .B(_0134_));
 sg13g2_o21ai_1 _1084_ (.B1(net145),
    .Y(_0144_),
    .A1(_0110_),
    .A2(_0111_));
 sg13g2_xnor2_1 _1085_ (.Y(_0145_),
    .A(_0005_),
    .B(_0144_));
 sg13g2_a221oi_1 _1086_ (.B2(_0115_),
    .C1(_0142_),
    .B1(_0145_),
    .A1(net143),
    .Y(_0146_),
    .A2(_0134_));
 sg13g2_o21ai_1 _1087_ (.B1(net145),
    .Y(_0147_),
    .A1(_0105_),
    .A2(_0138_));
 sg13g2_xor2_1 _1088_ (.B(_0147_),
    .A(_0005_),
    .X(_0148_));
 sg13g2_o21ai_1 _1089_ (.B1(_0146_),
    .Y(_0149_),
    .A1(_0118_),
    .A2(_0148_));
 sg13g2_nor3_1 _1090_ (.A(_0094_),
    .B(_0103_),
    .C(_0139_),
    .Y(_0150_));
 sg13g2_xnor2_1 _1091_ (.Y(_0151_),
    .A(_0006_),
    .B(_0131_));
 sg13g2_a22oi_1 _1092_ (.Y(_0152_),
    .B1(_0151_),
    .B2(_0115_),
    .A2(_0134_),
    .A1(_0110_));
 sg13g2_or2_1 _1093_ (.X(_0153_),
    .B(_0152_),
    .A(_0150_));
 sg13g2_and4_1 _1094_ (.A(_0126_),
    .B(_0141_),
    .C(_0149_),
    .D(_0153_),
    .X(_0154_));
 sg13g2_nand4_1 _1095_ (.B(_0141_),
    .C(_0149_),
    .A(_0126_),
    .Y(_0155_),
    .D(_0153_));
 sg13g2_nor3_1 _1096_ (.A(_0146_),
    .B(_0150_),
    .C(_0152_),
    .Y(_0156_));
 sg13g2_a21oi_2 _1097_ (.B1(_0156_),
    .Y(_0157_),
    .A2(_0149_),
    .A1(_0141_));
 sg13g2_a221oi_1 _1098_ (.B2(_0126_),
    .C1(_0156_),
    .B1(_0153_),
    .A1(_0141_),
    .Y(_0158_),
    .A2(_0149_));
 sg13g2_or2_1 _1099_ (.X(_0159_),
    .B(_0158_),
    .A(_0154_));
 sg13g2_or3_1 _1100_ (.A(_0130_),
    .B(_0154_),
    .C(_0158_),
    .X(_0160_));
 sg13g2_and2_1 _1101_ (.A(_0149_),
    .B(_0157_),
    .X(_0161_));
 sg13g2_mux2_1 _1102_ (.A0(_0141_),
    .A1(_0161_),
    .S(_0160_),
    .X(_0162_));
 sg13g2_and2_1 _1103_ (.A(_0141_),
    .B(_0155_),
    .X(_0163_));
 sg13g2_a21oi_2 _1104_ (.B1(_0161_),
    .Y(_0164_),
    .A2(_0163_),
    .A1(_0160_));
 sg13g2_xor2_1 _1105_ (.B(_0164_),
    .A(_0130_),
    .X(_0165_));
 sg13g2_or2_1 _1106_ (.X(_0166_),
    .B(_0118_),
    .A(_0085_));
 sg13g2_nand2_1 _1107_ (.Y(_0167_),
    .A(_0111_),
    .B(_0115_));
 sg13g2_nand3_1 _1108_ (.B(_0089_),
    .C(_0125_),
    .A(_0009_),
    .Y(_0168_));
 sg13g2_nand3_1 _1109_ (.B(_0167_),
    .C(_0168_),
    .A(_0166_),
    .Y(_0169_));
 sg13g2_xor2_1 _1110_ (.B(_0169_),
    .A(net148),
    .X(_0170_));
 sg13g2_nand2b_1 _1111_ (.Y(_0171_),
    .B(_0161_),
    .A_N(_0160_));
 sg13g2_o21ai_1 _1112_ (.B1(_0159_),
    .Y(_0172_),
    .A1(_0130_),
    .A2(_0164_));
 sg13g2_a22oi_1 _1113_ (.Y(_0173_),
    .B1(_0171_),
    .B2(_0172_),
    .A2(_0170_),
    .A1(_0165_));
 sg13g2_nor2_2 _1114_ (.A(_0162_),
    .B(_0173_),
    .Y(_0174_));
 sg13g2_nor2_1 _1115_ (.A(net150),
    .B(\top.controller.s2[1] ),
    .Y(_0175_));
 sg13g2_nor4_1 _1116_ (.A(_0108_),
    .B(_0111_),
    .C(_0114_),
    .D(_0175_),
    .Y(_0176_));
 sg13g2_o21ai_1 _1117_ (.B1(_0118_),
    .Y(_0177_),
    .A1(_0009_),
    .A2(_0115_));
 sg13g2_o21ai_1 _1118_ (.B1(_0166_),
    .Y(_0178_),
    .A1(_0176_),
    .A2(_0177_));
 sg13g2_nor2_1 _1119_ (.A(_0089_),
    .B(_0124_),
    .Y(_0179_));
 sg13g2_xor2_1 _1120_ (.B(_0179_),
    .A(_0178_),
    .X(_0180_));
 sg13g2_or2_1 _1121_ (.X(_0181_),
    .B(_0180_),
    .A(_0170_));
 sg13g2_o21ai_1 _1122_ (.B1(_0181_),
    .Y(_0182_),
    .A1(_0162_),
    .A2(_0173_));
 sg13g2_a21oi_1 _1123_ (.A1(_0170_),
    .A2(_0180_),
    .Y(_0183_),
    .B1(_0165_));
 sg13g2_nand3_1 _1124_ (.B(_0165_),
    .C(_0170_),
    .A(_0159_),
    .Y(_0184_));
 sg13g2_nand2b_1 _1125_ (.Y(_0185_),
    .B(_0184_),
    .A_N(_0162_));
 sg13g2_a21oi_2 _1126_ (.B1(_0185_),
    .Y(_0186_),
    .A2(_0183_),
    .A1(_0182_));
 sg13g2_a21o_1 _1127_ (.A2(_0183_),
    .A1(_0182_),
    .B1(_0185_),
    .X(_0187_));
 sg13g2_o21ai_1 _1128_ (.B1(_0095_),
    .Y(_0188_),
    .A1(_0103_),
    .A2(_0186_));
 sg13g2_nor2_2 _1129_ (.A(\top.controller.s1[6] ),
    .B(\top.controller.s1[7] ),
    .Y(_0189_));
 sg13g2_or2_2 _1130_ (.X(_0190_),
    .B(\top.controller.s1[7] ),
    .A(\top.controller.s1[6] ));
 sg13g2_nor2_2 _1131_ (.A(\top.controller.s1[0] ),
    .B(\top.controller.s1[1] ),
    .Y(_0191_));
 sg13g2_nor2_1 _1132_ (.A(net154),
    .B(net156),
    .Y(_0192_));
 sg13g2_or4_1 _1133_ (.A(net154),
    .B(net155),
    .C(\top.controller.s1[0] ),
    .D(net157),
    .X(_0193_));
 sg13g2_nand2_1 _1134_ (.Y(_0194_),
    .A(net152),
    .B(_0193_));
 sg13g2_nor2_1 _1135_ (.A(net151),
    .B(\top.controller.s1[7] ),
    .Y(_0195_));
 sg13g2_or2_1 _1136_ (.X(_0196_),
    .B(\top.controller.s1[7] ),
    .A(net151));
 sg13g2_a21oi_2 _1137_ (.B1(_0196_),
    .Y(_0197_),
    .A2(_0193_),
    .A1(net153));
 sg13g2_nor2_2 _1138_ (.A(_0189_),
    .B(_0197_),
    .Y(_0198_));
 sg13g2_o21ai_1 _1139_ (.B1(net156),
    .Y(_0199_),
    .A1(\top.controller.s1[0] ),
    .A2(net157));
 sg13g2_nand2_1 _1140_ (.Y(_0200_),
    .A(_0082_),
    .B(_0199_));
 sg13g2_nor2b_1 _1141_ (.A(\top.controller.s1[7] ),
    .B_N(\top.controller.s1[6] ),
    .Y(_0201_));
 sg13g2_nor2b_1 _1142_ (.A(net153),
    .B_N(net151),
    .Y(_0202_));
 sg13g2_nand4_1 _1143_ (.B(_0199_),
    .C(_0201_),
    .A(_0082_),
    .Y(_0203_),
    .D(_0202_));
 sg13g2_a21o_1 _1144_ (.A2(_0084_),
    .A1(\top.controller.s1[6] ),
    .B1(\top.controller.s1[7] ),
    .X(_0204_));
 sg13g2_and2_2 _1145_ (.A(_0203_),
    .B(_0204_),
    .X(_0205_));
 sg13g2_nand2_1 _1146_ (.Y(_0206_),
    .A(_0083_),
    .B(_0189_));
 sg13g2_a21oi_2 _1147_ (.B1(_0206_),
    .Y(_0207_),
    .A2(_0200_),
    .A1(net153));
 sg13g2_nor2_2 _1148_ (.A(net154),
    .B(net152),
    .Y(_0208_));
 sg13g2_or2_1 _1149_ (.X(_0209_),
    .B(net152),
    .A(net154));
 sg13g2_nand2b_1 _1150_ (.Y(_0210_),
    .B(_0191_),
    .A_N(net155));
 sg13g2_o21ai_1 _1151_ (.B1(_0207_),
    .Y(_0211_),
    .A1(_0209_),
    .A2(_0210_));
 sg13g2_a221oi_1 _1152_ (.B2(_0204_),
    .C1(_0189_),
    .B1(_0203_),
    .A1(_0194_),
    .Y(_0212_),
    .A2(_0195_));
 sg13g2_o21ai_1 _1153_ (.B1(net151),
    .Y(_0213_),
    .A1(net155),
    .A2(_0209_));
 sg13g2_nand2_1 _1154_ (.Y(_0214_),
    .A(_0212_),
    .B(_0213_));
 sg13g2_nor2b_1 _1155_ (.A(net152),
    .B_N(net154),
    .Y(_0215_));
 sg13g2_o21ai_1 _1156_ (.B1(_0189_),
    .Y(_0216_),
    .A1(_0083_),
    .A2(_0208_));
 sg13g2_nand2_1 _1157_ (.Y(_0217_),
    .A(_0189_),
    .B(_0215_));
 sg13g2_o21ai_1 _1158_ (.B1(_0216_),
    .Y(_0218_),
    .A1(_0210_),
    .A2(_0217_));
 sg13g2_nor2b_2 _1159_ (.A(_0207_),
    .B_N(_0218_),
    .Y(_0219_));
 sg13g2_nand3_1 _1160_ (.B(_0215_),
    .C(_0218_),
    .A(net151),
    .Y(_0220_));
 sg13g2_nand2b_1 _1161_ (.Y(_0221_),
    .B(net156),
    .A_N(_0001_));
 sg13g2_nand2_1 _1162_ (.Y(_0222_),
    .A(_0208_),
    .B(_0221_));
 sg13g2_nor2_1 _1163_ (.A(net151),
    .B(_0222_),
    .Y(_0223_));
 sg13g2_xnor2_1 _1164_ (.Y(_0224_),
    .A(_0002_),
    .B(_0223_));
 sg13g2_xnor2_1 _1165_ (.Y(_0225_),
    .A(_0214_),
    .B(_0224_));
 sg13g2_xnor2_1 _1166_ (.Y(_0226_),
    .A(_0220_),
    .B(_0225_));
 sg13g2_nand2_1 _1167_ (.Y(_0227_),
    .A(_0211_),
    .B(_0226_));
 sg13g2_nand2b_1 _1168_ (.Y(_0228_),
    .B(_0207_),
    .A_N(_0194_));
 sg13g2_nand2_1 _1169_ (.Y(_0229_),
    .A(_0082_),
    .B(_0221_));
 sg13g2_a21oi_1 _1170_ (.A1(net155),
    .A2(_0212_),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_xor2_1 _1171_ (.B(_0230_),
    .A(_0003_),
    .X(_0231_));
 sg13g2_nor2_1 _1172_ (.A(_0219_),
    .B(_0231_),
    .Y(_0232_));
 sg13g2_and2_1 _1173_ (.A(net154),
    .B(net152),
    .X(_0233_));
 sg13g2_o21ai_1 _1174_ (.B1(_0219_),
    .Y(_0234_),
    .A1(_0208_),
    .A2(_0233_));
 sg13g2_nand2_1 _1175_ (.Y(_0235_),
    .A(_0211_),
    .B(_0234_));
 sg13g2_o21ai_1 _1176_ (.B1(_0228_),
    .Y(_0236_),
    .A1(_0232_),
    .A2(_0235_));
 sg13g2_xnor2_1 _1177_ (.Y(_0237_),
    .A(_0084_),
    .B(_0222_));
 sg13g2_mux2_1 _1178_ (.A0(_0237_),
    .A1(_0213_),
    .S(_0212_),
    .X(_0238_));
 sg13g2_o21ai_1 _1179_ (.B1(_0220_),
    .Y(_0239_),
    .A1(_0219_),
    .A2(_0238_));
 sg13g2_nand2_1 _1180_ (.Y(_0240_),
    .A(_0211_),
    .B(_0239_));
 sg13g2_o21ai_1 _1181_ (.B1(\top.controller.s1[6] ),
    .Y(_0241_),
    .A1(net151),
    .A2(_0222_));
 sg13g2_xnor2_1 _1182_ (.Y(_0242_),
    .A(_0010_),
    .B(_0241_));
 sg13g2_xnor2_1 _1183_ (.Y(_0243_),
    .A(_0214_),
    .B(_0242_));
 sg13g2_o21ai_1 _1184_ (.B1(_0220_),
    .Y(_0244_),
    .A1(_0219_),
    .A2(_0243_));
 sg13g2_nand2b_1 _1185_ (.Y(_0245_),
    .B(_0226_),
    .A_N(_0240_));
 sg13g2_nand2b_2 _1186_ (.Y(_0246_),
    .B(_0245_),
    .A_N(_0244_));
 sg13g2_nor3_1 _1187_ (.A(_0226_),
    .B(_0240_),
    .C(_0244_),
    .Y(_0247_));
 sg13g2_or3_1 _1188_ (.A(_0226_),
    .B(_0240_),
    .C(_0244_),
    .X(_0248_));
 sg13g2_nand2_1 _1189_ (.Y(_0249_),
    .A(_0240_),
    .B(_0244_));
 sg13g2_nand2_1 _1190_ (.Y(_0250_),
    .A(_0248_),
    .B(_0249_));
 sg13g2_nand3_1 _1191_ (.B(_0248_),
    .C(_0249_),
    .A(_0236_),
    .Y(_0251_));
 sg13g2_nor2_2 _1192_ (.A(_0244_),
    .B(_0245_),
    .Y(_0252_));
 sg13g2_mux2_1 _1193_ (.A0(_0227_),
    .A1(_0252_),
    .S(_0251_),
    .X(_0253_));
 sg13g2_a221oi_1 _1194_ (.B2(_0249_),
    .C1(_0247_),
    .B1(_0236_),
    .A1(_0211_),
    .Y(_0254_),
    .A2(_0226_));
 sg13g2_nor2_2 _1195_ (.A(_0252_),
    .B(_0254_),
    .Y(_0255_));
 sg13g2_o21ai_1 _1196_ (.B1(_0236_),
    .Y(_0256_),
    .A1(_0252_),
    .A2(_0254_));
 sg13g2_or3_1 _1197_ (.A(_0236_),
    .B(_0252_),
    .C(_0254_),
    .X(_0257_));
 sg13g2_nand2_1 _1198_ (.Y(_0258_),
    .A(_0256_),
    .B(_0257_));
 sg13g2_o21ai_1 _1199_ (.B1(net155),
    .Y(_0259_),
    .A1(net157),
    .A2(_0212_));
 sg13g2_a21oi_1 _1200_ (.A1(_0004_),
    .A2(_0191_),
    .Y(_0260_),
    .B1(_0211_));
 sg13g2_a21oi_1 _1201_ (.A1(_0211_),
    .A2(_0259_),
    .Y(_0261_),
    .B1(_0219_));
 sg13g2_nor2b_1 _1202_ (.A(_0260_),
    .B_N(_0261_),
    .Y(_0262_));
 sg13g2_xnor2_1 _1203_ (.Y(_0263_),
    .A(net154),
    .B(_0262_));
 sg13g2_nand3b_1 _1204_ (.B(_0257_),
    .C(_0256_),
    .Y(_0264_),
    .A_N(_0263_));
 sg13g2_xnor2_1 _1205_ (.Y(_0265_),
    .A(_0250_),
    .B(_0256_));
 sg13g2_a21oi_2 _1206_ (.B1(_0253_),
    .Y(_0266_),
    .A2(_0265_),
    .A1(_0264_));
 sg13g2_a21o_1 _1207_ (.A2(_0265_),
    .A1(_0264_),
    .B1(_0253_),
    .X(_0267_));
 sg13g2_nand2_1 _1208_ (.Y(_0268_),
    .A(_0199_),
    .B(_0210_));
 sg13g2_or3_1 _1209_ (.A(net155),
    .B(net157),
    .C(_0212_),
    .X(_0269_));
 sg13g2_and2_1 _1210_ (.A(_0259_),
    .B(_0269_),
    .X(_0270_));
 sg13g2_o21ai_1 _1211_ (.B1(_0211_),
    .Y(_0271_),
    .A1(_0219_),
    .A2(_0270_));
 sg13g2_a21o_1 _1212_ (.A2(_0219_),
    .A1(_0004_),
    .B1(_0271_),
    .X(_0272_));
 sg13g2_o21ai_1 _1213_ (.B1(_0272_),
    .Y(_0273_),
    .A1(_0211_),
    .A2(_0268_));
 sg13g2_nand2_1 _1214_ (.Y(_0274_),
    .A(_0263_),
    .B(_0273_));
 sg13g2_o21ai_1 _1215_ (.B1(_0258_),
    .Y(_0275_),
    .A1(_0263_),
    .A2(_0273_));
 sg13g2_a21oi_2 _1216_ (.B1(_0275_),
    .Y(_0276_),
    .A2(_0274_),
    .A1(_0267_));
 sg13g2_a21o_1 _1217_ (.A2(_0274_),
    .A1(_0267_),
    .B1(_0275_),
    .X(_0277_));
 sg13g2_nand2b_1 _1218_ (.Y(_0278_),
    .B(_0250_),
    .A_N(_0264_));
 sg13g2_nor2b_1 _1219_ (.A(_0253_),
    .B_N(_0278_),
    .Y(_0279_));
 sg13g2_nand2b_1 _1220_ (.Y(_0280_),
    .B(_0278_),
    .A_N(_0253_));
 sg13g2_nor2_1 _1221_ (.A(_0276_),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_o21ai_1 _1222_ (.B1(_0198_),
    .Y(_0282_),
    .A1(_0205_),
    .A2(_0281_));
 sg13g2_or2_1 _1223_ (.X(_0283_),
    .B(_0199_),
    .A(_0082_));
 sg13g2_nand2_1 _1224_ (.Y(_0284_),
    .A(net152),
    .B(\top.controller.s1[5] ));
 sg13g2_nor3_2 _1225_ (.A(_0082_),
    .B(_0199_),
    .C(_0284_),
    .Y(_0285_));
 sg13g2_mux2_2 _1226_ (.A0(_0197_),
    .A1(_0285_),
    .S(_0189_),
    .X(_0286_));
 sg13g2_inv_1 _1227_ (.Y(_0287_),
    .A(_0286_));
 sg13g2_and3_1 _1228_ (.X(_0288_),
    .A(_0200_),
    .B(_0283_),
    .C(_0286_));
 sg13g2_nand2_2 _1229_ (.Y(_0289_),
    .A(\top.controller.s1[0] ),
    .B(net157));
 sg13g2_nor2_1 _1230_ (.A(_0004_),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_xnor2_1 _1231_ (.Y(_0291_),
    .A(_0082_),
    .B(_0290_));
 sg13g2_a21oi_1 _1232_ (.A1(_0287_),
    .A2(_0291_),
    .Y(_0292_),
    .B1(_0288_));
 sg13g2_inv_1 _1233_ (.Y(_0293_),
    .A(_0292_));
 sg13g2_nand3_1 _1234_ (.B(\top.controller.s1[0] ),
    .C(net157),
    .A(net155),
    .Y(_0294_));
 sg13g2_xor2_1 _1235_ (.B(_0289_),
    .A(net155),
    .X(_0295_));
 sg13g2_nor2_1 _1236_ (.A(_0286_),
    .B(_0295_),
    .Y(_0296_));
 sg13g2_xor2_1 _1237_ (.B(_0191_),
    .A(_0004_),
    .X(_0297_));
 sg13g2_a21oi_1 _1238_ (.A1(_0286_),
    .A2(_0297_),
    .Y(_0298_),
    .B1(_0296_));
 sg13g2_nand2_1 _1239_ (.Y(_0299_),
    .A(_0292_),
    .B(_0298_));
 sg13g2_nor2_1 _1240_ (.A(net153),
    .B(net151),
    .Y(_0300_));
 sg13g2_nand4_1 _1241_ (.B(net156),
    .C(\top.controller.s1[0] ),
    .A(net154),
    .Y(_0301_),
    .D(net157));
 sg13g2_a21o_1 _1242_ (.A2(_0301_),
    .A1(_0083_),
    .B1(_0300_),
    .X(_0302_));
 sg13g2_nand2_1 _1243_ (.Y(_0303_),
    .A(_0002_),
    .B(_0302_));
 sg13g2_xor2_1 _1244_ (.B(_0302_),
    .A(_0002_),
    .X(_0304_));
 sg13g2_inv_1 _1245_ (.Y(_0305_),
    .A(_0304_));
 sg13g2_nor3_1 _1246_ (.A(_0082_),
    .B(_0003_),
    .C(_0199_),
    .Y(_0306_));
 sg13g2_xnor2_1 _1247_ (.Y(_0307_),
    .A(\top.controller.s1[5] ),
    .B(_0306_));
 sg13g2_nor2_1 _1248_ (.A(_0003_),
    .B(_0301_),
    .Y(_0308_));
 sg13g2_xnor2_1 _1249_ (.Y(_0309_),
    .A(_0000_),
    .B(_0308_));
 sg13g2_mux2_2 _1250_ (.A0(_0309_),
    .A1(_0307_),
    .S(_0286_),
    .X(_0310_));
 sg13g2_nor2_1 _1251_ (.A(_0304_),
    .B(_0310_),
    .Y(_0311_));
 sg13g2_xor2_1 _1252_ (.B(_0303_),
    .A(_0010_),
    .X(_0312_));
 sg13g2_nor3_1 _1253_ (.A(_0304_),
    .B(_0310_),
    .C(_0312_),
    .Y(_0313_));
 sg13g2_nor2_1 _1254_ (.A(_0311_),
    .B(_0312_),
    .Y(_0314_));
 sg13g2_nor3_1 _1255_ (.A(_0305_),
    .B(_0310_),
    .C(_0312_),
    .Y(_0315_));
 sg13g2_o21ai_1 _1256_ (.B1(_0304_),
    .Y(_0316_),
    .A1(_0310_),
    .A2(_0312_));
 sg13g2_nand2b_1 _1257_ (.Y(_0317_),
    .B(_0316_),
    .A_N(_0313_));
 sg13g2_mux2_1 _1258_ (.A0(_0301_),
    .A1(_0283_),
    .S(_0286_),
    .X(_0318_));
 sg13g2_xor2_1 _1259_ (.B(_0318_),
    .A(net152),
    .X(_0319_));
 sg13g2_xnor2_1 _1260_ (.Y(_0320_),
    .A(net152),
    .B(_0318_));
 sg13g2_nand2_1 _1261_ (.Y(_0321_),
    .A(_0316_),
    .B(_0319_));
 sg13g2_nand2_1 _1262_ (.Y(_0322_),
    .A(_0310_),
    .B(_0312_));
 sg13g2_nand3b_1 _1263_ (.B(_0320_),
    .C(_0322_),
    .Y(_0323_),
    .A_N(_0313_));
 sg13g2_nand2_1 _1264_ (.Y(_0324_),
    .A(_0321_),
    .B(_0323_));
 sg13g2_nand2_2 _1265_ (.Y(_0325_),
    .A(_0317_),
    .B(_0323_));
 sg13g2_and2_1 _1266_ (.A(_0317_),
    .B(_0324_),
    .X(_0326_));
 sg13g2_mux2_1 _1267_ (.A0(_0317_),
    .A1(_0325_),
    .S(_0320_),
    .X(_0327_));
 sg13g2_nand2_1 _1268_ (.Y(_0328_),
    .A(_0313_),
    .B(_0320_));
 sg13g2_nor2b_1 _1269_ (.A(_0315_),
    .B_N(_0322_),
    .Y(_0329_));
 sg13g2_inv_1 _1270_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_o21ai_1 _1271_ (.B1(_0330_),
    .Y(_0331_),
    .A1(_0319_),
    .A2(_0325_));
 sg13g2_a22oi_1 _1272_ (.Y(_0332_),
    .B1(_0328_),
    .B2(_0331_),
    .A2(_0327_),
    .A1(_0293_));
 sg13g2_nor2_1 _1273_ (.A(_0326_),
    .B(_0332_),
    .Y(_0333_));
 sg13g2_o21ai_1 _1274_ (.B1(_0299_),
    .Y(_0334_),
    .A1(_0326_),
    .A2(_0332_));
 sg13g2_nor2_1 _1275_ (.A(_0292_),
    .B(_0298_),
    .Y(_0335_));
 sg13g2_nor2_1 _1276_ (.A(_0327_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_nand3_1 _1277_ (.B(_0327_),
    .C(_0330_),
    .A(_0293_),
    .Y(_0337_));
 sg13g2_nand2b_1 _1278_ (.Y(_0338_),
    .B(_0337_),
    .A_N(_0326_));
 sg13g2_a21oi_2 _1279_ (.B1(_0338_),
    .Y(_0339_),
    .A2(_0336_),
    .A1(_0334_));
 sg13g2_nand2b_1 _1280_ (.Y(_0340_),
    .B(_0339_),
    .A_N(_0198_));
 sg13g2_nor2_1 _1281_ (.A(_0097_),
    .B(_0116_),
    .Y(_0341_));
 sg13g2_nand2_1 _1282_ (.Y(_0342_),
    .A(net146),
    .B(_0341_));
 sg13g2_nand2_1 _1283_ (.Y(_0343_),
    .A(net143),
    .B(_0342_));
 sg13g2_o21ai_1 _1284_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0190_),
    .A2(_0285_));
 sg13g2_o21ai_1 _1285_ (.B1(_0123_),
    .Y(_0345_),
    .A1(_0112_),
    .A2(_0116_));
 sg13g2_nand3_1 _1286_ (.B(_0107_),
    .C(_0345_),
    .A(net143),
    .Y(_0346_));
 sg13g2_nor2_1 _1287_ (.A(_0106_),
    .B(_0346_),
    .Y(_0347_));
 sg13g2_nor2_1 _1288_ (.A(_0089_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_nor3_1 _1289_ (.A(_0009_),
    .B(_0089_),
    .C(_0347_),
    .Y(_0349_));
 sg13g2_xnor2_1 _1290_ (.Y(_0350_),
    .A(net148),
    .B(_0349_));
 sg13g2_xnor2_1 _1291_ (.Y(_0351_),
    .A(net150),
    .B(_0348_));
 sg13g2_nand2_1 _1292_ (.Y(_0352_),
    .A(_0350_),
    .B(_0351_));
 sg13g2_nand3_1 _1293_ (.B(_0342_),
    .C(_0346_),
    .A(_0007_),
    .Y(_0353_));
 sg13g2_a21o_1 _1294_ (.A2(_0346_),
    .A1(_0342_),
    .B1(_0007_),
    .X(_0354_));
 sg13g2_nand2_1 _1295_ (.Y(_0355_),
    .A(_0353_),
    .B(_0354_));
 sg13g2_nand2b_1 _1296_ (.Y(_0356_),
    .B(\top.controller.s2[3] ),
    .A_N(_0008_));
 sg13g2_nor2_1 _1297_ (.A(_0097_),
    .B(_0356_),
    .Y(_0357_));
 sg13g2_xor2_1 _1298_ (.B(_0357_),
    .A(net146),
    .X(_0358_));
 sg13g2_xnor2_1 _1299_ (.Y(_0359_),
    .A(net146),
    .B(_0357_));
 sg13g2_nor2_1 _1300_ (.A(_0112_),
    .B(_0356_),
    .Y(_0360_));
 sg13g2_xor2_1 _1301_ (.B(_0360_),
    .A(_0006_),
    .X(_0361_));
 sg13g2_xnor2_1 _1302_ (.Y(_0362_),
    .A(_0006_),
    .B(_0360_));
 sg13g2_mux2_1 _1303_ (.A0(_0361_),
    .A1(_0358_),
    .S(_0346_),
    .X(_0363_));
 sg13g2_mux2_1 _1304_ (.A0(_0362_),
    .A1(_0359_),
    .S(_0346_),
    .X(_0364_));
 sg13g2_a21oi_1 _1305_ (.A1(_0353_),
    .A2(_0354_),
    .Y(_0365_),
    .B1(_0364_));
 sg13g2_xnor2_1 _1306_ (.Y(_0366_),
    .A(_0005_),
    .B(_0353_));
 sg13g2_xor2_1 _1307_ (.B(_0353_),
    .A(_0005_),
    .X(_0367_));
 sg13g2_nor2_1 _1308_ (.A(_0365_),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_and4_1 _1309_ (.A(_0005_),
    .B(_0353_),
    .C(_0354_),
    .D(_0363_),
    .X(_0369_));
 sg13g2_nor2_2 _1310_ (.A(_0355_),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_and2_1 _1311_ (.A(_0365_),
    .B(_0366_),
    .X(_0371_));
 sg13g2_inv_1 _1312_ (.Y(_0372_),
    .A(_0371_));
 sg13g2_xnor2_1 _1313_ (.Y(_0373_),
    .A(net150),
    .B(_0106_));
 sg13g2_nor2_1 _1314_ (.A(_0346_),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_a21oi_1 _1315_ (.A1(net148),
    .A2(_0098_),
    .Y(_0375_),
    .B1(net147));
 sg13g2_nor3_2 _1316_ (.A(_0341_),
    .B(_0374_),
    .C(_0375_),
    .Y(_0376_));
 sg13g2_o21ai_1 _1317_ (.B1(_0376_),
    .Y(_0377_),
    .A1(_0363_),
    .A2(_0366_));
 sg13g2_a21oi_2 _1318_ (.B1(_0371_),
    .Y(_0378_),
    .A2(_0377_),
    .A1(_0370_));
 sg13g2_a21o_1 _1319_ (.A2(_0377_),
    .A1(_0370_),
    .B1(_0371_),
    .X(_0379_));
 sg13g2_nor2_1 _1320_ (.A(_0370_),
    .B(_0376_),
    .Y(_0380_));
 sg13g2_and2_1 _1321_ (.A(_0371_),
    .B(_0380_),
    .X(_0381_));
 sg13g2_a21o_1 _1322_ (.A2(_0378_),
    .A1(_0370_),
    .B1(_0381_),
    .X(_0382_));
 sg13g2_nand2_1 _1323_ (.Y(_0383_),
    .A(_0376_),
    .B(_0379_));
 sg13g2_a21oi_1 _1324_ (.A1(_0364_),
    .A2(_0367_),
    .Y(_0384_),
    .B1(_0369_));
 sg13g2_a21o_1 _1325_ (.A2(_0379_),
    .A1(_0376_),
    .B1(_0384_),
    .X(_0385_));
 sg13g2_nand3_1 _1326_ (.B(_0379_),
    .C(_0384_),
    .A(_0376_),
    .Y(_0386_));
 sg13g2_nand2_1 _1327_ (.Y(_0387_),
    .A(_0385_),
    .B(_0386_));
 sg13g2_nand2_1 _1328_ (.Y(_0388_),
    .A(_0372_),
    .B(_0380_));
 sg13g2_a221oi_1 _1329_ (.B2(_0372_),
    .C1(_0350_),
    .B1(_0380_),
    .A1(_0376_),
    .Y(_0389_),
    .A2(_0379_));
 sg13g2_a21oi_1 _1330_ (.A1(_0385_),
    .A2(_0386_),
    .Y(_0390_),
    .B1(_0389_));
 sg13g2_nor2_1 _1331_ (.A(_0382_),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_o21ai_1 _1332_ (.B1(_0352_),
    .Y(_0392_),
    .A1(_0382_),
    .A2(_0390_));
 sg13g2_nor2_1 _1333_ (.A(_0350_),
    .B(_0351_),
    .Y(_0393_));
 sg13g2_a21oi_1 _1334_ (.A1(_0383_),
    .A2(_0388_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_a221oi_1 _1335_ (.B2(_0394_),
    .C1(_0382_),
    .B1(_0392_),
    .A1(_0387_),
    .Y(_0395_),
    .A2(_0391_));
 sg13g2_a21oi_1 _1336_ (.A1(_0096_),
    .A2(_0395_),
    .Y(_0396_),
    .B1(_0344_));
 sg13g2_nand4_1 _1337_ (.B(_0282_),
    .C(_0340_),
    .A(_0188_),
    .Y(_0397_),
    .D(_0396_));
 sg13g2_o21ai_1 _1338_ (.B1(_0198_),
    .Y(_0398_),
    .A1(_0205_),
    .A2(_0266_));
 sg13g2_nor3_1 _1339_ (.A(_0198_),
    .B(_0326_),
    .C(_0332_),
    .Y(_0399_));
 sg13g2_a21oi_1 _1340_ (.A1(_0096_),
    .A2(_0391_),
    .Y(_0400_),
    .B1(_0344_));
 sg13g2_nor2b_1 _1341_ (.A(_0399_),
    .B_N(_0400_),
    .Y(_0401_));
 sg13g2_o21ai_1 _1342_ (.B1(_0095_),
    .Y(_0402_),
    .A1(_0103_),
    .A2(_0174_));
 sg13g2_nand3_1 _1343_ (.B(_0401_),
    .C(_0402_),
    .A(_0398_),
    .Y(_0403_));
 sg13g2_nand2_1 _1344_ (.Y(_0404_),
    .A(net137),
    .B(_0403_));
 sg13g2_xor2_1 _1345_ (.B(_0403_),
    .A(net137),
    .X(_0405_));
 sg13g2_nand2_1 _1346_ (.Y(_0406_),
    .A(_0109_),
    .B(_0186_));
 sg13g2_nand4_1 _1347_ (.B(_0195_),
    .C(_0208_),
    .A(\top.controller.s1[6] ),
    .Y(_0407_),
    .D(_0294_));
 sg13g2_o21ai_1 _1348_ (.B1(_0407_),
    .Y(_0408_),
    .A1(_0190_),
    .A2(_0302_));
 sg13g2_nand3b_1 _1349_ (.B(_0345_),
    .C(_0408_),
    .Y(_0409_),
    .A_N(_0114_));
 sg13g2_a21oi_2 _1350_ (.B1(_0284_),
    .Y(_0410_),
    .A2(_0289_),
    .A1(_0192_));
 sg13g2_nor2_2 _1351_ (.A(_0190_),
    .B(_0410_),
    .Y(_0411_));
 sg13g2_nand2b_2 _1352_ (.Y(_0412_),
    .B(_0189_),
    .A_N(_0410_));
 sg13g2_a221oi_1 _1353_ (.B2(_0339_),
    .C1(_0409_),
    .B1(_0411_),
    .A1(net142),
    .Y(_0413_),
    .A2(_0395_));
 sg13g2_nor3_2 _1354_ (.A(_0276_),
    .B(_0280_),
    .C(_0411_),
    .Y(_0414_));
 sg13g2_nand3_1 _1355_ (.B(_0279_),
    .C(_0412_),
    .A(_0277_),
    .Y(_0415_));
 sg13g2_nand3_1 _1356_ (.B(_0413_),
    .C(_0415_),
    .A(_0406_),
    .Y(_0416_));
 sg13g2_nor3_1 _1357_ (.A(_0206_),
    .B(_0209_),
    .C(_0210_),
    .Y(_0417_));
 sg13g2_a21oi_1 _1358_ (.A1(_0122_),
    .A2(_0123_),
    .Y(_0418_),
    .B1(_0417_));
 sg13g2_nand4_1 _1359_ (.B(net149),
    .C(_0100_),
    .A(_0085_),
    .Y(_0419_),
    .D(net143));
 sg13g2_o21ai_1 _1360_ (.B1(_0143_),
    .Y(_0420_),
    .A1(_0090_),
    .A2(_0419_));
 sg13g2_nand3_1 _1361_ (.B(_0418_),
    .C(_0420_),
    .A(_0218_),
    .Y(_0421_));
 sg13g2_nor2_1 _1362_ (.A(_0174_),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_nor3_2 _1363_ (.A(_0174_),
    .B(_0266_),
    .C(_0421_),
    .Y(_0423_));
 sg13g2_inv_2 _1364_ (.Y(_0424_),
    .A(_0423_));
 sg13g2_o21ai_1 _1365_ (.B1(_0413_),
    .Y(_0425_),
    .A1(net142),
    .A2(_0187_));
 sg13g2_nor2_2 _1366_ (.A(_0414_),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_o21ai_1 _1367_ (.B1(_0424_),
    .Y(_0427_),
    .A1(_0414_),
    .A2(_0425_));
 sg13g2_nand2_1 _1368_ (.Y(_0428_),
    .A(_0405_),
    .B(_0427_));
 sg13g2_nand3_1 _1369_ (.B(_0413_),
    .C(_0415_),
    .A(_0406_),
    .Y(_0429_));
 sg13g2_xor2_1 _1370_ (.B(_0427_),
    .A(_0405_),
    .X(_0430_));
 sg13g2_o21ai_1 _1371_ (.B1(_0422_),
    .Y(_0431_),
    .A1(_0276_),
    .A2(_0280_));
 sg13g2_o21ai_1 _1372_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0397_),
    .A2(_0426_));
 sg13g2_a21oi_2 _1373_ (.B1(_0432_),
    .Y(_0433_),
    .A2(_0426_),
    .A1(net137));
 sg13g2_inv_2 _1374_ (.Y(_0434_),
    .A(_0433_));
 sg13g2_a221oi_1 _1375_ (.B2(_0333_),
    .C1(_0409_),
    .B1(_0411_),
    .A1(net142),
    .Y(_0435_),
    .A2(_0391_));
 sg13g2_o21ai_1 _1376_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0267_),
    .A2(_0411_));
 sg13g2_a21oi_2 _1377_ (.B1(_0436_),
    .Y(_0437_),
    .A2(_0174_),
    .A1(_0109_));
 sg13g2_nand2b_1 _1378_ (.Y(_0438_),
    .B(_0437_),
    .A_N(_0403_));
 sg13g2_nor3_2 _1379_ (.A(_0164_),
    .B(_0255_),
    .C(_0421_),
    .Y(_0439_));
 sg13g2_inv_2 _1380_ (.Y(_0440_),
    .A(_0439_));
 sg13g2_o21ai_1 _1381_ (.B1(_0198_),
    .Y(_0441_),
    .A1(_0205_),
    .A2(_0255_));
 sg13g2_o21ai_1 _1382_ (.B1(_0095_),
    .Y(_0442_),
    .A1(_0103_),
    .A2(_0164_));
 sg13g2_nand2b_1 _1383_ (.Y(_0443_),
    .B(_0325_),
    .A_N(_0198_));
 sg13g2_a21oi_1 _1384_ (.A1(_0096_),
    .A2(_0378_),
    .Y(_0444_),
    .B1(_0344_));
 sg13g2_nand4_1 _1385_ (.B(_0442_),
    .C(_0443_),
    .A(_0441_),
    .Y(_0445_),
    .D(_0444_));
 sg13g2_nand2_1 _1386_ (.Y(_0446_),
    .A(net142),
    .B(_0379_));
 sg13g2_o21ai_1 _1387_ (.B1(_0446_),
    .Y(_0447_),
    .A1(net142),
    .A2(_0164_));
 sg13g2_nand2_1 _1388_ (.Y(_0448_),
    .A(_0325_),
    .B(_0411_));
 sg13g2_a21oi_1 _1389_ (.A1(_0325_),
    .A2(_0411_),
    .Y(_0449_),
    .B1(_0409_));
 sg13g2_nand2_1 _1390_ (.Y(_0450_),
    .A(_0255_),
    .B(_0412_));
 sg13g2_nand3_1 _1391_ (.B(_0449_),
    .C(_0450_),
    .A(_0447_),
    .Y(_0451_));
 sg13g2_nand2_1 _1392_ (.Y(_0452_),
    .A(_0109_),
    .B(_0164_));
 sg13g2_nand2_1 _1393_ (.Y(_0453_),
    .A(net142),
    .B(_0378_));
 sg13g2_a21oi_1 _1394_ (.A1(net142),
    .A2(_0378_),
    .Y(_0454_),
    .B1(_0409_));
 sg13g2_nand4_1 _1395_ (.B(_0450_),
    .C(_0452_),
    .A(_0448_),
    .Y(_0455_),
    .D(_0454_));
 sg13g2_nand4_1 _1396_ (.B(_0450_),
    .C(_0452_),
    .A(_0449_),
    .Y(_0456_),
    .D(_0453_));
 sg13g2_xnor2_1 _1397_ (.Y(_0457_),
    .A(_0445_),
    .B(_0455_));
 sg13g2_or2_1 _1398_ (.X(_0458_),
    .B(_0457_),
    .A(_0440_));
 sg13g2_xnor2_1 _1399_ (.Y(_0459_),
    .A(_0440_),
    .B(_0457_));
 sg13g2_or2_1 _1400_ (.X(_0460_),
    .B(_0459_),
    .A(_0438_));
 sg13g2_xnor2_1 _1401_ (.Y(_0461_),
    .A(_0438_),
    .B(_0459_));
 sg13g2_xor2_1 _1402_ (.B(_0437_),
    .A(_0403_),
    .X(_0462_));
 sg13g2_and2_1 _1403_ (.A(_0424_),
    .B(_0462_),
    .X(_0463_));
 sg13g2_nand2_1 _1404_ (.Y(_0464_),
    .A(_0424_),
    .B(_0462_));
 sg13g2_or3_1 _1405_ (.A(net137),
    .B(_0416_),
    .C(_0463_),
    .X(_0465_));
 sg13g2_nand3b_1 _1406_ (.B(_0426_),
    .C(_0464_),
    .Y(_0466_),
    .A_N(_0397_));
 sg13g2_xnor2_1 _1407_ (.Y(_0467_),
    .A(_0461_),
    .B(_0466_));
 sg13g2_inv_4 _1408_ (.A(net134),
    .Y(_0468_));
 sg13g2_nand2b_1 _1409_ (.Y(_0469_),
    .B(_0418_),
    .A_N(_0143_));
 sg13g2_or3_2 _1410_ (.A(_0216_),
    .B(_0246_),
    .C(_0469_),
    .X(_0470_));
 sg13g2_inv_2 _1411_ (.Y(_0471_),
    .A(_0470_));
 sg13g2_o21ai_1 _1412_ (.B1(_0198_),
    .Y(_0472_),
    .A1(_0205_),
    .A2(_0246_));
 sg13g2_nor2_1 _1413_ (.A(_0198_),
    .B(_0314_),
    .Y(_0473_));
 sg13g2_nor2_1 _1414_ (.A(_0095_),
    .B(_0368_),
    .Y(_0474_));
 sg13g2_nor3_1 _1415_ (.A(_0344_),
    .B(_0473_),
    .C(_0474_),
    .Y(_0475_));
 sg13g2_o21ai_1 _1416_ (.B1(_0095_),
    .Y(_0476_),
    .A1(_0103_),
    .A2(_0157_));
 sg13g2_nand3_1 _1417_ (.B(_0475_),
    .C(_0476_),
    .A(_0472_),
    .Y(_0477_));
 sg13g2_nor2_1 _1418_ (.A(_0246_),
    .B(_0411_),
    .Y(_0478_));
 sg13g2_a21oi_1 _1419_ (.A1(_0314_),
    .A2(_0411_),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_nand2_1 _1420_ (.Y(_0480_),
    .A(_0109_),
    .B(_0157_));
 sg13g2_o21ai_1 _1421_ (.B1(net142),
    .Y(_0481_),
    .A1(_0365_),
    .A2(_0367_));
 sg13g2_nand3b_1 _1422_ (.B(_0480_),
    .C(_0481_),
    .Y(_0482_),
    .A_N(_0409_));
 sg13g2_nand2_1 _1423_ (.Y(_0483_),
    .A(_0246_),
    .B(_0412_));
 sg13g2_nor2_1 _1424_ (.A(_0314_),
    .B(_0412_),
    .Y(_0484_));
 sg13g2_nor2_1 _1425_ (.A(_0409_),
    .B(_0484_),
    .Y(_0485_));
 sg13g2_and4_2 _1426_ (.A(_0480_),
    .B(_0481_),
    .C(_0483_),
    .D(_0485_),
    .X(_0486_));
 sg13g2_or3_1 _1427_ (.A(_0477_),
    .B(_0479_),
    .C(_0482_),
    .X(_0487_));
 sg13g2_nor2b_1 _1428_ (.A(_0477_),
    .B_N(_0486_),
    .Y(_0488_));
 sg13g2_xor2_1 _1429_ (.B(_0486_),
    .A(_0477_),
    .X(_0489_));
 sg13g2_or2_1 _1430_ (.X(_0490_),
    .B(_0489_),
    .A(_0470_));
 sg13g2_xnor2_1 _1431_ (.Y(_0491_),
    .A(_0471_),
    .B(_0489_));
 sg13g2_o21ai_1 _1432_ (.B1(_0458_),
    .Y(_0492_),
    .A1(_0445_),
    .A2(_0451_));
 sg13g2_o21ai_1 _1433_ (.B1(_0458_),
    .Y(_0493_),
    .A1(_0445_),
    .A2(_0455_));
 sg13g2_nand2_1 _1434_ (.Y(_0494_),
    .A(_0491_),
    .B(_0492_));
 sg13g2_xor2_1 _1435_ (.B(_0493_),
    .A(_0491_),
    .X(_0495_));
 sg13g2_o21ai_1 _1436_ (.B1(_0460_),
    .Y(_0496_),
    .A1(_0461_),
    .A2(_0465_));
 sg13g2_nand2_1 _1437_ (.Y(_0497_),
    .A(_0495_),
    .B(_0496_));
 sg13g2_nand4_1 _1438_ (.B(_0490_),
    .C(_0494_),
    .A(_0487_),
    .Y(_0498_),
    .D(_0497_));
 sg13g2_nand2_1 _1439_ (.Y(_0499_),
    .A(_0431_),
    .B(_0445_));
 sg13g2_nor2_1 _1440_ (.A(_0404_),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_inv_1 _1441_ (.Y(_0501_),
    .A(_0500_));
 sg13g2_xnor2_1 _1442_ (.Y(_0502_),
    .A(_0404_),
    .B(_0499_));
 sg13g2_and2_1 _1443_ (.A(_0437_),
    .B(_0439_),
    .X(_0503_));
 sg13g2_inv_1 _1444_ (.Y(_0504_),
    .A(_0503_));
 sg13g2_xnor2_1 _1445_ (.Y(_0505_),
    .A(_0437_),
    .B(_0439_));
 sg13g2_or2_1 _1446_ (.X(_0506_),
    .B(_0505_),
    .A(_0502_));
 sg13g2_or3_2 _1447_ (.A(_0414_),
    .B(_0425_),
    .C(_0455_),
    .X(_0507_));
 sg13g2_o21ai_1 _1448_ (.B1(_0455_),
    .Y(_0508_),
    .A1(_0414_),
    .A2(_0425_));
 sg13g2_xor2_1 _1449_ (.B(_0456_),
    .A(_0429_),
    .X(_0509_));
 sg13g2_a21oi_2 _1450_ (.B1(_0471_),
    .Y(_0510_),
    .A2(_0508_),
    .A1(_0507_));
 sg13g2_and3_1 _1451_ (.X(_0511_),
    .A(_0471_),
    .B(_0507_),
    .C(_0508_));
 sg13g2_nand3_1 _1452_ (.B(_0507_),
    .C(_0508_),
    .A(_0471_),
    .Y(_0512_));
 sg13g2_nor3_2 _1453_ (.A(_0504_),
    .B(_0510_),
    .C(_0511_),
    .Y(_0513_));
 sg13g2_nand3b_1 _1454_ (.B(_0512_),
    .C(_0503_),
    .Y(_0514_),
    .A_N(_0510_));
 sg13g2_o21ai_1 _1455_ (.B1(_0504_),
    .Y(_0515_),
    .A1(_0510_),
    .A2(_0511_));
 sg13g2_nor2b_1 _1456_ (.A(_0423_),
    .B_N(_0477_),
    .Y(_0516_));
 sg13g2_nor2b_1 _1457_ (.A(_0431_),
    .B_N(_0516_),
    .Y(_0517_));
 sg13g2_inv_1 _1458_ (.Y(_0518_),
    .A(_0517_));
 sg13g2_xnor2_1 _1459_ (.Y(_0519_),
    .A(_0431_),
    .B(_0516_));
 sg13g2_a21oi_1 _1460_ (.A1(_0514_),
    .A2(_0515_),
    .Y(_0520_),
    .B1(_0519_));
 sg13g2_nand3_1 _1461_ (.B(_0515_),
    .C(_0519_),
    .A(_0514_),
    .Y(_0521_));
 sg13g2_nand2b_1 _1462_ (.Y(_0522_),
    .B(_0521_),
    .A_N(_0520_));
 sg13g2_a21oi_2 _1463_ (.B1(_0522_),
    .Y(_0523_),
    .A2(_0506_),
    .A1(_0501_));
 sg13g2_nand2_2 _1464_ (.Y(_0524_),
    .A(_0431_),
    .B(_0440_));
 sg13g2_nor2_1 _1465_ (.A(_0424_),
    .B(_0524_),
    .Y(_0525_));
 sg13g2_nand2_1 _1466_ (.Y(_0526_),
    .A(_0424_),
    .B(_0524_));
 sg13g2_nand2b_1 _1467_ (.Y(_0527_),
    .B(_0526_),
    .A_N(_0525_));
 sg13g2_nand2_1 _1468_ (.Y(_0528_),
    .A(_0437_),
    .B(_0486_));
 sg13g2_xor2_1 _1469_ (.B(_0486_),
    .A(_0437_),
    .X(_0529_));
 sg13g2_inv_1 _1470_ (.Y(_0530_),
    .A(_0529_));
 sg13g2_nor2_1 _1471_ (.A(_0507_),
    .B(_0530_),
    .Y(_0531_));
 sg13g2_nand2b_1 _1472_ (.Y(_0532_),
    .B(_0529_),
    .A_N(_0507_));
 sg13g2_xnor2_1 _1473_ (.Y(_0533_),
    .A(_0507_),
    .B(_0529_));
 sg13g2_nand3_1 _1474_ (.B(_0509_),
    .C(_0529_),
    .A(_0471_),
    .Y(_0534_));
 sg13g2_mux2_1 _1475_ (.A0(_0530_),
    .A1(_0533_),
    .S(_0512_),
    .X(_0535_));
 sg13g2_xor2_1 _1476_ (.B(_0535_),
    .A(_0527_),
    .X(_0536_));
 sg13g2_a21oi_1 _1477_ (.A1(_0518_),
    .A2(_0521_),
    .Y(_0537_),
    .B1(_0536_));
 sg13g2_a21o_1 _1478_ (.A2(_0521_),
    .A1(_0518_),
    .B1(_0536_),
    .X(_0538_));
 sg13g2_nand3_1 _1479_ (.B(_0521_),
    .C(_0536_),
    .A(_0518_),
    .Y(_0539_));
 sg13g2_a21oi_1 _1480_ (.A1(_0538_),
    .A2(_0539_),
    .Y(_0540_),
    .B1(_0513_));
 sg13g2_nand3_1 _1481_ (.B(_0538_),
    .C(_0539_),
    .A(_0513_),
    .Y(_0541_));
 sg13g2_nor2b_1 _1482_ (.A(_0540_),
    .B_N(_0541_),
    .Y(_0542_));
 sg13g2_nand3b_1 _1483_ (.B(_0541_),
    .C(_0523_),
    .Y(_0543_),
    .A_N(_0540_));
 sg13g2_a21oi_2 _1484_ (.B1(_0537_),
    .Y(_0544_),
    .A2(_0539_),
    .A1(_0513_));
 sg13g2_nand2_1 _1485_ (.Y(_0545_),
    .A(_0423_),
    .B(_0470_));
 sg13g2_xnor2_1 _1486_ (.Y(_0546_),
    .A(_0423_),
    .B(_0471_));
 sg13g2_or2_1 _1487_ (.X(_0547_),
    .B(_0546_),
    .A(_0524_));
 sg13g2_and2_1 _1488_ (.A(_0524_),
    .B(_0546_),
    .X(_0548_));
 sg13g2_xor2_1 _1489_ (.B(_0546_),
    .A(_0524_),
    .X(_0549_));
 sg13g2_and4_1 _1490_ (.A(_0437_),
    .B(_0486_),
    .C(_0507_),
    .D(_0508_),
    .X(_0550_));
 sg13g2_a22oi_1 _1491_ (.Y(_0551_),
    .B1(_0507_),
    .B2(_0508_),
    .A2(_0486_),
    .A1(_0437_));
 sg13g2_o21ai_1 _1492_ (.B1(_0532_),
    .Y(_0552_),
    .A1(_0550_),
    .A2(_0551_));
 sg13g2_xnor2_1 _1493_ (.Y(_0553_),
    .A(_0549_),
    .B(_0552_));
 sg13g2_a21o_1 _1494_ (.A2(_0535_),
    .A1(_0526_),
    .B1(_0525_),
    .X(_0554_));
 sg13g2_nor2b_1 _1495_ (.A(_0553_),
    .B_N(_0554_),
    .Y(_0555_));
 sg13g2_xor2_1 _1496_ (.B(_0554_),
    .A(_0553_),
    .X(_0556_));
 sg13g2_or2_1 _1497_ (.X(_0557_),
    .B(_0556_),
    .A(_0534_));
 sg13g2_xor2_1 _1498_ (.B(_0556_),
    .A(_0534_),
    .X(_0558_));
 sg13g2_inv_1 _1499_ (.Y(_0559_),
    .A(_0558_));
 sg13g2_xor2_1 _1500_ (.B(_0558_),
    .A(_0544_),
    .X(_0560_));
 sg13g2_nor2_1 _1501_ (.A(_0543_),
    .B(_0560_),
    .Y(_0561_));
 sg13g2_or2_1 _1502_ (.X(_0562_),
    .B(_0550_),
    .A(_0533_));
 sg13g2_nor2_1 _1503_ (.A(_0424_),
    .B(_0470_),
    .Y(_0563_));
 sg13g2_nor3_2 _1504_ (.A(_0533_),
    .B(_0550_),
    .C(_0563_),
    .Y(_0564_));
 sg13g2_nand2b_1 _1505_ (.Y(_0565_),
    .B(_0549_),
    .A_N(_0564_));
 sg13g2_xnor2_1 _1506_ (.Y(_0566_),
    .A(_0549_),
    .B(_0564_));
 sg13g2_a21oi_1 _1507_ (.A1(_0549_),
    .A2(_0552_),
    .Y(_0567_),
    .B1(_0548_));
 sg13g2_nand2b_1 _1508_ (.Y(_0568_),
    .B(_0566_),
    .A_N(_0567_));
 sg13g2_xnor2_1 _1509_ (.Y(_0569_),
    .A(_0566_),
    .B(_0567_));
 sg13g2_o21ai_1 _1510_ (.B1(_0557_),
    .Y(_0570_),
    .A1(_0555_),
    .A2(_0569_));
 sg13g2_o21ai_1 _1511_ (.B1(_0570_),
    .Y(_0571_),
    .A1(_0544_),
    .A2(_0559_));
 sg13g2_nor3_1 _1512_ (.A(_0543_),
    .B(_0560_),
    .C(_0570_),
    .Y(_0572_));
 sg13g2_a21o_1 _1513_ (.A2(_0565_),
    .A1(_0547_),
    .B1(_0553_),
    .X(_0573_));
 sg13g2_nand3_1 _1514_ (.B(_0553_),
    .C(_0565_),
    .A(_0547_),
    .Y(_0574_));
 sg13g2_nand2_1 _1515_ (.Y(_0575_),
    .A(_0573_),
    .B(_0574_));
 sg13g2_and3_1 _1516_ (.X(_0576_),
    .A(_0557_),
    .B(_0568_),
    .C(_0575_));
 sg13g2_nor2_1 _1517_ (.A(net128),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_o21ai_1 _1518_ (.B1(_0460_),
    .Y(_0578_),
    .A1(_0461_),
    .A2(_0466_));
 sg13g2_nand2_1 _1519_ (.Y(_0579_),
    .A(_0495_),
    .B(_0578_));
 sg13g2_xor2_1 _1520_ (.B(_0578_),
    .A(_0495_),
    .X(_0580_));
 sg13g2_inv_1 _1521_ (.Y(_0581_),
    .A(_0580_));
 sg13g2_nor2_1 _1522_ (.A(_0423_),
    .B(_0439_),
    .Y(_0582_));
 sg13g2_inv_1 _1523_ (.Y(_0583_),
    .A(_0582_));
 sg13g2_nor2b_1 _1524_ (.A(_0431_),
    .B_N(_0545_),
    .Y(_0584_));
 sg13g2_a21oi_1 _1525_ (.A1(_0424_),
    .A2(_0471_),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_o21ai_1 _1526_ (.B1(net137),
    .Y(_0586_),
    .A1(_0583_),
    .A2(_0585_));
 sg13g2_a21o_1 _1527_ (.A2(_0585_),
    .A1(_0583_),
    .B1(_0586_),
    .X(_0587_));
 sg13g2_a22oi_1 _1528_ (.Y(_0588_),
    .B1(_0549_),
    .B2(_0552_),
    .A2(_0470_),
    .A1(_0439_));
 sg13g2_nor2_1 _1529_ (.A(_0587_),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_xnor2_1 _1530_ (.Y(_0590_),
    .A(_0587_),
    .B(_0588_));
 sg13g2_nor2_1 _1531_ (.A(_0573_),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_xor2_1 _1532_ (.B(_0590_),
    .A(_0573_),
    .X(_0592_));
 sg13g2_a21oi_1 _1533_ (.A1(_0562_),
    .A2(_0592_),
    .Y(_0593_),
    .B1(_0591_));
 sg13g2_o21ai_1 _1534_ (.B1(_0403_),
    .Y(_0594_),
    .A1(_0439_),
    .A2(_0546_));
 sg13g2_a21o_1 _1535_ (.A2(_0470_),
    .A1(_0439_),
    .B1(_0594_),
    .X(_0595_));
 sg13g2_nor2b_1 _1536_ (.A(_0595_),
    .B_N(_0586_),
    .Y(_0596_));
 sg13g2_xnor2_1 _1537_ (.Y(_0597_),
    .A(_0586_),
    .B(_0595_));
 sg13g2_and2_1 _1538_ (.A(_0589_),
    .B(_0597_),
    .X(_0598_));
 sg13g2_xor2_1 _1539_ (.B(_0597_),
    .A(_0589_),
    .X(_0599_));
 sg13g2_a21oi_2 _1540_ (.B1(_0531_),
    .Y(_0600_),
    .A2(_0528_),
    .A1(_0455_));
 sg13g2_xor2_1 _1541_ (.B(_0600_),
    .A(_0599_),
    .X(_0601_));
 sg13g2_nor2b_1 _1542_ (.A(_0593_),
    .B_N(_0601_),
    .Y(_0602_));
 sg13g2_nand2_1 _1543_ (.Y(_0603_),
    .A(_0403_),
    .B(_0545_));
 sg13g2_nand3_1 _1544_ (.B(_0445_),
    .C(_0470_),
    .A(_0440_),
    .Y(_0604_));
 sg13g2_nor2_1 _1545_ (.A(_0603_),
    .B(_0604_),
    .Y(_0605_));
 sg13g2_xnor2_1 _1546_ (.Y(_0606_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_xor2_1 _1547_ (.B(_0606_),
    .A(_0596_),
    .X(_0607_));
 sg13g2_nor2_1 _1548_ (.A(_0486_),
    .B(_0531_),
    .Y(_0608_));
 sg13g2_nor2b_1 _1549_ (.A(_0608_),
    .B_N(_0607_),
    .Y(_0609_));
 sg13g2_xnor2_1 _1550_ (.Y(_0610_),
    .A(_0607_),
    .B(_0608_));
 sg13g2_a21oi_1 _1551_ (.A1(_0599_),
    .A2(_0600_),
    .Y(_0611_),
    .B1(_0598_));
 sg13g2_nand2b_1 _1552_ (.Y(_0612_),
    .B(_0610_),
    .A_N(_0611_));
 sg13g2_xnor2_1 _1553_ (.Y(_0613_),
    .A(_0610_),
    .B(_0611_));
 sg13g2_o21ai_1 _1554_ (.B1(_0613_),
    .Y(_0614_),
    .A1(net128),
    .A2(_0602_));
 sg13g2_or3_1 _1555_ (.A(net128),
    .B(_0602_),
    .C(_0613_),
    .X(_0615_));
 sg13g2_and2_1 _1556_ (.A(_0614_),
    .B(_0615_),
    .X(_0616_));
 sg13g2_inv_1 _1557_ (.Y(_0617_),
    .A(_0616_));
 sg13g2_and3_1 _1558_ (.X(_0618_),
    .A(net130),
    .B(_0614_),
    .C(_0615_));
 sg13g2_nand2_1 _1559_ (.Y(_0619_),
    .A(net130),
    .B(_0616_));
 sg13g2_a21oi_1 _1560_ (.A1(_0614_),
    .A2(_0615_),
    .Y(_0620_),
    .B1(net130));
 sg13g2_nor2_1 _1561_ (.A(_0618_),
    .B(_0620_),
    .Y(_0621_));
 sg13g2_nor2b_1 _1562_ (.A(_0601_),
    .B_N(_0593_),
    .Y(_0622_));
 sg13g2_nor3_2 _1563_ (.A(net128),
    .B(_0602_),
    .C(_0622_),
    .Y(_0623_));
 sg13g2_nor2_1 _1564_ (.A(net135),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_o21ai_1 _1565_ (.B1(_0463_),
    .Y(_0625_),
    .A1(net137),
    .A2(_0416_));
 sg13g2_and2_1 _1566_ (.A(_0466_),
    .B(_0625_),
    .X(_0626_));
 sg13g2_nand2_2 _1567_ (.Y(_0627_),
    .A(_0466_),
    .B(_0625_));
 sg13g2_xnor2_1 _1568_ (.Y(_0628_),
    .A(_0562_),
    .B(_0592_));
 sg13g2_nor2_1 _1569_ (.A(net128),
    .B(_0628_),
    .Y(_0629_));
 sg13g2_nor3_1 _1570_ (.A(net128),
    .B(net132),
    .C(_0628_),
    .Y(_0630_));
 sg13g2_o21ai_1 _1571_ (.B1(net132),
    .Y(_0631_),
    .A1(net128),
    .A2(_0628_));
 sg13g2_nand2b_1 _1572_ (.Y(_0632_),
    .B(_0631_),
    .A_N(_0630_));
 sg13g2_o21ai_1 _1573_ (.B1(_0434_),
    .Y(_0633_),
    .A1(net128),
    .A2(_0576_));
 sg13g2_a21oi_1 _1574_ (.A1(_0631_),
    .A2(_0633_),
    .Y(_0634_),
    .B1(_0630_));
 sg13g2_a221oi_1 _1575_ (.B2(_0633_),
    .C1(_0630_),
    .B1(_0631_),
    .A1(net135),
    .Y(_0635_),
    .A2(_0623_));
 sg13g2_nor2_1 _1576_ (.A(_0624_),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_or4_1 _1577_ (.A(_0618_),
    .B(_0620_),
    .C(_0624_),
    .D(_0635_),
    .X(_0637_));
 sg13g2_a21oi_1 _1578_ (.A1(_0596_),
    .A2(_0606_),
    .Y(_0638_),
    .B1(_0609_));
 sg13g2_xnor2_1 _1579_ (.Y(_0639_),
    .A(_0477_),
    .B(_0605_));
 sg13g2_xnor2_1 _1580_ (.Y(_0640_),
    .A(_0638_),
    .B(_0639_));
 sg13g2_a21o_1 _1581_ (.A2(_0614_),
    .A1(_0612_),
    .B1(_0640_),
    .X(_0641_));
 sg13g2_nand3_1 _1582_ (.B(_0614_),
    .C(_0640_),
    .A(_0612_),
    .Y(_0642_));
 sg13g2_and2_1 _1583_ (.A(_0641_),
    .B(_0642_),
    .X(_0643_));
 sg13g2_a21oi_1 _1584_ (.A1(_0491_),
    .A2(_0493_),
    .Y(_0644_),
    .B1(_0488_));
 sg13g2_and3_2 _1585_ (.X(_0645_),
    .A(_0490_),
    .B(_0579_),
    .C(_0644_));
 sg13g2_inv_2 _1586_ (.Y(_0646_),
    .A(net129));
 sg13g2_a21o_1 _1587_ (.A2(_0642_),
    .A1(_0641_),
    .B1(_0646_),
    .X(_0647_));
 sg13g2_nand3_1 _1588_ (.B(_0641_),
    .C(_0642_),
    .A(_0498_),
    .Y(_0648_));
 sg13g2_and4_1 _1589_ (.A(_0619_),
    .B(_0637_),
    .C(_0647_),
    .D(_0648_),
    .X(_0649_));
 sg13g2_a22oi_1 _1590_ (.Y(_0650_),
    .B1(_0647_),
    .B2(_0648_),
    .A2(_0637_),
    .A1(_0619_));
 sg13g2_or2_2 _1591_ (.X(_0651_),
    .B(_0650_),
    .A(_0649_));
 sg13g2_nor3_1 _1592_ (.A(net136),
    .B(_0649_),
    .C(_0650_),
    .Y(_0652_));
 sg13g2_xor2_1 _1593_ (.B(_0652_),
    .A(_0577_),
    .X(_0653_));
 sg13g2_xnor2_1 _1594_ (.Y(_0654_),
    .A(_0468_),
    .B(_0623_));
 sg13g2_xnor2_1 _1595_ (.Y(_0655_),
    .A(_0634_),
    .B(_0654_));
 sg13g2_mux2_1 _1596_ (.A0(_0655_),
    .A1(_0623_),
    .S(_0651_),
    .X(_0656_));
 sg13g2_inv_1 _1597_ (.Y(_0657_),
    .A(_0656_));
 sg13g2_nand2_1 _1598_ (.Y(_0658_),
    .A(_0629_),
    .B(_0651_));
 sg13g2_xor2_1 _1599_ (.B(_0633_),
    .A(_0632_),
    .X(_0659_));
 sg13g2_o21ai_1 _1600_ (.B1(_0658_),
    .Y(_0660_),
    .A1(_0651_),
    .A2(_0659_));
 sg13g2_and2_1 _1601_ (.A(net135),
    .B(_0660_),
    .X(_0661_));
 sg13g2_xnor2_1 _1602_ (.Y(_0662_),
    .A(_0468_),
    .B(_0660_));
 sg13g2_nand2_1 _1603_ (.Y(_0663_),
    .A(_0627_),
    .B(_0653_));
 sg13g2_xnor2_1 _1604_ (.Y(_0664_),
    .A(_0627_),
    .B(_0653_));
 sg13g2_xnor2_1 _1605_ (.Y(_0665_),
    .A(_0561_),
    .B(_0571_));
 sg13g2_inv_1 _1606_ (.Y(_0666_),
    .A(_0665_));
 sg13g2_nand2_1 _1607_ (.Y(_0667_),
    .A(_0434_),
    .B(_0665_));
 sg13g2_inv_1 _1608_ (.Y(_0668_),
    .A(_0667_));
 sg13g2_o21ai_1 _1609_ (.B1(_0663_),
    .Y(_0669_),
    .A1(_0664_),
    .A2(_0668_));
 sg13g2_a21oi_1 _1610_ (.A1(_0662_),
    .A2(_0669_),
    .Y(_0670_),
    .B1(_0661_));
 sg13g2_a221oi_1 _1611_ (.B2(_0669_),
    .C1(_0661_),
    .B1(_0662_),
    .A1(net130),
    .Y(_0671_),
    .A2(_0656_));
 sg13g2_nand2_1 _1612_ (.Y(_0672_),
    .A(net131),
    .B(_0657_));
 sg13g2_xnor2_1 _1613_ (.Y(_0673_),
    .A(_0621_),
    .B(_0636_));
 sg13g2_a21oi_1 _1614_ (.A1(_0617_),
    .A2(_0651_),
    .Y(_0674_),
    .B1(_0673_));
 sg13g2_o21ai_1 _1615_ (.B1(_0672_),
    .Y(_0675_),
    .A1(net129),
    .A2(_0674_));
 sg13g2_nor2b_1 _1616_ (.A(_0643_),
    .B_N(_0651_),
    .Y(_0676_));
 sg13g2_a21oi_1 _1617_ (.A1(net129),
    .A2(_0674_),
    .Y(_0677_),
    .B1(_0676_));
 sg13g2_o21ai_1 _1618_ (.B1(_0677_),
    .Y(_0678_),
    .A1(_0671_),
    .A2(_0675_));
 sg13g2_xnor2_1 _1619_ (.Y(_0679_),
    .A(_0664_),
    .B(_0667_));
 sg13g2_mux2_2 _1620_ (.A0(_0653_),
    .A1(_0679_),
    .S(_0678_),
    .X(_0680_));
 sg13g2_xnor2_1 _1621_ (.Y(_0681_),
    .A(_0543_),
    .B(_0560_));
 sg13g2_nand3_1 _1622_ (.B(_0506_),
    .C(_0522_),
    .A(_0501_),
    .Y(_0682_));
 sg13g2_nand2b_1 _1623_ (.Y(_0683_),
    .B(_0682_),
    .A_N(_0523_));
 sg13g2_xnor2_1 _1624_ (.Y(_0684_),
    .A(_0502_),
    .B(_0505_));
 sg13g2_xnor2_1 _1625_ (.Y(_0685_),
    .A(_0523_),
    .B(_0542_));
 sg13g2_nor2_1 _1626_ (.A(_0428_),
    .B(_0684_),
    .Y(_0686_));
 sg13g2_nand2b_1 _1627_ (.Y(_0687_),
    .B(_0686_),
    .A_N(_0683_));
 sg13g2_o21ai_1 _1628_ (.B1(_0681_),
    .Y(_0688_),
    .A1(_0685_),
    .A2(_0687_));
 sg13g2_nand2b_1 _1629_ (.Y(_0689_),
    .B(_0434_),
    .A_N(_0688_));
 sg13g2_inv_1 _1630_ (.Y(_0690_),
    .A(_0689_));
 sg13g2_xnor2_1 _1631_ (.Y(_0691_),
    .A(net136),
    .B(_0665_));
 sg13g2_xnor2_1 _1632_ (.Y(_0692_),
    .A(_0434_),
    .B(_0665_));
 sg13g2_mux2_1 _1633_ (.A0(_0665_),
    .A1(_0691_),
    .S(_0678_),
    .X(_0693_));
 sg13g2_mux2_1 _1634_ (.A0(_0666_),
    .A1(_0692_),
    .S(_0678_),
    .X(_0694_));
 sg13g2_nor2_1 _1635_ (.A(net132),
    .B(_0693_),
    .Y(_0695_));
 sg13g2_xnor2_1 _1636_ (.Y(_0696_),
    .A(_0627_),
    .B(_0693_));
 sg13g2_xnor2_1 _1637_ (.Y(_0697_),
    .A(net132),
    .B(_0693_));
 sg13g2_a22oi_1 _1638_ (.Y(_0698_),
    .B1(_0694_),
    .B2(_0627_),
    .A2(_0680_),
    .A1(net135));
 sg13g2_o21ai_1 _1639_ (.B1(_0698_),
    .Y(_0699_),
    .A1(_0690_),
    .A2(_0697_));
 sg13g2_nor2_1 _1640_ (.A(net135),
    .B(_0680_),
    .Y(_0700_));
 sg13g2_inv_1 _1641_ (.Y(_0701_),
    .A(_0700_));
 sg13g2_and2_1 _1642_ (.A(_0699_),
    .B(_0701_),
    .X(_0702_));
 sg13g2_xor2_1 _1643_ (.B(_0669_),
    .A(_0662_),
    .X(_0703_));
 sg13g2_mux2_1 _1644_ (.A0(_0660_),
    .A1(_0703_),
    .S(_0678_),
    .X(_0704_));
 sg13g2_and2_1 _1645_ (.A(net130),
    .B(_0704_),
    .X(_0705_));
 sg13g2_xnor2_1 _1646_ (.Y(_0706_),
    .A(net131),
    .B(_0704_));
 sg13g2_xnor2_1 _1647_ (.Y(_0707_),
    .A(net130),
    .B(_0656_));
 sg13g2_xnor2_1 _1648_ (.Y(_0708_),
    .A(_0670_),
    .B(_0707_));
 sg13g2_mux2_1 _1649_ (.A0(_0657_),
    .A1(_0708_),
    .S(_0678_),
    .X(_0709_));
 sg13g2_inv_1 _1650_ (.Y(_0710_),
    .A(_0709_));
 sg13g2_or2_1 _1651_ (.X(_0711_),
    .B(_0709_),
    .A(_0646_));
 sg13g2_nand2_1 _1652_ (.Y(_0712_),
    .A(_0646_),
    .B(_0709_));
 sg13g2_and3_1 _1653_ (.X(_0713_),
    .A(_0706_),
    .B(_0711_),
    .C(_0712_));
 sg13g2_and3_1 _1654_ (.X(_0714_),
    .A(_0699_),
    .B(_0701_),
    .C(_0713_));
 sg13g2_nand3_1 _1655_ (.B(_0701_),
    .C(_0713_),
    .A(_0699_),
    .Y(_0715_));
 sg13g2_nand2b_1 _1656_ (.Y(_0716_),
    .B(_0711_),
    .A_N(_0676_));
 sg13g2_a21oi_2 _1657_ (.B1(_0716_),
    .Y(_0717_),
    .A2(_0712_),
    .A1(_0705_));
 sg13g2_a21o_2 _1658_ (.A2(_0712_),
    .A1(_0705_),
    .B1(_0716_),
    .X(_0718_));
 sg13g2_nor2_2 _1659_ (.A(_0714_),
    .B(_0718_),
    .Y(_0719_));
 sg13g2_xnor2_1 _1660_ (.Y(_0720_),
    .A(_0468_),
    .B(_0680_));
 sg13g2_a21oi_1 _1661_ (.A1(_0689_),
    .A2(_0696_),
    .Y(_0721_),
    .B1(_0695_));
 sg13g2_xnor2_1 _1662_ (.Y(_0722_),
    .A(_0720_),
    .B(_0721_));
 sg13g2_nand3_1 _1663_ (.B(_0715_),
    .C(_0717_),
    .A(_0680_),
    .Y(_0723_));
 sg13g2_o21ai_1 _1664_ (.B1(_0722_),
    .Y(_0724_),
    .A1(_0714_),
    .A2(_0718_));
 sg13g2_and2_1 _1665_ (.A(_0723_),
    .B(_0724_),
    .X(_0725_));
 sg13g2_inv_1 _1666_ (.Y(_0726_),
    .A(_0725_));
 sg13g2_xnor2_1 _1667_ (.Y(_0727_),
    .A(net136),
    .B(_0688_));
 sg13g2_o21ai_1 _1668_ (.B1(_0727_),
    .Y(_0728_),
    .A1(_0714_),
    .A2(_0718_));
 sg13g2_nand3_1 _1669_ (.B(_0715_),
    .C(_0717_),
    .A(_0688_),
    .Y(_0729_));
 sg13g2_nand2_1 _1670_ (.Y(_0730_),
    .A(_0728_),
    .B(_0729_));
 sg13g2_nand3_1 _1671_ (.B(_0728_),
    .C(_0729_),
    .A(net132),
    .Y(_0731_));
 sg13g2_a21oi_1 _1672_ (.A1(_0728_),
    .A2(_0729_),
    .Y(_0732_),
    .B1(net132));
 sg13g2_xor2_1 _1673_ (.B(_0687_),
    .A(_0685_),
    .X(_0733_));
 sg13g2_nor2_1 _1674_ (.A(net136),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_inv_1 _1675_ (.Y(_0735_),
    .A(_0734_));
 sg13g2_a21oi_2 _1676_ (.B1(_0732_),
    .Y(_0736_),
    .A2(_0735_),
    .A1(_0731_));
 sg13g2_xnor2_1 _1677_ (.Y(_0737_),
    .A(_0690_),
    .B(_0696_));
 sg13g2_nand3_1 _1678_ (.B(_0715_),
    .C(_0717_),
    .A(_0694_),
    .Y(_0738_));
 sg13g2_o21ai_1 _1679_ (.B1(_0737_),
    .Y(_0739_),
    .A1(_0714_),
    .A2(_0718_));
 sg13g2_and2_1 _1680_ (.A(_0738_),
    .B(_0739_),
    .X(_0740_));
 sg13g2_a21oi_1 _1681_ (.A1(_0738_),
    .A2(_0739_),
    .Y(_0741_),
    .B1(_0468_));
 sg13g2_a21o_1 _1682_ (.A2(_0739_),
    .A1(_0738_),
    .B1(_0468_),
    .X(_0742_));
 sg13g2_nand3_1 _1683_ (.B(_0738_),
    .C(_0739_),
    .A(_0468_),
    .Y(_0743_));
 sg13g2_nand2_1 _1684_ (.Y(_0744_),
    .A(_0742_),
    .B(_0743_));
 sg13g2_nand3_1 _1685_ (.B(_0723_),
    .C(_0724_),
    .A(net131),
    .Y(_0745_));
 sg13g2_a21oi_1 _1686_ (.A1(_0723_),
    .A2(_0724_),
    .Y(_0746_),
    .B1(net131));
 sg13g2_a21o_1 _1687_ (.A2(_0724_),
    .A1(_0723_),
    .B1(net131),
    .X(_0747_));
 sg13g2_nand2_1 _1688_ (.Y(_0748_),
    .A(_0745_),
    .B(_0747_));
 sg13g2_nand4_1 _1689_ (.B(_0743_),
    .C(_0745_),
    .A(_0742_),
    .Y(_0749_),
    .D(_0747_));
 sg13g2_a21oi_1 _1690_ (.A1(_0741_),
    .A2(_0745_),
    .Y(_0750_),
    .B1(_0746_));
 sg13g2_o21ai_1 _1691_ (.B1(_0750_),
    .Y(_0751_),
    .A1(_0736_),
    .A2(_0749_));
 sg13g2_nor2_1 _1692_ (.A(_0702_),
    .B(_0706_),
    .Y(_0752_));
 sg13g2_nand2_1 _1693_ (.Y(_0753_),
    .A(_0702_),
    .B(_0706_));
 sg13g2_nor2_1 _1694_ (.A(_0717_),
    .B(_0752_),
    .Y(_0754_));
 sg13g2_a22oi_1 _1695_ (.Y(_0755_),
    .B1(_0753_),
    .B2(_0754_),
    .A2(_0719_),
    .A1(_0704_));
 sg13g2_xnor2_1 _1696_ (.Y(_0756_),
    .A(net129),
    .B(_0755_));
 sg13g2_nand2b_1 _1697_ (.Y(_0757_),
    .B(_0753_),
    .A_N(_0705_));
 sg13g2_a22oi_1 _1698_ (.Y(_0758_),
    .B1(_0757_),
    .B2(_0716_),
    .A2(_0719_),
    .A1(_0710_));
 sg13g2_o21ai_1 _1699_ (.B1(_0758_),
    .Y(_0759_),
    .A1(_0646_),
    .A2(_0755_));
 sg13g2_a21oi_2 _1700_ (.B1(_0759_),
    .Y(_0760_),
    .A2(_0756_),
    .A1(_0751_));
 sg13g2_o21ai_1 _1701_ (.B1(_0742_),
    .Y(_0761_),
    .A1(_0736_),
    .A2(_0744_));
 sg13g2_xnor2_1 _1702_ (.Y(_0762_),
    .A(_0748_),
    .B(_0761_));
 sg13g2_mux2_1 _1703_ (.A0(_0762_),
    .A1(_0726_),
    .S(_0760_),
    .X(_0763_));
 sg13g2_inv_1 _1704_ (.Y(_0764_),
    .A(_0763_));
 sg13g2_and2_1 _1705_ (.A(net129),
    .B(_0763_),
    .X(_0765_));
 sg13g2_nand2_1 _1706_ (.Y(_0766_),
    .A(_0498_),
    .B(_0764_));
 sg13g2_xnor2_1 _1707_ (.Y(_0767_),
    .A(net129),
    .B(_0763_));
 sg13g2_xnor2_1 _1708_ (.Y(_0768_),
    .A(_0736_),
    .B(_0744_));
 sg13g2_mux2_1 _1709_ (.A0(_0768_),
    .A1(_0740_),
    .S(_0760_),
    .X(_0769_));
 sg13g2_nor2_1 _1710_ (.A(net131),
    .B(_0769_),
    .Y(_0770_));
 sg13g2_xnor2_1 _1711_ (.Y(_0771_),
    .A(net131),
    .B(_0769_));
 sg13g2_or2_1 _1712_ (.X(_0772_),
    .B(_0771_),
    .A(_0767_));
 sg13g2_nand2_1 _1713_ (.Y(_0773_),
    .A(_0730_),
    .B(_0760_));
 sg13g2_xnor2_1 _1714_ (.Y(_0774_),
    .A(net132),
    .B(_0730_));
 sg13g2_xnor2_1 _1715_ (.Y(_0775_),
    .A(_0735_),
    .B(_0774_));
 sg13g2_o21ai_1 _1716_ (.B1(_0773_),
    .Y(_0776_),
    .A1(_0760_),
    .A2(_0775_));
 sg13g2_and2_1 _1717_ (.A(net135),
    .B(_0776_),
    .X(_0777_));
 sg13g2_nor2_1 _1718_ (.A(_0467_),
    .B(_0776_),
    .Y(_0778_));
 sg13g2_or2_1 _1719_ (.X(_0779_),
    .B(_0776_),
    .A(net135));
 sg13g2_xnor2_1 _1720_ (.Y(_0780_),
    .A(net136),
    .B(_0733_));
 sg13g2_mux2_1 _1721_ (.A0(_0780_),
    .A1(_0733_),
    .S(_0760_),
    .X(_0781_));
 sg13g2_and2_1 _1722_ (.A(_0627_),
    .B(_0781_),
    .X(_0782_));
 sg13g2_xnor2_1 _1723_ (.Y(_0783_),
    .A(_0683_),
    .B(_0686_));
 sg13g2_nor2_1 _1724_ (.A(_0433_),
    .B(_0783_),
    .Y(_0784_));
 sg13g2_inv_1 _1725_ (.Y(_0785_),
    .A(_0784_));
 sg13g2_nand2b_1 _1726_ (.Y(_0786_),
    .B(net133),
    .A_N(_0781_));
 sg13g2_nand2b_1 _1727_ (.Y(_0787_),
    .B(_0786_),
    .A_N(_0782_));
 sg13g2_a21o_1 _1728_ (.A2(_0786_),
    .A1(_0785_),
    .B1(_0782_),
    .X(_0788_));
 sg13g2_a21oi_1 _1729_ (.A1(_0779_),
    .A2(_0788_),
    .Y(_0789_),
    .B1(_0777_));
 sg13g2_a221oi_1 _1730_ (.B2(_0786_),
    .C1(_0782_),
    .B1(_0785_),
    .A1(_0467_),
    .Y(_0790_),
    .A2(_0776_));
 sg13g2_nor3_1 _1731_ (.A(_0772_),
    .B(_0778_),
    .C(_0790_),
    .Y(_0791_));
 sg13g2_or3_1 _1732_ (.A(_0772_),
    .B(_0778_),
    .C(_0790_),
    .X(_0792_));
 sg13g2_or2_1 _1733_ (.X(_0793_),
    .B(_0756_),
    .A(_0751_));
 sg13g2_a22oi_1 _1734_ (.Y(_0794_),
    .B1(_0758_),
    .B2(_0755_),
    .A2(_0756_),
    .A1(_0751_));
 sg13g2_a21o_1 _1735_ (.A2(_0794_),
    .A1(_0793_),
    .B1(_0765_),
    .X(_0795_));
 sg13g2_a21oi_2 _1736_ (.B1(_0795_),
    .Y(_0796_),
    .A2(_0770_),
    .A1(_0766_));
 sg13g2_a21o_1 _1737_ (.A2(_0770_),
    .A1(_0766_),
    .B1(_0795_),
    .X(_0797_));
 sg13g2_nand2_2 _1738_ (.Y(_0798_),
    .A(_0792_),
    .B(_0796_));
 sg13g2_xnor2_1 _1739_ (.Y(_0799_),
    .A(_0433_),
    .B(_0783_));
 sg13g2_a21oi_2 _1740_ (.B1(_0799_),
    .Y(_0800_),
    .A2(_0796_),
    .A1(_0792_));
 sg13g2_nor3_1 _1741_ (.A(_0783_),
    .B(_0791_),
    .C(_0797_),
    .Y(_0801_));
 sg13g2_nor2_1 _1742_ (.A(_0800_),
    .B(_0801_),
    .Y(_0802_));
 sg13g2_nor2_1 _1743_ (.A(_0777_),
    .B(_0778_),
    .Y(_0803_));
 sg13g2_xor2_1 _1744_ (.B(_0803_),
    .A(_0788_),
    .X(_0804_));
 sg13g2_mux2_1 _1745_ (.A0(_0776_),
    .A1(_0804_),
    .S(_0798_),
    .X(_0805_));
 sg13g2_nand2b_1 _1746_ (.Y(_0806_),
    .B(_0580_),
    .A_N(_0805_));
 sg13g2_nor3_1 _1747_ (.A(_0781_),
    .B(_0791_),
    .C(_0797_),
    .Y(_0807_));
 sg13g2_xnor2_1 _1748_ (.Y(_0808_),
    .A(_0784_),
    .B(_0787_));
 sg13g2_a21oi_2 _1749_ (.B1(_0807_),
    .Y(_0809_),
    .A2(_0808_),
    .A1(_0798_));
 sg13g2_xnor2_1 _1750_ (.Y(_0810_),
    .A(net134),
    .B(_0809_));
 sg13g2_nor3_1 _1751_ (.A(net133),
    .B(_0800_),
    .C(_0801_),
    .Y(_0811_));
 sg13g2_xor2_1 _1752_ (.B(_0684_),
    .A(_0428_),
    .X(_0812_));
 sg13g2_nor2_1 _1753_ (.A(net136),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_inv_1 _1754_ (.Y(_0814_),
    .A(_0813_));
 sg13g2_o21ai_1 _1755_ (.B1(net133),
    .Y(_0815_),
    .A1(_0800_),
    .A2(_0801_));
 sg13g2_nor2b_1 _1756_ (.A(_0811_),
    .B_N(_0815_),
    .Y(_0816_));
 sg13g2_a21oi_2 _1757_ (.B1(_0811_),
    .Y(_0817_),
    .A2(_0815_),
    .A1(_0814_));
 sg13g2_nor2_1 _1758_ (.A(_0810_),
    .B(_0817_),
    .Y(_0818_));
 sg13g2_a22oi_1 _1759_ (.Y(_0819_),
    .B1(_0809_),
    .B2(net134),
    .A2(_0805_),
    .A1(net130));
 sg13g2_o21ai_1 _1760_ (.B1(_0819_),
    .Y(_0820_),
    .A1(_0810_),
    .A2(_0817_));
 sg13g2_nand2_1 _1761_ (.Y(_0821_),
    .A(_0806_),
    .B(_0820_));
 sg13g2_nor2_1 _1762_ (.A(_0769_),
    .B(_0798_),
    .Y(_0822_));
 sg13g2_nor2_1 _1763_ (.A(_0771_),
    .B(_0789_),
    .Y(_0823_));
 sg13g2_xor2_1 _1764_ (.B(_0789_),
    .A(_0771_),
    .X(_0824_));
 sg13g2_a21oi_2 _1765_ (.B1(_0822_),
    .Y(_0825_),
    .A2(_0824_),
    .A1(_0798_));
 sg13g2_xnor2_1 _1766_ (.Y(_0826_),
    .A(_0645_),
    .B(_0825_));
 sg13g2_and3_1 _1767_ (.X(_0827_),
    .A(_0806_),
    .B(_0820_),
    .C(_0826_));
 sg13g2_nand3_1 _1768_ (.B(_0820_),
    .C(_0826_),
    .A(_0806_),
    .Y(_0828_));
 sg13g2_nand3_1 _1769_ (.B(_0792_),
    .C(_0796_),
    .A(_0763_),
    .Y(_0829_));
 sg13g2_o21ai_1 _1770_ (.B1(_0829_),
    .Y(_0830_),
    .A1(_0646_),
    .A2(_0825_));
 sg13g2_nor2_1 _1771_ (.A(_0770_),
    .B(_0823_),
    .Y(_0831_));
 sg13g2_xor2_1 _1772_ (.B(_0831_),
    .A(_0767_),
    .X(_0832_));
 sg13g2_a21oi_2 _1773_ (.B1(_0830_),
    .Y(_0833_),
    .A2(_0832_),
    .A1(_0798_));
 sg13g2_a21o_1 _1774_ (.A2(_0832_),
    .A1(_0798_),
    .B1(_0830_),
    .X(_0834_));
 sg13g2_nor2_2 _1775_ (.A(_0827_),
    .B(_0834_),
    .Y(_0835_));
 sg13g2_xnor2_1 _1776_ (.Y(_0836_),
    .A(_0813_),
    .B(_0816_));
 sg13g2_mux2_1 _1777_ (.A0(_0836_),
    .A1(_0802_),
    .S(_0835_),
    .X(_0837_));
 sg13g2_nor2_1 _1778_ (.A(net134),
    .B(_0837_),
    .Y(_0838_));
 sg13g2_xnor2_1 _1779_ (.Y(_0839_),
    .A(net136),
    .B(_0812_));
 sg13g2_a21oi_1 _1780_ (.A1(_0828_),
    .A2(_0833_),
    .Y(_0840_),
    .B1(_0839_));
 sg13g2_nor3_2 _1781_ (.A(_0812_),
    .B(_0827_),
    .C(_0834_),
    .Y(_0841_));
 sg13g2_nor2_1 _1782_ (.A(_0840_),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_nor3_1 _1783_ (.A(net133),
    .B(_0840_),
    .C(_0841_),
    .Y(_0843_));
 sg13g2_o21ai_1 _1784_ (.B1(net133),
    .Y(_0844_),
    .A1(_0840_),
    .A2(_0841_));
 sg13g2_nor2b_1 _1785_ (.A(_0843_),
    .B_N(_0844_),
    .Y(_0845_));
 sg13g2_or2_1 _1786_ (.X(_0846_),
    .B(net136),
    .A(_0430_));
 sg13g2_a21oi_1 _1787_ (.A1(_0844_),
    .A2(_0846_),
    .Y(_0847_),
    .B1(_0843_));
 sg13g2_a221oi_1 _1788_ (.B2(_0846_),
    .C1(_0843_),
    .B1(_0844_),
    .A1(net134),
    .Y(_0848_),
    .A2(_0837_));
 sg13g2_nor2_1 _1789_ (.A(_0838_),
    .B(_0848_),
    .Y(_0849_));
 sg13g2_nand3_1 _1790_ (.B(_0828_),
    .C(_0833_),
    .A(_0809_),
    .Y(_0850_));
 sg13g2_xnor2_1 _1791_ (.Y(_0851_),
    .A(_0810_),
    .B(_0817_));
 sg13g2_o21ai_1 _1792_ (.B1(_0850_),
    .Y(_0852_),
    .A1(_0835_),
    .A2(_0851_));
 sg13g2_xnor2_1 _1793_ (.Y(_0853_),
    .A(_0581_),
    .B(_0852_));
 sg13g2_xnor2_1 _1794_ (.Y(_0854_),
    .A(net131),
    .B(_0805_));
 sg13g2_a21oi_1 _1795_ (.A1(net134),
    .A2(_0809_),
    .Y(_0855_),
    .B1(_0818_));
 sg13g2_xnor2_1 _1796_ (.Y(_0856_),
    .A(_0854_),
    .B(_0855_));
 sg13g2_mux2_2 _1797_ (.A0(_0856_),
    .A1(_0805_),
    .S(_0835_),
    .X(_0857_));
 sg13g2_nor2_1 _1798_ (.A(_0645_),
    .B(_0857_),
    .Y(_0858_));
 sg13g2_xnor2_1 _1799_ (.Y(_0859_),
    .A(net129),
    .B(_0857_));
 sg13g2_nor4_2 _1800_ (.A(_0838_),
    .B(_0848_),
    .C(_0853_),
    .Y(_0860_),
    .D(_0859_));
 sg13g2_a21o_1 _1801_ (.A2(_0833_),
    .A1(_0825_),
    .B1(_0827_),
    .X(_0861_));
 sg13g2_a21o_1 _1802_ (.A2(_0834_),
    .A1(_0821_),
    .B1(_0861_),
    .X(_0862_));
 sg13g2_a22oi_1 _1803_ (.Y(_0863_),
    .B1(_0857_),
    .B2(net129),
    .A2(_0852_),
    .A1(_0581_));
 sg13g2_o21ai_1 _1804_ (.B1(_0862_),
    .Y(_0864_),
    .A1(_0858_),
    .A2(_0863_));
 sg13g2_nor2_2 _1805_ (.A(_0860_),
    .B(_0864_),
    .Y(_0865_));
 sg13g2_o21ai_1 _1806_ (.B1(_0434_),
    .Y(_0866_),
    .A1(_0860_),
    .A2(_0864_));
 sg13g2_xnor2_1 _1807_ (.Y(_0867_),
    .A(_0430_),
    .B(_0866_));
 sg13g2_nand3_1 _1808_ (.B(_0426_),
    .C(_0464_),
    .A(net137),
    .Y(_0868_));
 sg13g2_xor2_1 _1809_ (.B(_0846_),
    .A(_0845_),
    .X(_0869_));
 sg13g2_mux2_1 _1810_ (.A0(_0869_),
    .A1(_0842_),
    .S(_0865_),
    .X(_0870_));
 sg13g2_a21oi_1 _1811_ (.A1(net137),
    .A2(_0426_),
    .Y(_0871_),
    .B1(net132));
 sg13g2_a221oi_1 _1812_ (.B2(net134),
    .C1(_0871_),
    .B1(_0870_),
    .A1(_0867_),
    .Y(_0872_),
    .A2(_0868_));
 sg13g2_xnor2_1 _1813_ (.Y(_0873_),
    .A(_0468_),
    .B(_0837_));
 sg13g2_xnor2_1 _1814_ (.Y(_0874_),
    .A(_0847_),
    .B(_0873_));
 sg13g2_mux2_1 _1815_ (.A0(_0874_),
    .A1(_0837_),
    .S(_0865_),
    .X(_0875_));
 sg13g2_nor2_1 _1816_ (.A(net130),
    .B(_0875_),
    .Y(_0876_));
 sg13g2_nor2_1 _1817_ (.A(net134),
    .B(_0870_),
    .Y(_0877_));
 sg13g2_nor3_1 _1818_ (.A(_0872_),
    .B(_0876_),
    .C(_0877_),
    .Y(_0878_));
 sg13g2_xnor2_1 _1819_ (.Y(_0879_),
    .A(_0849_),
    .B(_0853_));
 sg13g2_mux2_1 _1820_ (.A0(_0879_),
    .A1(_0852_),
    .S(_0865_),
    .X(_0880_));
 sg13g2_xor2_1 _1821_ (.B(_0880_),
    .A(_0498_),
    .X(_0881_));
 sg13g2_a21o_1 _1822_ (.A2(_0875_),
    .A1(_0581_),
    .B1(_0881_),
    .X(_0882_));
 sg13g2_nand2b_2 _1823_ (.Y(_0883_),
    .B(\top.controller.ef1 ),
    .A_N(_0572_));
 sg13g2_inv_1 _1824_ (.Y(_0884_),
    .A(_0883_));
 sg13g2_nand2_1 _1825_ (.Y(_0885_),
    .A(_0498_),
    .B(_0862_));
 sg13g2_a21oi_1 _1826_ (.A1(_0857_),
    .A2(_0865_),
    .Y(_0886_),
    .B1(_0885_));
 sg13g2_nor2b_1 _1827_ (.A(_0880_),
    .B_N(_0886_),
    .Y(_0887_));
 sg13g2_nor2_1 _1828_ (.A(_0883_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_o21ai_1 _1829_ (.B1(_0888_),
    .Y(_0889_),
    .A1(_0878_),
    .A2(_0882_));
 sg13g2_a21oi_1 _1830_ (.A1(_0088_),
    .A2(_0889_),
    .Y(_0014_),
    .B1(_0081_));
 sg13g2_nor2_1 _1831_ (.A(_0865_),
    .B(_0883_),
    .Y(_0890_));
 sg13g2_a21oi_1 _1832_ (.A1(net144),
    .A2(net116),
    .Y(_0891_),
    .B1(_0890_));
 sg13g2_nor2_1 _1833_ (.A(net158),
    .B(net117),
    .Y(_0015_));
 sg13g2_nor2_1 _1834_ (.A(_0835_),
    .B(_0883_),
    .Y(_0892_));
 sg13g2_a21oi_1 _1835_ (.A1(_0079_),
    .A2(net100),
    .Y(_0893_),
    .B1(_0892_));
 sg13g2_nor2_1 _1836_ (.A(net158),
    .B(net101),
    .Y(_0016_));
 sg13g2_a22oi_1 _1837_ (.Y(_0894_),
    .B1(_0798_),
    .B2(_0884_),
    .A2(net109),
    .A1(net144));
 sg13g2_nor2_1 _1838_ (.A(net158),
    .B(net110),
    .Y(_0017_));
 sg13g2_nor2_1 _1839_ (.A(_0760_),
    .B(_0883_),
    .Y(_0895_));
 sg13g2_a21oi_1 _1840_ (.A1(net144),
    .A2(net105),
    .Y(_0896_),
    .B1(_0895_));
 sg13g2_nor2_1 _1841_ (.A(net158),
    .B(net106),
    .Y(_0018_));
 sg13g2_nor2_1 _1842_ (.A(_0719_),
    .B(_0883_),
    .Y(_0897_));
 sg13g2_a21oi_1 _1843_ (.A1(net144),
    .A2(net114),
    .Y(_0898_),
    .B1(_0897_));
 sg13g2_nor2_1 _1844_ (.A(net158),
    .B(net115),
    .Y(_0019_));
 sg13g2_a22oi_1 _1845_ (.Y(_0899_),
    .B1(_0678_),
    .B2(_0884_),
    .A2(net118),
    .A1(net144));
 sg13g2_nor2_1 _1846_ (.A(net158),
    .B(net119),
    .Y(_0020_));
 sg13g2_nor2_1 _1847_ (.A(_0651_),
    .B(_0883_),
    .Y(_0900_));
 sg13g2_a21oi_1 _1848_ (.A1(net94),
    .A2(net144),
    .Y(_0901_),
    .B1(_0900_));
 sg13g2_nor2_1 _1849_ (.A(net158),
    .B(net95),
    .Y(_0021_));
 sg13g2_nor4_1 _1850_ (.A(\top.controller.r2[3] ),
    .B(\top.controller.r2[2] ),
    .C(\top.controller.r2[1] ),
    .D(\top.controller.r2[0] ),
    .Y(_0902_));
 sg13g2_nor4_1 _1851_ (.A(\top.controller.r2[7] ),
    .B(\top.controller.r2[6] ),
    .C(\top.controller.r2[5] ),
    .D(\top.controller.r2[4] ),
    .Y(_0903_));
 sg13g2_nor4_1 _1852_ (.A(\top.controller.r1[3] ),
    .B(\top.controller.r1[2] ),
    .C(\top.controller.r1[1] ),
    .D(\top.controller.r1[0] ),
    .Y(_0904_));
 sg13g2_nor4_1 _1853_ (.A(\top.controller.r1[7] ),
    .B(\top.controller.r1[6] ),
    .C(\top.controller.r1[5] ),
    .D(\top.controller.r1[4] ),
    .Y(_0905_));
 sg13g2_a22oi_1 _1854_ (.Y(_0906_),
    .B1(_0904_),
    .B2(_0905_),
    .A2(_0903_),
    .A1(_0902_));
 sg13g2_nand2_1 _1855_ (.Y(_0907_),
    .A(net166),
    .B(_0906_));
 sg13g2_or2_1 _1856_ (.X(_0908_),
    .B(_0907_),
    .A(_0087_));
 sg13g2_nand2_1 _1857_ (.Y(_0909_),
    .A(net97),
    .B(net139));
 sg13g2_o21ai_1 _1858_ (.B1(_0909_),
    .Y(_0022_),
    .A1(_0078_),
    .A2(net139));
 sg13g2_nand2_1 _1859_ (.Y(_0910_),
    .A(net157),
    .B(net141));
 sg13g2_o21ai_1 _1860_ (.B1(_0910_),
    .Y(_0023_),
    .A1(_0077_),
    .A2(net141));
 sg13g2_nand2_1 _1861_ (.Y(_0911_),
    .A(net156),
    .B(net139));
 sg13g2_o21ai_1 _1862_ (.B1(_0911_),
    .Y(_0024_),
    .A1(_0076_),
    .A2(net139));
 sg13g2_nor2_1 _1863_ (.A(net85),
    .B(net139),
    .Y(_0912_));
 sg13g2_a21oi_1 _1864_ (.A1(_0082_),
    .A2(net139),
    .Y(_0025_),
    .B1(_0912_));
 sg13g2_nand2_1 _1865_ (.Y(_0913_),
    .A(net153),
    .B(net138));
 sg13g2_o21ai_1 _1866_ (.B1(_0913_),
    .Y(_0026_),
    .A1(_0074_),
    .A2(net138));
 sg13g2_nor2_1 _1867_ (.A(net72),
    .B(net138),
    .Y(_0914_));
 sg13g2_a21oi_1 _1868_ (.A1(_0083_),
    .A2(net138),
    .Y(_0027_),
    .B1(_0914_));
 sg13g2_nand2_1 _1869_ (.Y(_0915_),
    .A(net84),
    .B(net138));
 sg13g2_o21ai_1 _1870_ (.B1(_0915_),
    .Y(_0028_),
    .A1(_0072_),
    .A2(net138));
 sg13g2_nand2_1 _1871_ (.Y(_0916_),
    .A(net93),
    .B(net138));
 sg13g2_o21ai_1 _1872_ (.B1(_0916_),
    .Y(_0029_),
    .A1(_0071_),
    .A2(net138));
 sg13g2_o21ai_1 _1873_ (.B1(net164),
    .Y(_0917_),
    .A1(net163),
    .A2(net1));
 sg13g2_a21oi_1 _1874_ (.A1(net162),
    .A2(_0078_),
    .Y(_0030_),
    .B1(_0917_));
 sg13g2_o21ai_1 _1875_ (.B1(net164),
    .Y(_0918_),
    .A1(net161),
    .A2(net2));
 sg13g2_a21oi_1 _1876_ (.A1(net163),
    .A2(_0077_),
    .Y(_0031_),
    .B1(_0918_));
 sg13g2_o21ai_1 _1877_ (.B1(net164),
    .Y(_0919_),
    .A1(net161),
    .A2(net3));
 sg13g2_a21oi_1 _1878_ (.A1(net161),
    .A2(_0076_),
    .Y(_0032_),
    .B1(_0919_));
 sg13g2_o21ai_1 _1879_ (.B1(net164),
    .Y(_0920_),
    .A1(net161),
    .A2(net4));
 sg13g2_a21oi_1 _1880_ (.A1(net163),
    .A2(_0075_),
    .Y(_0033_),
    .B1(_0920_));
 sg13g2_o21ai_1 _1881_ (.B1(net165),
    .Y(_0921_),
    .A1(net159),
    .A2(net5));
 sg13g2_a21oi_1 _1882_ (.A1(net159),
    .A2(_0074_),
    .Y(_0034_),
    .B1(_0921_));
 sg13g2_o21ai_1 _1883_ (.B1(net165),
    .Y(_0922_),
    .A1(net159),
    .A2(net6));
 sg13g2_a21oi_1 _1884_ (.A1(net159),
    .A2(_0073_),
    .Y(_0035_),
    .B1(_0922_));
 sg13g2_o21ai_1 _1885_ (.B1(net166),
    .Y(_0923_),
    .A1(net159),
    .A2(net7));
 sg13g2_a21oi_1 _1886_ (.A1(net159),
    .A2(_0072_),
    .Y(_0036_),
    .B1(_0923_));
 sg13g2_o21ai_1 _1887_ (.B1(net166),
    .Y(_0924_),
    .A1(net8),
    .A2(net159));
 sg13g2_a21oi_1 _1888_ (.A1(net159),
    .A2(_0071_),
    .Y(_0037_),
    .B1(_0924_));
 sg13g2_o21ai_1 _1889_ (.B1(net165),
    .Y(_0925_),
    .A1(net162),
    .A2(net82));
 sg13g2_a21oi_1 _1890_ (.A1(net162),
    .A2(_0070_),
    .Y(_0038_),
    .B1(_0925_));
 sg13g2_o21ai_1 _1891_ (.B1(net164),
    .Y(_0926_),
    .A1(net163),
    .A2(net77));
 sg13g2_a21oi_1 _1892_ (.A1(net162),
    .A2(_0069_),
    .Y(_0039_),
    .B1(_0926_));
 sg13g2_o21ai_1 _1893_ (.B1(net164),
    .Y(_0055_),
    .A1(net162),
    .A2(net104));
 sg13g2_a21oi_1 _1894_ (.A1(net162),
    .A2(_0068_),
    .Y(_0040_),
    .B1(_0055_));
 sg13g2_o21ai_1 _1895_ (.B1(net164),
    .Y(_0056_),
    .A1(net162),
    .A2(net89));
 sg13g2_a21oi_1 _1896_ (.A1(net162),
    .A2(_0067_),
    .Y(_0041_),
    .B1(_0056_));
 sg13g2_o21ai_1 _1897_ (.B1(net164),
    .Y(_0057_),
    .A1(net161),
    .A2(net108));
 sg13g2_a21oi_1 _1898_ (.A1(net161),
    .A2(_0066_),
    .Y(_0042_),
    .B1(_0057_));
 sg13g2_o21ai_1 _1899_ (.B1(net165),
    .Y(_0058_),
    .A1(net161),
    .A2(net86));
 sg13g2_a21oi_1 _1900_ (.A1(net161),
    .A2(_0065_),
    .Y(_0043_),
    .B1(_0058_));
 sg13g2_o21ai_1 _1901_ (.B1(net165),
    .Y(_0059_),
    .A1(net160),
    .A2(net112));
 sg13g2_a21oi_1 _1902_ (.A1(net160),
    .A2(_0064_),
    .Y(_0044_),
    .B1(_0059_));
 sg13g2_o21ai_1 _1903_ (.B1(net165),
    .Y(_0060_),
    .A1(net102),
    .A2(net160));
 sg13g2_a21oi_1 _1904_ (.A1(_0063_),
    .A2(net160),
    .Y(_0045_),
    .B1(_0060_));
 sg13g2_mux2_1 _1905_ (.A0(net82),
    .A1(\top.controller.s2[0] ),
    .S(net140),
    .X(_0046_));
 sg13g2_mux2_1 _1906_ (.A0(net77),
    .A1(\top.controller.s2[1] ),
    .S(net141),
    .X(_0047_));
 sg13g2_nor2_1 _1907_ (.A(net104),
    .B(net139),
    .Y(_0061_));
 sg13g2_a21oi_1 _1908_ (.A1(_0085_),
    .A2(net140),
    .Y(_0048_),
    .B1(_0061_));
 sg13g2_mux2_1 _1909_ (.A0(net89),
    .A1(net149),
    .S(net140),
    .X(_0049_));
 sg13g2_nor2_1 _1910_ (.A(net108),
    .B(net139),
    .Y(_0062_));
 sg13g2_a21oi_1 _1911_ (.A1(_0086_),
    .A2(net140),
    .Y(_0050_),
    .B1(_0062_));
 sg13g2_mux2_1 _1912_ (.A0(net86),
    .A1(net146),
    .S(net140),
    .X(_0051_));
 sg13g2_mux2_1 _1913_ (.A0(net112),
    .A1(net145),
    .S(net140),
    .X(_0052_));
 sg13g2_mux2_1 _1914_ (.A0(net102),
    .A1(\top.controller.s2[7] ),
    .S(net140),
    .X(_0053_));
 sg13g2_a22oi_1 _1915_ (.Y(_0054_),
    .B1(_0907_),
    .B2(net144),
    .A2(_0087_),
    .A1(net166));
 sg13g2_dfrbp_1 _1916_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net61),
    .D(net69),
    .Q_N(_0011_),
    .Q(\top.controller.count[0] ));
 sg13g2_dfrbp_1 _1917_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net54),
    .D(net71),
    .Q_N(_0957_),
    .Q(\top.controller.count[1] ));
 sg13g2_dfrbp_1 _1918_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net53),
    .D(net81),
    .Q_N(_0956_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1919_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(_0015_),
    .Q_N(_0955_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1920_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net49),
    .D(_0016_),
    .Q_N(_0954_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1921_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net47),
    .D(_0017_),
    .Q_N(_0953_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1922_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net45),
    .D(_0018_),
    .Q_N(_0952_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1923_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net43),
    .D(_0019_),
    .Q_N(_0951_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1924_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net41),
    .D(_0020_),
    .Q_N(_0950_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1925_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net39),
    .D(_0021_),
    .Q_N(_0949_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1926_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net37),
    .D(_0022_),
    .Q_N(_0948_),
    .Q(\top.controller.s1[0] ));
 sg13g2_dfrbp_1 _1927_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net36),
    .D(_0023_),
    .Q_N(_0001_),
    .Q(\top.controller.s1[1] ));
 sg13g2_dfrbp_1 _1928_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net35),
    .D(_0024_),
    .Q_N(_0004_),
    .Q(\top.controller.s1[2] ));
 sg13g2_dfrbp_1 _1929_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net34),
    .D(_0025_),
    .Q_N(_0947_),
    .Q(\top.controller.s1[3] ));
 sg13g2_dfrbp_1 _1930_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net33),
    .D(_0026_),
    .Q_N(_0003_),
    .Q(\top.controller.s1[4] ));
 sg13g2_dfrbp_1 _1931_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net32),
    .D(_0027_),
    .Q_N(_0000_),
    .Q(\top.controller.s1[5] ));
 sg13g2_dfrbp_1 _1932_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net31),
    .D(_0028_),
    .Q_N(_0002_),
    .Q(\top.controller.s1[6] ));
 sg13g2_dfrbp_1 _1933_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net30),
    .D(_0029_),
    .Q_N(_0010_),
    .Q(\top.controller.s1[7] ));
 sg13g2_dfrbp_1 _1934_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net29),
    .D(_0030_),
    .Q_N(_0946_),
    .Q(\top.controller.r1[0] ));
 sg13g2_dfrbp_1 _1935_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net27),
    .D(_0031_),
    .Q_N(_0945_),
    .Q(\top.controller.r1[1] ));
 sg13g2_dfrbp_1 _1936_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net25),
    .D(_0032_),
    .Q_N(_0944_),
    .Q(\top.controller.r1[2] ));
 sg13g2_dfrbp_1 _1937_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net66),
    .D(_0033_),
    .Q_N(_0943_),
    .Q(\top.controller.r1[3] ));
 sg13g2_dfrbp_1 _1938_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net64),
    .D(_0034_),
    .Q_N(_0942_),
    .Q(\top.controller.r1[4] ));
 sg13g2_dfrbp_1 _1939_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net62),
    .D(_0035_),
    .Q_N(_0941_),
    .Q(\top.controller.r1[5] ));
 sg13g2_dfrbp_1 _1940_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net60),
    .D(_0036_),
    .Q_N(_0940_),
    .Q(\top.controller.r1[6] ));
 sg13g2_dfrbp_1 _1941_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net58),
    .D(_0037_),
    .Q_N(_0939_),
    .Q(\top.controller.r1[7] ));
 sg13g2_dfrbp_1 _1942_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net56),
    .D(_0038_),
    .Q_N(_0938_),
    .Q(\top.controller.r2[0] ));
 sg13g2_dfrbp_1 _1943_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net52),
    .D(_0039_),
    .Q_N(_0937_),
    .Q(\top.controller.r2[1] ));
 sg13g2_dfrbp_1 _1944_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net48),
    .D(_0040_),
    .Q_N(_0936_),
    .Q(\top.controller.r2[2] ));
 sg13g2_dfrbp_1 _1945_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net44),
    .D(_0041_),
    .Q_N(_0935_),
    .Q(\top.controller.r2[3] ));
 sg13g2_dfrbp_1 _1946_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net40),
    .D(_0042_),
    .Q_N(_0934_),
    .Q(\top.controller.r2[4] ));
 sg13g2_dfrbp_1 _1947_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net28),
    .D(_0043_),
    .Q_N(_0933_),
    .Q(\top.controller.r2[5] ));
 sg13g2_dfrbp_1 _1948_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net67),
    .D(_0044_),
    .Q_N(_0932_),
    .Q(\top.controller.r2[6] ));
 sg13g2_dfrbp_1 _1949_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net63),
    .D(_0045_),
    .Q_N(_0931_),
    .Q(\top.controller.r2[7] ));
 sg13g2_dfrbp_1 _1950_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net59),
    .D(net83),
    .Q_N(_0930_),
    .Q(\top.controller.s2[0] ));
 sg13g2_dfrbp_1 _1951_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net57),
    .D(net78),
    .Q_N(_0929_),
    .Q(\top.controller.s2[1] ));
 sg13g2_dfrbp_1 _1952_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net55),
    .D(_0048_),
    .Q_N(_0009_),
    .Q(\top.controller.s2[2] ));
 sg13g2_dfrbp_1 _1953_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net50),
    .D(net90),
    .Q_N(_0928_),
    .Q(\top.controller.s2[3] ));
 sg13g2_dfrbp_1 _1954_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net46),
    .D(_0050_),
    .Q_N(_0008_),
    .Q(\top.controller.s2[4] ));
 sg13g2_dfrbp_1 _1955_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net42),
    .D(net87),
    .Q_N(_0006_),
    .Q(\top.controller.s2[5] ));
 sg13g2_dfrbp_1 _1956_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net38),
    .D(net113),
    .Q_N(_0007_),
    .Q(\top.controller.s2[6] ));
 sg13g2_dfrbp_1 _1957_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net26),
    .D(net103),
    .Q_N(_0005_),
    .Q(\top.controller.s2[7] ));
 sg13g2_dfrbp_1 _1958_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net65),
    .D(net99),
    .Q_N(_0927_),
    .Q(\top.controller.ef1 ));
 sg13g2_tiehi _1957__26 (.L_HI(net26));
 sg13g2_tiehi _1935__27 (.L_HI(net27));
 sg13g2_tiehi _1947__28 (.L_HI(net28));
 sg13g2_tiehi _1934__29 (.L_HI(net29));
 sg13g2_tiehi _1933__30 (.L_HI(net30));
 sg13g2_tiehi _1932__31 (.L_HI(net31));
 sg13g2_tiehi _1931__32 (.L_HI(net32));
 sg13g2_tiehi _1930__33 (.L_HI(net33));
 sg13g2_tiehi _1929__34 (.L_HI(net34));
 sg13g2_tiehi _1928__35 (.L_HI(net35));
 sg13g2_tiehi _1927__36 (.L_HI(net36));
 sg13g2_tiehi _1926__37 (.L_HI(net37));
 sg13g2_tiehi _1956__38 (.L_HI(net38));
 sg13g2_tiehi _1925__39 (.L_HI(net39));
 sg13g2_tiehi _1946__40 (.L_HI(net40));
 sg13g2_tiehi _1924__41 (.L_HI(net41));
 sg13g2_tiehi _1955__42 (.L_HI(net42));
 sg13g2_tiehi _1923__43 (.L_HI(net43));
 sg13g2_tiehi _1945__44 (.L_HI(net44));
 sg13g2_tiehi _1922__45 (.L_HI(net45));
 sg13g2_tiehi _1954__46 (.L_HI(net46));
 sg13g2_tiehi _1921__47 (.L_HI(net47));
 sg13g2_tiehi _1944__48 (.L_HI(net48));
 sg13g2_tiehi _1920__49 (.L_HI(net49));
 sg13g2_tiehi _1953__50 (.L_HI(net50));
 sg13g2_tiehi _1919__51 (.L_HI(net51));
 sg13g2_tiehi _1943__52 (.L_HI(net52));
 sg13g2_tiehi _1918__53 (.L_HI(net53));
 sg13g2_tiehi _1917__54 (.L_HI(net54));
 sg13g2_tiehi _1952__55 (.L_HI(net55));
 sg13g2_tiehi _1942__56 (.L_HI(net56));
 sg13g2_tiehi _1951__57 (.L_HI(net57));
 sg13g2_tiehi _1941__58 (.L_HI(net58));
 sg13g2_tiehi _1950__59 (.L_HI(net59));
 sg13g2_tiehi _1940__60 (.L_HI(net60));
 sg13g2_tiehi _1916__61 (.L_HI(net61));
 sg13g2_tiehi _1939__62 (.L_HI(net62));
 sg13g2_tiehi _1949__63 (.L_HI(net63));
 sg13g2_tiehi _1938__64 (.L_HI(net64));
 sg13g2_tiehi _1958__65 (.L_HI(net65));
 sg13g2_tiehi _1937__66 (.L_HI(net66));
 sg13g2_tiehi _1948__67 (.L_HI(net67));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_resfuzzy_10 (.L_LO(net10));
 sg13g2_tielo tt_um_resfuzzy_11 (.L_LO(net11));
 sg13g2_tielo tt_um_resfuzzy_12 (.L_LO(net12));
 sg13g2_tielo tt_um_resfuzzy_13 (.L_LO(net13));
 sg13g2_tielo tt_um_resfuzzy_14 (.L_LO(net14));
 sg13g2_tielo tt_um_resfuzzy_15 (.L_LO(net15));
 sg13g2_tielo tt_um_resfuzzy_16 (.L_LO(net16));
 sg13g2_tielo tt_um_resfuzzy_17 (.L_LO(net17));
 sg13g2_tielo tt_um_resfuzzy_18 (.L_LO(net18));
 sg13g2_tielo tt_um_resfuzzy_19 (.L_LO(net19));
 sg13g2_tielo tt_um_resfuzzy_20 (.L_LO(net20));
 sg13g2_tielo tt_um_resfuzzy_21 (.L_LO(net21));
 sg13g2_tielo tt_um_resfuzzy_22 (.L_LO(net22));
 sg13g2_tielo tt_um_resfuzzy_23 (.L_LO(net23));
 sg13g2_tielo tt_um_resfuzzy_24 (.L_LO(net24));
 sg13g2_tiehi _1936__25 (.L_HI(net25));
 sg13g2_buf_2 fanout128 (.A(_0572_),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(_0645_));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_0581_));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(_0580_));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(_0626_));
 sg13g2_buf_1 fanout133 (.A(_0626_),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net135));
 sg13g2_buf_2 fanout135 (.A(_0467_),
    .X(net135));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(_0433_));
 sg13g2_buf_2 fanout137 (.A(_0397_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net141),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(net141));
 sg13g2_buf_2 fanout141 (.A(_0908_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_0108_),
    .X(net142));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(_0104_));
 sg13g2_buf_2 fanout144 (.A(_0079_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(\top.controller.s2[6] ),
    .X(net145));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(\top.controller.s2[5] ));
 sg13g2_buf_2 fanout147 (.A(\top.controller.s2[4] ),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net149));
 sg13g2_buf_2 fanout149 (.A(\top.controller.s2[3] ),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(net120),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(\top.controller.s1[5] ),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net75),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(\top.controller.s1[3] ),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(\top.controller.s1[2] ),
    .X(net155));
 sg13g2_buf_1 fanout156 (.A(net96),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(net111),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_0081_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(uio_in[0]),
    .X(net159));
 sg13g2_buf_1 fanout160 (.A(uio_in[0]),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(net163),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(net163),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(uio_in[0]),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net165),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(rst_n),
    .X(net166));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_resfuzzy_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0011_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0012_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold3 (.A(\top.controller.count[0] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0013_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold5 (.A(\top.controller.r1[5] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold6 (.A(\top.controller.r1[4] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold7 (.A(\top.controller.s1[5] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold8 (.A(\top.controller.s1[4] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold9 (.A(\top.controller.r1[7] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold10 (.A(\top.controller.r2[1] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0047_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold12 (.A(\top.controller.r1[6] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold13 (.A(uo_out[0]),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0014_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold15 (.A(\top.controller.r2[0] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0046_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold17 (.A(\top.controller.s1[6] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold18 (.A(\top.controller.r1[3] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold19 (.A(\top.controller.r2[5] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0051_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold21 (.A(\top.controller.r1[2] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold22 (.A(\top.controller.r2[3] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0049_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold24 (.A(\top.controller.s1[3] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold25 (.A(\top.controller.r1[0] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold26 (.A(\top.controller.s1[7] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold27 (.A(uo_out[7]),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0901_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold29 (.A(\top.controller.s1[2] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold30 (.A(\top.controller.s1[0] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold31 (.A(\top.controller.count[1] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0054_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold33 (.A(uo_out[2]),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0893_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold35 (.A(\top.controller.r2[7] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0053_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold37 (.A(\top.controller.r2[2] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold38 (.A(uo_out[4]),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0896_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold40 (.A(\top.controller.r1[1] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold41 (.A(\top.controller.r2[4] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold42 (.A(uo_out[3]),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0894_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold44 (.A(\top.controller.s1[1] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold45 (.A(\top.controller.r2[6] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0052_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold47 (.A(uo_out[5]),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0898_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold49 (.A(uo_out[1]),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0891_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold51 (.A(uo_out[6]),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0899_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold53 (.A(\top.controller.s2[2] ),
    .X(net120));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_70 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_decap_8 FILLER_13_78 ();
 sg13g2_decap_8 FILLER_13_85 ();
 sg13g2_decap_8 FILLER_13_92 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_decap_4 FILLER_13_116 ();
 sg13g2_fill_1 FILLER_13_120 ();
 sg13g2_decap_8 FILLER_13_125 ();
 sg13g2_decap_8 FILLER_13_132 ();
 sg13g2_fill_2 FILLER_13_139 ();
 sg13g2_fill_2 FILLER_13_145 ();
 sg13g2_fill_1 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_fill_2 FILLER_14_63 ();
 sg13g2_decap_4 FILLER_14_86 ();
 sg13g2_fill_1 FILLER_14_111 ();
 sg13g2_decap_4 FILLER_14_132 ();
 sg13g2_decap_4 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_decap_8 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_decap_8 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_fill_2 FILLER_14_271 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_4 FILLER_14_328 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_decap_4 FILLER_14_356 ();
 sg13g2_fill_2 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_35 ();
 sg13g2_fill_2 FILLER_15_49 ();
 sg13g2_fill_1 FILLER_15_51 ();
 sg13g2_decap_4 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_111 ();
 sg13g2_fill_2 FILLER_15_118 ();
 sg13g2_fill_1 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_125 ();
 sg13g2_decap_8 FILLER_15_132 ();
 sg13g2_fill_2 FILLER_15_149 ();
 sg13g2_fill_2 FILLER_15_157 ();
 sg13g2_fill_1 FILLER_15_168 ();
 sg13g2_decap_4 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_194 ();
 sg13g2_decap_8 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_208 ();
 sg13g2_decap_4 FILLER_15_215 ();
 sg13g2_fill_2 FILLER_15_219 ();
 sg13g2_decap_4 FILLER_15_230 ();
 sg13g2_fill_1 FILLER_15_234 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_314 ();
 sg13g2_fill_2 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_decap_4 FILLER_15_347 ();
 sg13g2_fill_2 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_50 ();
 sg13g2_fill_1 FILLER_16_57 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_decap_8 FILLER_16_75 ();
 sg13g2_fill_2 FILLER_16_82 ();
 sg13g2_decap_4 FILLER_16_97 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_fill_1 FILLER_16_131 ();
 sg13g2_fill_1 FILLER_16_151 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_fill_2 FILLER_16_179 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_299 ();
 sg13g2_decap_4 FILLER_16_306 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_333 ();
 sg13g2_fill_1 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_fill_2 FILLER_16_360 ();
 sg13g2_fill_2 FILLER_16_367 ();
 sg13g2_fill_2 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_51 ();
 sg13g2_decap_8 FILLER_17_78 ();
 sg13g2_decap_8 FILLER_17_85 ();
 sg13g2_decap_4 FILLER_17_92 ();
 sg13g2_fill_1 FILLER_17_109 ();
 sg13g2_decap_8 FILLER_17_141 ();
 sg13g2_fill_2 FILLER_17_148 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_fill_1 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_fill_2 FILLER_17_270 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_323 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_fill_2 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_45 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_58 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_113 ();
 sg13g2_fill_2 FILLER_18_120 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_fill_2 FILLER_18_151 ();
 sg13g2_fill_1 FILLER_18_153 ();
 sg13g2_decap_8 FILLER_18_169 ();
 sg13g2_decap_4 FILLER_18_176 ();
 sg13g2_fill_2 FILLER_18_180 ();
 sg13g2_decap_8 FILLER_18_191 ();
 sg13g2_decap_4 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_257 ();
 sg13g2_fill_1 FILLER_18_259 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_fill_2 FILLER_18_280 ();
 sg13g2_decap_4 FILLER_18_304 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_314 ();
 sg13g2_decap_4 FILLER_18_321 ();
 sg13g2_fill_1 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_fill_1 FILLER_18_363 ();
 sg13g2_decap_4 FILLER_18_374 ();
 sg13g2_fill_2 FILLER_18_394 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_16 ();
 sg13g2_fill_2 FILLER_19_23 ();
 sg13g2_decap_8 FILLER_19_33 ();
 sg13g2_fill_2 FILLER_19_40 ();
 sg13g2_fill_1 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_55 ();
 sg13g2_fill_1 FILLER_19_59 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_70 ();
 sg13g2_decap_4 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_89 ();
 sg13g2_decap_4 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_decap_4 FILLER_19_162 ();
 sg13g2_fill_1 FILLER_19_166 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_fill_2 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_219 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_decap_4 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_281 ();
 sg13g2_decap_4 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_296 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_fill_2 FILLER_19_383 ();
 sg13g2_fill_1 FILLER_19_385 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_4 ();
 sg13g2_fill_2 FILLER_20_36 ();
 sg13g2_fill_1 FILLER_20_38 ();
 sg13g2_fill_1 FILLER_20_64 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_143 ();
 sg13g2_fill_1 FILLER_20_150 ();
 sg13g2_decap_4 FILLER_20_163 ();
 sg13g2_fill_2 FILLER_20_177 ();
 sg13g2_decap_8 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_220 ();
 sg13g2_decap_8 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_244 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_262 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_fill_1 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_fill_2 FILLER_20_325 ();
 sg13g2_fill_1 FILLER_20_327 ();
 sg13g2_decap_4 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_fill_2 FILLER_20_354 ();
 sg13g2_fill_1 FILLER_20_356 ();
 sg13g2_decap_4 FILLER_20_374 ();
 sg13g2_fill_1 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_22 ();
 sg13g2_decap_4 FILLER_21_29 ();
 sg13g2_fill_1 FILLER_21_33 ();
 sg13g2_fill_2 FILLER_21_64 ();
 sg13g2_fill_2 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_fill_2 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_decap_4 FILLER_21_113 ();
 sg13g2_fill_1 FILLER_21_117 ();
 sg13g2_decap_8 FILLER_21_134 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_decap_4 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_227 ();
 sg13g2_fill_2 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_282 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_358 ();
 sg13g2_fill_1 FILLER_21_360 ();
 sg13g2_decap_4 FILLER_21_366 ();
 sg13g2_decap_4 FILLER_21_377 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_22 ();
 sg13g2_fill_1 FILLER_22_34 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_decap_8 FILLER_22_75 ();
 sg13g2_decap_4 FILLER_22_82 ();
 sg13g2_fill_2 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_decap_4 FILLER_22_136 ();
 sg13g2_fill_2 FILLER_22_166 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_decap_4 FILLER_22_189 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_decap_4 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_233 ();
 sg13g2_fill_1 FILLER_22_235 ();
 sg13g2_decap_4 FILLER_22_256 ();
 sg13g2_fill_2 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_276 ();
 sg13g2_decap_8 FILLER_22_283 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_decap_4 FILLER_22_317 ();
 sg13g2_decap_4 FILLER_22_332 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_4 FILLER_22_381 ();
 sg13g2_fill_2 FILLER_22_401 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_23 ();
 sg13g2_fill_1 FILLER_23_30 ();
 sg13g2_fill_2 FILLER_23_39 ();
 sg13g2_fill_1 FILLER_23_41 ();
 sg13g2_decap_8 FILLER_23_50 ();
 sg13g2_decap_8 FILLER_23_57 ();
 sg13g2_decap_8 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_94 ();
 sg13g2_fill_1 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_decap_4 FILLER_23_117 ();
 sg13g2_fill_1 FILLER_23_121 ();
 sg13g2_fill_2 FILLER_23_125 ();
 sg13g2_fill_1 FILLER_23_127 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_4 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_decap_4 FILLER_23_151 ();
 sg13g2_fill_2 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_277 ();
 sg13g2_fill_2 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_decap_8 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_4 FILLER_23_341 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_351 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_decap_4 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_30 ();
 sg13g2_decap_8 FILLER_24_44 ();
 sg13g2_decap_4 FILLER_24_51 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_fill_1 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_104 ();
 sg13g2_fill_1 FILLER_24_106 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_decap_4 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_160 ();
 sg13g2_fill_2 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_169 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_234 ();
 sg13g2_fill_2 FILLER_24_241 ();
 sg13g2_decap_8 FILLER_24_248 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_9 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_fill_2 FILLER_25_32 ();
 sg13g2_fill_2 FILLER_25_55 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_79 ();
 sg13g2_decap_4 FILLER_25_86 ();
 sg13g2_fill_1 FILLER_25_90 ();
 sg13g2_decap_8 FILLER_25_99 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_decap_8 FILLER_25_120 ();
 sg13g2_fill_2 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_139 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_decap_4 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_231 ();
 sg13g2_decap_4 FILLER_25_240 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_fill_2 FILLER_25_254 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_fill_2 FILLER_25_265 ();
 sg13g2_decap_4 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_decap_4 FILLER_25_312 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_decap_4 FILLER_25_376 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_30 ();
 sg13g2_decap_4 FILLER_26_52 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_4 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_225 ();
 sg13g2_decap_4 FILLER_26_241 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_4 FILLER_26_287 ();
 sg13g2_fill_2 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_310 ();
 sg13g2_fill_2 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_367 ();
 sg13g2_decap_4 FILLER_26_379 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_16 ();
 sg13g2_fill_1 FILLER_27_26 ();
 sg13g2_fill_2 FILLER_27_30 ();
 sg13g2_fill_1 FILLER_27_32 ();
 sg13g2_decap_4 FILLER_27_47 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_decap_8 FILLER_27_60 ();
 sg13g2_fill_1 FILLER_27_67 ();
 sg13g2_decap_4 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_110 ();
 sg13g2_decap_8 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_4 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_2 FILLER_27_156 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_decap_8 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_2 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_241 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_fill_2 FILLER_27_285 ();
 sg13g2_decap_4 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_314 ();
 sg13g2_fill_2 FILLER_27_335 ();
 sg13g2_fill_2 FILLER_27_356 ();
 sg13g2_fill_2 FILLER_27_388 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_38 ();
 sg13g2_fill_1 FILLER_28_40 ();
 sg13g2_decap_8 FILLER_28_54 ();
 sg13g2_decap_4 FILLER_28_61 ();
 sg13g2_fill_2 FILLER_28_65 ();
 sg13g2_decap_4 FILLER_28_78 ();
 sg13g2_fill_2 FILLER_28_82 ();
 sg13g2_fill_1 FILLER_28_89 ();
 sg13g2_decap_4 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_118 ();
 sg13g2_decap_4 FILLER_28_125 ();
 sg13g2_decap_4 FILLER_28_134 ();
 sg13g2_fill_2 FILLER_28_138 ();
 sg13g2_decap_8 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_4 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_209 ();
 sg13g2_decap_4 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_236 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_decap_8 FILLER_28_284 ();
 sg13g2_decap_4 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_decap_4 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_4 ();
 sg13g2_fill_2 FILLER_29_23 ();
 sg13g2_fill_2 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_37 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_195 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_decap_8 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_fill_2 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_fill_1 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_27 ();
 sg13g2_fill_1 FILLER_30_29 ();
 sg13g2_fill_2 FILLER_30_46 ();
 sg13g2_decap_8 FILLER_30_57 ();
 sg13g2_decap_4 FILLER_30_81 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_decap_8 FILLER_30_94 ();
 sg13g2_fill_2 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_decap_4 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_decap_4 FILLER_30_178 ();
 sg13g2_decap_8 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_fill_2 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_fill_2 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_282 ();
 sg13g2_decap_4 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_293 ();
 sg13g2_fill_1 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_45 ();
 sg13g2_decap_4 FILLER_31_52 ();
 sg13g2_fill_1 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_4 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_decap_4 FILLER_31_250 ();
 sg13g2_decap_4 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_fill_1 FILLER_31_335 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_18 ();
 sg13g2_fill_2 FILLER_32_31 ();
 sg13g2_fill_1 FILLER_32_33 ();
 sg13g2_fill_2 FILLER_32_60 ();
 sg13g2_fill_1 FILLER_32_62 ();
 sg13g2_fill_2 FILLER_32_78 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_fill_2 FILLER_32_134 ();
 sg13g2_fill_2 FILLER_32_158 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_decap_4 FILLER_32_181 ();
 sg13g2_fill_1 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_196 ();
 sg13g2_decap_4 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_209 ();
 sg13g2_decap_4 FILLER_32_246 ();
 sg13g2_fill_2 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_2 FILLER_32_322 ();
 sg13g2_fill_1 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_2 FILLER_33_25 ();
 sg13g2_fill_2 FILLER_33_32 ();
 sg13g2_fill_1 FILLER_33_34 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_fill_2 FILLER_33_102 ();
 sg13g2_fill_1 FILLER_33_104 ();
 sg13g2_decap_4 FILLER_33_122 ();
 sg13g2_fill_1 FILLER_33_126 ();
 sg13g2_decap_4 FILLER_33_136 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_170 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_decap_8 FILLER_33_278 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_decap_4 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_30 ();
 sg13g2_decap_4 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_decap_8 FILLER_34_44 ();
 sg13g2_fill_2 FILLER_34_83 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_decap_8 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_269 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_372 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_4 FILLER_35_42 ();
 sg13g2_fill_1 FILLER_35_46 ();
 sg13g2_fill_2 FILLER_35_64 ();
 sg13g2_fill_2 FILLER_35_80 ();
 sg13g2_fill_2 FILLER_35_134 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_fill_1 FILLER_35_159 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_194 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_4 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_39 ();
 sg13g2_fill_2 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_69 ();
 sg13g2_decap_8 FILLER_36_83 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_142 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_236 ();
 sg13g2_fill_1 FILLER_36_240 ();
 sg13g2_fill_2 FILLER_36_251 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_fill_1 FILLER_36_258 ();
 sg13g2_decap_4 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_285 ();
 sg13g2_decap_4 FILLER_36_297 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_71 ();
 sg13g2_decap_8 FILLER_37_76 ();
 sg13g2_decap_8 FILLER_37_83 ();
 sg13g2_decap_8 FILLER_37_90 ();
 sg13g2_decap_8 FILLER_37_97 ();
 sg13g2_decap_4 FILLER_37_104 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_decap_8 FILLER_37_113 ();
 sg13g2_decap_8 FILLER_37_124 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_decap_8 FILLER_37_143 ();
 sg13g2_decap_4 FILLER_37_150 ();
 sg13g2_decap_8 FILLER_37_167 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_decap_4 FILLER_37_188 ();
 sg13g2_fill_2 FILLER_37_222 ();
 sg13g2_decap_4 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_fill_2 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_214 ();
 sg13g2_fill_1 FILLER_38_218 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_decap_4 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_283 ();
 sg13g2_fill_2 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

module tt_um_nyan (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire \gfx.bitmap_x[0] ;
 wire \gfx.bitmap_x[1] ;
 wire \gfx.bitmap_x[2] ;
 wire \gfx.bitmap_x[3] ;
 wire \gfx.bitmap_y[0] ;
 wire \gfx.bitmap_y[1] ;
 wire \gfx.bitmap_y[2] ;
 wire \gfx.bitmap_y[3] ;
 wire \gfx.frame_counter[0] ;
 wire \gfx.frame_counter[1] ;
 wire \gfx.frame_counter[2] ;
 wire \gfx.frame_counter[3] ;
 wire \gfx.frame_counter[4] ;
 wire \gfx.hsync ;
 wire \gfx.pixel_x[0] ;
 wire \gfx.pixel_x[1] ;
 wire \gfx.pixel_x[2] ;
 wire \gfx.pixel_x[7] ;
 wire \gfx.pixel_x[8] ;
 wire \gfx.pixel_x[9] ;
 wire \gfx.pixel_y[0] ;
 wire \gfx.pixel_y[1] ;
 wire \gfx.pixel_y[2] ;
 wire \gfx.pixel_y[7] ;
 wire \gfx.pixel_y[8] ;
 wire \gfx.pixel_y[9] ;
 wire \gfx.vsync ;
 wire \music.do_note ;
 wire \music.extended_sample[0] ;
 wire \music.extended_sample[10] ;
 wire \music.extended_sample[11] ;
 wire \music.extended_sample[12] ;
 wire \music.extended_sample[13] ;
 wire \music.extended_sample[14] ;
 wire \music.extended_sample[1] ;
 wire \music.extended_sample[2] ;
 wire \music.extended_sample[3] ;
 wire \music.extended_sample[4] ;
 wire \music.extended_sample[5] ;
 wire \music.extended_sample[6] ;
 wire \music.extended_sample[7] ;
 wire \music.extended_sample[8] ;
 wire \music.extended_sample[9] ;
 wire \music.melody_pos[0] ;
 wire \music.melody_pos[1] ;
 wire \music.melody_pos[2] ;
 wire \music.melody_pos[3] ;
 wire \music.melody_pos[4] ;
 wire \music.note[0] ;
 wire \music.note[1] ;
 wire \music.note[2] ;
 wire \music.note_length ;
 wire \music.note_pos[0] ;
 wire \music.note_pos[10] ;
 wire \music.note_pos[11] ;
 wire \music.note_pos[12] ;
 wire \music.note_pos[13] ;
 wire \music.note_pos[14] ;
 wire \music.note_pos[15] ;
 wire \music.note_pos[1] ;
 wire \music.note_pos[2] ;
 wire \music.note_pos[3] ;
 wire \music.note_pos[4] ;
 wire \music.note_pos[5] ;
 wire \music.note_pos[6] ;
 wire \music.note_pos[7] ;
 wire \music.note_pos[8] ;
 wire \music.note_pos[9] ;
 wire \music.pwm ;
 wire \music.pwm_pos[0] ;
 wire \music.pwm_pos[10] ;
 wire \music.pwm_pos[11] ;
 wire \music.pwm_pos[12] ;
 wire \music.pwm_pos[13] ;
 wire \music.pwm_pos[14] ;
 wire \music.pwm_pos[1] ;
 wire \music.pwm_pos[2] ;
 wire \music.pwm_pos[3] ;
 wire \music.pwm_pos[4] ;
 wire \music.pwm_pos[5] ;
 wire \music.pwm_pos[6] ;
 wire \music.pwm_pos[7] ;
 wire \music.pwm_pos[8] ;
 wire \music.pwm_pos[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net1;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;

 sg13g2_inv_1 _1454_ (.Y(_0513_),
    .A(net215));
 sg13g2_inv_1 _1455_ (.Y(_0514_),
    .A(net151));
 sg13g2_inv_1 _1456_ (.Y(_0515_),
    .A(net238));
 sg13g2_inv_1 _1457_ (.Y(_0516_),
    .A(\music.note_pos[5] ));
 sg13g2_inv_1 _1458_ (.Y(_0517_),
    .A(\music.pwm_pos[3] ));
 sg13g2_inv_1 _1459_ (.Y(_0518_),
    .A(\music.pwm_pos[2] ));
 sg13g2_inv_1 _1460_ (.Y(_0519_),
    .A(\music.pwm_pos[5] ));
 sg13g2_inv_1 _1461_ (.Y(_0520_),
    .A(\music.pwm_pos[6] ));
 sg13g2_inv_1 _1462_ (.Y(_0521_),
    .A(net587));
 sg13g2_inv_1 _1463_ (.Y(_0522_),
    .A(net117));
 sg13g2_inv_1 _1464_ (.Y(_0523_),
    .A(net574));
 sg13g2_inv_1 _1465_ (.Y(_0524_),
    .A(net567));
 sg13g2_inv_1 _1466_ (.Y(_0525_),
    .A(net577));
 sg13g2_inv_1 _1467_ (.Y(_0526_),
    .A(net226));
 sg13g2_inv_1 _1468_ (.Y(_0527_),
    .A(\music.extended_sample[10] ));
 sg13g2_inv_1 _1469_ (.Y(_0528_),
    .A(net208));
 sg13g2_inv_1 _1470_ (.Y(_0529_),
    .A(net126));
 sg13g2_inv_1 _1471_ (.Y(_0530_),
    .A(net563));
 sg13g2_inv_2 _1472_ (.Y(_0531_),
    .A(_0011_));
 sg13g2_inv_1 _1473_ (.Y(_0532_),
    .A(_0009_));
 sg13g2_inv_1 _1474_ (.Y(_0533_),
    .A(net110));
 sg13g2_inv_1 _1475_ (.Y(_0534_),
    .A(\music.note[2] ));
 sg13g2_inv_1 _1476_ (.Y(_0535_),
    .A(net157));
 sg13g2_inv_1 _1477_ (.Y(_0536_),
    .A(\music.extended_sample[5] ));
 sg13g2_inv_1 _1478_ (.Y(_0537_),
    .A(net105));
 sg13g2_inv_1 _1479_ (.Y(_0538_),
    .A(net213));
 sg13g2_inv_1 _1480_ (.Y(_0539_),
    .A(net196));
 sg13g2_inv_1 _1481_ (.Y(_0540_),
    .A(net211));
 sg13g2_o21ai_1 _1482_ (.B1(\music.pwm_pos[0] ),
    .Y(_0541_),
    .A1(\music.pwm_pos[1] ),
    .A2(_0526_));
 sg13g2_a22oi_1 _1483_ (.Y(_0542_),
    .B1(_0527_),
    .B2(\music.pwm_pos[2] ),
    .A2(_0526_),
    .A1(\music.pwm_pos[1] ));
 sg13g2_o21ai_1 _1484_ (.B1(_0542_),
    .Y(_0543_),
    .A1(\music.extended_sample[8] ),
    .A2(_0541_));
 sg13g2_a22oi_1 _1485_ (.Y(_0544_),
    .B1(\music.extended_sample[10] ),
    .B2(_0518_),
    .A2(\music.extended_sample[11] ),
    .A1(_0517_));
 sg13g2_a22oi_1 _1486_ (.Y(_0545_),
    .B1(_0543_),
    .B2(_0544_),
    .A2(_0529_),
    .A1(\music.pwm_pos[4] ));
 sg13g2_o21ai_1 _1487_ (.B1(_0545_),
    .Y(_0546_),
    .A1(_0517_),
    .A2(\music.extended_sample[11] ));
 sg13g2_nand2b_1 _1488_ (.Y(_0547_),
    .B(\music.extended_sample[12] ),
    .A_N(\music.pwm_pos[4] ));
 sg13g2_a22oi_1 _1489_ (.Y(_0548_),
    .B1(_0546_),
    .B2(_0547_),
    .A2(_0528_),
    .A1(\music.pwm_pos[5] ));
 sg13g2_a221oi_1 _1490_ (.B2(_0519_),
    .C1(_0548_),
    .B1(\music.extended_sample[13] ),
    .A1(_0520_),
    .Y(_0549_),
    .A2(\music.extended_sample[14] ));
 sg13g2_nor3_1 _1491_ (.A(\music.pwm_pos[13] ),
    .B(\music.pwm_pos[12] ),
    .C(\music.pwm_pos[14] ),
    .Y(_0550_));
 sg13g2_nor4_1 _1492_ (.A(\music.pwm_pos[9] ),
    .B(\music.pwm_pos[8] ),
    .C(\music.pwm_pos[11] ),
    .D(\music.pwm_pos[10] ),
    .Y(_0551_));
 sg13g2_nand2_2 _1493_ (.Y(_0552_),
    .A(_0550_),
    .B(_0551_));
 sg13g2_nor2_1 _1494_ (.A(_0520_),
    .B(\music.extended_sample[14] ),
    .Y(_0553_));
 sg13g2_nor4_1 _1495_ (.A(\music.pwm_pos[7] ),
    .B(_0549_),
    .C(_0552_),
    .D(_0553_),
    .Y(\music.pwm ));
 sg13g2_nor3_1 _1496_ (.A(\music.pwm_pos[5] ),
    .B(\music.pwm_pos[4] ),
    .C(\music.pwm_pos[6] ),
    .Y(_0554_));
 sg13g2_nand2_1 _1497_ (.Y(_0555_),
    .A(\music.pwm_pos[7] ),
    .B(_0554_));
 sg13g2_or4_1 _1498_ (.A(\music.pwm_pos[1] ),
    .B(\music.pwm_pos[0] ),
    .C(\music.pwm_pos[3] ),
    .D(\music.pwm_pos[2] ),
    .X(_0556_));
 sg13g2_nor3_2 _1499_ (.A(_0552_),
    .B(_0555_),
    .C(_0556_),
    .Y(_0557_));
 sg13g2_nor2b_1 _1500_ (.A(\music.note_pos[13] ),
    .B_N(\music.note_pos[12] ),
    .Y(_0558_));
 sg13g2_nor2_1 _1501_ (.A(\music.note_pos[1] ),
    .B(\music.note_pos[0] ),
    .Y(_0559_));
 sg13g2_nand2_1 _1502_ (.Y(_0560_),
    .A(_0516_),
    .B(\music.note_pos[4] ));
 sg13g2_nand4_1 _1503_ (.B(\music.note_pos[4] ),
    .C(_0558_),
    .A(_0516_),
    .Y(_0561_),
    .D(_0559_));
 sg13g2_nor2_1 _1504_ (.A(\music.note_pos[11] ),
    .B(\music.note_pos[9] ),
    .Y(_0562_));
 sg13g2_nand3_1 _1505_ (.B(\music.note_pos[8] ),
    .C(_0562_),
    .A(\music.note_pos[10] ),
    .Y(_0563_));
 sg13g2_nor4_1 _1506_ (.A(\music.do_note ),
    .B(\music.note_pos[15] ),
    .C(\music.note_pos[14] ),
    .D(\music.note_pos[7] ),
    .Y(_0564_));
 sg13g2_nand4_1 _1507_ (.B(\music.note_pos[3] ),
    .C(\music.note_pos[2] ),
    .A(\music.note_pos[6] ),
    .Y(_0565_),
    .D(_0564_));
 sg13g2_nor3_2 _1508_ (.A(_0561_),
    .B(_0563_),
    .C(_0565_),
    .Y(_0566_));
 sg13g2_nand2_2 _1509_ (.Y(_0567_),
    .A(_0557_),
    .B(_0566_));
 sg13g2_inv_1 _1510_ (.Y(_0568_),
    .A(_0567_));
 sg13g2_nor3_1 _1511_ (.A(_0552_),
    .B(_0555_),
    .C(_0556_),
    .Y(_0569_));
 sg13g2_nor2_2 _1512_ (.A(net583),
    .B(_0568_),
    .Y(_0570_));
 sg13g2_nand2_2 _1513_ (.Y(_0571_),
    .A(net586),
    .B(_0567_));
 sg13g2_nand2_1 _1514_ (.Y(_0572_),
    .A(\music.melody_pos[1] ),
    .B(\music.melody_pos[0] ));
 sg13g2_xor2_1 _1515_ (.B(_0572_),
    .A(_0007_),
    .X(_0573_));
 sg13g2_or2_1 _1516_ (.X(_0574_),
    .B(\music.melody_pos[0] ),
    .A(\music.melody_pos[1] ));
 sg13g2_nor3_1 _1517_ (.A(_0514_),
    .B(\music.melody_pos[2] ),
    .C(_0574_),
    .Y(_0575_));
 sg13g2_a21oi_1 _1518_ (.A1(\music.melody_pos[3] ),
    .A2(_0575_),
    .Y(_0576_),
    .B1(_0567_));
 sg13g2_nand2_1 _1519_ (.Y(_0577_),
    .A(net586),
    .B(_0576_));
 sg13g2_inv_1 _1520_ (.Y(_0578_),
    .A(_0577_));
 sg13g2_a22oi_1 _1521_ (.Y(_0579_),
    .B1(_0573_),
    .B2(_0578_),
    .A2(_0570_),
    .A1(\music.melody_pos[2] ));
 sg13g2_inv_1 _1522_ (.Y(_0096_),
    .A(_0579_));
 sg13g2_nand3_1 _1523_ (.B(_0572_),
    .C(_0574_),
    .A(_0568_),
    .Y(_0580_));
 sg13g2_o21ai_1 _1524_ (.B1(_0580_),
    .Y(_0581_),
    .A1(net245),
    .A2(_0568_));
 sg13g2_nand2_1 _1525_ (.Y(_0582_),
    .A(net112),
    .B(_0576_));
 sg13g2_o21ai_1 _1526_ (.B1(_0582_),
    .Y(_0583_),
    .A1(_0006_),
    .A2(_0568_));
 sg13g2_nand2_1 _1527_ (.Y(_0584_),
    .A(net586),
    .B(_0583_));
 sg13g2_nor2_1 _1528_ (.A(_0581_),
    .B(_0584_),
    .Y(_0585_));
 sg13g2_nor2_1 _1529_ (.A(_0579_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_nand3_1 _1530_ (.B(_0579_),
    .C(_0583_),
    .A(net586),
    .Y(_0587_));
 sg13g2_xnor2_1 _1531_ (.Y(_0588_),
    .A(_0096_),
    .B(_0585_));
 sg13g2_nand2_1 _1532_ (.Y(_0589_),
    .A(net586),
    .B(_0581_));
 sg13g2_or2_1 _1533_ (.X(_0590_),
    .B(_0589_),
    .A(_0583_));
 sg13g2_nand2_1 _1534_ (.Y(_0591_),
    .A(_0588_),
    .B(_0590_));
 sg13g2_nand3_1 _1535_ (.B(\music.melody_pos[1] ),
    .C(\music.melody_pos[0] ),
    .A(\music.melody_pos[2] ),
    .Y(_0592_));
 sg13g2_nand4_1 _1536_ (.B(\music.melody_pos[2] ),
    .C(\music.melody_pos[1] ),
    .A(\music.melody_pos[3] ),
    .Y(_0593_),
    .D(\music.melody_pos[0] ));
 sg13g2_xor2_1 _1537_ (.B(_0593_),
    .A(_0008_),
    .X(_0594_));
 sg13g2_nand2_1 _1538_ (.Y(_0595_),
    .A(_0578_),
    .B(_0594_));
 sg13g2_o21ai_1 _1539_ (.B1(_0595_),
    .Y(_0596_),
    .A1(net243),
    .A2(_0571_));
 sg13g2_inv_1 _1540_ (.Y(_0597_),
    .A(_0596_));
 sg13g2_nand2_1 _1541_ (.Y(_0598_),
    .A(net242),
    .B(_0570_));
 sg13g2_xor2_1 _1542_ (.B(_0592_),
    .A(\music.melody_pos[3] ),
    .X(_0599_));
 sg13g2_o21ai_1 _1543_ (.B1(_0598_),
    .Y(_0097_),
    .A1(_0577_),
    .A2(_0599_));
 sg13g2_nand2b_1 _1544_ (.Y(_0600_),
    .B(_0596_),
    .A_N(_0097_));
 sg13g2_or2_1 _1545_ (.X(_0601_),
    .B(_0583_),
    .A(_0579_));
 sg13g2_nor2_1 _1546_ (.A(_0579_),
    .B(_0590_),
    .Y(_0602_));
 sg13g2_nor2_1 _1547_ (.A(_0600_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_nor2_1 _1548_ (.A(_0097_),
    .B(_0602_),
    .Y(_0604_));
 sg13g2_a221oi_1 _1549_ (.B2(_0587_),
    .C1(_0596_),
    .B1(_0604_),
    .A1(_0588_),
    .Y(_0605_),
    .A2(_0097_));
 sg13g2_a21oi_1 _1550_ (.A1(_0591_),
    .A2(_0603_),
    .Y(_0000_),
    .B1(_0605_));
 sg13g2_nor2_1 _1551_ (.A(_0586_),
    .B(_0097_),
    .Y(_0606_));
 sg13g2_nand2_1 _1552_ (.Y(_0607_),
    .A(_0579_),
    .B(_0589_));
 sg13g2_and3_1 _1553_ (.X(_0608_),
    .A(_0581_),
    .B(_0097_),
    .C(_0601_));
 sg13g2_a21oi_1 _1554_ (.A1(_0606_),
    .A2(_0607_),
    .Y(_0609_),
    .B1(_0608_));
 sg13g2_a21oi_1 _1555_ (.A1(_0579_),
    .A2(_0590_),
    .Y(_0610_),
    .B1(_0600_));
 sg13g2_nand2b_1 _1556_ (.Y(_0611_),
    .B(_0610_),
    .A_N(_0586_));
 sg13g2_o21ai_1 _1557_ (.B1(_0611_),
    .Y(_0001_),
    .A1(_0596_),
    .A2(_0609_));
 sg13g2_a21oi_1 _1558_ (.A1(_0597_),
    .A2(_0608_),
    .Y(_0002_),
    .B1(_0606_));
 sg13g2_nand2_1 _1559_ (.Y(_0612_),
    .A(_0096_),
    .B(_0589_));
 sg13g2_a21oi_1 _1560_ (.A1(_0590_),
    .A2(_0612_),
    .Y(_0613_),
    .B1(_0608_));
 sg13g2_and4_1 _1561_ (.A(_0581_),
    .B(_0590_),
    .C(_0097_),
    .D(_0612_),
    .X(_0614_));
 sg13g2_nor3_1 _1562_ (.A(_0596_),
    .B(_0613_),
    .C(_0614_),
    .Y(_0019_));
 sg13g2_nand2b_1 _1563_ (.Y(_0615_),
    .B(net587),
    .A_N(_0557_));
 sg13g2_nor2_1 _1564_ (.A(_0537_),
    .B(net542),
    .Y(_0020_));
 sg13g2_xnor2_1 _1565_ (.Y(_0616_),
    .A(\music.pwm_pos[1] ),
    .B(net197));
 sg13g2_nor2_1 _1566_ (.A(net542),
    .B(net198),
    .Y(_0021_));
 sg13g2_and3_1 _1567_ (.X(_0617_),
    .A(\music.pwm_pos[1] ),
    .B(\music.pwm_pos[0] ),
    .C(net143));
 sg13g2_a21oi_1 _1568_ (.A1(\music.pwm_pos[1] ),
    .A2(\music.pwm_pos[0] ),
    .Y(_0618_),
    .B1(net143));
 sg13g2_nor3_1 _1569_ (.A(net542),
    .B(_0617_),
    .C(net144),
    .Y(_0022_));
 sg13g2_and2_1 _1570_ (.A(net177),
    .B(_0617_),
    .X(_0619_));
 sg13g2_nor2_1 _1571_ (.A(net177),
    .B(_0617_),
    .Y(_0620_));
 sg13g2_nor3_1 _1572_ (.A(net542),
    .B(_0619_),
    .C(net178),
    .Y(_0023_));
 sg13g2_and2_1 _1573_ (.A(net199),
    .B(_0619_),
    .X(_0621_));
 sg13g2_nor2_1 _1574_ (.A(net199),
    .B(_0619_),
    .Y(_0622_));
 sg13g2_nor3_1 _1575_ (.A(net542),
    .B(_0621_),
    .C(_0622_),
    .Y(_0024_));
 sg13g2_and2_1 _1576_ (.A(net190),
    .B(_0621_),
    .X(_0623_));
 sg13g2_nor2_1 _1577_ (.A(net190),
    .B(_0621_),
    .Y(_0624_));
 sg13g2_nor3_1 _1578_ (.A(net542),
    .B(_0623_),
    .C(net191),
    .Y(_0025_));
 sg13g2_xnor2_1 _1579_ (.Y(_0625_),
    .A(net214),
    .B(_0623_));
 sg13g2_nor2_1 _1580_ (.A(net542),
    .B(_0625_),
    .Y(_0026_));
 sg13g2_a21oi_1 _1581_ (.A1(\music.pwm_pos[6] ),
    .A2(_0623_),
    .Y(_0626_),
    .B1(net172));
 sg13g2_and3_1 _1582_ (.X(_0627_),
    .A(\music.pwm_pos[6] ),
    .B(net172),
    .C(_0623_));
 sg13g2_nor3_1 _1583_ (.A(net542),
    .B(net173),
    .C(_0627_),
    .Y(_0027_));
 sg13g2_nor2_1 _1584_ (.A(net186),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_and2_1 _1585_ (.A(net186),
    .B(_0627_),
    .X(_0629_));
 sg13g2_nor3_1 _1586_ (.A(net543),
    .B(net187),
    .C(_0629_),
    .Y(_0028_));
 sg13g2_xnor2_1 _1587_ (.Y(_0630_),
    .A(net212),
    .B(_0629_));
 sg13g2_nor2_1 _1588_ (.A(net543),
    .B(_0630_),
    .Y(_0029_));
 sg13g2_a21oi_1 _1589_ (.A1(\music.pwm_pos[9] ),
    .A2(_0629_),
    .Y(_0631_),
    .B1(net138));
 sg13g2_and3_1 _1590_ (.X(_0632_),
    .A(\music.pwm_pos[9] ),
    .B(net138),
    .C(_0629_));
 sg13g2_nor3_1 _1591_ (.A(net543),
    .B(net139),
    .C(_0632_),
    .Y(_0030_));
 sg13g2_nor2_1 _1592_ (.A(net182),
    .B(_0632_),
    .Y(_0633_));
 sg13g2_and2_1 _1593_ (.A(net182),
    .B(_0632_),
    .X(_0634_));
 sg13g2_nor3_1 _1594_ (.A(net543),
    .B(net183),
    .C(_0634_),
    .Y(_0031_));
 sg13g2_nor2_1 _1595_ (.A(net162),
    .B(_0634_),
    .Y(_0635_));
 sg13g2_and2_1 _1596_ (.A(net162),
    .B(_0634_),
    .X(_0636_));
 sg13g2_nor3_1 _1597_ (.A(net543),
    .B(net163),
    .C(_0636_),
    .Y(_0032_));
 sg13g2_nor2_1 _1598_ (.A(net167),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_and2_1 _1599_ (.A(net167),
    .B(_0636_),
    .X(_0638_));
 sg13g2_nor3_1 _1600_ (.A(net543),
    .B(_0637_),
    .C(_0638_),
    .Y(_0033_));
 sg13g2_a21oi_1 _1601_ (.A1(net189),
    .A2(_0638_),
    .Y(_0639_),
    .B1(net543));
 sg13g2_o21ai_1 _1602_ (.B1(_0639_),
    .Y(_0640_),
    .A1(net189),
    .A2(_0638_));
 sg13g2_inv_1 _1603_ (.Y(_0034_),
    .A(_0640_));
 sg13g2_and2_1 _1604_ (.A(net565),
    .B(\gfx.bitmap_y[3] ),
    .X(_0641_));
 sg13g2_nand3_1 _1605_ (.B(net184),
    .C(_0641_),
    .A(net566),
    .Y(_0642_));
 sg13g2_nor4_1 _1606_ (.A(\gfx.pixel_y[0] ),
    .B(net569),
    .C(\gfx.pixel_y[9] ),
    .D(_0642_),
    .Y(_0643_));
 sg13g2_nor3_1 _1607_ (.A(_0522_),
    .B(_0523_),
    .C(\gfx.pixel_y[2] ),
    .Y(_0644_));
 sg13g2_a21oi_1 _1608_ (.A1(_0643_),
    .A2(_0644_),
    .Y(_0645_),
    .B1(net146));
 sg13g2_and4_1 _1609_ (.A(_0522_),
    .B(net575),
    .C(\gfx.pixel_y[2] ),
    .D(_0643_),
    .X(_0646_));
 sg13g2_o21ai_1 _1610_ (.B1(net588),
    .Y(_0035_),
    .A1(net147),
    .A2(_0646_));
 sg13g2_nor3_1 _1611_ (.A(\gfx.bitmap_x[0] ),
    .B(\gfx.pixel_x[2] ),
    .C(\gfx.pixel_x[8] ),
    .Y(_0647_));
 sg13g2_nand2_1 _1612_ (.Y(_0648_),
    .A(\gfx.pixel_x[9] ),
    .B(_0647_));
 sg13g2_nor3_1 _1613_ (.A(\gfx.pixel_x[1] ),
    .B(\gfx.pixel_x[0] ),
    .C(_0648_),
    .Y(_0649_));
 sg13g2_nor2b_2 _1614_ (.A(net578),
    .B_N(net577),
    .Y(_0650_));
 sg13g2_nor2b_1 _1615_ (.A(\gfx.bitmap_x[2] ),
    .B_N(net581),
    .Y(_0651_));
 sg13g2_nand3_1 _1616_ (.B(_0650_),
    .C(_0651_),
    .A(_0649_),
    .Y(_0652_));
 sg13g2_nand2b_1 _1617_ (.Y(_0653_),
    .B(_0652_),
    .A_N(net231));
 sg13g2_and2_1 _1618_ (.A(net582),
    .B(\gfx.bitmap_x[2] ),
    .X(_0654_));
 sg13g2_nand2_1 _1619_ (.Y(_0655_),
    .A(net581),
    .B(net580));
 sg13g2_nand4_1 _1620_ (.B(net579),
    .C(_0649_),
    .A(net153),
    .Y(_0656_),
    .D(_0654_));
 sg13g2_a21o_1 _1621_ (.A2(_0656_),
    .A1(_0653_),
    .B1(net584),
    .X(_0036_));
 sg13g2_nor2b_1 _1622_ (.A(net588),
    .B_N(net235),
    .Y(_0657_));
 sg13g2_nand2_2 _1623_ (.Y(_0658_),
    .A(net568),
    .B(net566));
 sg13g2_nor2_1 _1624_ (.A(net565),
    .B(\gfx.bitmap_y[3] ),
    .Y(_0659_));
 sg13g2_nand2_1 _1625_ (.Y(_0660_),
    .A(_0658_),
    .B(_0659_));
 sg13g2_and2_1 _1626_ (.A(_0010_),
    .B(_0660_),
    .X(_0661_));
 sg13g2_nand2_2 _1627_ (.Y(_0662_),
    .A(_0010_),
    .B(_0660_));
 sg13g2_and3_1 _1628_ (.X(_0663_),
    .A(_0525_),
    .B(net578),
    .C(_0651_));
 sg13g2_nor2_2 _1629_ (.A(net581),
    .B(net580),
    .Y(_0664_));
 sg13g2_nor2_1 _1630_ (.A(_0654_),
    .B(_0664_),
    .Y(_0665_));
 sg13g2_xnor2_1 _1631_ (.Y(_0666_),
    .A(net582),
    .B(net580));
 sg13g2_nor2_1 _1632_ (.A(net578),
    .B(_0666_),
    .Y(_0667_));
 sg13g2_or3_2 _1633_ (.A(net581),
    .B(net580),
    .C(net579),
    .X(_0668_));
 sg13g2_a22oi_1 _1634_ (.Y(_0669_),
    .B1(_0668_),
    .B2(_0525_),
    .A2(_0664_),
    .A1(_0650_));
 sg13g2_a221oi_1 _1635_ (.B2(_0525_),
    .C1(net581),
    .B1(_0668_),
    .A1(_0650_),
    .Y(_0670_),
    .A2(_0664_));
 sg13g2_nor2b_1 _1636_ (.A(net577),
    .B_N(net581),
    .Y(_0671_));
 sg13g2_nor2_1 _1637_ (.A(_0670_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_or2_1 _1638_ (.X(_0673_),
    .B(_0671_),
    .A(_0670_));
 sg13g2_a21oi_1 _1639_ (.A1(_0667_),
    .A2(_0672_),
    .Y(_0674_),
    .B1(_0663_));
 sg13g2_xor2_1 _1640_ (.B(_0664_),
    .A(net578),
    .X(_0675_));
 sg13g2_nor2_1 _1641_ (.A(_0672_),
    .B(_0675_),
    .Y(_0676_));
 sg13g2_or2_1 _1642_ (.X(_0677_),
    .B(net576),
    .A(net577));
 sg13g2_nand2_1 _1643_ (.Y(_0678_),
    .A(net577),
    .B(net576));
 sg13g2_xor2_1 _1644_ (.B(net576),
    .A(net577),
    .X(_0679_));
 sg13g2_a21oi_2 _1645_ (.B1(_0679_),
    .Y(_0680_),
    .A2(_0664_),
    .A1(_0650_));
 sg13g2_a21o_1 _1646_ (.A2(_0664_),
    .A1(_0650_),
    .B1(_0679_),
    .X(_0681_));
 sg13g2_nand3b_1 _1647_ (.B(_0650_),
    .C(_0664_),
    .Y(_0682_),
    .A_N(net576));
 sg13g2_nand2_1 _1648_ (.Y(_0683_),
    .A(_0681_),
    .B(_0682_));
 sg13g2_nand2_1 _1649_ (.Y(_0684_),
    .A(_0666_),
    .B(_0683_));
 sg13g2_and3_1 _1650_ (.X(_0685_),
    .A(_0666_),
    .B(_0681_),
    .C(_0682_));
 sg13g2_nor3_2 _1651_ (.A(_0654_),
    .B(_0664_),
    .C(_0679_),
    .Y(_0686_));
 sg13g2_nand2_1 _1652_ (.Y(_0687_),
    .A(_0014_),
    .B(_0669_));
 sg13g2_o21ai_1 _1653_ (.B1(_0687_),
    .Y(_0688_),
    .A1(_0685_),
    .A2(_0686_));
 sg13g2_or3_1 _1654_ (.A(_0685_),
    .B(_0686_),
    .C(_0687_),
    .X(_0689_));
 sg13g2_and3_1 _1655_ (.X(_0690_),
    .A(_0676_),
    .B(_0688_),
    .C(_0689_));
 sg13g2_nand3_1 _1656_ (.B(_0688_),
    .C(_0689_),
    .A(_0676_),
    .Y(_0691_));
 sg13g2_a21oi_1 _1657_ (.A1(_0688_),
    .A2(_0689_),
    .Y(_0692_),
    .B1(_0676_));
 sg13g2_or3_1 _1658_ (.A(_0674_),
    .B(_0690_),
    .C(_0692_),
    .X(_0693_));
 sg13g2_o21ai_1 _1659_ (.B1(_0674_),
    .Y(_0694_),
    .A1(_0690_),
    .A2(_0692_));
 sg13g2_and3_1 _1660_ (.X(_0695_),
    .A(net555),
    .B(_0693_),
    .C(_0694_));
 sg13g2_nand3_1 _1661_ (.B(_0693_),
    .C(_0694_),
    .A(net555),
    .Y(_0696_));
 sg13g2_nand2_2 _1662_ (.Y(_0697_),
    .A(_0011_),
    .B(_0658_));
 sg13g2_xor2_1 _1663_ (.B(_0697_),
    .A(net565),
    .X(_0698_));
 sg13g2_xnor2_1 _1664_ (.Y(_0699_),
    .A(\gfx.pixel_y[7] ),
    .B(_0697_));
 sg13g2_or2_1 _1665_ (.X(_0700_),
    .B(_0675_),
    .A(_0667_));
 sg13g2_nor4_1 _1666_ (.A(_0667_),
    .B(_0670_),
    .C(_0671_),
    .D(_0675_),
    .Y(_0701_));
 sg13g2_a221oi_1 _1667_ (.B2(_0700_),
    .C1(_0701_),
    .B1(_0673_),
    .A1(net578),
    .Y(_0702_),
    .A2(_0651_));
 sg13g2_or3_2 _1668_ (.A(_0663_),
    .B(net551),
    .C(_0702_),
    .X(_0703_));
 sg13g2_xnor2_1 _1669_ (.Y(_0704_),
    .A(_0531_),
    .B(_0658_));
 sg13g2_xnor2_1 _1670_ (.Y(_0705_),
    .A(_0011_),
    .B(_0658_));
 sg13g2_xnor2_1 _1671_ (.Y(_0706_),
    .A(net582),
    .B(net578));
 sg13g2_xnor2_1 _1672_ (.Y(_0707_),
    .A(net568),
    .B(net566));
 sg13g2_nand2_1 _1673_ (.Y(_0708_),
    .A(net580),
    .B(net559));
 sg13g2_xor2_1 _1674_ (.B(net559),
    .A(net580),
    .X(_0709_));
 sg13g2_xnor2_1 _1675_ (.Y(_0710_),
    .A(net580),
    .B(net559));
 sg13g2_nand2_2 _1676_ (.Y(_0711_),
    .A(net570),
    .B(net582));
 sg13g2_o21ai_1 _1677_ (.B1(_0708_),
    .Y(_0712_),
    .A1(_0710_),
    .A2(_0711_));
 sg13g2_xnor2_1 _1678_ (.Y(_0713_),
    .A(_0705_),
    .B(_0706_));
 sg13g2_nand2b_1 _1679_ (.Y(_0714_),
    .B(_0712_),
    .A_N(_0713_));
 sg13g2_o21ai_1 _1680_ (.B1(_0714_),
    .Y(_0715_),
    .A1(_0705_),
    .A2(_0706_));
 sg13g2_o21ai_1 _1681_ (.B1(net551),
    .Y(_0716_),
    .A1(_0663_),
    .A2(_0702_));
 sg13g2_nand2_1 _1682_ (.Y(_0717_),
    .A(_0703_),
    .B(_0716_));
 sg13g2_and3_2 _1683_ (.X(_0718_),
    .A(_0703_),
    .B(_0715_),
    .C(_0716_));
 sg13g2_nand3_1 _1684_ (.B(_0715_),
    .C(_0716_),
    .A(_0703_),
    .Y(_0719_));
 sg13g2_and2_1 _1685_ (.A(_0703_),
    .B(net515),
    .X(_0720_));
 sg13g2_nand2_1 _1686_ (.Y(_0721_),
    .A(_0703_),
    .B(net515));
 sg13g2_a21oi_1 _1687_ (.A1(_0693_),
    .A2(_0694_),
    .Y(_0722_),
    .B1(net555));
 sg13g2_a21o_1 _1688_ (.A2(_0694_),
    .A1(_0693_),
    .B1(net555),
    .X(_0723_));
 sg13g2_nor3_1 _1689_ (.A(_0695_),
    .B(_0720_),
    .C(_0722_),
    .Y(_0724_));
 sg13g2_nand3_1 _1690_ (.B(_0721_),
    .C(_0723_),
    .A(_0696_),
    .Y(_0725_));
 sg13g2_o21ai_1 _1691_ (.B1(_0696_),
    .Y(_0726_),
    .A1(_0720_),
    .A2(_0722_));
 sg13g2_o21ai_1 _1692_ (.B1(_0691_),
    .Y(_0727_),
    .A1(_0674_),
    .A2(_0692_));
 sg13g2_o21ai_1 _1693_ (.B1(_0014_),
    .Y(_0728_),
    .A1(_0685_),
    .A2(_0686_));
 sg13g2_nand2_1 _1694_ (.Y(_0729_),
    .A(_0669_),
    .B(_0728_));
 sg13g2_nor2_1 _1695_ (.A(_0675_),
    .B(_0679_),
    .Y(_0730_));
 sg13g2_a21oi_1 _1696_ (.A1(_0675_),
    .A2(_0681_),
    .Y(_0731_),
    .B1(_0730_));
 sg13g2_xor2_1 _1697_ (.B(_0731_),
    .A(_0684_),
    .X(_0732_));
 sg13g2_nor2_1 _1698_ (.A(_0729_),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_xor2_1 _1699_ (.B(_0732_),
    .A(_0729_),
    .X(_0734_));
 sg13g2_xnor2_1 _1700_ (.Y(_0735_),
    .A(_0727_),
    .B(_0734_));
 sg13g2_nor2_1 _1701_ (.A(net554),
    .B(_0735_),
    .Y(_0736_));
 sg13g2_nand2_1 _1702_ (.Y(_0737_),
    .A(net554),
    .B(_0735_));
 sg13g2_xnor2_1 _1703_ (.Y(_0738_),
    .A(net555),
    .B(_0735_));
 sg13g2_xor2_1 _1704_ (.B(_0738_),
    .A(_0726_),
    .X(_0739_));
 sg13g2_xnor2_1 _1705_ (.Y(_0740_),
    .A(_0726_),
    .B(_0738_));
 sg13g2_a21oi_1 _1706_ (.A1(_0696_),
    .A2(_0723_),
    .Y(_0741_),
    .B1(_0721_));
 sg13g2_o21ai_1 _1707_ (.B1(_0720_),
    .Y(_0742_),
    .A1(_0695_),
    .A2(_0722_));
 sg13g2_nor2_1 _1708_ (.A(net492),
    .B(net480),
    .Y(_0743_));
 sg13g2_nand2_1 _1709_ (.Y(_0744_),
    .A(net485),
    .B(net476));
 sg13g2_xnor2_1 _1710_ (.Y(_0745_),
    .A(_0712_),
    .B(_0713_));
 sg13g2_xor2_1 _1711_ (.B(_0713_),
    .A(_0712_),
    .X(_0746_));
 sg13g2_xor2_1 _1712_ (.B(net582),
    .A(net570),
    .X(_0747_));
 sg13g2_xnor2_1 _1713_ (.Y(_0748_),
    .A(_0709_),
    .B(_0711_));
 sg13g2_xnor2_1 _1714_ (.Y(_0749_),
    .A(_0710_),
    .B(_0711_));
 sg13g2_nor2_1 _1715_ (.A(net571),
    .B(net547),
    .Y(_0750_));
 sg13g2_nand2b_1 _1716_ (.Y(_0751_),
    .B(net545),
    .A_N(net557));
 sg13g2_nor2_2 _1717_ (.A(net571),
    .B(net558),
    .Y(_0752_));
 sg13g2_or2_2 _1718_ (.X(_0753_),
    .B(net558),
    .A(net571));
 sg13g2_nor2_2 _1719_ (.A(net548),
    .B(_0753_),
    .Y(_0754_));
 sg13g2_nand2_2 _1720_ (.Y(_0755_),
    .A(net545),
    .B(_0752_));
 sg13g2_nand2_2 _1721_ (.Y(_0756_),
    .A(net540),
    .B(_0755_));
 sg13g2_inv_2 _1722_ (.Y(_0757_),
    .A(_0756_));
 sg13g2_a21oi_2 _1723_ (.B1(_0715_),
    .Y(_0758_),
    .A2(_0716_),
    .A1(_0703_));
 sg13g2_a21o_2 _1724_ (.A2(_0716_),
    .A1(_0703_),
    .B1(_0715_),
    .X(_0759_));
 sg13g2_nand2_1 _1725_ (.Y(_0760_),
    .A(_0715_),
    .B(_0717_));
 sg13g2_or2_1 _1726_ (.X(_0761_),
    .B(_0717_),
    .A(_0715_));
 sg13g2_nor2_1 _1727_ (.A(_0718_),
    .B(_0758_),
    .Y(_0762_));
 sg13g2_nand2_1 _1728_ (.Y(_0763_),
    .A(net515),
    .B(_0759_));
 sg13g2_and2_2 _1729_ (.A(net571),
    .B(net558),
    .X(_0764_));
 sg13g2_nand2_2 _1730_ (.Y(_0765_),
    .A(net571),
    .B(net558));
 sg13g2_nor2_1 _1731_ (.A(_0710_),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_nand2_2 _1732_ (.Y(_0767_),
    .A(_0709_),
    .B(_0764_));
 sg13g2_nor2_1 _1733_ (.A(net537),
    .B(_0766_),
    .Y(_0768_));
 sg13g2_nand2_1 _1734_ (.Y(_0769_),
    .A(net531),
    .B(_0767_));
 sg13g2_a21oi_2 _1735_ (.B1(_0768_),
    .Y(_0770_),
    .A2(_0759_),
    .A1(net515));
 sg13g2_nand2_1 _1736_ (.Y(_0771_),
    .A(net499),
    .B(_0769_));
 sg13g2_a22oi_1 _1737_ (.Y(_0772_),
    .B1(_0756_),
    .B2(_0770_),
    .A2(net474),
    .A1(net487));
 sg13g2_nand2_2 _1738_ (.Y(_0773_),
    .A(_0709_),
    .B(net557));
 sg13g2_nor2_2 _1739_ (.A(net539),
    .B(_0773_),
    .Y(_0774_));
 sg13g2_inv_1 _1740_ (.Y(_0775_),
    .A(_0774_));
 sg13g2_and2_2 _1741_ (.A(net572),
    .B(net557),
    .X(_0776_));
 sg13g2_nand2_2 _1742_ (.Y(_0777_),
    .A(net572),
    .B(net557));
 sg13g2_nand2_2 _1743_ (.Y(_0778_),
    .A(_0709_),
    .B(_0776_));
 sg13g2_nand2_1 _1744_ (.Y(_0779_),
    .A(net573),
    .B(_0774_));
 sg13g2_nor2_1 _1745_ (.A(net501),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_or3_1 _1746_ (.A(net491),
    .B(net479),
    .C(_0780_),
    .X(_0781_));
 sg13g2_nand3b_1 _1747_ (.B(_0781_),
    .C(net564),
    .Y(_0782_),
    .A_N(_0772_));
 sg13g2_a21oi_2 _1748_ (.B1(net512),
    .Y(_0783_),
    .A2(net475),
    .A1(net487));
 sg13g2_nor2_1 _1749_ (.A(net557),
    .B(net545),
    .Y(_0784_));
 sg13g2_nand2b_2 _1750_ (.Y(_0785_),
    .B(net547),
    .A_N(net557));
 sg13g2_nor2_2 _1751_ (.A(net572),
    .B(net557),
    .Y(_0786_));
 sg13g2_or2_2 _1752_ (.X(_0787_),
    .B(net557),
    .A(net572));
 sg13g2_nor2_1 _1753_ (.A(_0749_),
    .B(_0787_),
    .Y(_0788_));
 sg13g2_nand2_2 _1754_ (.Y(_0789_),
    .A(net548),
    .B(_0786_));
 sg13g2_nand2_2 _1755_ (.Y(_0790_),
    .A(_0778_),
    .B(_0789_));
 sg13g2_nand2_1 _1756_ (.Y(_0791_),
    .A(net528),
    .B(_0790_));
 sg13g2_inv_1 _1757_ (.Y(_0792_),
    .A(_0791_));
 sg13g2_nor3_2 _1758_ (.A(net490),
    .B(net478),
    .C(net497),
    .Y(_0793_));
 sg13g2_nor2_1 _1759_ (.A(net546),
    .B(_0753_),
    .Y(_0794_));
 sg13g2_nand2_2 _1760_ (.Y(_0795_),
    .A(net548),
    .B(_0752_));
 sg13g2_nor2_1 _1761_ (.A(net540),
    .B(_0795_),
    .Y(_0796_));
 sg13g2_nand2_1 _1762_ (.Y(_0797_),
    .A(net527),
    .B(_0794_));
 sg13g2_a22oi_1 _1763_ (.Y(_0798_),
    .B1(_0793_),
    .B2(_0796_),
    .A2(_0792_),
    .A1(_0783_));
 sg13g2_o21ai_1 _1764_ (.B1(_0782_),
    .Y(_0799_),
    .A1(net564),
    .A2(_0798_));
 sg13g2_a21oi_1 _1765_ (.A1(_0727_),
    .A2(_0734_),
    .Y(_0800_),
    .B1(_0733_));
 sg13g2_o21ai_1 _1766_ (.B1(_0683_),
    .Y(_0801_),
    .A1(_0665_),
    .A2(_0731_));
 sg13g2_nand2b_1 _1767_ (.Y(_0802_),
    .B(_0668_),
    .A_N(_0678_));
 sg13g2_or2_1 _1768_ (.X(_0803_),
    .B(_0678_),
    .A(_0675_));
 sg13g2_o21ai_1 _1769_ (.B1(_0803_),
    .Y(_0804_),
    .A1(_0669_),
    .A2(_0730_));
 sg13g2_nor2_1 _1770_ (.A(_0801_),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_xnor2_1 _1771_ (.Y(_0806_),
    .A(_0801_),
    .B(_0804_));
 sg13g2_xor2_1 _1772_ (.B(_0806_),
    .A(_0800_),
    .X(_0807_));
 sg13g2_nand2_1 _1773_ (.Y(_0808_),
    .A(net555),
    .B(_0807_));
 sg13g2_nor2_1 _1774_ (.A(net555),
    .B(_0807_),
    .Y(_0809_));
 sg13g2_xnor2_1 _1775_ (.Y(_0810_),
    .A(net554),
    .B(_0807_));
 sg13g2_o21ai_1 _1776_ (.B1(_0737_),
    .Y(_0811_),
    .A1(_0726_),
    .A2(_0736_));
 sg13g2_xnor2_1 _1777_ (.Y(_0812_),
    .A(_0810_),
    .B(_0811_));
 sg13g2_xor2_1 _1778_ (.B(_0811_),
    .A(_0810_),
    .X(_0813_));
 sg13g2_nor2_2 _1779_ (.A(net536),
    .B(net548),
    .Y(_0814_));
 sg13g2_nand2_2 _1780_ (.Y(_0815_),
    .A(net529),
    .B(_0749_));
 sg13g2_nor3_1 _1781_ (.A(_0718_),
    .B(_0758_),
    .C(_0815_),
    .Y(_0816_));
 sg13g2_nand2_1 _1782_ (.Y(_0817_),
    .A(net511),
    .B(_0814_));
 sg13g2_a21oi_1 _1783_ (.A1(net486),
    .A2(net474),
    .Y(_0818_),
    .B1(net500));
 sg13g2_nor2_2 _1784_ (.A(net530),
    .B(_0773_),
    .Y(_0819_));
 sg13g2_inv_1 _1785_ (.Y(_0820_),
    .A(_0819_));
 sg13g2_a21oi_1 _1786_ (.A1(net487),
    .A2(net474),
    .Y(_0821_),
    .B1(_0819_));
 sg13g2_o21ai_1 _1787_ (.B1(_0817_),
    .Y(_0822_),
    .A1(net451),
    .A2(_0821_));
 sg13g2_nor2_2 _1788_ (.A(_0748_),
    .B(_0764_),
    .Y(_0823_));
 sg13g2_nand2_2 _1789_ (.Y(_0824_),
    .A(net546),
    .B(_0765_));
 sg13g2_nor2_2 _1790_ (.A(net531),
    .B(_0823_),
    .Y(_0825_));
 sg13g2_nand2_1 _1791_ (.Y(_0826_),
    .A(net540),
    .B(_0824_));
 sg13g2_nand2_1 _1792_ (.Y(_0827_),
    .A(net512),
    .B(_0824_));
 sg13g2_nor3_2 _1793_ (.A(_0718_),
    .B(_0758_),
    .C(_0826_),
    .Y(_0828_));
 sg13g2_nor4_2 _1794_ (.A(net491),
    .B(net479),
    .C(_0780_),
    .Y(_0829_),
    .D(_0828_));
 sg13g2_a21oi_2 _1795_ (.B1(_0814_),
    .Y(_0830_),
    .A2(_0759_),
    .A1(_0719_));
 sg13g2_nor2_1 _1796_ (.A(net511),
    .B(_0825_),
    .Y(_0831_));
 sg13g2_nand2_1 _1797_ (.Y(_0832_),
    .A(net501),
    .B(_0826_));
 sg13g2_o21ai_1 _1798_ (.B1(_0829_),
    .Y(_0833_),
    .A1(_0814_),
    .A2(_0832_));
 sg13g2_a21o_1 _1799_ (.A2(_0833_),
    .A1(_0822_),
    .B1(net564),
    .X(_0834_));
 sg13g2_nor2_2 _1800_ (.A(net531),
    .B(_0749_),
    .Y(_0835_));
 sg13g2_nand2_2 _1801_ (.Y(_0836_),
    .A(net536),
    .B(net547));
 sg13g2_nor2_1 _1802_ (.A(net545),
    .B(_0752_),
    .Y(_0837_));
 sg13g2_nor2_1 _1803_ (.A(_0752_),
    .B(_0836_),
    .Y(_0838_));
 sg13g2_nand2_2 _1804_ (.Y(_0839_),
    .A(net540),
    .B(net522));
 sg13g2_nor2_1 _1805_ (.A(net530),
    .B(net524),
    .Y(_0840_));
 sg13g2_nor2_2 _1806_ (.A(net528),
    .B(_0755_),
    .Y(_0841_));
 sg13g2_nand2_1 _1807_ (.Y(_0842_),
    .A(net539),
    .B(_0754_));
 sg13g2_nand2_1 _1808_ (.Y(_0843_),
    .A(_0839_),
    .B(_0842_));
 sg13g2_and2_1 _1809_ (.A(net529),
    .B(_0773_),
    .X(_0844_));
 sg13g2_nand2_2 _1810_ (.Y(_0845_),
    .A(net530),
    .B(_0773_));
 sg13g2_a221oi_1 _1811_ (.B2(_0761_),
    .C1(_0845_),
    .B1(_0760_),
    .A1(net483),
    .Y(_0846_),
    .A2(net471));
 sg13g2_nand2_2 _1812_ (.Y(_0847_),
    .A(net500),
    .B(_0839_));
 sg13g2_nor3_1 _1813_ (.A(net491),
    .B(net479),
    .C(_0847_),
    .Y(_0848_));
 sg13g2_nor2_1 _1814_ (.A(net562),
    .B(_0846_),
    .Y(_0849_));
 sg13g2_a22oi_1 _1815_ (.Y(_0850_),
    .B1(_0845_),
    .B2(_0848_),
    .A2(_0843_),
    .A1(_0793_));
 sg13g2_a21oi_1 _1816_ (.A1(_0849_),
    .A2(_0850_),
    .Y(_0851_),
    .B1(net463));
 sg13g2_a221oi_1 _1817_ (.B2(_0851_),
    .C1(_0812_),
    .B1(_0834_),
    .A1(net463),
    .Y(_0852_),
    .A2(_0799_));
 sg13g2_nor2_1 _1818_ (.A(net540),
    .B(_0764_),
    .Y(_0853_));
 sg13g2_nor2_1 _1819_ (.A(net541),
    .B(_0824_),
    .Y(_0854_));
 sg13g2_a21oi_2 _1820_ (.B1(_0854_),
    .Y(_0855_),
    .A2(_0759_),
    .A1(_0719_));
 sg13g2_and2_2 _1821_ (.A(_0710_),
    .B(net558),
    .X(_0856_));
 sg13g2_nand2_1 _1822_ (.Y(_0857_),
    .A(_0710_),
    .B(_0764_));
 sg13g2_nand2_1 _1823_ (.Y(_0858_),
    .A(net533),
    .B(_0856_));
 sg13g2_nor2_2 _1824_ (.A(net525),
    .B(net544),
    .Y(_0859_));
 sg13g2_nor2_1 _1825_ (.A(net526),
    .B(net523),
    .Y(_0860_));
 sg13g2_nand2_2 _1826_ (.Y(_0861_),
    .A(net537),
    .B(_0794_));
 sg13g2_nor2_2 _1827_ (.A(_0859_),
    .B(_0860_),
    .Y(_0862_));
 sg13g2_a21oi_1 _1828_ (.A1(net523),
    .A2(net544),
    .Y(_0863_),
    .B1(net527));
 sg13g2_and2_2 _1829_ (.A(_0012_),
    .B(_0819_),
    .X(_0864_));
 sg13g2_nor4_2 _1830_ (.A(_0718_),
    .B(_0758_),
    .C(_0841_),
    .Y(_0865_),
    .D(_0864_));
 sg13g2_nand2_1 _1831_ (.Y(_0866_),
    .A(net528),
    .B(net522));
 sg13g2_a22oi_1 _1832_ (.Y(_0867_),
    .B1(_0865_),
    .B2(_0866_),
    .A2(_0862_),
    .A1(_0855_));
 sg13g2_nor2_1 _1833_ (.A(net456),
    .B(_0867_),
    .Y(_0868_));
 sg13g2_nand2_2 _1834_ (.Y(_0869_),
    .A(net541),
    .B(_0767_));
 sg13g2_nand2b_2 _1835_ (.Y(_0870_),
    .B(net525),
    .A_N(net524));
 sg13g2_nor2_2 _1836_ (.A(net538),
    .B(_0755_),
    .Y(_0871_));
 sg13g2_nand2_2 _1837_ (.Y(_0872_),
    .A(net530),
    .B(_0754_));
 sg13g2_nand4_1 _1838_ (.B(_0775_),
    .C(_0869_),
    .A(net497),
    .Y(_0873_),
    .D(_0872_));
 sg13g2_or2_2 _1839_ (.X(_0874_),
    .B(net522),
    .A(net540));
 sg13g2_nor2_1 _1840_ (.A(net535),
    .B(net521),
    .Y(_0875_));
 sg13g2_nand4_1 _1841_ (.B(net470),
    .C(net504),
    .A(net482),
    .Y(_0876_),
    .D(_0875_));
 sg13g2_o21ai_1 _1842_ (.B1(_0876_),
    .Y(_0877_),
    .A1(_0744_),
    .A2(_0873_));
 sg13g2_o21ai_1 _1843_ (.B1(net463),
    .Y(_0878_),
    .A1(_0868_),
    .A2(_0877_));
 sg13g2_nand2_1 _1844_ (.Y(_0879_),
    .A(_0831_),
    .B(_0874_));
 sg13g2_a21oi_1 _1845_ (.A1(net486),
    .A2(net474),
    .Y(_0880_),
    .B1(_0828_));
 sg13g2_nand2_2 _1846_ (.Y(_0881_),
    .A(_0755_),
    .B(_0768_));
 sg13g2_nor2_2 _1847_ (.A(net499),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_a21oi_1 _1848_ (.A1(net499),
    .A2(_0871_),
    .Y(_0883_),
    .B1(_0882_));
 sg13g2_a221oi_1 _1849_ (.B2(net456),
    .C1(net461),
    .B1(_0883_),
    .A1(_0879_),
    .Y(_0884_),
    .A2(_0880_));
 sg13g2_nor2_1 _1850_ (.A(net560),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_nand2_1 _1851_ (.Y(_0886_),
    .A(_0777_),
    .B(_0787_));
 sg13g2_nand3_1 _1852_ (.B(net546),
    .C(_0886_),
    .A(net534),
    .Y(_0887_));
 sg13g2_and2_1 _1853_ (.A(_0872_),
    .B(_0887_),
    .X(_0888_));
 sg13g2_a221oi_1 _1854_ (.B2(_0815_),
    .C1(net454),
    .B1(_0839_),
    .A1(net512),
    .Y(_0889_),
    .A2(_0824_));
 sg13g2_nor2_1 _1855_ (.A(net546),
    .B(_0764_),
    .Y(_0890_));
 sg13g2_nand2_2 _1856_ (.Y(_0891_),
    .A(net547),
    .B(_0765_));
 sg13g2_nand2_1 _1857_ (.Y(_0892_),
    .A(_0767_),
    .B(_0824_));
 sg13g2_nand2_1 _1858_ (.Y(_0893_),
    .A(net538),
    .B(_0790_));
 sg13g2_o21ai_1 _1859_ (.B1(_0893_),
    .Y(_0894_),
    .A1(net540),
    .A2(_0892_));
 sg13g2_nor2_2 _1860_ (.A(net534),
    .B(_0823_),
    .Y(_0895_));
 sg13g2_nor2_1 _1861_ (.A(_0757_),
    .B(_0854_),
    .Y(_0896_));
 sg13g2_nand2_1 _1862_ (.Y(_0897_),
    .A(net512),
    .B(_0874_));
 sg13g2_nor2_1 _1863_ (.A(net509),
    .B(_0864_),
    .Y(_0898_));
 sg13g2_or2_1 _1864_ (.X(_0899_),
    .B(_0864_),
    .A(net508));
 sg13g2_nand4_1 _1865_ (.B(net473),
    .C(_0897_),
    .A(net486),
    .Y(_0900_),
    .D(_0899_));
 sg13g2_o21ai_1 _1866_ (.B1(net560),
    .Y(_0901_),
    .A1(net461),
    .A2(_0900_));
 sg13g2_mux2_1 _1867_ (.A0(_0888_),
    .A1(_0896_),
    .S(net466),
    .X(_0902_));
 sg13g2_a221oi_1 _1868_ (.B2(_0783_),
    .C1(_0901_),
    .B1(_0902_),
    .A1(net461),
    .Y(_0903_),
    .A2(_0889_));
 sg13g2_nor3_1 _1869_ (.A(net462),
    .B(_0869_),
    .C(_0896_),
    .Y(_0904_));
 sg13g2_nor2_1 _1870_ (.A(net466),
    .B(_0894_),
    .Y(_0905_));
 sg13g2_o21ai_1 _1871_ (.B1(net451),
    .Y(_0906_),
    .A1(_0904_),
    .A2(_0905_));
 sg13g2_a221oi_1 _1872_ (.B2(_0906_),
    .C1(_0813_),
    .B1(_0903_),
    .A1(_0878_),
    .Y(_0907_),
    .A2(_0885_));
 sg13g2_o21ai_1 _1873_ (.B1(_0808_),
    .Y(_0908_),
    .A1(_0809_),
    .A2(_0811_));
 sg13g2_o21ai_1 _1874_ (.B1(_0802_),
    .Y(_0909_),
    .A1(net576),
    .A2(_0668_));
 sg13g2_nor2_1 _1875_ (.A(_0805_),
    .B(_0909_),
    .Y(_0910_));
 sg13g2_o21ai_1 _1876_ (.B1(_0910_),
    .Y(_0911_),
    .A1(_0800_),
    .A2(_0806_));
 sg13g2_xnor2_1 _1877_ (.Y(_0912_),
    .A(net555),
    .B(_0911_));
 sg13g2_xnor2_1 _1878_ (.Y(_0913_),
    .A(_0908_),
    .B(_0912_));
 sg13g2_nor3_1 _1879_ (.A(_0852_),
    .B(_0907_),
    .C(net448),
    .Y(_0914_));
 sg13g2_nand2_1 _1880_ (.Y(_0915_),
    .A(\gfx.pixel_y[8] ),
    .B(_0660_));
 sg13g2_nor2_1 _1881_ (.A(net565),
    .B(\gfx.pixel_y[8] ),
    .Y(_0916_));
 sg13g2_nor3_1 _1882_ (.A(\gfx.pixel_y[9] ),
    .B(\gfx.pixel_x[9] ),
    .C(_0916_),
    .Y(_0917_));
 sg13g2_nand2_1 _1883_ (.Y(_0918_),
    .A(_0915_),
    .B(_0917_));
 sg13g2_nor2_1 _1884_ (.A(_0680_),
    .B(_0918_),
    .Y(_0919_));
 sg13g2_inv_1 _1885_ (.Y(_0920_),
    .A(net516));
 sg13g2_nor2_1 _1886_ (.A(_0755_),
    .B(net501),
    .Y(_0921_));
 sg13g2_nor3_2 _1887_ (.A(net491),
    .B(net479),
    .C(_0921_),
    .Y(_0922_));
 sg13g2_and2_2 _1888_ (.A(net533),
    .B(net524),
    .X(_0923_));
 sg13g2_nand2_2 _1889_ (.Y(_0924_),
    .A(net535),
    .B(net524));
 sg13g2_nand2_1 _1890_ (.Y(_0925_),
    .A(net501),
    .B(_0825_));
 sg13g2_nor2_2 _1891_ (.A(net506),
    .B(_0874_),
    .Y(_0926_));
 sg13g2_a21oi_2 _1892_ (.B1(_0926_),
    .Y(_0927_),
    .A2(net471),
    .A1(net483));
 sg13g2_nor2_1 _1893_ (.A(net501),
    .B(_0825_),
    .Y(_0928_));
 sg13g2_nand2_1 _1894_ (.Y(_0929_),
    .A(_0845_),
    .B(_0928_));
 sg13g2_nand2_1 _1895_ (.Y(_0930_),
    .A(net495),
    .B(_0835_));
 sg13g2_a221oi_1 _1896_ (.B2(_0924_),
    .C1(_0926_),
    .B1(net506),
    .A1(net483),
    .Y(_0931_),
    .A2(net472));
 sg13g2_nand2_2 _1897_ (.Y(_0932_),
    .A(_0757_),
    .B(_0892_));
 sg13g2_nand2_1 _1898_ (.Y(_0933_),
    .A(_0765_),
    .B(net522));
 sg13g2_nand4_1 _1899_ (.B(_0828_),
    .C(net544),
    .A(_0757_),
    .Y(_0934_),
    .D(_0891_));
 sg13g2_nand2_1 _1900_ (.Y(_0935_),
    .A(_0755_),
    .B(net495));
 sg13g2_or3_1 _1901_ (.A(net527),
    .B(net521),
    .C(_0935_),
    .X(_0936_));
 sg13g2_nand3_1 _1902_ (.B(_0934_),
    .C(_0936_),
    .A(net455),
    .Y(_0937_));
 sg13g2_nand2_1 _1903_ (.Y(_0938_),
    .A(_0767_),
    .B(_0825_));
 sg13g2_a221oi_1 _1904_ (.B2(net456),
    .C1(net511),
    .B1(_0938_),
    .A1(_0769_),
    .Y(_0939_),
    .A2(_0821_));
 sg13g2_nand3_1 _1905_ (.B(_0827_),
    .C(_0847_),
    .A(net456),
    .Y(_0940_));
 sg13g2_nand2_2 _1906_ (.Y(_0941_),
    .A(_0012_),
    .B(net548));
 sg13g2_nand2_2 _1907_ (.Y(_0942_),
    .A(net531),
    .B(_0941_));
 sg13g2_nand3_1 _1908_ (.B(_0839_),
    .C(_0942_),
    .A(net512),
    .Y(_0943_));
 sg13g2_a22oi_1 _1909_ (.Y(_0944_),
    .B1(_0881_),
    .B2(_0943_),
    .A2(net475),
    .A1(net486));
 sg13g2_nand2b_1 _1910_ (.Y(_0945_),
    .B(_0944_),
    .A_N(_0882_));
 sg13g2_a21oi_1 _1911_ (.A1(_0940_),
    .A2(_0945_),
    .Y(_0946_),
    .B1(net560));
 sg13g2_a22oi_1 _1912_ (.Y(_0947_),
    .B1(_0927_),
    .B2(_0929_),
    .A2(_0925_),
    .A1(_0922_));
 sg13g2_a21o_1 _1913_ (.A2(_0947_),
    .A1(net561),
    .B1(net462),
    .X(_0948_));
 sg13g2_a21o_1 _1914_ (.A2(_0836_),
    .A1(net450),
    .B1(_0939_),
    .X(_0949_));
 sg13g2_a21oi_1 _1915_ (.A1(_0930_),
    .A2(_0931_),
    .Y(_0950_),
    .B1(net564));
 sg13g2_a221oi_1 _1916_ (.B2(_0937_),
    .C1(net465),
    .B1(_0950_),
    .A1(net564),
    .Y(_0951_),
    .A2(_0949_));
 sg13g2_o21ai_1 _1917_ (.B1(net447),
    .Y(_0952_),
    .A1(_0946_),
    .A2(_0948_));
 sg13g2_o21ai_1 _1918_ (.B1(net516),
    .Y(_0953_),
    .A1(_0951_),
    .A2(_0952_));
 sg13g2_nor2_1 _1919_ (.A(_0677_),
    .B(_0918_),
    .Y(_0954_));
 sg13g2_and2_2 _1920_ (.A(net579),
    .B(_0954_),
    .X(_0955_));
 sg13g2_nor2_1 _1921_ (.A(_0523_),
    .B(net568),
    .Y(_0956_));
 sg13g2_nand2b_2 _1922_ (.Y(_0957_),
    .B(net574),
    .A_N(net568));
 sg13g2_nand2_1 _1923_ (.Y(_0958_),
    .A(_0707_),
    .B(_0957_));
 sg13g2_nor2_1 _1924_ (.A(_0705_),
    .B(_0958_),
    .Y(_0959_));
 sg13g2_nand2_1 _1925_ (.Y(_0960_),
    .A(net549),
    .B(_0959_));
 sg13g2_nor2b_2 _1926_ (.A(net574),
    .B_N(net568),
    .Y(_0961_));
 sg13g2_nor2_2 _1927_ (.A(net559),
    .B(_0961_),
    .Y(_0962_));
 sg13g2_nor2_1 _1928_ (.A(net556),
    .B(net552),
    .Y(_0963_));
 sg13g2_a21oi_1 _1929_ (.A1(net552),
    .A2(_0962_),
    .Y(_0964_),
    .B1(net556));
 sg13g2_nor2_1 _1930_ (.A(_0531_),
    .B(_0957_),
    .Y(_0965_));
 sg13g2_nor3_1 _1931_ (.A(net549),
    .B(_0959_),
    .C(_0965_),
    .Y(_0966_));
 sg13g2_nor2_1 _1932_ (.A(_0524_),
    .B(_0957_),
    .Y(_0967_));
 sg13g2_nand2_2 _1933_ (.Y(_0968_),
    .A(net567),
    .B(_0956_));
 sg13g2_o21ai_1 _1934_ (.B1(_0705_),
    .Y(_0969_),
    .A1(net574),
    .A2(_0658_));
 sg13g2_o21ai_1 _1935_ (.B1(_0966_),
    .Y(_0970_),
    .A1(_0967_),
    .A2(_0969_));
 sg13g2_o21ai_1 _1936_ (.B1(net556),
    .Y(_0971_),
    .A1(net552),
    .A2(_0969_));
 sg13g2_o21ai_1 _1937_ (.B1(_0971_),
    .Y(_0972_),
    .A1(_0662_),
    .A2(_0968_));
 sg13g2_a22oi_1 _1938_ (.Y(_0973_),
    .B1(_0970_),
    .B2(_0972_),
    .A2(_0964_),
    .A1(_0960_));
 sg13g2_nor3_1 _1939_ (.A(net574),
    .B(net568),
    .C(net567),
    .Y(_0974_));
 sg13g2_nor2_2 _1940_ (.A(_0697_),
    .B(_0974_),
    .Y(_0975_));
 sg13g2_nor2_1 _1941_ (.A(net553),
    .B(_0975_),
    .Y(_0976_));
 sg13g2_nor2_1 _1942_ (.A(_0662_),
    .B(_0976_),
    .Y(_0977_));
 sg13g2_nor2_1 _1943_ (.A(_0705_),
    .B(_0962_),
    .Y(_0978_));
 sg13g2_nand2b_1 _1944_ (.Y(_0979_),
    .B(_0704_),
    .A_N(_0962_));
 sg13g2_o21ai_1 _1945_ (.B1(net553),
    .Y(_0980_),
    .A1(\gfx.pixel_y[7] ),
    .A2(_0978_));
 sg13g2_nand2_1 _1946_ (.Y(_0981_),
    .A(_0977_),
    .B(_0980_));
 sg13g2_nor2_1 _1947_ (.A(net549),
    .B(_0968_),
    .Y(_0982_));
 sg13g2_a21oi_1 _1948_ (.A1(net549),
    .A2(_0978_),
    .Y(_0983_),
    .B1(_0982_));
 sg13g2_o21ai_1 _1949_ (.B1(_0981_),
    .Y(_0984_),
    .A1(net556),
    .A2(_0983_));
 sg13g2_nand2_1 _1950_ (.Y(_0985_),
    .A(net561),
    .B(_0984_));
 sg13g2_a21oi_1 _1951_ (.A1(net563),
    .A2(_0973_),
    .Y(_0986_),
    .B1(net516));
 sg13g2_a21oi_1 _1952_ (.A1(_0985_),
    .A2(_0986_),
    .Y(_0987_),
    .B1(_0955_));
 sg13g2_o21ai_1 _1953_ (.B1(_0987_),
    .Y(_0988_),
    .A1(_0914_),
    .A2(_0953_));
 sg13g2_and2_1 _1954_ (.A(net563),
    .B(_0955_),
    .X(_0989_));
 sg13g2_and2_1 _1955_ (.A(net561),
    .B(_0955_),
    .X(_0990_));
 sg13g2_a22oi_1 _1956_ (.Y(_0991_),
    .B1(_0990_),
    .B2(_0973_),
    .A2(_0989_),
    .A1(_0984_));
 sg13g2_and2_1 _1957_ (.A(_0988_),
    .B(_0991_),
    .X(_0992_));
 sg13g2_nand2_2 _1958_ (.Y(_0993_),
    .A(_0988_),
    .B(_0991_));
 sg13g2_nor3_1 _1959_ (.A(net508),
    .B(_0844_),
    .C(_0864_),
    .Y(_0994_));
 sg13g2_nor3_2 _1960_ (.A(net490),
    .B(net480),
    .C(_0994_),
    .Y(_0995_));
 sg13g2_nand2_1 _1961_ (.Y(_0996_),
    .A(net529),
    .B(_0789_));
 sg13g2_a21oi_1 _1962_ (.A1(net573),
    .A2(net546),
    .Y(_0997_),
    .B1(_0996_));
 sg13g2_or3_1 _1963_ (.A(net498),
    .B(_0840_),
    .C(_0997_),
    .X(_0998_));
 sg13g2_nor2_2 _1964_ (.A(net548),
    .B(_0752_),
    .Y(_0999_));
 sg13g2_and2_2 _1965_ (.A(net534),
    .B(_0999_),
    .X(_1000_));
 sg13g2_a21o_1 _1966_ (.A2(_1000_),
    .A1(net499),
    .B1(_0828_),
    .X(_1001_));
 sg13g2_a22oi_1 _1967_ (.Y(_1002_),
    .B1(_1001_),
    .B2(net454),
    .A2(_0998_),
    .A1(_0995_));
 sg13g2_nor2_1 _1968_ (.A(net529),
    .B(_0941_),
    .Y(_1003_));
 sg13g2_a21oi_1 _1969_ (.A1(net451),
    .A2(_1003_),
    .Y(_1004_),
    .B1(net461));
 sg13g2_nand2_1 _1970_ (.Y(_1005_),
    .A(net527),
    .B(_0766_));
 sg13g2_nand2_1 _1971_ (.Y(_1006_),
    .A(_0765_),
    .B(_0923_));
 sg13g2_a221oi_1 _1972_ (.B2(_1006_),
    .C1(net507),
    .B1(_1005_),
    .A1(net483),
    .Y(_1007_),
    .A2(net471));
 sg13g2_nand2_1 _1973_ (.Y(_1008_),
    .A(net572),
    .B(_0748_));
 sg13g2_nor2_2 _1974_ (.A(net526),
    .B(_1008_),
    .Y(_1009_));
 sg13g2_nand2_2 _1975_ (.Y(_1010_),
    .A(net573),
    .B(_0835_));
 sg13g2_a22oi_1 _1976_ (.Y(_1011_),
    .B1(_0814_),
    .B2(net573),
    .A2(_0774_),
    .A1(net571));
 sg13g2_nand2_1 _1977_ (.Y(_1012_),
    .A(_1010_),
    .B(_1011_));
 sg13g2_nor4_1 _1978_ (.A(net493),
    .B(net481),
    .C(net501),
    .D(_1012_),
    .Y(_1013_));
 sg13g2_nor2_2 _1979_ (.A(net538),
    .B(_0789_),
    .Y(_1014_));
 sg13g2_nor4_1 _1980_ (.A(net491),
    .B(net479),
    .C(_0847_),
    .D(_1014_),
    .Y(_1015_));
 sg13g2_nor4_2 _1981_ (.A(_0846_),
    .B(_1007_),
    .C(_1013_),
    .Y(_1016_),
    .D(_1015_));
 sg13g2_nor2b_1 _1982_ (.A(_1003_),
    .B_N(_0830_),
    .Y(_1017_));
 sg13g2_nor3_1 _1983_ (.A(net490),
    .B(net478),
    .C(_1017_),
    .Y(_1018_));
 sg13g2_nor2_2 _1984_ (.A(net547),
    .B(_0776_),
    .Y(_1019_));
 sg13g2_nand2_1 _1985_ (.Y(_1020_),
    .A(net545),
    .B(_0777_));
 sg13g2_nor2_1 _1986_ (.A(_0786_),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_nand2_2 _1987_ (.Y(_1022_),
    .A(_0787_),
    .B(_1019_));
 sg13g2_a21oi_1 _1988_ (.A1(net529),
    .A2(_1022_),
    .Y(_1023_),
    .B1(net498));
 sg13g2_nor4_1 _1989_ (.A(net492),
    .B(net478),
    .C(_1017_),
    .D(_1023_),
    .Y(_1024_));
 sg13g2_a221oi_1 _1990_ (.B2(_0751_),
    .C1(_0771_),
    .B1(net539),
    .A1(net488),
    .Y(_1025_),
    .A2(net476));
 sg13g2_nor3_1 _1991_ (.A(net466),
    .B(_1024_),
    .C(_1025_),
    .Y(_1026_));
 sg13g2_nand2_1 _1992_ (.Y(_1027_),
    .A(_0757_),
    .B(net450));
 sg13g2_a21oi_2 _1993_ (.B1(net529),
    .Y(_1028_),
    .A2(net546),
    .A1(net573));
 sg13g2_a221oi_1 _1994_ (.B2(_1028_),
    .C1(net498),
    .B1(net523),
    .A1(net529),
    .Y(_1029_),
    .A2(net546));
 sg13g2_nor2_2 _1995_ (.A(net526),
    .B(_0786_),
    .Y(_1030_));
 sg13g2_nor3_1 _1996_ (.A(net510),
    .B(_1014_),
    .C(_1030_),
    .Y(_1031_));
 sg13g2_or3_1 _1997_ (.A(net457),
    .B(_1029_),
    .C(_1031_),
    .X(_1032_));
 sg13g2_a21oi_1 _1998_ (.A1(net530),
    .A2(net548),
    .Y(_1033_),
    .B1(_0823_));
 sg13g2_nor2_2 _1999_ (.A(_0709_),
    .B(_0777_),
    .Y(_1034_));
 sg13g2_nand2_2 _2000_ (.Y(_1035_),
    .A(_0710_),
    .B(_0776_));
 sg13g2_nor2_2 _2001_ (.A(net528),
    .B(_1034_),
    .Y(_1036_));
 sg13g2_nand2_1 _2002_ (.Y(_1037_),
    .A(net523),
    .B(_1036_));
 sg13g2_o21ai_1 _2003_ (.B1(_1037_),
    .Y(_1038_),
    .A1(_0754_),
    .A2(_0996_));
 sg13g2_nand2_1 _2004_ (.Y(_1039_),
    .A(net508),
    .B(_1038_));
 sg13g2_o21ai_1 _2005_ (.B1(_1039_),
    .Y(_1040_),
    .A1(net508),
    .A2(_1033_));
 sg13g2_a21oi_1 _2006_ (.A1(net457),
    .A2(_1040_),
    .Y(_1041_),
    .B1(net461));
 sg13g2_a221oi_1 _2007_ (.B2(_1016_),
    .C1(net560),
    .B1(_1004_),
    .A1(net461),
    .Y(_1042_),
    .A2(_1002_));
 sg13g2_a221oi_1 _2008_ (.B2(_1041_),
    .C1(net563),
    .B1(_1032_),
    .A1(_1026_),
    .Y(_1043_),
    .A2(_1027_));
 sg13g2_or2_1 _2009_ (.X(_1044_),
    .B(_1043_),
    .A(_1042_));
 sg13g2_nor3_2 _2010_ (.A(net525),
    .B(_0776_),
    .C(net521),
    .Y(_1045_));
 sg13g2_and3_1 _2011_ (.X(_1046_),
    .A(net455),
    .B(net496),
    .C(_1045_));
 sg13g2_a21oi_1 _2012_ (.A1(_0891_),
    .A2(_1020_),
    .Y(_1047_),
    .B1(net535));
 sg13g2_nor3_1 _2013_ (.A(net497),
    .B(_0788_),
    .C(_1047_),
    .Y(_1048_));
 sg13g2_a221oi_1 _2014_ (.B2(_0831_),
    .C1(_1048_),
    .B1(_0755_),
    .A1(net485),
    .Y(_1049_),
    .A2(net473));
 sg13g2_nor2_2 _2015_ (.A(net547),
    .B(_0787_),
    .Y(_1050_));
 sg13g2_nor2_2 _2016_ (.A(net525),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_nor2_1 _2017_ (.A(_0895_),
    .B(_1051_),
    .Y(_1052_));
 sg13g2_nor2b_1 _2018_ (.A(_1052_),
    .B_N(_0793_),
    .Y(_1053_));
 sg13g2_or4_1 _2019_ (.A(net464),
    .B(_1046_),
    .C(_1049_),
    .D(_1053_),
    .X(_1054_));
 sg13g2_nand2_1 _2020_ (.Y(_1055_),
    .A(net528),
    .B(_1035_));
 sg13g2_o21ai_1 _2021_ (.B1(net528),
    .Y(_1056_),
    .A1(_0890_),
    .A2(_1021_));
 sg13g2_o21ai_1 _2022_ (.B1(_1056_),
    .Y(_1057_),
    .A1(net528),
    .A2(_0753_));
 sg13g2_a22oi_1 _2023_ (.Y(_1058_),
    .B1(_1057_),
    .B2(net497),
    .A2(_1055_),
    .A1(_0865_));
 sg13g2_a21oi_1 _2024_ (.A1(net454),
    .A2(_1058_),
    .Y(_1059_),
    .B1(net463));
 sg13g2_o21ai_1 _2025_ (.B1(_0793_),
    .Y(_1060_),
    .A1(_0792_),
    .A2(_1036_));
 sg13g2_nand3_1 _2026_ (.B(_0779_),
    .C(_0898_),
    .A(net456),
    .Y(_1061_));
 sg13g2_nand3_1 _2027_ (.B(_1060_),
    .C(_1061_),
    .A(_1059_),
    .Y(_1062_));
 sg13g2_a21o_1 _2028_ (.A2(_1062_),
    .A1(_1054_),
    .B1(net563),
    .X(_1063_));
 sg13g2_nor3_1 _2029_ (.A(net494),
    .B(_0814_),
    .C(_0859_),
    .Y(_1064_));
 sg13g2_nor3_1 _2030_ (.A(net494),
    .B(_0859_),
    .C(_0875_),
    .Y(_1065_));
 sg13g2_nor2_2 _2031_ (.A(net545),
    .B(_0776_),
    .Y(_1066_));
 sg13g2_nand2_2 _2032_ (.Y(_1067_),
    .A(net547),
    .B(_0777_));
 sg13g2_nor2_1 _2033_ (.A(_0786_),
    .B(_1067_),
    .Y(_1068_));
 sg13g2_nor3_1 _2034_ (.A(net504),
    .B(_0924_),
    .C(_1068_),
    .Y(_1069_));
 sg13g2_nand2_1 _2035_ (.Y(_1070_),
    .A(net526),
    .B(net523));
 sg13g2_nand2_1 _2036_ (.Y(_1071_),
    .A(_0865_),
    .B(_1070_));
 sg13g2_o21ai_1 _2037_ (.B1(net494),
    .Y(_1072_),
    .A1(_0895_),
    .A2(_1045_));
 sg13g2_nand2_1 _2038_ (.Y(_1073_),
    .A(net511),
    .B(_0861_));
 sg13g2_nand2_1 _2039_ (.Y(_1074_),
    .A(net536),
    .B(_1050_));
 sg13g2_nand4_1 _2040_ (.B(_0861_),
    .C(_0881_),
    .A(net506),
    .Y(_1075_),
    .D(_1074_));
 sg13g2_nand4_1 _2041_ (.B(net471),
    .C(_0935_),
    .A(net483),
    .Y(_1076_),
    .D(_1075_));
 sg13g2_nor2_2 _2042_ (.A(net534),
    .B(_1019_),
    .Y(_1077_));
 sg13g2_and2_1 _2043_ (.A(net535),
    .B(_0857_),
    .X(_1078_));
 sg13g2_a21oi_1 _2044_ (.A1(net515),
    .A2(_0759_),
    .Y(_1079_),
    .B1(_1078_));
 sg13g2_a22oi_1 _2045_ (.Y(_1080_),
    .B1(_1078_),
    .B2(_1067_),
    .A2(_1077_),
    .A1(_0753_));
 sg13g2_nor3_2 _2046_ (.A(_0718_),
    .B(_0758_),
    .C(_0796_),
    .Y(_1081_));
 sg13g2_nand2_1 _2047_ (.Y(_1082_),
    .A(net506),
    .B(_0797_));
 sg13g2_a22oi_1 _2048_ (.Y(_1083_),
    .B1(_1081_),
    .B2(_0938_),
    .A2(_1080_),
    .A1(net496));
 sg13g2_o21ai_1 _2049_ (.B1(_1083_),
    .Y(_1084_),
    .A1(net493),
    .A2(net481));
 sg13g2_a22oi_1 _2050_ (.Y(_1085_),
    .B1(_1071_),
    .B2(_1072_),
    .A2(net470),
    .A1(net482));
 sg13g2_nor4_1 _2051_ (.A(net489),
    .B(net477),
    .C(_1065_),
    .D(_1069_),
    .Y(_1086_));
 sg13g2_or3_1 _2052_ (.A(net464),
    .B(_1085_),
    .C(_1086_),
    .X(_1087_));
 sg13g2_nand3_1 _2053_ (.B(_1076_),
    .C(_1084_),
    .A(net464),
    .Y(_1088_));
 sg13g2_nand3_1 _2054_ (.B(_1087_),
    .C(_1088_),
    .A(net564),
    .Y(_1089_));
 sg13g2_and2_1 _2055_ (.A(_0812_),
    .B(_1089_),
    .X(_1090_));
 sg13g2_a221oi_1 _2056_ (.B2(_1090_),
    .C1(net447),
    .B1(_1063_),
    .A1(net449),
    .Y(_1091_),
    .A2(_1044_));
 sg13g2_nand2_2 _2057_ (.Y(_1092_),
    .A(_0753_),
    .B(_0823_));
 sg13g2_nor2b_1 _2058_ (.A(_0942_),
    .B_N(_1092_),
    .Y(_1093_));
 sg13g2_nor2_1 _2059_ (.A(net498),
    .B(_1093_),
    .Y(_1094_));
 sg13g2_a221oi_1 _2060_ (.B2(_0898_),
    .C1(_1094_),
    .B1(_0872_),
    .A1(net488),
    .Y(_1095_),
    .A2(net473));
 sg13g2_nor2_1 _2061_ (.A(net538),
    .B(_0790_),
    .Y(_1096_));
 sg13g2_nor3_1 _2062_ (.A(net509),
    .B(_0843_),
    .C(_1096_),
    .Y(_1097_));
 sg13g2_a21oi_1 _2063_ (.A1(net457),
    .A2(_1097_),
    .Y(_1098_),
    .B1(_1095_));
 sg13g2_a22oi_1 _2064_ (.Y(_1099_),
    .B1(_1022_),
    .B2(net539),
    .A2(_0844_),
    .A1(_0787_));
 sg13g2_nor2_1 _2065_ (.A(net508),
    .B(_1099_),
    .Y(_1100_));
 sg13g2_a221oi_1 _2066_ (.B2(_0924_),
    .C1(_1100_),
    .B1(net508),
    .A1(net485),
    .Y(_1101_),
    .A2(net476));
 sg13g2_nor4_1 _2067_ (.A(net528),
    .B(net497),
    .C(_0788_),
    .D(_1021_),
    .Y(_1102_));
 sg13g2_nor2_2 _2068_ (.A(net538),
    .B(net544),
    .Y(_1103_));
 sg13g2_nor2_2 _2069_ (.A(net532),
    .B(_0824_),
    .Y(_1104_));
 sg13g2_nor3_1 _2070_ (.A(_0790_),
    .B(_1103_),
    .C(_1104_),
    .Y(_1105_));
 sg13g2_nor2_1 _2071_ (.A(net508),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_nor4_1 _2072_ (.A(net490),
    .B(net478),
    .C(_1102_),
    .D(_1106_),
    .Y(_1107_));
 sg13g2_or3_1 _2073_ (.A(net466),
    .B(_1101_),
    .C(_1107_),
    .X(_1108_));
 sg13g2_o21ai_1 _2074_ (.B1(_1108_),
    .Y(_1109_),
    .A1(net461),
    .A2(_1098_));
 sg13g2_and3_1 _2075_ (.X(_1110_),
    .A(net498),
    .B(_0787_),
    .C(_1028_));
 sg13g2_o21ai_1 _2076_ (.B1(net454),
    .Y(_1111_),
    .A1(_0853_),
    .A2(_1110_));
 sg13g2_nand2_1 _2077_ (.Y(_1112_),
    .A(net536),
    .B(_1066_));
 sg13g2_and2_1 _2078_ (.A(net506),
    .B(_1112_),
    .X(_1113_));
 sg13g2_nor2_1 _2079_ (.A(_0766_),
    .B(_0794_),
    .Y(_1114_));
 sg13g2_nand2b_1 _2080_ (.Y(_1115_),
    .B(_1114_),
    .A_N(_0856_));
 sg13g2_nor2_1 _2081_ (.A(net538),
    .B(_0941_),
    .Y(_1116_));
 sg13g2_o21ai_1 _2082_ (.B1(_0942_),
    .Y(_1117_),
    .A1(net531),
    .A2(_1115_));
 sg13g2_a22oi_1 _2083_ (.Y(_1118_),
    .B1(_1117_),
    .B2(net499),
    .A2(_1113_),
    .A1(_0872_));
 sg13g2_a221oi_1 _2084_ (.B2(net456),
    .C1(net466),
    .B1(_1118_),
    .A1(net451),
    .Y(_1119_),
    .A2(_0836_));
 sg13g2_a21oi_1 _2085_ (.A1(_0753_),
    .A2(_1077_),
    .Y(_1120_),
    .B1(_0841_));
 sg13g2_nand3_1 _2086_ (.B(_0770_),
    .C(_0932_),
    .A(net456),
    .Y(_1121_));
 sg13g2_a221oi_1 _2087_ (.B2(_1120_),
    .C1(_0855_),
    .B1(net510),
    .A1(net485),
    .Y(_1122_),
    .A2(net473));
 sg13g2_nor2_1 _2088_ (.A(net463),
    .B(_1122_),
    .Y(_1123_));
 sg13g2_a221oi_1 _2089_ (.B2(_1123_),
    .C1(net560),
    .B1(_1121_),
    .A1(_1111_),
    .Y(_1124_),
    .A2(_1119_));
 sg13g2_a21oi_1 _2090_ (.A1(net560),
    .A2(_1109_),
    .Y(_1125_),
    .B1(_1124_));
 sg13g2_a21o_1 _2091_ (.A2(_1125_),
    .A1(net447),
    .B1(_0920_),
    .X(_1126_));
 sg13g2_nor2_1 _2092_ (.A(_0956_),
    .B(_0961_),
    .Y(_1127_));
 sg13g2_inv_1 _2093_ (.Y(_1128_),
    .A(_1127_));
 sg13g2_nand3_1 _2094_ (.B(_0957_),
    .C(_0962_),
    .A(net552),
    .Y(_1129_));
 sg13g2_nand3_1 _2095_ (.B(_0011_),
    .C(_0961_),
    .A(net567),
    .Y(_1130_));
 sg13g2_nand2_1 _2096_ (.Y(_1131_),
    .A(net549),
    .B(_1130_));
 sg13g2_nor3_1 _2097_ (.A(net568),
    .B(_0524_),
    .C(_0531_),
    .Y(_1132_));
 sg13g2_a21oi_1 _2098_ (.A1(_0011_),
    .A2(_0967_),
    .Y(_1133_),
    .B1(_1131_));
 sg13g2_a21oi_1 _2099_ (.A1(net571),
    .A2(net559),
    .Y(_1134_),
    .B1(_0704_));
 sg13g2_o21ai_1 _2100_ (.B1(net556),
    .Y(_1135_),
    .A1(net551),
    .A2(_1134_));
 sg13g2_nand3_1 _2101_ (.B(net559),
    .C(_1127_),
    .A(_0705_),
    .Y(_1136_));
 sg13g2_nand2_1 _2102_ (.Y(_1137_),
    .A(_0704_),
    .B(_0968_));
 sg13g2_nand3_1 _2103_ (.B(_0958_),
    .C(_0968_),
    .A(_0704_),
    .Y(_1138_));
 sg13g2_nand2_1 _2104_ (.Y(_1139_),
    .A(_1136_),
    .B(_1138_));
 sg13g2_nor2_1 _2105_ (.A(_1133_),
    .B(_1135_),
    .Y(_1140_));
 sg13g2_a22oi_1 _2106_ (.Y(_1141_),
    .B1(_1140_),
    .B2(_1129_),
    .A2(_1139_),
    .A1(_0963_));
 sg13g2_and2_1 _2107_ (.A(net549),
    .B(_0969_),
    .X(_1142_));
 sg13g2_nand3_1 _2108_ (.B(_0957_),
    .C(_0962_),
    .A(_0704_),
    .Y(_1143_));
 sg13g2_and3_1 _2109_ (.X(_1144_),
    .A(_0662_),
    .B(_1130_),
    .C(_1143_));
 sg13g2_nand2b_1 _2110_ (.Y(_1145_),
    .B(_0961_),
    .A_N(net567));
 sg13g2_nor2_1 _2111_ (.A(net567),
    .B(_1127_),
    .Y(_1146_));
 sg13g2_o21ai_1 _2112_ (.B1(net565),
    .Y(_1147_),
    .A1(net567),
    .A2(_1128_));
 sg13g2_a21oi_1 _2113_ (.A1(_1137_),
    .A2(_1147_),
    .Y(_1148_),
    .B1(net549));
 sg13g2_a21oi_1 _2114_ (.A1(_0011_),
    .A2(_0962_),
    .Y(_1149_),
    .B1(net553));
 sg13g2_nor3_1 _2115_ (.A(net554),
    .B(_1148_),
    .C(_1149_),
    .Y(_1150_));
 sg13g2_a21oi_1 _2116_ (.A1(_1142_),
    .A2(_1144_),
    .Y(_1151_),
    .B1(_1150_));
 sg13g2_nand2_1 _2117_ (.Y(_1152_),
    .A(net563),
    .B(_1151_));
 sg13g2_a21oi_1 _2118_ (.A1(net561),
    .A2(_1141_),
    .Y(_1153_),
    .B1(net516));
 sg13g2_a21oi_1 _2119_ (.A1(_1152_),
    .A2(_1153_),
    .Y(_1154_),
    .B1(_0955_));
 sg13g2_o21ai_1 _2120_ (.B1(_1154_),
    .Y(_1155_),
    .A1(_1091_),
    .A2(_1126_));
 sg13g2_and2_1 _2121_ (.A(_0989_),
    .B(_1141_),
    .X(_1156_));
 sg13g2_a21o_1 _2122_ (.A2(_1151_),
    .A1(_0990_),
    .B1(_1156_),
    .X(_1157_));
 sg13g2_inv_1 _2123_ (.Y(_1158_),
    .A(_1157_));
 sg13g2_and2_2 _2124_ (.A(_1155_),
    .B(_1158_),
    .X(_1159_));
 sg13g2_nand2_2 _2125_ (.Y(_1160_),
    .A(_1155_),
    .B(_1158_));
 sg13g2_nor3_1 _2126_ (.A(net533),
    .B(_0784_),
    .C(_1034_),
    .Y(_1161_));
 sg13g2_nor2_1 _2127_ (.A(_1051_),
    .B(_1161_),
    .Y(_1162_));
 sg13g2_nor2_1 _2128_ (.A(_0777_),
    .B(_0930_),
    .Y(_1163_));
 sg13g2_nand2_1 _2129_ (.Y(_1164_),
    .A(net458),
    .B(_1163_));
 sg13g2_a221oi_1 _2130_ (.B2(net525),
    .C1(_1050_),
    .B1(_1035_),
    .A1(_0765_),
    .Y(_1165_),
    .A2(net521));
 sg13g2_nand3_1 _2131_ (.B(_0795_),
    .C(net544),
    .A(net531),
    .Y(_1166_));
 sg13g2_nand4_1 _2132_ (.B(_0793_),
    .C(net523),
    .A(net526),
    .Y(_1167_),
    .D(net544));
 sg13g2_a22oi_1 _2133_ (.Y(_1168_),
    .B1(_1165_),
    .B2(net450),
    .A2(_1162_),
    .A1(_0783_));
 sg13g2_nand4_1 _2134_ (.B(_1164_),
    .C(_1167_),
    .A(net464),
    .Y(_1169_),
    .D(_1168_));
 sg13g2_o21ai_1 _2135_ (.B1(_0887_),
    .Y(_1170_),
    .A1(_0845_),
    .A2(_1050_));
 sg13g2_nand2_2 _2136_ (.Y(_1171_),
    .A(net547),
    .B(_0787_));
 sg13g2_nand2_1 _2137_ (.Y(_1172_),
    .A(_1036_),
    .B(_1171_));
 sg13g2_a22oi_1 _2138_ (.Y(_1173_),
    .B1(_1172_),
    .B2(_0830_),
    .A2(_1035_),
    .A1(_0816_));
 sg13g2_nor3_1 _2139_ (.A(net489),
    .B(net477),
    .C(_1173_),
    .Y(_1174_));
 sg13g2_nand2_1 _2140_ (.Y(_1175_),
    .A(net525),
    .B(_0778_));
 sg13g2_nor2b_1 _2141_ (.A(_1068_),
    .B_N(_1175_),
    .Y(_1176_));
 sg13g2_a221oi_1 _2142_ (.B2(net450),
    .C1(_1174_),
    .B1(_1176_),
    .A1(_0783_),
    .Y(_1177_),
    .A2(_1170_));
 sg13g2_a21oi_1 _2143_ (.A1(net459),
    .A2(_1177_),
    .Y(_1178_),
    .B1(net449));
 sg13g2_o21ai_1 _2144_ (.B1(net497),
    .Y(_1179_),
    .A1(_0869_),
    .A2(_1021_));
 sg13g2_a21oi_1 _2145_ (.A1(_1073_),
    .A2(_1179_),
    .Y(_1180_),
    .B1(_0781_));
 sg13g2_a21oi_1 _2146_ (.A1(net504),
    .A2(_1070_),
    .Y(_1181_),
    .B1(_0830_));
 sg13g2_a221oi_1 _2147_ (.B2(_0819_),
    .C1(_1181_),
    .B1(net494),
    .A1(net482),
    .Y(_1182_),
    .A2(net470));
 sg13g2_o21ai_1 _2148_ (.B1(net464),
    .Y(_1183_),
    .A1(_1180_),
    .A2(_1182_));
 sg13g2_o21ai_1 _2149_ (.B1(_0930_),
    .Y(_1184_),
    .A1(_0757_),
    .A2(_1082_));
 sg13g2_nor3_1 _2150_ (.A(net453),
    .B(_0926_),
    .C(_1184_),
    .Y(_1185_));
 sg13g2_nor2_1 _2151_ (.A(net533),
    .B(_1068_),
    .Y(_1186_));
 sg13g2_nor3_1 _2152_ (.A(net505),
    .B(_0819_),
    .C(_1186_),
    .Y(_1187_));
 sg13g2_a221oi_1 _2153_ (.B2(_0862_),
    .C1(_1187_),
    .B1(net504),
    .A1(net482),
    .Y(_1188_),
    .A2(net470));
 sg13g2_or4_1 _2154_ (.A(net465),
    .B(_0846_),
    .C(_1185_),
    .D(_1188_),
    .X(_1189_));
 sg13g2_nand3_1 _2155_ (.B(_1183_),
    .C(_1189_),
    .A(net449),
    .Y(_1190_));
 sg13g2_a21oi_1 _2156_ (.A1(_1169_),
    .A2(_1178_),
    .Y(_1191_),
    .B1(net564));
 sg13g2_nand2_1 _2157_ (.Y(_1192_),
    .A(net524),
    .B(_1175_));
 sg13g2_nand2_1 _2158_ (.Y(_1193_),
    .A(net505),
    .B(_1192_));
 sg13g2_nor4_1 _2159_ (.A(net527),
    .B(net495),
    .C(_0999_),
    .D(_1066_),
    .Y(_1194_));
 sg13g2_nor2_1 _2160_ (.A(_1110_),
    .B(_1194_),
    .Y(_1195_));
 sg13g2_a221oi_1 _2161_ (.B2(net455),
    .C1(net459),
    .B1(_1195_),
    .A1(_0927_),
    .Y(_1196_),
    .A2(_1193_));
 sg13g2_nand2_1 _2162_ (.Y(_1197_),
    .A(_0770_),
    .B(_0820_));
 sg13g2_nand3_1 _2163_ (.B(_0778_),
    .C(_0789_),
    .A(net524),
    .Y(_1198_));
 sg13g2_a221oi_1 _2164_ (.B2(net504),
    .C1(_0841_),
    .B1(_1198_),
    .A1(net526),
    .Y(_1199_),
    .A2(_0778_));
 sg13g2_a221oi_1 _2165_ (.B2(net453),
    .C1(net464),
    .B1(_1199_),
    .A1(_0829_),
    .Y(_1200_),
    .A2(_1197_));
 sg13g2_o21ai_1 _2166_ (.B1(net449),
    .Y(_1201_),
    .A1(_1196_),
    .A2(_1200_));
 sg13g2_nor4_2 _2167_ (.A(_0774_),
    .B(_0840_),
    .C(_0871_),
    .Y(_1202_),
    .D(_1009_));
 sg13g2_nand2_1 _2168_ (.Y(_1203_),
    .A(_0778_),
    .B(_1051_));
 sg13g2_nand2_1 _2169_ (.Y(_1204_),
    .A(net525),
    .B(_1171_));
 sg13g2_nor2_1 _2170_ (.A(_0863_),
    .B(_1077_),
    .Y(_1205_));
 sg13g2_mux4_1 _2171_ (.S0(net503),
    .A0(_1202_),
    .A1(_1204_),
    .A2(_1205_),
    .A3(_1203_),
    .S1(net452),
    .X(_1206_));
 sg13g2_a221oi_1 _2172_ (.B2(_0785_),
    .C1(net494),
    .B1(_1035_),
    .A1(net525),
    .Y(_1207_),
    .A2(net523));
 sg13g2_a21oi_1 _2173_ (.A1(_1079_),
    .A2(_1204_),
    .Y(_1208_),
    .B1(_1207_));
 sg13g2_or2_1 _2174_ (.X(_1209_),
    .B(_1208_),
    .A(net455));
 sg13g2_nor2_2 _2175_ (.A(net572),
    .B(_0870_),
    .Y(_1210_));
 sg13g2_nor2_1 _2176_ (.A(net504),
    .B(_1210_),
    .Y(_1211_));
 sg13g2_a21oi_1 _2177_ (.A1(net503),
    .A2(_1192_),
    .Y(_1212_),
    .B1(_1210_));
 sg13g2_a21oi_1 _2178_ (.A1(net503),
    .A2(_1210_),
    .Y(_1213_),
    .B1(_1212_));
 sg13g2_a21oi_1 _2179_ (.A1(net455),
    .A2(_1213_),
    .Y(_1214_),
    .B1(net459));
 sg13g2_a221oi_1 _2180_ (.B2(_1214_),
    .C1(net449),
    .B1(_1209_),
    .A1(net459),
    .Y(_1215_),
    .A2(_1206_));
 sg13g2_nor2_1 _2181_ (.A(net562),
    .B(_1215_),
    .Y(_1216_));
 sg13g2_a221oi_1 _2182_ (.B2(_1216_),
    .C1(net448),
    .B1(_1201_),
    .A1(_1190_),
    .Y(_1217_),
    .A2(_1191_));
 sg13g2_a21oi_2 _2183_ (.B1(net533),
    .Y(_1218_),
    .A2(net544),
    .A1(_0785_));
 sg13g2_nor3_2 _2184_ (.A(net510),
    .B(_0864_),
    .C(_1218_),
    .Y(_1219_));
 sg13g2_nor4_1 _2185_ (.A(net491),
    .B(net479),
    .C(_0828_),
    .D(_1219_),
    .Y(_1220_));
 sg13g2_nand2_2 _2186_ (.Y(_1221_),
    .A(net533),
    .B(_0785_));
 sg13g2_nor2_1 _2187_ (.A(_0856_),
    .B(_1221_),
    .Y(_1222_));
 sg13g2_and2_1 _2188_ (.A(_0830_),
    .B(_0839_),
    .X(_1223_));
 sg13g2_nor4_1 _2189_ (.A(net492),
    .B(net480),
    .C(_0828_),
    .D(_1223_),
    .Y(_1224_));
 sg13g2_nor2_2 _2190_ (.A(_1019_),
    .B(_1221_),
    .Y(_1225_));
 sg13g2_nand2b_2 _2191_ (.Y(_1226_),
    .B(net506),
    .A_N(_1225_));
 sg13g2_nor2_1 _2192_ (.A(_0835_),
    .B(_0997_),
    .Y(_1227_));
 sg13g2_a22oi_1 _2193_ (.Y(_1228_),
    .B1(_1226_),
    .B2(_1227_),
    .A2(net475),
    .A1(net486));
 sg13g2_nor2_1 _2194_ (.A(_0756_),
    .B(net512),
    .Y(_1229_));
 sg13g2_nor4_1 _2195_ (.A(net491),
    .B(net479),
    .C(_0921_),
    .D(_1229_),
    .Y(_1230_));
 sg13g2_a221oi_1 _2196_ (.B2(_0928_),
    .C1(_0926_),
    .B1(_0870_),
    .A1(net483),
    .Y(_1231_),
    .A2(net471));
 sg13g2_nand4_1 _2197_ (.B(net474),
    .C(_0827_),
    .A(net486),
    .Y(_1232_),
    .D(_0832_));
 sg13g2_o21ai_1 _2198_ (.B1(_0839_),
    .Y(_1233_),
    .A1(net540),
    .A2(_0753_));
 sg13g2_a221oi_1 _2199_ (.B2(_1233_),
    .C1(_0770_),
    .B1(net512),
    .A1(net486),
    .Y(_1234_),
    .A2(net474));
 sg13g2_o21ai_1 _2200_ (.B1(net462),
    .Y(_1235_),
    .A1(_1224_),
    .A2(_1228_));
 sg13g2_o21ai_1 _2201_ (.B1(net467),
    .Y(_1236_),
    .A1(_1230_),
    .A2(_1231_));
 sg13g2_nand3_1 _2202_ (.B(_1235_),
    .C(_1236_),
    .A(net561),
    .Y(_1237_));
 sg13g2_o21ai_1 _2203_ (.B1(_0791_),
    .Y(_1238_),
    .A1(_0856_),
    .A2(_1221_));
 sg13g2_o21ai_1 _2204_ (.B1(net497),
    .Y(_1239_),
    .A1(_1103_),
    .A2(_1238_));
 sg13g2_a22oi_1 _2205_ (.Y(_1240_),
    .B1(_1073_),
    .B2(_1239_),
    .A2(net474),
    .A1(net487));
 sg13g2_o21ai_1 _2206_ (.B1(net463),
    .Y(_1241_),
    .A1(_1220_),
    .A2(_1240_));
 sg13g2_nand3b_1 _2207_ (.B(net466),
    .C(_1232_),
    .Y(_1242_),
    .A_N(_1234_));
 sg13g2_nand3_1 _2208_ (.B(_1241_),
    .C(_1242_),
    .A(\gfx.frame_counter[4] ),
    .Y(_1243_));
 sg13g2_nand3_1 _2209_ (.B(_1237_),
    .C(_1243_),
    .A(net447),
    .Y(_1244_));
 sg13g2_nand2_1 _2210_ (.Y(_1245_),
    .A(net516),
    .B(_1244_));
 sg13g2_o21ai_1 _2211_ (.B1(_0964_),
    .Y(_1246_),
    .A1(net552),
    .A2(_0979_));
 sg13g2_o21ai_1 _2212_ (.B1(_1246_),
    .Y(_1247_),
    .A1(_0966_),
    .A2(_0971_));
 sg13g2_nand2_1 _2213_ (.Y(_1248_),
    .A(net563),
    .B(_1247_));
 sg13g2_o21ai_1 _2214_ (.B1(net554),
    .Y(_1249_),
    .A1(net549),
    .A2(_0967_));
 sg13g2_inv_1 _2215_ (.Y(_1250_),
    .A(_1249_));
 sg13g2_nand2_1 _2216_ (.Y(_1251_),
    .A(net550),
    .B(_1137_));
 sg13g2_o21ai_1 _2217_ (.B1(net552),
    .Y(_1252_),
    .A1(_0978_),
    .A2(_1132_));
 sg13g2_a22oi_1 _2218_ (.Y(_1253_),
    .B1(_1252_),
    .B2(_0977_),
    .A2(_1251_),
    .A1(_1250_));
 sg13g2_a21oi_1 _2219_ (.A1(net560),
    .A2(_1253_),
    .Y(_1254_),
    .B1(net516));
 sg13g2_a21oi_1 _2220_ (.A1(_1248_),
    .A2(_1254_),
    .Y(_1255_),
    .B1(_0955_));
 sg13g2_o21ai_1 _2221_ (.B1(_1255_),
    .Y(_1256_),
    .A1(_1217_),
    .A2(_1245_));
 sg13g2_a22oi_1 _2222_ (.Y(_1257_),
    .B1(_1253_),
    .B2(_0989_),
    .A2(_1247_),
    .A1(_0990_));
 sg13g2_and2_1 _2223_ (.A(net445),
    .B(net468),
    .X(_1258_));
 sg13g2_nand2_1 _2224_ (.Y(_1259_),
    .A(net445),
    .B(net468));
 sg13g2_and2_2 _2225_ (.A(\gfx.bitmap_x[0] ),
    .B(_0919_),
    .X(_1260_));
 sg13g2_nand2_2 _2226_ (.Y(_1261_),
    .A(\gfx.bitmap_x[0] ),
    .B(net516));
 sg13g2_nand2_1 _2227_ (.Y(_1262_),
    .A(_0755_),
    .B(net503));
 sg13g2_a221oi_1 _2228_ (.B2(net545),
    .C1(_1262_),
    .B1(net533),
    .A1(net482),
    .Y(_1263_),
    .A2(net470));
 sg13g2_nor2_1 _2229_ (.A(net524),
    .B(_1030_),
    .Y(_1264_));
 sg13g2_mux2_1 _2230_ (.A0(_1225_),
    .A1(_1264_),
    .S(net503),
    .X(_1265_));
 sg13g2_nor3_1 _2231_ (.A(net489),
    .B(net477),
    .C(_1265_),
    .Y(_1266_));
 sg13g2_a221oi_1 _2232_ (.B2(_0870_),
    .C1(net503),
    .B1(_0775_),
    .A1(net482),
    .Y(_1267_),
    .A2(net470));
 sg13g2_or3_1 _2233_ (.A(_1263_),
    .B(_1266_),
    .C(_1267_),
    .X(_1268_));
 sg13g2_nor2_1 _2234_ (.A(net503),
    .B(_0860_),
    .Y(_1269_));
 sg13g2_o21ai_1 _2235_ (.B1(_1269_),
    .Y(_1270_),
    .A1(_0845_),
    .A2(_0999_));
 sg13g2_nand3_1 _2236_ (.B(_0858_),
    .C(_1035_),
    .A(net503),
    .Y(_1271_));
 sg13g2_nand3_1 _2237_ (.B(_1270_),
    .C(_1271_),
    .A(net452),
    .Y(_1272_));
 sg13g2_a221oi_1 _2238_ (.B2(net533),
    .C1(_0784_),
    .B1(_1035_),
    .A1(net494),
    .Y(_1273_),
    .A2(_0778_));
 sg13g2_a21oi_1 _2239_ (.A1(net455),
    .A2(_1273_),
    .Y(_1274_),
    .B1(net459));
 sg13g2_a221oi_1 _2240_ (.B2(_1274_),
    .C1(net449),
    .B1(_1272_),
    .A1(net459),
    .Y(_1275_),
    .A2(_1268_));
 sg13g2_nand2_1 _2241_ (.Y(_1276_),
    .A(_0874_),
    .B(_0924_));
 sg13g2_nor3_1 _2242_ (.A(net495),
    .B(_0923_),
    .C(_1077_),
    .Y(_1277_));
 sg13g2_a21oi_1 _2243_ (.A1(_0797_),
    .A2(_1010_),
    .Y(_1278_),
    .B1(net507));
 sg13g2_or3_1 _2244_ (.A(net452),
    .B(_1277_),
    .C(_1278_),
    .X(_1279_));
 sg13g2_or3_1 _2245_ (.A(net527),
    .B(_0750_),
    .C(net521),
    .X(_1280_));
 sg13g2_a221oi_1 _2246_ (.B2(net450),
    .C1(net464),
    .B1(_1280_),
    .A1(_0783_),
    .Y(_1281_),
    .A2(_1276_));
 sg13g2_o21ai_1 _2247_ (.B1(_0858_),
    .Y(_1282_),
    .A1(_1050_),
    .A2(_1204_));
 sg13g2_or2_1 _2248_ (.X(_1283_),
    .B(_1282_),
    .A(net495));
 sg13g2_nor2_1 _2249_ (.A(_0838_),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_nor4_1 _2250_ (.A(net506),
    .B(_0819_),
    .C(_0895_),
    .D(_1000_),
    .Y(_1285_));
 sg13g2_nand4_1 _2251_ (.B(_0815_),
    .C(_0824_),
    .A(net511),
    .Y(_1286_),
    .D(_0861_));
 sg13g2_nand2_1 _2252_ (.Y(_1287_),
    .A(net544),
    .B(_1171_));
 sg13g2_nor2_1 _2253_ (.A(net538),
    .B(_1287_),
    .Y(_1288_));
 sg13g2_nor2_1 _2254_ (.A(_1051_),
    .B(_1288_),
    .Y(_1289_));
 sg13g2_o21ai_1 _2255_ (.B1(net455),
    .Y(_1290_),
    .A1(_1284_),
    .A2(_1285_));
 sg13g2_o21ai_1 _2256_ (.B1(_1286_),
    .Y(_1291_),
    .A1(_0847_),
    .A2(_1289_));
 sg13g2_a21oi_1 _2257_ (.A1(net452),
    .A2(_1291_),
    .Y(_0105_),
    .B1(net459));
 sg13g2_a221oi_1 _2258_ (.B2(_0105_),
    .C1(_0812_),
    .B1(_1290_),
    .A1(_1279_),
    .Y(_0106_),
    .A2(_1281_));
 sg13g2_or3_1 _2259_ (.A(net448),
    .B(_1275_),
    .C(_0106_),
    .X(_0107_));
 sg13g2_a21oi_1 _2260_ (.A1(net538),
    .A2(_0790_),
    .Y(_0108_),
    .B1(_1103_));
 sg13g2_nor3_1 _2261_ (.A(net489),
    .B(net477),
    .C(_0108_),
    .Y(_0109_));
 sg13g2_a221oi_1 _2262_ (.B2(net572),
    .C1(_0784_),
    .B1(net545),
    .A1(net482),
    .Y(_0110_),
    .A2(net470));
 sg13g2_or3_1 _2263_ (.A(net504),
    .B(_0109_),
    .C(_0110_),
    .X(_0111_));
 sg13g2_nor2_1 _2264_ (.A(_1034_),
    .B(_1221_),
    .Y(_0112_));
 sg13g2_and2_1 _2265_ (.A(net508),
    .B(_1028_),
    .X(_0113_));
 sg13g2_and2_1 _2266_ (.A(_1171_),
    .B(_0113_),
    .X(_0114_));
 sg13g2_a221oi_1 _2267_ (.B2(net458),
    .C1(net464),
    .B1(_0114_),
    .A1(net450),
    .Y(_0115_),
    .A2(_0112_));
 sg13g2_o21ai_1 _2268_ (.B1(_1092_),
    .Y(_0116_),
    .A1(net537),
    .A2(net558));
 sg13g2_a221oi_1 _2269_ (.B2(_0761_),
    .C1(_0116_),
    .B1(_0760_),
    .A1(net484),
    .Y(_0117_),
    .A2(net471));
 sg13g2_nand2_1 _2270_ (.Y(_0118_),
    .A(net522),
    .B(_0853_));
 sg13g2_a21oi_1 _2271_ (.A1(_0932_),
    .A2(_0118_),
    .Y(_0119_),
    .B1(net511));
 sg13g2_nor4_1 _2272_ (.A(net491),
    .B(net479),
    .C(_0921_),
    .D(_0119_),
    .Y(_0120_));
 sg13g2_a221oi_1 _2273_ (.B2(_1166_),
    .C1(net511),
    .B1(_0869_),
    .A1(net483),
    .Y(_0121_),
    .A2(net471));
 sg13g2_or3_1 _2274_ (.A(_0117_),
    .B(_0120_),
    .C(_0121_),
    .X(_0122_));
 sg13g2_a22oi_1 _2275_ (.Y(_0123_),
    .B1(_0122_),
    .B2(net465),
    .A2(_0115_),
    .A1(_0111_));
 sg13g2_a21oi_1 _2276_ (.A1(net448),
    .A2(_0123_),
    .Y(_0124_),
    .B1(net564));
 sg13g2_a21oi_1 _2277_ (.A1(net536),
    .A2(_0856_),
    .Y(_0125_),
    .B1(net521));
 sg13g2_nand4_1 _2278_ (.B(_0870_),
    .C(_0935_),
    .A(net455),
    .Y(_0126_),
    .D(_0125_));
 sg13g2_nor2_1 _2279_ (.A(_0856_),
    .B(_1066_),
    .Y(_0127_));
 sg13g2_a22oi_1 _2280_ (.Y(_0128_),
    .B1(_0127_),
    .B2(net536),
    .A2(_1077_),
    .A1(_0785_));
 sg13g2_a22oi_1 _2281_ (.Y(_0129_),
    .B1(_0128_),
    .B2(net495),
    .A2(_1112_),
    .A1(_1081_));
 sg13g2_a21oi_1 _2282_ (.A1(net452),
    .A2(_0129_),
    .Y(_0130_),
    .B1(net460));
 sg13g2_a22oi_1 _2283_ (.Y(_0131_),
    .B1(_0891_),
    .B2(net527),
    .A2(_0759_),
    .A1(net515));
 sg13g2_nor3_1 _2284_ (.A(net494),
    .B(_0895_),
    .C(_1222_),
    .Y(_0132_));
 sg13g2_a21o_1 _2285_ (.A2(_0131_),
    .A1(net524),
    .B1(_0132_),
    .X(_0133_));
 sg13g2_nor4_1 _2286_ (.A(net489),
    .B(net477),
    .C(_1064_),
    .D(_1269_),
    .Y(_0134_));
 sg13g2_a21oi_1 _2287_ (.A1(net452),
    .A2(_0133_),
    .Y(_0135_),
    .B1(_0134_));
 sg13g2_a221oi_1 _2288_ (.B2(net459),
    .C1(net449),
    .B1(_0135_),
    .A1(_0126_),
    .Y(_0136_),
    .A2(_0130_));
 sg13g2_a21oi_1 _2289_ (.A1(net572),
    .A2(_0814_),
    .Y(_0137_),
    .B1(_1066_));
 sg13g2_mux2_1 _2290_ (.A0(_1225_),
    .A1(_0137_),
    .S(net506),
    .X(_0138_));
 sg13g2_nor4_1 _2291_ (.A(net493),
    .B(net481),
    .C(_0926_),
    .D(_0138_),
    .Y(_0139_));
 sg13g2_nand2_1 _2292_ (.Y(_0140_),
    .A(_0845_),
    .B(_1010_));
 sg13g2_a22oi_1 _2293_ (.Y(_0141_),
    .B1(_0140_),
    .B2(net507),
    .A2(_0131_),
    .A1(_1006_));
 sg13g2_a21oi_1 _2294_ (.A1(net483),
    .A2(net471),
    .Y(_0142_),
    .B1(_0141_));
 sg13g2_or2_1 _2295_ (.X(_0143_),
    .B(_0142_),
    .A(_0139_));
 sg13g2_nand3_1 _2296_ (.B(_0778_),
    .C(_0820_),
    .A(net495),
    .Y(_0144_));
 sg13g2_a21o_1 _2297_ (.A2(_0144_),
    .A1(_1283_),
    .B1(net452),
    .X(_0145_));
 sg13g2_a22oi_1 _2298_ (.Y(_0146_),
    .B1(_1114_),
    .B2(_0828_),
    .A2(_0836_),
    .A1(_0770_));
 sg13g2_a21oi_1 _2299_ (.A1(net452),
    .A2(_0146_),
    .Y(_0147_),
    .B1(net465));
 sg13g2_a221oi_1 _2300_ (.B2(_0147_),
    .C1(_0812_),
    .B1(_0145_),
    .A1(net465),
    .Y(_0148_),
    .A2(_0143_));
 sg13g2_or3_1 _2301_ (.A(net448),
    .B(_0136_),
    .C(_0148_),
    .X(_0149_));
 sg13g2_nor2b_1 _2302_ (.A(_1051_),
    .B_N(_0770_),
    .Y(_0150_));
 sg13g2_nor2_1 _2303_ (.A(net496),
    .B(_1092_),
    .Y(_0151_));
 sg13g2_nor4_1 _2304_ (.A(net489),
    .B(net477),
    .C(_0150_),
    .D(_0151_),
    .Y(_0152_));
 sg13g2_nor3_1 _2305_ (.A(net536),
    .B(_0750_),
    .C(net521),
    .Y(_0153_));
 sg13g2_nor3_1 _2306_ (.A(net495),
    .B(_0863_),
    .C(_0153_),
    .Y(_0154_));
 sg13g2_a221oi_1 _2307_ (.B2(net453),
    .C1(_0152_),
    .B1(_0154_),
    .A1(_0783_),
    .Y(_0155_),
    .A2(_0118_));
 sg13g2_nor4_1 _2308_ (.A(net490),
    .B(net478),
    .C(_0899_),
    .D(_1014_),
    .Y(_0156_));
 sg13g2_nor3_1 _2309_ (.A(_0718_),
    .B(_0758_),
    .C(_1171_),
    .Y(_0157_));
 sg13g2_nand2_1 _2310_ (.Y(_0158_),
    .A(_0815_),
    .B(_1287_));
 sg13g2_a21o_1 _2311_ (.A2(_0158_),
    .A1(_0855_),
    .B1(_0157_),
    .X(_0159_));
 sg13g2_a221oi_1 _2312_ (.B2(_0924_),
    .C1(_0159_),
    .B1(net510),
    .A1(net482),
    .Y(_0160_),
    .A2(net470));
 sg13g2_nor3_1 _2313_ (.A(_0859_),
    .B(_1009_),
    .C(_1210_),
    .Y(_0161_));
 sg13g2_nor4_1 _2314_ (.A(net489),
    .B(net477),
    .C(net494),
    .D(_0161_),
    .Y(_0162_));
 sg13g2_or3_1 _2315_ (.A(_0156_),
    .B(_0160_),
    .C(_0162_),
    .X(_0163_));
 sg13g2_mux2_1 _2316_ (.A0(_0155_),
    .A1(_0163_),
    .S(net460),
    .X(_0164_));
 sg13g2_a21oi_1 _2317_ (.A1(net448),
    .A2(_0164_),
    .Y(_0165_),
    .B1(net562));
 sg13g2_a221oi_1 _2318_ (.B2(_0165_),
    .C1(_0920_),
    .B1(_0149_),
    .A1(_0107_),
    .Y(_0166_),
    .A2(_0124_));
 sg13g2_nor2_1 _2319_ (.A(net516),
    .B(_0955_),
    .Y(_0167_));
 sg13g2_a21oi_2 _2320_ (.B1(_0989_),
    .Y(_0168_),
    .A2(_0167_),
    .A1(net560));
 sg13g2_nand4_1 _2321_ (.B(_1130_),
    .C(_1136_),
    .A(net550),
    .Y(_0169_),
    .D(_1143_));
 sg13g2_nand2b_1 _2322_ (.Y(_0170_),
    .B(net559),
    .A_N(_0013_));
 sg13g2_nand3_1 _2323_ (.B(_1145_),
    .C(_0170_),
    .A(_0705_),
    .Y(_0171_));
 sg13g2_nand3_1 _2324_ (.B(_1143_),
    .C(_0171_),
    .A(net553),
    .Y(_0172_));
 sg13g2_a21oi_1 _2325_ (.A1(_0011_),
    .A2(_1146_),
    .Y(_0173_),
    .B1(_1131_));
 sg13g2_nor2_1 _2326_ (.A(net554),
    .B(_0173_),
    .Y(_0174_));
 sg13g2_a22oi_1 _2327_ (.Y(_0175_),
    .B1(_0172_),
    .B2(_0174_),
    .A2(_0169_),
    .A1(_1250_));
 sg13g2_a21o_1 _2328_ (.A2(_0167_),
    .A1(net563),
    .B1(_0990_),
    .X(_0176_));
 sg13g2_o21ai_1 _2329_ (.B1(_0975_),
    .Y(_0177_),
    .A1(net571),
    .A2(net559));
 sg13g2_a21oi_1 _2330_ (.A1(_0704_),
    .A2(_1146_),
    .Y(_0178_),
    .B1(net550));
 sg13g2_a221oi_1 _2331_ (.B2(_0178_),
    .C1(net554),
    .B1(_0177_),
    .A1(net550),
    .Y(_0179_),
    .A2(_1136_));
 sg13g2_nand4_1 _2332_ (.B(net567),
    .C(\gfx.pixel_y[7] ),
    .A(_0523_),
    .Y(_0180_),
    .D(_0531_));
 sg13g2_a21oi_1 _2333_ (.A1(_1129_),
    .A2(_0180_),
    .Y(_0181_),
    .B1(net556));
 sg13g2_o21ai_1 _2334_ (.B1(_0176_),
    .Y(_0182_),
    .A1(_0179_),
    .A2(_0181_));
 sg13g2_o21ai_1 _2335_ (.B1(_0182_),
    .Y(_0183_),
    .A1(_0168_),
    .A2(_0175_));
 sg13g2_nor2_2 _2336_ (.A(_0166_),
    .B(_0183_),
    .Y(_0184_));
 sg13g2_or2_2 _2337_ (.X(_0185_),
    .B(_0183_),
    .A(_0166_));
 sg13g2_nand2_2 _2338_ (.Y(_0186_),
    .A(net523),
    .B(_1022_));
 sg13g2_inv_1 _2339_ (.Y(_0187_),
    .A(_0186_));
 sg13g2_a221oi_1 _2340_ (.B2(_0187_),
    .C1(net510),
    .B1(_1055_),
    .A1(net485),
    .Y(_0188_),
    .A2(net473));
 sg13g2_nand2_1 _2341_ (.Y(_0189_),
    .A(_0815_),
    .B(_0865_));
 sg13g2_a22oi_1 _2342_ (.Y(_0190_),
    .B1(_0923_),
    .B2(_1008_),
    .A2(_0789_),
    .A1(net504));
 sg13g2_nor3_1 _2343_ (.A(net489),
    .B(net477),
    .C(_0190_),
    .Y(_0191_));
 sg13g2_a21oi_1 _2344_ (.A1(net485),
    .A2(net473),
    .Y(_0192_),
    .B1(_0189_));
 sg13g2_or3_1 _2345_ (.A(_0188_),
    .B(_0191_),
    .C(_0192_),
    .X(_0193_));
 sg13g2_or4_1 _2346_ (.A(net453),
    .B(_0882_),
    .C(_1051_),
    .D(_1211_),
    .X(_0194_));
 sg13g2_o21ai_1 _2347_ (.B1(net534),
    .Y(_0195_),
    .A1(_0890_),
    .A2(_1019_));
 sg13g2_a21oi_1 _2348_ (.A1(net505),
    .A2(_0195_),
    .Y(_0196_),
    .B1(_1079_));
 sg13g2_a21oi_1 _2349_ (.A1(net484),
    .A2(net472),
    .Y(_0197_),
    .B1(_0196_));
 sg13g2_a21oi_1 _2350_ (.A1(_1070_),
    .A2(_0197_),
    .Y(_0198_),
    .B1(net460));
 sg13g2_a221oi_1 _2351_ (.B2(_0198_),
    .C1(net449),
    .B1(_0194_),
    .A1(net463),
    .Y(_0199_),
    .A2(_0193_));
 sg13g2_or3_1 _2352_ (.A(net498),
    .B(_0997_),
    .C(_1104_),
    .X(_0200_));
 sg13g2_a22oi_1 _2353_ (.Y(_0201_),
    .B1(_1000_),
    .B2(net499),
    .A2(_0933_),
    .A1(_0828_));
 sg13g2_inv_1 _2354_ (.Y(_0202_),
    .A(_0201_));
 sg13g2_a22oi_1 _2355_ (.Y(_0203_),
    .B1(_0202_),
    .B2(net454),
    .A2(_0200_),
    .A1(_0995_));
 sg13g2_nand3_1 _2356_ (.B(_0898_),
    .C(_0942_),
    .A(_0842_),
    .Y(_0204_));
 sg13g2_a21oi_1 _2357_ (.A1(_0862_),
    .A2(_0874_),
    .Y(_0205_),
    .B1(net511));
 sg13g2_a21oi_1 _2358_ (.A1(_1011_),
    .A2(_1113_),
    .Y(_0206_),
    .B1(_0205_));
 sg13g2_mux2_1 _2359_ (.A0(_0204_),
    .A1(_0206_),
    .S(net457),
    .X(_0207_));
 sg13g2_a221oi_1 _2360_ (.B2(_1004_),
    .C1(_0812_),
    .B1(_0207_),
    .A1(net461),
    .Y(_0208_),
    .A2(_0203_));
 sg13g2_or3_1 _2361_ (.A(net447),
    .B(_0199_),
    .C(_0208_),
    .X(_0209_));
 sg13g2_o21ai_1 _2362_ (.B1(net451),
    .Y(_0210_),
    .A1(net522),
    .A2(_0924_));
 sg13g2_a221oi_1 _2363_ (.B2(_1067_),
    .C1(_0832_),
    .B1(_0824_),
    .A1(net486),
    .Y(_0211_),
    .A2(net475));
 sg13g2_a21oi_1 _2364_ (.A1(net515),
    .A2(_0759_),
    .Y(_0212_),
    .B1(_1104_));
 sg13g2_and2_1 _2365_ (.A(_1056_),
    .B(_0212_),
    .X(_0213_));
 sg13g2_o21ai_1 _2366_ (.B1(_1221_),
    .Y(_0214_),
    .A1(net539),
    .A2(_0754_));
 sg13g2_nor2_1 _2367_ (.A(net498),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_nor4_2 _2368_ (.A(net490),
    .B(net478),
    .C(_0213_),
    .Y(_0216_),
    .D(_0215_));
 sg13g2_nor3_1 _2369_ (.A(net467),
    .B(_0211_),
    .C(_0216_),
    .Y(_0217_));
 sg13g2_o21ai_1 _2370_ (.B1(_0922_),
    .Y(_0218_),
    .A1(_0771_),
    .A2(_0186_));
 sg13g2_a21o_1 _2371_ (.A2(_1115_),
    .A1(net531),
    .B1(_1104_),
    .X(_0219_));
 sg13g2_o21ai_1 _2372_ (.B1(net499),
    .Y(_0220_),
    .A1(_0754_),
    .A2(_0874_));
 sg13g2_o21ai_1 _2373_ (.B1(_0220_),
    .Y(_0221_),
    .A1(net500),
    .A2(_0219_));
 sg13g2_a21oi_1 _2374_ (.A1(net454),
    .A2(_0221_),
    .Y(_0222_),
    .B1(net462));
 sg13g2_a22oi_1 _2375_ (.Y(_0223_),
    .B1(_0218_),
    .B2(_0222_),
    .A2(_0217_),
    .A1(_0210_));
 sg13g2_a21oi_1 _2376_ (.A1(net447),
    .A2(_0223_),
    .Y(_0224_),
    .B1(_0009_));
 sg13g2_nand3_1 _2377_ (.B(_0891_),
    .C(_1022_),
    .A(net534),
    .Y(_0225_));
 sg13g2_o21ai_1 _2378_ (.B1(net534),
    .Y(_0226_),
    .A1(net521),
    .A2(_0856_));
 sg13g2_o21ai_1 _2379_ (.B1(_0226_),
    .Y(_0227_),
    .A1(_0999_),
    .A2(_1204_));
 sg13g2_a22oi_1 _2380_ (.Y(_0228_),
    .B1(_0227_),
    .B2(net510),
    .A2(_0225_),
    .A1(_0855_));
 sg13g2_nor3_1 _2381_ (.A(net490),
    .B(net478),
    .C(_0228_),
    .Y(_0229_));
 sg13g2_a221oi_1 _2382_ (.B2(_1028_),
    .C1(net498),
    .B1(_0795_),
    .A1(net485),
    .Y(_0230_),
    .A2(net473));
 sg13g2_a221oi_1 _2383_ (.B2(_0942_),
    .C1(net509),
    .B1(_0839_),
    .A1(net485),
    .Y(_0231_),
    .A2(net473));
 sg13g2_or3_1 _2384_ (.A(_0229_),
    .B(_0230_),
    .C(_0231_),
    .X(_0232_));
 sg13g2_nor2_1 _2385_ (.A(net529),
    .B(_0186_),
    .Y(_0233_));
 sg13g2_a22oi_1 _2386_ (.Y(_0234_),
    .B1(_0233_),
    .B2(net451),
    .A2(_1018_),
    .A1(_0841_));
 sg13g2_a221oi_1 _2387_ (.B2(_1026_),
    .C1(_0812_),
    .B1(_0234_),
    .A1(net466),
    .Y(_0235_),
    .A2(_0232_));
 sg13g2_nor2_1 _2388_ (.A(_1047_),
    .B(_1051_),
    .Y(_0236_));
 sg13g2_a221oi_1 _2389_ (.B2(net531),
    .C1(_1000_),
    .B1(_1035_),
    .A1(net573),
    .Y(_0237_),
    .A2(_0835_));
 sg13g2_a22oi_1 _2390_ (.Y(_0238_),
    .B1(_0237_),
    .B2(net450),
    .A2(_1116_),
    .A1(_0793_));
 sg13g2_a221oi_1 _2391_ (.B2(_0783_),
    .C1(net460),
    .B1(_0236_),
    .A1(net458),
    .Y(_0239_),
    .A2(_1163_));
 sg13g2_a21oi_1 _2392_ (.A1(net497),
    .A2(_1037_),
    .Y(_0240_),
    .B1(_1103_));
 sg13g2_nor3_1 _2393_ (.A(net490),
    .B(net478),
    .C(_0240_),
    .Y(_0241_));
 sg13g2_nor3_1 _2394_ (.A(net536),
    .B(_0856_),
    .C(_1066_),
    .Y(_0242_));
 sg13g2_o21ai_1 _2395_ (.B1(net450),
    .Y(_0243_),
    .A1(_0838_),
    .A2(_0242_));
 sg13g2_nand2_1 _2396_ (.Y(_0244_),
    .A(_0881_),
    .B(_1092_));
 sg13g2_a221oi_1 _2397_ (.B2(net515),
    .C1(_0244_),
    .B1(_0759_),
    .A1(net487),
    .Y(_0245_),
    .A2(net474));
 sg13g2_nor3_1 _2398_ (.A(net466),
    .B(_0241_),
    .C(_0245_),
    .Y(_0246_));
 sg13g2_a221oi_1 _2399_ (.B2(_0246_),
    .C1(_0813_),
    .B1(_0243_),
    .A1(_0238_),
    .Y(_0247_),
    .A2(_0239_));
 sg13g2_or3_1 _2400_ (.A(net447),
    .B(_0235_),
    .C(_0247_),
    .X(_0248_));
 sg13g2_nand3_1 _2401_ (.B(_0842_),
    .C(_0996_),
    .A(net509),
    .Y(_0249_));
 sg13g2_nand2b_1 _2402_ (.Y(_0250_),
    .B(_0855_),
    .A_N(_0864_));
 sg13g2_nand2_1 _2403_ (.Y(_0251_),
    .A(_0249_),
    .B(_0250_));
 sg13g2_a21oi_1 _2404_ (.A1(_0756_),
    .A2(_0797_),
    .Y(_0252_),
    .B1(_0819_));
 sg13g2_nand2b_1 _2405_ (.Y(_0253_),
    .B(_1211_),
    .A_N(_0252_));
 sg13g2_o21ai_1 _2406_ (.B1(_0253_),
    .Y(_0254_),
    .A1(net499),
    .A2(_1104_));
 sg13g2_nor3_1 _2407_ (.A(_0841_),
    .B(_0899_),
    .C(_1096_),
    .Y(_0255_));
 sg13g2_a21oi_1 _2408_ (.A1(_0933_),
    .A2(_0113_),
    .Y(_0256_),
    .B1(_0255_));
 sg13g2_nand3_1 _2409_ (.B(_0874_),
    .C(_0932_),
    .A(net500),
    .Y(_0257_));
 sg13g2_mux4_1 _2410_ (.S0(net462),
    .A0(_0251_),
    .A1(_0254_),
    .A2(_0257_),
    .A3(_0256_),
    .S1(net456),
    .X(_0258_));
 sg13g2_a21oi_1 _2411_ (.A1(net447),
    .A2(_0258_),
    .Y(_0259_),
    .B1(_0532_));
 sg13g2_a221oi_1 _2412_ (.B2(_0259_),
    .C1(_0920_),
    .B1(_0248_),
    .A1(_0209_),
    .Y(_0260_),
    .A2(_0224_));
 sg13g2_mux2_1 _2413_ (.A0(_0013_),
    .A1(net566),
    .S(net574),
    .X(_0261_));
 sg13g2_nand2_1 _2414_ (.Y(_0262_),
    .A(_0705_),
    .B(_0261_));
 sg13g2_nand3_1 _2415_ (.B(_0979_),
    .C(_0262_),
    .A(net552),
    .Y(_0263_));
 sg13g2_nand3_1 _2416_ (.B(_0968_),
    .C(_0975_),
    .A(net550),
    .Y(_0264_));
 sg13g2_nand3_1 _2417_ (.B(_0263_),
    .C(_0264_),
    .A(net556),
    .Y(_0265_));
 sg13g2_nand3_1 _2418_ (.B(_1142_),
    .C(_1145_),
    .A(_0957_),
    .Y(_0266_));
 sg13g2_nand2b_1 _2419_ (.Y(_0267_),
    .B(_0266_),
    .A_N(_0982_));
 sg13g2_o21ai_1 _2420_ (.B1(_0265_),
    .Y(_0268_),
    .A1(net556),
    .A2(_0267_));
 sg13g2_nand2_1 _2421_ (.Y(_0269_),
    .A(_0176_),
    .B(_0268_));
 sg13g2_nand2b_1 _2422_ (.Y(_0270_),
    .B(_1137_),
    .A_N(_0974_));
 sg13g2_a221oi_1 _2423_ (.B2(net552),
    .C1(net554),
    .B1(_0270_),
    .A1(_1130_),
    .Y(_0271_),
    .A2(_1149_));
 sg13g2_a21o_1 _2424_ (.A2(_1144_),
    .A1(_0976_),
    .B1(_0271_),
    .X(_0272_));
 sg13g2_o21ai_1 _2425_ (.B1(_0269_),
    .Y(_0273_),
    .A1(_0168_),
    .A2(_0272_));
 sg13g2_nor2_1 _2426_ (.A(_0260_),
    .B(_0273_),
    .Y(_0274_));
 sg13g2_or2_2 _2427_ (.X(_0275_),
    .B(_0273_),
    .A(_0260_));
 sg13g2_a21oi_1 _2428_ (.A1(_0185_),
    .A2(net444),
    .Y(_0276_),
    .B1(_1261_));
 sg13g2_nand2_1 _2429_ (.Y(_0277_),
    .A(_0184_),
    .B(_0275_));
 sg13g2_or2_1 _2430_ (.X(_0278_),
    .B(_0276_),
    .A(_1258_));
 sg13g2_a21oi_1 _2431_ (.A1(_0276_),
    .A2(_0277_),
    .Y(_0279_),
    .B1(_1258_));
 sg13g2_a221oi_1 _2432_ (.B2(_0277_),
    .C1(_1160_),
    .B1(_0276_),
    .A1(net445),
    .Y(_0280_),
    .A2(net468));
 sg13g2_o21ai_1 _2433_ (.B1(_1260_),
    .Y(_0281_),
    .A1(_0166_),
    .A2(_0183_));
 sg13g2_a22oi_1 _2434_ (.Y(_0282_),
    .B1(_1260_),
    .B2(_0185_),
    .A2(_1158_),
    .A1(_1155_));
 sg13g2_nand2_1 _2435_ (.Y(_0283_),
    .A(_1160_),
    .B(_0281_));
 sg13g2_and3_1 _2436_ (.X(_0284_),
    .A(net446),
    .B(net469),
    .C(_0281_));
 sg13g2_nand3_1 _2437_ (.B(net468),
    .C(_0281_),
    .A(net445),
    .Y(_0285_));
 sg13g2_nand3_1 _2438_ (.B(net468),
    .C(_0275_),
    .A(net445),
    .Y(_0286_));
 sg13g2_nand3b_1 _2439_ (.B(_0285_),
    .C(_0286_),
    .Y(_0287_),
    .A_N(_0282_));
 sg13g2_o21ai_1 _2440_ (.B1(_0993_),
    .Y(_0288_),
    .A1(_0280_),
    .A2(_0287_));
 sg13g2_a22oi_1 _2441_ (.Y(_0289_),
    .B1(_1260_),
    .B2(_0274_),
    .A2(net469),
    .A1(net446));
 sg13g2_o21ai_1 _2442_ (.B1(_1261_),
    .Y(_0290_),
    .A1(_0260_),
    .A2(_0273_));
 sg13g2_a22oi_1 _2443_ (.Y(_0291_),
    .B1(_0275_),
    .B2(_0281_),
    .A2(net469),
    .A1(net446));
 sg13g2_o21ai_1 _2444_ (.B1(net444),
    .Y(_0292_),
    .A1(_1260_),
    .A2(_0185_));
 sg13g2_a21o_1 _2445_ (.A2(_0292_),
    .A1(_0291_),
    .B1(_1160_),
    .X(_0293_));
 sg13g2_and4_1 _2446_ (.A(net445),
    .B(net468),
    .C(_1260_),
    .D(net444),
    .X(_0294_));
 sg13g2_o21ai_1 _2447_ (.B1(_0992_),
    .Y(_0295_),
    .A1(_1159_),
    .A2(_0294_));
 sg13g2_o21ai_1 _2448_ (.B1(_0293_),
    .Y(_0296_),
    .A1(_1159_),
    .A2(_0184_));
 sg13g2_o21ai_1 _2449_ (.B1(_0288_),
    .Y(_0297_),
    .A1(_0295_),
    .A2(_0296_));
 sg13g2_nor2_1 _2450_ (.A(_0919_),
    .B(_0954_),
    .Y(_0298_));
 sg13g2_a21oi_1 _2451_ (.A1(_0677_),
    .A2(_0680_),
    .Y(_0299_),
    .B1(_0918_));
 sg13g2_nand2_1 _2452_ (.Y(_0300_),
    .A(net588),
    .B(_0299_));
 sg13g2_inv_1 _2453_ (.Y(_0301_),
    .A(_0300_));
 sg13g2_a21o_1 _2454_ (.A2(_0301_),
    .A1(_0297_),
    .B1(_0657_),
    .X(_0037_));
 sg13g2_nand4_1 _2455_ (.B(net468),
    .C(net444),
    .A(net445),
    .Y(_0302_),
    .D(_0281_));
 sg13g2_nor3_2 _2456_ (.A(_1261_),
    .B(_0166_),
    .C(_0183_),
    .Y(_0303_));
 sg13g2_a21oi_1 _2457_ (.A1(net446),
    .A2(net469),
    .Y(_0304_),
    .B1(_0303_));
 sg13g2_nor2_1 _2458_ (.A(_1160_),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_a21o_1 _2459_ (.A2(_0305_),
    .A1(_0302_),
    .B1(_0295_),
    .X(_0306_));
 sg13g2_a21oi_1 _2460_ (.A1(_0288_),
    .A2(_0306_),
    .Y(_0307_),
    .B1(_0300_));
 sg13g2_a21o_1 _2461_ (.A2(net207),
    .A1(net584),
    .B1(_0307_),
    .X(_0038_));
 sg13g2_nand4_1 _2462_ (.B(\gfx.pixel_x[0] ),
    .C(\gfx.bitmap_x[0] ),
    .A(\gfx.pixel_x[1] ),
    .Y(_0308_),
    .D(net247));
 sg13g2_nor2_1 _2463_ (.A(net577),
    .B(net579),
    .Y(_0309_));
 sg13g2_o21ai_1 _2464_ (.B1(_0309_),
    .Y(_0310_),
    .A1(_0655_),
    .A2(_0308_));
 sg13g2_nand3_1 _2465_ (.B(\gfx.pixel_x[9] ),
    .C(_0310_),
    .A(net576),
    .Y(_0311_));
 sg13g2_and2_1 _2466_ (.A(net587),
    .B(_0311_),
    .X(_0312_));
 sg13g2_a22oi_1 _2467_ (.Y(_0313_),
    .B1(_0312_),
    .B2(net106),
    .A2(\gfx.pixel_x[0] ),
    .A1(net583));
 sg13g2_inv_1 _2468_ (.Y(_0039_),
    .A(net107));
 sg13g2_nor2b_1 _2469_ (.A(net587),
    .B_N(net239),
    .Y(_0314_));
 sg13g2_xor2_1 _2470_ (.B(\gfx.pixel_x[0] ),
    .A(net239),
    .X(_0315_));
 sg13g2_a21o_1 _2471_ (.A2(_0315_),
    .A1(_0312_),
    .B1(_0314_),
    .X(_0040_));
 sg13g2_nor2_1 _2472_ (.A(net584),
    .B(_0311_),
    .Y(_0316_));
 sg13g2_nand3_1 _2473_ (.B(\gfx.pixel_x[1] ),
    .C(\gfx.pixel_x[0] ),
    .A(net587),
    .Y(_0317_));
 sg13g2_nand4_1 _2474_ (.B(\gfx.pixel_x[1] ),
    .C(\gfx.pixel_x[0] ),
    .A(net587),
    .Y(_0318_),
    .D(net216));
 sg13g2_xor2_1 _2475_ (.B(_0317_),
    .A(net216),
    .X(_0319_));
 sg13g2_nor2_1 _2476_ (.A(net519),
    .B(net217),
    .Y(_0041_));
 sg13g2_nor2_1 _2477_ (.A(net584),
    .B(_0308_),
    .Y(_0320_));
 sg13g2_nor2b_1 _2478_ (.A(net220),
    .B_N(_0318_),
    .Y(_0321_));
 sg13g2_nor3_1 _2479_ (.A(net519),
    .B(_0320_),
    .C(net221),
    .Y(_0042_));
 sg13g2_xor2_1 _2480_ (.B(_0308_),
    .A(net224),
    .X(_0322_));
 sg13g2_a22oi_1 _2481_ (.Y(_0323_),
    .B1(_0312_),
    .B2(net225),
    .A2(net581),
    .A1(net585));
 sg13g2_inv_1 _2482_ (.Y(_0043_),
    .A(_0323_));
 sg13g2_nor3_1 _2483_ (.A(net585),
    .B(_0655_),
    .C(_0308_),
    .Y(_0324_));
 sg13g2_a21oi_1 _2484_ (.A1(net581),
    .A2(_0320_),
    .Y(_0325_),
    .B1(net580));
 sg13g2_nor3_1 _2485_ (.A(net519),
    .B(_0324_),
    .C(_0325_),
    .Y(_0044_));
 sg13g2_and2_1 _2486_ (.A(net578),
    .B(_0324_),
    .X(_0326_));
 sg13g2_nor2_1 _2487_ (.A(net578),
    .B(_0324_),
    .Y(_0327_));
 sg13g2_nor3_1 _2488_ (.A(net519),
    .B(_0326_),
    .C(_0327_),
    .Y(_0045_));
 sg13g2_nor2_1 _2489_ (.A(net153),
    .B(_0326_),
    .Y(_0328_));
 sg13g2_and2_1 _2490_ (.A(net577),
    .B(_0326_),
    .X(_0329_));
 sg13g2_nor3_1 _2491_ (.A(net519),
    .B(_0328_),
    .C(_0329_),
    .Y(_0046_));
 sg13g2_xnor2_1 _2492_ (.Y(_0330_),
    .A(net576),
    .B(_0329_));
 sg13g2_nor2_1 _2493_ (.A(net519),
    .B(_0330_),
    .Y(_0047_));
 sg13g2_a21oi_1 _2494_ (.A1(net576),
    .A2(_0329_),
    .Y(_0331_),
    .B1(net194));
 sg13g2_nor2_1 _2495_ (.A(net519),
    .B(net195),
    .Y(_0048_));
 sg13g2_and3_1 _2496_ (.X(_0332_),
    .A(net446),
    .B(net469),
    .C(_0290_));
 sg13g2_a21oi_1 _2497_ (.A1(_0281_),
    .A2(_0332_),
    .Y(_0333_),
    .B1(_1160_));
 sg13g2_or3_1 _2498_ (.A(_0185_),
    .B(_0289_),
    .C(_0332_),
    .X(_0334_));
 sg13g2_a22oi_1 _2499_ (.Y(_0335_),
    .B1(_0334_),
    .B2(_1160_),
    .A2(_0333_),
    .A1(_0278_));
 sg13g2_and3_1 _2500_ (.X(_0336_),
    .A(net446),
    .B(net469),
    .C(_0303_));
 sg13g2_nand2_1 _2501_ (.Y(_0337_),
    .A(_1259_),
    .B(_0281_));
 sg13g2_a221oi_1 _2502_ (.B2(_0185_),
    .C1(net444),
    .B1(_1260_),
    .A1(net446),
    .Y(_0338_),
    .A2(net469));
 sg13g2_o21ai_1 _2503_ (.B1(_1160_),
    .Y(_0339_),
    .A1(_0336_),
    .A2(_0338_));
 sg13g2_and3_1 _2504_ (.X(_0340_),
    .A(_1155_),
    .B(_1158_),
    .C(_0275_));
 sg13g2_a21oi_1 _2505_ (.A1(_0284_),
    .A2(_0340_),
    .Y(_0341_),
    .B1(_0993_));
 sg13g2_a21oi_1 _2506_ (.A1(_0339_),
    .A2(_0341_),
    .Y(_0342_),
    .B1(_0298_));
 sg13g2_o21ai_1 _2507_ (.B1(_0342_),
    .Y(_0343_),
    .A1(_0992_),
    .A2(_0335_));
 sg13g2_nand2b_1 _2508_ (.Y(_0344_),
    .B(_0642_),
    .A_N(\gfx.pixel_y[9] ));
 sg13g2_a21oi_1 _2509_ (.A1(\gfx.pixel_x[9] ),
    .A2(_0677_),
    .Y(_0345_),
    .B1(_0344_));
 sg13g2_a21oi_2 _2510_ (.B1(net584),
    .Y(_0346_),
    .A2(_0345_),
    .A1(_0298_));
 sg13g2_a22oi_1 _2511_ (.Y(_0049_),
    .B1(_0343_),
    .B2(_0346_),
    .A2(_0538_),
    .A1(net585));
 sg13g2_nand3_1 _2512_ (.B(_0991_),
    .C(net444),
    .A(_0988_),
    .Y(_0347_));
 sg13g2_o21ai_1 _2513_ (.B1(_0295_),
    .Y(_0348_),
    .A1(_0337_),
    .A2(_0347_));
 sg13g2_nand2_1 _2514_ (.Y(_0349_),
    .A(_0184_),
    .B(_0290_));
 sg13g2_a22oi_1 _2515_ (.Y(_0350_),
    .B1(_0184_),
    .B2(_0290_),
    .A2(net468),
    .A1(net445));
 sg13g2_nand3b_1 _2516_ (.B(_1159_),
    .C(_0285_),
    .Y(_0351_),
    .A_N(_0350_));
 sg13g2_o21ai_1 _2517_ (.B1(_0282_),
    .Y(_0352_),
    .A1(_0289_),
    .A2(_0332_));
 sg13g2_a21o_1 _2518_ (.A2(_0286_),
    .A1(_0285_),
    .B1(_1160_),
    .X(_0353_));
 sg13g2_nand3b_1 _2519_ (.B(_0352_),
    .C(_0353_),
    .Y(_0354_),
    .A_N(_0280_));
 sg13g2_a22oi_1 _2520_ (.Y(_0355_),
    .B1(_0354_),
    .B2(_0993_),
    .A2(_0351_),
    .A1(_0348_));
 sg13g2_nand2_1 _2521_ (.Y(_0356_),
    .A(net584),
    .B(net171));
 sg13g2_o21ai_1 _2522_ (.B1(_0356_),
    .Y(_0050_),
    .A1(_0300_),
    .A2(_0355_));
 sg13g2_a21oi_1 _2523_ (.A1(net575),
    .A2(\gfx.pixel_y[2] ),
    .Y(_0357_),
    .B1(\gfx.pixel_y[8] ));
 sg13g2_nor4_1 _2524_ (.A(net569),
    .B(net566),
    .C(net565),
    .D(\gfx.bitmap_y[3] ),
    .Y(_0358_));
 sg13g2_nand2_1 _2525_ (.Y(_0359_),
    .A(\gfx.pixel_y[9] ),
    .B(net520));
 sg13g2_a21oi_1 _2526_ (.A1(_0357_),
    .A2(_0358_),
    .Y(_0360_),
    .B1(_0359_));
 sg13g2_inv_1 _2527_ (.Y(_0361_),
    .A(net513));
 sg13g2_nand2b_1 _2528_ (.Y(_0362_),
    .B(net520),
    .A_N(net149));
 sg13g2_o21ai_1 _2529_ (.B1(_0362_),
    .Y(_0363_),
    .A1(\gfx.pixel_y[0] ),
    .A2(net519));
 sg13g2_nor2_1 _2530_ (.A(net514),
    .B(net150),
    .Y(_0051_));
 sg13g2_a21oi_1 _2531_ (.A1(\gfx.pixel_y[0] ),
    .A2(net520),
    .Y(_0364_),
    .B1(net117));
 sg13g2_and3_1 _2532_ (.X(_0365_),
    .A(\gfx.pixel_y[0] ),
    .B(net117),
    .C(net520));
 sg13g2_nor3_1 _2533_ (.A(net514),
    .B(net118),
    .C(_0365_),
    .Y(_0052_));
 sg13g2_nor2_1 _2534_ (.A(net200),
    .B(_0365_),
    .Y(_0366_));
 sg13g2_and2_1 _2535_ (.A(net200),
    .B(_0365_),
    .X(_0367_));
 sg13g2_nor3_1 _2536_ (.A(net513),
    .B(net201),
    .C(_0367_),
    .Y(_0053_));
 sg13g2_nor2_1 _2537_ (.A(net574),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_and2_1 _2538_ (.A(net574),
    .B(_0367_),
    .X(_0369_));
 sg13g2_nor3_1 _2539_ (.A(net513),
    .B(_0368_),
    .C(_0369_),
    .Y(_0054_));
 sg13g2_and2_1 _2540_ (.A(net569),
    .B(_0369_),
    .X(_0370_));
 sg13g2_o21ai_1 _2541_ (.B1(_0361_),
    .Y(_0371_),
    .A1(net569),
    .A2(_0369_));
 sg13g2_nor2_1 _2542_ (.A(_0370_),
    .B(_0371_),
    .Y(_0055_));
 sg13g2_nor2b_1 _2543_ (.A(net202),
    .B_N(_0369_),
    .Y(_0372_));
 sg13g2_xnor2_1 _2544_ (.Y(_0373_),
    .A(net566),
    .B(_0372_));
 sg13g2_nor2_1 _2545_ (.A(net513),
    .B(net203),
    .Y(_0056_));
 sg13g2_and2_1 _2546_ (.A(net566),
    .B(_0370_),
    .X(_0374_));
 sg13g2_a21oi_1 _2547_ (.A1(net219),
    .A2(_0374_),
    .Y(_0375_),
    .B1(net513));
 sg13g2_o21ai_1 _2548_ (.B1(_0375_),
    .Y(_0376_),
    .A1(net219),
    .A2(_0374_));
 sg13g2_inv_1 _2549_ (.Y(_0057_),
    .A(_0376_));
 sg13g2_and4_1 _2550_ (.A(net568),
    .B(net566),
    .C(_0531_),
    .D(_0369_),
    .X(_0377_));
 sg13g2_o21ai_1 _2551_ (.B1(_0361_),
    .Y(_0378_),
    .A1(net565),
    .A2(_0377_));
 sg13g2_a21oi_1 _2552_ (.A1(net565),
    .A2(_0377_),
    .Y(_0058_),
    .B1(_0378_));
 sg13g2_a21oi_1 _2553_ (.A1(_0641_),
    .A2(_0374_),
    .Y(_0379_),
    .B1(net184));
 sg13g2_nor2b_1 _2554_ (.A(_0642_),
    .B_N(_0370_),
    .Y(_0380_));
 sg13g2_nor3_1 _2555_ (.A(net513),
    .B(net185),
    .C(_0380_),
    .Y(_0059_));
 sg13g2_nor2_1 _2556_ (.A(net192),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_nor2_1 _2557_ (.A(net513),
    .B(_0381_),
    .Y(_0060_));
 sg13g2_nand2_1 _2558_ (.Y(_0382_),
    .A(_1159_),
    .B(_0349_));
 sg13g2_nand2_1 _2559_ (.Y(_0383_),
    .A(_0185_),
    .B(_0275_));
 sg13g2_nand3_1 _2560_ (.B(_0349_),
    .C(_0383_),
    .A(_1159_),
    .Y(_0384_));
 sg13g2_a21oi_1 _2561_ (.A1(_0283_),
    .A2(_0384_),
    .Y(_0385_),
    .B1(_0993_));
 sg13g2_a21oi_1 _2562_ (.A1(_1155_),
    .A2(_1158_),
    .Y(_0386_),
    .B1(net444));
 sg13g2_a221oi_1 _2563_ (.B2(net444),
    .C1(_0386_),
    .B1(_1260_),
    .A1(_0988_),
    .Y(_0387_),
    .A2(_0991_));
 sg13g2_a21o_1 _2564_ (.A2(_0387_),
    .A1(_0382_),
    .B1(_1258_),
    .X(_0388_));
 sg13g2_a21oi_1 _2565_ (.A1(_0988_),
    .A2(_0991_),
    .Y(_0389_),
    .B1(_0303_));
 sg13g2_a221oi_1 _2566_ (.B2(_0340_),
    .C1(_1259_),
    .B1(_0389_),
    .A1(_0303_),
    .Y(_0390_),
    .A2(_0386_));
 sg13g2_nor2_1 _2567_ (.A(_0298_),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_o21ai_1 _2568_ (.B1(_0391_),
    .Y(_0392_),
    .A1(_0385_),
    .A2(_0388_));
 sg13g2_a22oi_1 _2569_ (.Y(_0061_),
    .B1(_0346_),
    .B2(_0392_),
    .A2(_0539_),
    .A1(net584));
 sg13g2_nand2_1 _2570_ (.Y(_0393_),
    .A(_0993_),
    .B(_0286_));
 sg13g2_nand3b_1 _2571_ (.B(_0992_),
    .C(_0302_),
    .Y(_0394_),
    .A_N(_0350_));
 sg13g2_o21ai_1 _2572_ (.B1(_0394_),
    .Y(_0395_),
    .A1(_0279_),
    .A2(_0393_));
 sg13g2_a221oi_1 _2573_ (.B2(_0347_),
    .C1(_1259_),
    .B1(_0277_),
    .A1(_0992_),
    .Y(_0396_),
    .A2(_1261_));
 sg13g2_a21o_1 _2574_ (.A2(_0281_),
    .A1(_1259_),
    .B1(_1159_),
    .X(_0397_));
 sg13g2_o21ai_1 _2575_ (.B1(_0299_),
    .Y(_0398_),
    .A1(_0396_),
    .A2(_0397_));
 sg13g2_a21o_1 _2576_ (.A2(_0395_),
    .A1(_1159_),
    .B1(_0398_),
    .X(_0399_));
 sg13g2_a22oi_1 _2577_ (.Y(_0062_),
    .B1(_0346_),
    .B2(_0399_),
    .A2(_0540_),
    .A1(net584));
 sg13g2_nand2_1 _2578_ (.Y(_0400_),
    .A(\music.do_note ),
    .B(_0562_));
 sg13g2_nand3b_1 _2579_ (.B(\music.note_pos[2] ),
    .C(_0559_),
    .Y(_0401_),
    .A_N(\music.note_pos[3] ));
 sg13g2_nor4_1 _2580_ (.A(\music.note_pos[8] ),
    .B(\music.note_pos[7] ),
    .C(\music.note_pos[6] ),
    .D(\music.note_length ),
    .Y(_0402_));
 sg13g2_nor4_1 _2581_ (.A(_0515_),
    .B(\music.note_pos[13] ),
    .C(\music.note_pos[12] ),
    .D(\music.note_pos[10] ),
    .Y(_0403_));
 sg13g2_nand3b_1 _2582_ (.B(_0402_),
    .C(_0403_),
    .Y(_0404_),
    .A_N(_0401_));
 sg13g2_nor4_1 _2583_ (.A(\music.note_pos[15] ),
    .B(_0560_),
    .C(_0400_),
    .D(_0404_),
    .Y(_0405_));
 sg13g2_and2_1 _2584_ (.A(\music.do_note ),
    .B(\music.note_pos[15] ),
    .X(_0406_));
 sg13g2_nand4_1 _2585_ (.B(\music.note_pos[7] ),
    .C(_0558_),
    .A(_0515_),
    .Y(_0407_),
    .D(_0406_));
 sg13g2_nor3_1 _2586_ (.A(\music.note_pos[6] ),
    .B(\music.note_pos[5] ),
    .C(\music.note_pos[4] ),
    .Y(_0408_));
 sg13g2_nand2_1 _2587_ (.Y(_0409_),
    .A(\music.note_length ),
    .B(_0408_));
 sg13g2_nor4_1 _2588_ (.A(_0563_),
    .B(_0401_),
    .C(_0407_),
    .D(_0409_),
    .Y(_0410_));
 sg13g2_nand2b_1 _2589_ (.Y(_0411_),
    .B(_0557_),
    .A_N(_0410_));
 sg13g2_nor3_1 _2590_ (.A(_0566_),
    .B(_0405_),
    .C(_0411_),
    .Y(_0412_));
 sg13g2_nor2_1 _2591_ (.A(net188),
    .B(_0412_),
    .Y(_0413_));
 sg13g2_and2_1 _2592_ (.A(net188),
    .B(_0557_),
    .X(_0414_));
 sg13g2_nor3_1 _2593_ (.A(net583),
    .B(_0413_),
    .C(_0414_),
    .Y(_0063_));
 sg13g2_xnor2_1 _2594_ (.Y(_0415_),
    .A(net205),
    .B(_0414_));
 sg13g2_nor2_1 _2595_ (.A(net583),
    .B(_0415_),
    .Y(_0064_));
 sg13g2_and3_1 _2596_ (.X(_0416_),
    .A(net164),
    .B(\music.note_pos[1] ),
    .C(_0414_));
 sg13g2_a21oi_1 _2597_ (.A1(\music.note_pos[1] ),
    .A2(_0414_),
    .Y(_0417_),
    .B1(net164));
 sg13g2_nand2_1 _2598_ (.Y(_0418_),
    .A(_0557_),
    .B(_0410_));
 sg13g2_nand2_1 _2599_ (.Y(_0419_),
    .A(net586),
    .B(_0418_));
 sg13g2_and4_1 _2600_ (.A(net164),
    .B(net205),
    .C(net188),
    .D(_0569_),
    .X(_0420_));
 sg13g2_nand2_1 _2601_ (.Y(_0421_),
    .A(_0557_),
    .B(_0405_));
 sg13g2_nand3_1 _2602_ (.B(_0418_),
    .C(_0421_),
    .A(_0567_),
    .Y(_0422_));
 sg13g2_nor4_1 _2603_ (.A(net583),
    .B(_0416_),
    .C(net165),
    .D(_0422_),
    .Y(_0065_));
 sg13g2_and2_1 _2604_ (.A(net210),
    .B(_0416_),
    .X(_0423_));
 sg13g2_nor2_1 _2605_ (.A(net210),
    .B(_0420_),
    .Y(_0424_));
 sg13g2_nor3_1 _2606_ (.A(_0571_),
    .B(_0423_),
    .C(_0424_),
    .Y(_0066_));
 sg13g2_or2_1 _2607_ (.X(_0425_),
    .B(_0423_),
    .A(net234));
 sg13g2_nand2_1 _2608_ (.Y(_0426_),
    .A(net234),
    .B(_0423_));
 sg13g2_nand4_1 _2609_ (.B(_0421_),
    .C(_0425_),
    .A(_0570_),
    .Y(_0427_),
    .D(_0426_));
 sg13g2_inv_1 _2610_ (.Y(_0067_),
    .A(_0427_));
 sg13g2_a21oi_1 _2611_ (.A1(\music.note_pos[4] ),
    .A2(_0423_),
    .Y(_0428_),
    .B1(net141));
 sg13g2_and4_2 _2612_ (.A(net141),
    .B(net248),
    .C(net210),
    .D(_0420_),
    .X(_0429_));
 sg13g2_nor3_1 _2613_ (.A(net583),
    .B(net142),
    .C(_0429_),
    .Y(_0068_));
 sg13g2_xnor2_1 _2614_ (.Y(_0430_),
    .A(net222),
    .B(_0429_));
 sg13g2_nor2_1 _2615_ (.A(_0571_),
    .B(net223),
    .Y(_0069_));
 sg13g2_a21oi_1 _2616_ (.A1(\music.note_pos[6] ),
    .A2(_0429_),
    .Y(_0431_),
    .B1(net179));
 sg13g2_and3_1 _2617_ (.X(_0432_),
    .A(net179),
    .B(net246),
    .C(_0429_));
 sg13g2_nor3_1 _2618_ (.A(_0419_),
    .B(net180),
    .C(_0432_),
    .Y(_0070_));
 sg13g2_nor2_1 _2619_ (.A(net206),
    .B(_0432_),
    .Y(_0433_));
 sg13g2_nand2_1 _2620_ (.Y(_0434_),
    .A(_0570_),
    .B(_0418_));
 sg13g2_and2_1 _2621_ (.A(net206),
    .B(_0432_),
    .X(_0435_));
 sg13g2_nor3_1 _2622_ (.A(_0433_),
    .B(_0434_),
    .C(_0435_),
    .Y(_0071_));
 sg13g2_o21ai_1 _2623_ (.B1(net586),
    .Y(_0436_),
    .A1(net136),
    .A2(_0435_));
 sg13g2_a21oi_1 _2624_ (.A1(net136),
    .A2(_0435_),
    .Y(_0072_),
    .B1(_0436_));
 sg13g2_a21oi_1 _2625_ (.A1(net136),
    .A2(_0435_),
    .Y(_0437_),
    .B1(net155));
 sg13g2_and3_1 _2626_ (.X(_0438_),
    .A(net155),
    .B(net136),
    .C(_0435_));
 sg13g2_nor3_1 _2627_ (.A(_0434_),
    .B(net156),
    .C(_0438_),
    .Y(_0073_));
 sg13g2_and2_1 _2628_ (.A(net193),
    .B(_0438_),
    .X(_0439_));
 sg13g2_o21ai_1 _2629_ (.B1(net588),
    .Y(_0440_),
    .A1(net193),
    .A2(_0438_));
 sg13g2_nor2_1 _2630_ (.A(_0439_),
    .B(_0440_),
    .Y(_0074_));
 sg13g2_xnor2_1 _2631_ (.Y(_0441_),
    .A(net204),
    .B(_0439_));
 sg13g2_nor2_1 _2632_ (.A(_0434_),
    .B(_0441_),
    .Y(_0075_));
 sg13g2_a21oi_1 _2633_ (.A1(\music.note_pos[12] ),
    .A2(_0439_),
    .Y(_0442_),
    .B1(net132));
 sg13g2_nand3_1 _2634_ (.B(net204),
    .C(_0439_),
    .A(net132),
    .Y(_0443_));
 sg13g2_nand2_1 _2635_ (.Y(_0444_),
    .A(net587),
    .B(_0443_));
 sg13g2_nor2_1 _2636_ (.A(net133),
    .B(_0444_),
    .Y(_0076_));
 sg13g2_nand2_1 _2637_ (.Y(_0445_),
    .A(_0515_),
    .B(_0443_));
 sg13g2_or2_1 _2638_ (.X(_0446_),
    .B(_0443_),
    .A(_0515_));
 sg13g2_and4_1 _2639_ (.A(net588),
    .B(_0421_),
    .C(_0445_),
    .D(_0446_),
    .X(_0077_));
 sg13g2_xor2_1 _2640_ (.B(_0446_),
    .A(net218),
    .X(_0447_));
 sg13g2_nor2_1 _2641_ (.A(_0419_),
    .B(_0447_),
    .Y(_0078_));
 sg13g2_nor2_1 _2642_ (.A(\music.note[0] ),
    .B(\music.note[1] ),
    .Y(_0448_));
 sg13g2_or2_1 _2643_ (.X(_0449_),
    .B(\music.note[1] ),
    .A(\music.note[0] ));
 sg13g2_a21oi_1 _2644_ (.A1(_0534_),
    .A2(\music.note[1] ),
    .Y(_0450_),
    .B1(\music.note[0] ));
 sg13g2_and3_1 _2645_ (.X(_0451_),
    .A(\music.do_note ),
    .B(net586),
    .C(_0557_));
 sg13g2_inv_1 _2646_ (.Y(_0452_),
    .A(net517));
 sg13g2_nand2_1 _2647_ (.Y(_0453_),
    .A(_0450_),
    .B(net518));
 sg13g2_xnor2_1 _2648_ (.Y(_0079_),
    .A(net122),
    .B(_0453_));
 sg13g2_nor2_1 _2649_ (.A(\music.note[0] ),
    .B(\music.note[2] ),
    .Y(_0454_));
 sg13g2_nand2_1 _2650_ (.Y(_0455_),
    .A(\music.extended_sample[1] ),
    .B(_0454_));
 sg13g2_xor2_1 _2651_ (.B(_0454_),
    .A(\music.extended_sample[1] ),
    .X(_0456_));
 sg13g2_nand3_1 _2652_ (.B(_0450_),
    .C(_0456_),
    .A(\music.extended_sample[0] ),
    .Y(_0457_));
 sg13g2_a21o_1 _2653_ (.A2(_0450_),
    .A1(\music.extended_sample[0] ),
    .B1(_0456_),
    .X(_0458_));
 sg13g2_and2_1 _2654_ (.A(_0457_),
    .B(_0458_),
    .X(_0459_));
 sg13g2_mux2_1 _2655_ (.A0(net175),
    .A1(_0459_),
    .S(net518),
    .X(_0080_));
 sg13g2_nor2_1 _2656_ (.A(net161),
    .B(net518),
    .Y(_0460_));
 sg13g2_nand2b_1 _2657_ (.Y(_0461_),
    .B(\music.note[0] ),
    .A_N(\music.note[1] ));
 sg13g2_mux2_1 _2658_ (.A0(\music.note[0] ),
    .A1(_0461_),
    .S(_0534_),
    .X(_0462_));
 sg13g2_nor2b_1 _2659_ (.A(_0462_),
    .B_N(\music.extended_sample[2] ),
    .Y(_0463_));
 sg13g2_xor2_1 _2660_ (.B(_0462_),
    .A(\music.extended_sample[2] ),
    .X(_0464_));
 sg13g2_a21oi_1 _2661_ (.A1(_0455_),
    .A2(_0457_),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_and3_1 _2662_ (.X(_0466_),
    .A(_0455_),
    .B(_0457_),
    .C(_0464_));
 sg13g2_o21ai_1 _2663_ (.B1(net518),
    .Y(_0467_),
    .A1(_0465_),
    .A2(_0466_));
 sg13g2_nor2b_1 _2664_ (.A(_0460_),
    .B_N(_0467_),
    .Y(_0081_));
 sg13g2_nand2_1 _2665_ (.Y(_0468_),
    .A(_0004_),
    .B(_0461_));
 sg13g2_nand2_1 _2666_ (.Y(_0469_),
    .A(\music.extended_sample[3] ),
    .B(_0468_));
 sg13g2_xnor2_1 _2667_ (.Y(_0470_),
    .A(_0535_),
    .B(_0468_));
 sg13g2_or3_1 _2668_ (.A(_0463_),
    .B(_0465_),
    .C(_0470_),
    .X(_0471_));
 sg13g2_o21ai_1 _2669_ (.B1(_0470_),
    .Y(_0472_),
    .A1(_0463_),
    .A2(_0465_));
 sg13g2_a21oi_1 _2670_ (.A1(_0471_),
    .A2(_0472_),
    .Y(_0473_),
    .B1(_0452_));
 sg13g2_a21oi_1 _2671_ (.A1(_0535_),
    .A2(_0452_),
    .Y(_0082_),
    .B1(_0473_));
 sg13g2_nand2_1 _2672_ (.Y(_0474_),
    .A(net124),
    .B(_0452_));
 sg13g2_a21oi_1 _2673_ (.A1(_0004_),
    .A2(_0449_),
    .Y(_0475_),
    .B1(net124));
 sg13g2_nand3_1 _2674_ (.B(net124),
    .C(_0449_),
    .A(_0004_),
    .Y(_0476_));
 sg13g2_nor2b_1 _2675_ (.A(_0475_),
    .B_N(_0476_),
    .Y(_0477_));
 sg13g2_nand2_1 _2676_ (.Y(_0478_),
    .A(_0469_),
    .B(_0472_));
 sg13g2_and2_1 _2677_ (.A(_0477_),
    .B(_0478_),
    .X(_0479_));
 sg13g2_inv_1 _2678_ (.Y(_0480_),
    .A(_0479_));
 sg13g2_o21ai_1 _2679_ (.B1(net517),
    .Y(_0481_),
    .A1(_0477_),
    .A2(_0478_));
 sg13g2_o21ai_1 _2680_ (.B1(_0474_),
    .Y(_0083_),
    .A1(_0479_),
    .A2(_0481_));
 sg13g2_nor2_1 _2681_ (.A(net168),
    .B(net517),
    .Y(_0482_));
 sg13g2_nand2_1 _2682_ (.Y(_0483_),
    .A(_0476_),
    .B(_0480_));
 sg13g2_nor2_1 _2683_ (.A(\music.note[2] ),
    .B(_0449_),
    .Y(_0484_));
 sg13g2_nand2_1 _2684_ (.Y(_0485_),
    .A(_0536_),
    .B(_0484_));
 sg13g2_xnor2_1 _2685_ (.Y(_0486_),
    .A(net168),
    .B(_0484_));
 sg13g2_xnor2_1 _2686_ (.Y(_0487_),
    .A(_0483_),
    .B(_0486_));
 sg13g2_a21oi_1 _2687_ (.A1(net517),
    .A2(_0487_),
    .Y(_0084_),
    .B1(_0482_));
 sg13g2_nor2_1 _2688_ (.A(net135),
    .B(net517),
    .Y(_0488_));
 sg13g2_a21oi_1 _2689_ (.A1(_0004_),
    .A2(_0448_),
    .Y(_0489_),
    .B1(\music.extended_sample[6] ));
 sg13g2_and3_1 _2690_ (.X(_0490_),
    .A(_0004_),
    .B(\music.extended_sample[6] ),
    .C(_0448_));
 sg13g2_or2_1 _2691_ (.X(_0491_),
    .B(_0490_),
    .A(_0489_));
 sg13g2_o21ai_1 _2692_ (.B1(_0476_),
    .Y(_0492_),
    .A1(_0536_),
    .A2(_0484_));
 sg13g2_a21oi_1 _2693_ (.A1(_0479_),
    .A2(_0485_),
    .Y(_0493_),
    .B1(_0492_));
 sg13g2_nor2_1 _2694_ (.A(_0491_),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_xnor2_1 _2695_ (.Y(_0495_),
    .A(_0491_),
    .B(_0493_));
 sg13g2_a21oi_1 _2696_ (.A1(net517),
    .A2(_0495_),
    .Y(_0085_),
    .B1(_0488_));
 sg13g2_nor2_1 _2697_ (.A(_0490_),
    .B(_0494_),
    .Y(_0496_));
 sg13g2_nor3_2 _2698_ (.A(_0005_),
    .B(_0452_),
    .C(_0496_),
    .Y(_0497_));
 sg13g2_nor2_1 _2699_ (.A(net120),
    .B(net517),
    .Y(_0498_));
 sg13g2_and3_1 _2700_ (.X(_0499_),
    .A(_0005_),
    .B(net517),
    .C(_0496_));
 sg13g2_nor3_1 _2701_ (.A(_0497_),
    .B(_0498_),
    .C(_0499_),
    .Y(_0086_));
 sg13g2_and2_1 _2702_ (.A(net130),
    .B(_0497_),
    .X(_0500_));
 sg13g2_xor2_1 _2703_ (.B(_0497_),
    .A(net130),
    .X(_0087_));
 sg13g2_xnor2_1 _2704_ (.Y(_0088_),
    .A(_0526_),
    .B(_0500_));
 sg13g2_a21oi_1 _2705_ (.A1(\music.extended_sample[9] ),
    .A2(_0500_),
    .Y(_0501_),
    .B1(net158));
 sg13g2_nand3_1 _2706_ (.B(net158),
    .C(_0500_),
    .A(\music.extended_sample[9] ),
    .Y(_0502_));
 sg13g2_nor2b_1 _2707_ (.A(net159),
    .B_N(_0502_),
    .Y(_0089_));
 sg13g2_nand4_1 _2708_ (.B(net169),
    .C(net158),
    .A(\music.extended_sample[9] ),
    .Y(_0503_),
    .D(_0500_));
 sg13g2_xnor2_1 _2709_ (.Y(_0090_),
    .A(net169),
    .B(_0502_));
 sg13g2_nor2_1 _2710_ (.A(_0529_),
    .B(_0503_),
    .Y(_0504_));
 sg13g2_xnor2_1 _2711_ (.Y(_0091_),
    .A(net126),
    .B(_0503_));
 sg13g2_nor3_1 _2712_ (.A(_0528_),
    .B(_0529_),
    .C(_0503_),
    .Y(_0505_));
 sg13g2_xnor2_1 _2713_ (.Y(_0092_),
    .A(_0528_),
    .B(_0504_));
 sg13g2_xor2_1 _2714_ (.B(_0505_),
    .A(net128),
    .X(_0093_));
 sg13g2_nand2_1 _2715_ (.Y(_0506_),
    .A(\music.melody_pos[0] ),
    .B(_0570_));
 sg13g2_o21ai_1 _2716_ (.B1(_0506_),
    .Y(_0094_),
    .A1(net583),
    .A2(net113));
 sg13g2_nand2_1 _2717_ (.Y(_0507_),
    .A(net236),
    .B(_0567_));
 sg13g2_a21o_1 _2718_ (.A2(_0507_),
    .A1(_0580_),
    .B1(net583),
    .X(_0508_));
 sg13g2_inv_1 _2719_ (.Y(_0095_),
    .A(_0508_));
 sg13g2_o21ai_1 _2720_ (.B1(_0595_),
    .Y(_0098_),
    .A1(_0514_),
    .A2(_0571_));
 sg13g2_mux2_1 _2721_ (.A0(\gfx.frame_counter[0] ),
    .A1(net108),
    .S(net514),
    .X(_0099_));
 sg13g2_nand3_1 _2722_ (.B(net228),
    .C(net514),
    .A(\gfx.frame_counter[0] ),
    .Y(_0509_));
 sg13g2_a21o_1 _2723_ (.A2(net514),
    .A1(\gfx.frame_counter[0] ),
    .B1(net228),
    .X(_0510_));
 sg13g2_and2_1 _2724_ (.A(_0509_),
    .B(net229),
    .X(_0100_));
 sg13g2_nand4_1 _2725_ (.B(net228),
    .C(net115),
    .A(net233),
    .Y(_0511_),
    .D(net513));
 sg13g2_xnor2_1 _2726_ (.Y(_0101_),
    .A(net115),
    .B(_0509_));
 sg13g2_nor2_2 _2727_ (.A(_0533_),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_xnor2_1 _2728_ (.Y(_0102_),
    .A(net110),
    .B(_0511_));
 sg13g2_xnor2_1 _2729_ (.Y(_0103_),
    .A(net562),
    .B(_0512_));
 sg13g2_o21ai_1 _2730_ (.B1(_0570_),
    .Y(_0104_),
    .A1(_0513_),
    .A2(_0422_));
 sg13g2_dfrbp_1 _2731_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net33),
    .D(_0019_),
    .Q_N(_1361_),
    .Q(\music.note_length ));
 sg13g2_dfrbp_1 _2732_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net62),
    .D(_0020_),
    .Q_N(_0018_),
    .Q(\music.pwm_pos[0] ));
 sg13g2_dfrbp_1 _2733_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net61),
    .D(_0021_),
    .Q_N(_1360_),
    .Q(\music.pwm_pos[1] ));
 sg13g2_dfrbp_1 _2734_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net60),
    .D(net145),
    .Q_N(_1359_),
    .Q(\music.pwm_pos[2] ));
 sg13g2_dfrbp_1 _2735_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net59),
    .D(_0023_),
    .Q_N(_1358_),
    .Q(\music.pwm_pos[3] ));
 sg13g2_dfrbp_1 _2736_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net58),
    .D(_0024_),
    .Q_N(_1357_),
    .Q(\music.pwm_pos[4] ));
 sg13g2_dfrbp_1 _2737_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net57),
    .D(_0025_),
    .Q_N(_1356_),
    .Q(\music.pwm_pos[5] ));
 sg13g2_dfrbp_1 _2738_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net56),
    .D(_0026_),
    .Q_N(_1355_),
    .Q(\music.pwm_pos[6] ));
 sg13g2_dfrbp_1 _2739_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net55),
    .D(net174),
    .Q_N(_1354_),
    .Q(\music.pwm_pos[7] ));
 sg13g2_dfrbp_1 _2740_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net54),
    .D(_0028_),
    .Q_N(_1353_),
    .Q(\music.pwm_pos[8] ));
 sg13g2_dfrbp_1 _2741_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net53),
    .D(_0029_),
    .Q_N(_1352_),
    .Q(\music.pwm_pos[9] ));
 sg13g2_dfrbp_1 _2742_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net52),
    .D(net140),
    .Q_N(_1351_),
    .Q(\music.pwm_pos[10] ));
 sg13g2_dfrbp_1 _2743_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net51),
    .D(_0031_),
    .Q_N(_1350_),
    .Q(\music.pwm_pos[11] ));
 sg13g2_dfrbp_1 _2744_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net50),
    .D(_0032_),
    .Q_N(_1349_),
    .Q(\music.pwm_pos[12] ));
 sg13g2_dfrbp_1 _2745_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net49),
    .D(_0033_),
    .Q_N(_1348_),
    .Q(\music.pwm_pos[13] ));
 sg13g2_dfrbp_1 _2746_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(_0034_),
    .Q_N(_1347_),
    .Q(\music.pwm_pos[14] ));
 sg13g2_dfrbp_1 _2747_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net47),
    .D(net148),
    .Q_N(_1346_),
    .Q(\gfx.vsync ));
 sg13g2_dfrbp_1 _2748_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net34),
    .D(net232),
    .Q_N(_1362_),
    .Q(\gfx.hsync ));
 sg13g2_dfrbp_1 _2749_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net35),
    .D(_0000_),
    .Q_N(_1363_),
    .Q(\music.note[0] ));
 sg13g2_dfrbp_1 _2750_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net29),
    .D(_0001_),
    .Q_N(_1364_),
    .Q(\music.note[1] ));
 sg13g2_dfrbp_1 _2751_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net45),
    .D(_0002_),
    .Q_N(_0004_),
    .Q(\music.note[2] ));
 sg13g2_dfrbp_1 _2752_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net43),
    .D(_0037_),
    .Q_N(_1345_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2753_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net42),
    .D(_0038_),
    .Q_N(_1344_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _2754_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net41),
    .D(_0039_),
    .Q_N(_0017_),
    .Q(\gfx.pixel_x[0] ));
 sg13g2_dfrbp_1 _2755_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net39),
    .D(net240),
    .Q_N(_1343_),
    .Q(\gfx.pixel_x[1] ));
 sg13g2_dfrbp_1 _2756_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net37),
    .D(_0041_),
    .Q_N(_1342_),
    .Q(\gfx.pixel_x[2] ));
 sg13g2_dfrbp_1 _2757_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net32),
    .D(_0042_),
    .Q_N(_1341_),
    .Q(\gfx.bitmap_x[0] ));
 sg13g2_dfrbp_1 _2758_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net30),
    .D(_0043_),
    .Q_N(_0014_),
    .Q(\gfx.bitmap_x[1] ));
 sg13g2_dfrbp_1 _2759_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net28),
    .D(_0044_),
    .Q_N(_1340_),
    .Q(\gfx.bitmap_x[2] ));
 sg13g2_dfrbp_1 _2760_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net26),
    .D(_0045_),
    .Q_N(_1339_),
    .Q(\gfx.bitmap_x[3] ));
 sg13g2_dfrbp_1 _2761_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net24),
    .D(net154),
    .Q_N(_1338_),
    .Q(\gfx.pixel_x[7] ));
 sg13g2_dfrbp_1 _2762_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net22),
    .D(_0047_),
    .Q_N(_1337_),
    .Q(\gfx.pixel_x[8] ));
 sg13g2_dfrbp_1 _2763_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net20),
    .D(_0048_),
    .Q_N(_1336_),
    .Q(\gfx.pixel_x[9] ));
 sg13g2_dfrbp_1 _2764_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net18),
    .D(_0049_),
    .Q_N(_1335_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2765_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net17),
    .D(_0050_),
    .Q_N(_1334_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2766_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net16),
    .D(_0051_),
    .Q_N(_0016_),
    .Q(\gfx.pixel_y[0] ));
 sg13g2_dfrbp_1 _2767_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net103),
    .D(net119),
    .Q_N(_1333_),
    .Q(\gfx.pixel_y[1] ));
 sg13g2_dfrbp_1 _2768_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net101),
    .D(_0053_),
    .Q_N(_1332_),
    .Q(\gfx.pixel_y[2] ));
 sg13g2_dfrbp_1 _2769_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net99),
    .D(_0054_),
    .Q_N(_0012_),
    .Q(\gfx.bitmap_y[0] ));
 sg13g2_dfrbp_1 _2770_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net97),
    .D(_0055_),
    .Q_N(_0013_),
    .Q(\gfx.bitmap_y[1] ));
 sg13g2_dfrbp_1 _2771_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net95),
    .D(_0056_),
    .Q_N(_1331_),
    .Q(\gfx.bitmap_y[2] ));
 sg13g2_dfrbp_1 _2772_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net93),
    .D(_0057_),
    .Q_N(_0011_),
    .Q(\gfx.bitmap_y[3] ));
 sg13g2_dfrbp_1 _2773_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net91),
    .D(_0058_),
    .Q_N(_0010_),
    .Q(\gfx.pixel_y[7] ));
 sg13g2_dfrbp_1 _2774_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net89),
    .D(_0059_),
    .Q_N(_1330_),
    .Q(\gfx.pixel_y[8] ));
 sg13g2_dfrbp_1 _2775_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net87),
    .D(_0060_),
    .Q_N(_1329_),
    .Q(\gfx.pixel_y[9] ));
 sg13g2_dfrbp_1 _2776_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net85),
    .D(_0061_),
    .Q_N(_1328_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2777_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net84),
    .D(_0062_),
    .Q_N(_1327_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _2778_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net83),
    .D(_0063_),
    .Q_N(_1326_),
    .Q(\music.note_pos[0] ));
 sg13g2_dfrbp_1 _2779_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net81),
    .D(_0064_),
    .Q_N(_1325_),
    .Q(\music.note_pos[1] ));
 sg13g2_dfrbp_1 _2780_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net79),
    .D(net166),
    .Q_N(_1324_),
    .Q(\music.note_pos[2] ));
 sg13g2_dfrbp_1 _2781_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net77),
    .D(_0066_),
    .Q_N(_1323_),
    .Q(\music.note_pos[3] ));
 sg13g2_dfrbp_1 _2782_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net75),
    .D(_0067_),
    .Q_N(_1322_),
    .Q(\music.note_pos[4] ));
 sg13g2_dfrbp_1 _2783_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net73),
    .D(_0068_),
    .Q_N(_1321_),
    .Q(\music.note_pos[5] ));
 sg13g2_dfrbp_1 _2784_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net71),
    .D(_0069_),
    .Q_N(_1320_),
    .Q(\music.note_pos[6] ));
 sg13g2_dfrbp_1 _2785_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net69),
    .D(net181),
    .Q_N(_1319_),
    .Q(\music.note_pos[7] ));
 sg13g2_dfrbp_1 _2786_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net67),
    .D(_0071_),
    .Q_N(_1318_),
    .Q(\music.note_pos[8] ));
 sg13g2_dfrbp_1 _2787_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net65),
    .D(net137),
    .Q_N(_1317_),
    .Q(\music.note_pos[9] ));
 sg13g2_dfrbp_1 _2788_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net63),
    .D(_0073_),
    .Q_N(_1316_),
    .Q(\music.note_pos[10] ));
 sg13g2_dfrbp_1 _2789_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net44),
    .D(_0074_),
    .Q_N(_1315_),
    .Q(\music.note_pos[11] ));
 sg13g2_dfrbp_1 _2790_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net38),
    .D(_0075_),
    .Q_N(_1314_),
    .Q(\music.note_pos[12] ));
 sg13g2_dfrbp_1 _2791_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net31),
    .D(net134),
    .Q_N(_1313_),
    .Q(\music.note_pos[13] ));
 sg13g2_dfrbp_1 _2792_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net27),
    .D(_0077_),
    .Q_N(_1312_),
    .Q(\music.note_pos[14] ));
 sg13g2_dfrbp_1 _2793_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net23),
    .D(_0078_),
    .Q_N(_1311_),
    .Q(\music.note_pos[15] ));
 sg13g2_dfrbp_1 _2794_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net19),
    .D(net123),
    .Q_N(_1310_),
    .Q(\music.extended_sample[0] ));
 sg13g2_dfrbp_1 _2795_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net15),
    .D(net176),
    .Q_N(_1309_),
    .Q(\music.extended_sample[1] ));
 sg13g2_dfrbp_1 _2796_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net102),
    .D(_0081_),
    .Q_N(_1308_),
    .Q(\music.extended_sample[2] ));
 sg13g2_dfrbp_1 _2797_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net100),
    .D(_0082_),
    .Q_N(_1307_),
    .Q(\music.extended_sample[3] ));
 sg13g2_dfrbp_1 _2798_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net98),
    .D(net125),
    .Q_N(_1306_),
    .Q(\music.extended_sample[4] ));
 sg13g2_dfrbp_1 _2799_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net96),
    .D(_0084_),
    .Q_N(_1305_),
    .Q(\music.extended_sample[5] ));
 sg13g2_dfrbp_1 _2800_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net94),
    .D(_0085_),
    .Q_N(_1304_),
    .Q(\music.extended_sample[6] ));
 sg13g2_dfrbp_1 _2801_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net92),
    .D(net121),
    .Q_N(_0005_),
    .Q(\music.extended_sample[7] ));
 sg13g2_dfrbp_1 _2802_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net90),
    .D(net131),
    .Q_N(_1303_),
    .Q(\music.extended_sample[8] ));
 sg13g2_dfrbp_1 _2803_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net88),
    .D(net227),
    .Q_N(_1302_),
    .Q(\music.extended_sample[9] ));
 sg13g2_dfrbp_1 _2804_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net86),
    .D(net160),
    .Q_N(_1301_),
    .Q(\music.extended_sample[10] ));
 sg13g2_dfrbp_1 _2805_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net82),
    .D(net170),
    .Q_N(_1300_),
    .Q(\music.extended_sample[11] ));
 sg13g2_dfrbp_1 _2806_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net80),
    .D(net127),
    .Q_N(_1299_),
    .Q(\music.extended_sample[12] ));
 sg13g2_dfrbp_1 _2807_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net78),
    .D(net209),
    .Q_N(_1298_),
    .Q(\music.extended_sample[13] ));
 sg13g2_dfrbp_1 _2808_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net76),
    .D(net129),
    .Q_N(_1297_),
    .Q(\music.extended_sample[14] ));
 sg13g2_dfrbp_1 _2809_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net74),
    .D(net114),
    .Q_N(_0006_),
    .Q(\music.melody_pos[0] ));
 sg13g2_dfrbp_1 _2810_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net70),
    .D(_0095_),
    .Q_N(_0003_),
    .Q(\music.melody_pos[1] ));
 sg13g2_dfrbp_1 _2811_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net66),
    .D(_0096_),
    .Q_N(_0007_),
    .Q(\music.melody_pos[2] ));
 sg13g2_dfrbp_1 _2812_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net46),
    .D(_0097_),
    .Q_N(_1296_),
    .Q(\music.melody_pos[3] ));
 sg13g2_dfrbp_1 _2813_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net36),
    .D(net152),
    .Q_N(_0008_),
    .Q(\music.melody_pos[4] ));
 sg13g2_dfrbp_1 _2814_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net25),
    .D(net109),
    .Q_N(_0015_),
    .Q(\gfx.frame_counter[0] ));
 sg13g2_dfrbp_1 _2815_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net21),
    .D(net230),
    .Q_N(_1295_),
    .Q(\gfx.frame_counter[1] ));
 sg13g2_dfrbp_1 _2816_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net72),
    .D(net116),
    .Q_N(_1294_),
    .Q(\gfx.frame_counter[2] ));
 sg13g2_dfrbp_1 _2817_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net68),
    .D(net111),
    .Q_N(_1293_),
    .Q(\gfx.frame_counter[3] ));
 sg13g2_dfrbp_1 _2818_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net64),
    .D(_0103_),
    .Q_N(_0009_),
    .Q(\gfx.frame_counter[4] ));
 sg13g2_dfrbp_1 _2819_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net40),
    .D(_0104_),
    .Q_N(_1292_),
    .Q(\music.do_note ));
 sg13g2_tiehi _2766__16 (.L_HI(net16));
 sg13g2_tiehi _2765__17 (.L_HI(net17));
 sg13g2_tiehi _2764__18 (.L_HI(net18));
 sg13g2_tiehi _2794__19 (.L_HI(net19));
 sg13g2_tiehi _2763__20 (.L_HI(net20));
 sg13g2_tiehi _2815__21 (.L_HI(net21));
 sg13g2_tiehi _2762__22 (.L_HI(net22));
 sg13g2_tiehi _2793__23 (.L_HI(net23));
 sg13g2_tiehi _2761__24 (.L_HI(net24));
 sg13g2_tiehi _2814__25 (.L_HI(net25));
 sg13g2_tiehi _2760__26 (.L_HI(net26));
 sg13g2_tiehi _2792__27 (.L_HI(net27));
 sg13g2_tiehi _2759__28 (.L_HI(net28));
 sg13g2_tiehi _2750__29 (.L_HI(net29));
 sg13g2_tiehi _2758__30 (.L_HI(net30));
 sg13g2_tiehi _2791__31 (.L_HI(net31));
 sg13g2_tiehi _2757__32 (.L_HI(net32));
 sg13g2_tiehi _2731__33 (.L_HI(net33));
 sg13g2_tiehi _2748__34 (.L_HI(net34));
 sg13g2_tiehi _2749__35 (.L_HI(net35));
 sg13g2_tiehi _2813__36 (.L_HI(net36));
 sg13g2_tiehi _2756__37 (.L_HI(net37));
 sg13g2_tiehi _2790__38 (.L_HI(net38));
 sg13g2_tiehi _2755__39 (.L_HI(net39));
 sg13g2_tiehi _2819__40 (.L_HI(net40));
 sg13g2_tiehi _2754__41 (.L_HI(net41));
 sg13g2_tiehi _2753__42 (.L_HI(net42));
 sg13g2_tiehi _2752__43 (.L_HI(net43));
 sg13g2_tiehi _2789__44 (.L_HI(net44));
 sg13g2_tiehi _2751__45 (.L_HI(net45));
 sg13g2_tiehi _2812__46 (.L_HI(net46));
 sg13g2_tiehi _2747__47 (.L_HI(net47));
 sg13g2_tiehi _2746__48 (.L_HI(net48));
 sg13g2_tiehi _2745__49 (.L_HI(net49));
 sg13g2_tiehi _2744__50 (.L_HI(net50));
 sg13g2_tiehi _2743__51 (.L_HI(net51));
 sg13g2_tiehi _2742__52 (.L_HI(net52));
 sg13g2_tiehi _2741__53 (.L_HI(net53));
 sg13g2_tiehi _2740__54 (.L_HI(net54));
 sg13g2_tiehi _2739__55 (.L_HI(net55));
 sg13g2_tiehi _2738__56 (.L_HI(net56));
 sg13g2_tiehi _2737__57 (.L_HI(net57));
 sg13g2_tiehi _2736__58 (.L_HI(net58));
 sg13g2_tiehi _2735__59 (.L_HI(net59));
 sg13g2_tiehi _2734__60 (.L_HI(net60));
 sg13g2_tiehi _2733__61 (.L_HI(net61));
 sg13g2_tiehi _2732__62 (.L_HI(net62));
 sg13g2_tiehi _2788__63 (.L_HI(net63));
 sg13g2_tiehi _2818__64 (.L_HI(net64));
 sg13g2_tiehi _2787__65 (.L_HI(net65));
 sg13g2_tiehi _2811__66 (.L_HI(net66));
 sg13g2_tiehi _2786__67 (.L_HI(net67));
 sg13g2_tiehi _2817__68 (.L_HI(net68));
 sg13g2_tiehi _2785__69 (.L_HI(net69));
 sg13g2_tiehi _2810__70 (.L_HI(net70));
 sg13g2_tiehi _2784__71 (.L_HI(net71));
 sg13g2_tiehi _2816__72 (.L_HI(net72));
 sg13g2_tiehi _2783__73 (.L_HI(net73));
 sg13g2_tiehi _2809__74 (.L_HI(net74));
 sg13g2_tiehi _2782__75 (.L_HI(net75));
 sg13g2_tiehi _2808__76 (.L_HI(net76));
 sg13g2_tiehi _2781__77 (.L_HI(net77));
 sg13g2_tiehi _2807__78 (.L_HI(net78));
 sg13g2_tiehi _2780__79 (.L_HI(net79));
 sg13g2_tiehi _2806__80 (.L_HI(net80));
 sg13g2_tiehi _2779__81 (.L_HI(net81));
 sg13g2_tiehi _2805__82 (.L_HI(net82));
 sg13g2_tiehi _2778__83 (.L_HI(net83));
 sg13g2_tiehi _2777__84 (.L_HI(net84));
 sg13g2_tiehi _2776__85 (.L_HI(net85));
 sg13g2_tiehi _2804__86 (.L_HI(net86));
 sg13g2_tiehi _2775__87 (.L_HI(net87));
 sg13g2_tiehi _2803__88 (.L_HI(net88));
 sg13g2_tiehi _2774__89 (.L_HI(net89));
 sg13g2_tiehi _2802__90 (.L_HI(net90));
 sg13g2_tiehi _2773__91 (.L_HI(net91));
 sg13g2_tiehi _2801__92 (.L_HI(net92));
 sg13g2_tiehi _2772__93 (.L_HI(net93));
 sg13g2_tiehi _2800__94 (.L_HI(net94));
 sg13g2_tiehi _2771__95 (.L_HI(net95));
 sg13g2_tiehi _2799__96 (.L_HI(net96));
 sg13g2_tiehi _2770__97 (.L_HI(net97));
 sg13g2_tiehi _2798__98 (.L_HI(net98));
 sg13g2_tiehi _2769__99 (.L_HI(net99));
 sg13g2_tiehi _2797__100 (.L_HI(net100));
 sg13g2_tiehi _2768__101 (.L_HI(net101));
 sg13g2_tiehi _2796__102 (.L_HI(net102));
 sg13g2_tiehi _2767__103 (.L_HI(net103));
 sg13g2_tiehi tt_um_nyan_104 (.L_HI(net104));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_nyan_2 (.L_LO(net2));
 sg13g2_tielo tt_um_nyan_3 (.L_LO(net3));
 sg13g2_tielo tt_um_nyan_4 (.L_LO(net4));
 sg13g2_tielo tt_um_nyan_5 (.L_LO(net5));
 sg13g2_tielo tt_um_nyan_6 (.L_LO(net6));
 sg13g2_tielo tt_um_nyan_7 (.L_LO(net7));
 sg13g2_tielo tt_um_nyan_8 (.L_LO(net8));
 sg13g2_tielo tt_um_nyan_9 (.L_LO(net9));
 sg13g2_tielo tt_um_nyan_10 (.L_LO(net10));
 sg13g2_tielo tt_um_nyan_11 (.L_LO(net11));
 sg13g2_tielo tt_um_nyan_12 (.L_LO(net12));
 sg13g2_tielo tt_um_nyan_13 (.L_LO(net13));
 sg13g2_tielo tt_um_nyan_14 (.L_LO(net14));
 sg13g2_tiehi _2795__15 (.L_HI(net15));
 sg13g2_buf_1 _2924_ (.A(\music.pwm ),
    .X(uio_out[7]));
 sg13g2_buf_1 _2925_ (.A(\gfx.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2926_ (.A(\gfx.hsync ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout444 (.A(_0274_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(net446),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_1256_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_0913_),
    .X(net448));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(_0813_));
 sg13g2_buf_4 fanout450 (.X(net450),
    .A(_0818_));
 sg13g2_buf_2 fanout451 (.A(_0818_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(net454),
    .X(net452));
 sg13g2_buf_1 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(_0744_));
 sg13g2_buf_2 fanout455 (.A(net458),
    .X(net455));
 sg13g2_buf_4 fanout456 (.X(net456),
    .A(net458));
 sg13g2_buf_1 fanout457 (.A(net458),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_0743_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(net460),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_0740_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_0740_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(net463),
    .X(net462));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(_0740_));
 sg13g2_buf_2 fanout464 (.A(net467),
    .X(net464));
 sg13g2_buf_1 fanout465 (.A(net467),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net467),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_0739_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(net469),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_1257_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(net472),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_1 fanout472 (.A(_0742_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(net476),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net476),
    .X(net474));
 sg13g2_buf_1 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_0742_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(net481),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(net480),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(net481),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_0741_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net484),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(net484),
    .X(net483));
 sg13g2_buf_1 fanout484 (.A(_0725_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net488),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(net487),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_0725_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(net493),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net492),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(net492),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(net493),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_0724_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(net496),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net496),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(net502),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net502),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net502),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(net501),
    .X(net499));
 sg13g2_buf_1 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(net502),
    .X(net501));
 sg13g2_buf_1 fanout502 (.A(_0763_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(net505),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(net505),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(net507),
    .X(net505));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(net507));
 sg13g2_buf_2 fanout507 (.A(_0762_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net510),
    .X(net508));
 sg13g2_buf_1 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(_0762_));
 sg13g2_buf_2 fanout511 (.A(net512),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_0762_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_0360_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_0360_),
    .X(net514));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(_0719_));
 sg13g2_buf_2 fanout516 (.A(_0919_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_0451_),
    .X(net517));
 sg13g2_buf_1 fanout518 (.A(_0451_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_0316_),
    .X(net519));
 sg13g2_buf_1 fanout520 (.A(_0316_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_0837_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_0837_),
    .X(net522));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(_0795_));
 sg13g2_buf_2 fanout524 (.A(_0751_),
    .X(net524));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(net526));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(net527));
 sg13g2_buf_2 fanout527 (.A(net532),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net530),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(net532),
    .X(net530));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(net532));
 sg13g2_buf_2 fanout532 (.A(_0746_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net537),
    .X(net534));
 sg13g2_buf_1 fanout535 (.A(net537),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_0745_),
    .X(net537));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(net541));
 sg13g2_buf_2 fanout539 (.A(net541),
    .X(net539));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(net541));
 sg13g2_buf_2 fanout541 (.A(_0745_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_0615_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_0615_),
    .X(net543));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(_0857_));
 sg13g2_buf_4 fanout545 (.X(net545),
    .A(net546));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(_0749_));
 sg13g2_buf_4 fanout547 (.X(net547),
    .A(net548));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(_0748_));
 sg13g2_buf_2 fanout549 (.A(net551),
    .X(net549));
 sg13g2_buf_1 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_0699_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_0698_),
    .X(net552));
 sg13g2_buf_1 fanout553 (.A(_0698_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_0662_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_0661_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_0661_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_0747_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_0747_),
    .X(net558));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(_0707_));
 sg13g2_buf_2 fanout560 (.A(net562),
    .X(net560));
 sg13g2_buf_1 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_0530_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(\gfx.frame_counter[4] ),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(\gfx.frame_counter[4] ),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(net244),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(\gfx.bitmap_y[2] ),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(\gfx.bitmap_y[2] ),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net570),
    .X(net568));
 sg13g2_buf_1 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(\gfx.bitmap_y[1] ),
    .X(net570));
 sg13g2_buf_4 fanout571 (.X(net571),
    .A(_0012_));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(net575));
 sg13g2_buf_2 fanout573 (.A(net575),
    .X(net573));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(net575));
 sg13g2_buf_2 fanout575 (.A(\gfx.bitmap_y[0] ),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net241),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(\gfx.pixel_x[7] ),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(\gfx.bitmap_x[3] ),
    .X(net579));
 sg13g2_buf_4 fanout580 (.X(net580),
    .A(net237));
 sg13g2_buf_2 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(\gfx.bitmap_x[1] ),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(net585),
    .X(net583));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(net585));
 sg13g2_buf_2 fanout585 (.A(_0521_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(rst_n));
 sg13g2_tielo tt_um_nyan_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0018_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0017_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0313_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0015_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0099_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold6 (.A(\gfx.frame_counter[3] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0102_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0006_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0582_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0094_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold11 (.A(\gfx.frame_counter[2] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0101_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold13 (.A(\gfx.pixel_y[1] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0364_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0052_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold16 (.A(\music.extended_sample[7] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0086_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold18 (.A(\music.extended_sample[0] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0079_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold20 (.A(\music.extended_sample[4] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0083_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold22 (.A(\music.extended_sample[12] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0091_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold24 (.A(\music.extended_sample[14] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0093_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold26 (.A(\music.extended_sample[8] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0087_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold28 (.A(\music.note_pos[13] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0442_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0076_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold31 (.A(\music.extended_sample[6] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold32 (.A(\music.note_pos[9] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0072_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold34 (.A(\music.pwm_pos[10] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0631_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0030_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold37 (.A(\music.note_pos[5] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0428_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold39 (.A(\music.pwm_pos[2] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0618_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0022_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold42 (.A(\gfx.vsync ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0645_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0035_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0016_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0363_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold47 (.A(\music.melody_pos[4] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0098_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold49 (.A(\gfx.pixel_x[7] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0046_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold51 (.A(\music.note_pos[10] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0437_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold53 (.A(\music.extended_sample[3] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold54 (.A(\music.extended_sample[10] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0501_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0089_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold57 (.A(\music.extended_sample[2] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold58 (.A(\music.pwm_pos[12] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0635_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold60 (.A(\music.note_pos[2] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0417_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0065_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold63 (.A(\music.pwm_pos[13] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold64 (.A(\music.extended_sample[5] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold65 (.A(\music.extended_sample[11] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0090_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold67 (.A(uo_out[1]),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold68 (.A(\music.pwm_pos[7] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0626_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0027_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold71 (.A(\music.extended_sample[1] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0080_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold73 (.A(\music.pwm_pos[3] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0620_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold75 (.A(\music.note_pos[7] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0431_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0070_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold78 (.A(\music.pwm_pos[11] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0633_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold80 (.A(\gfx.pixel_y[8] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0379_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold82 (.A(\music.pwm_pos[8] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0628_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold84 (.A(\music.note_pos[0] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold85 (.A(\music.pwm_pos[14] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold86 (.A(\music.pwm_pos[5] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0624_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold88 (.A(\gfx.pixel_y[9] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold89 (.A(\music.note_pos[11] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold90 (.A(\gfx.pixel_x[9] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0331_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold92 (.A(uo_out[6]),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold93 (.A(\music.pwm_pos[0] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0616_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold95 (.A(\music.pwm_pos[4] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold96 (.A(\gfx.pixel_y[2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0366_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0013_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0373_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold100 (.A(\music.note_pos[12] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold101 (.A(\music.note_pos[1] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold102 (.A(\music.note_pos[8] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold103 (.A(uo_out[0]),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold104 (.A(\music.extended_sample[13] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0092_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold106 (.A(\music.note_pos[3] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold107 (.A(uo_out[2]),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold108 (.A(\music.pwm_pos[9] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold109 (.A(uo_out[5]),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold110 (.A(\music.pwm_pos[6] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold111 (.A(\music.do_note ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold112 (.A(\gfx.pixel_x[2] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0319_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold114 (.A(\music.note_pos[15] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold115 (.A(\gfx.bitmap_y[3] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold116 (.A(\gfx.bitmap_x[0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0321_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold118 (.A(\music.note_pos[6] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0430_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0014_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0322_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold122 (.A(\music.extended_sample[9] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0088_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold124 (.A(\gfx.frame_counter[1] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0510_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0100_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold127 (.A(\gfx.hsync ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0036_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold129 (.A(\gfx.frame_counter[0] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold130 (.A(\music.note_pos[4] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold131 (.A(uo_out[4]),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold132 (.A(\music.melody_pos[1] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold133 (.A(\gfx.bitmap_x[2] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold134 (.A(\music.note_pos[14] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold135 (.A(\gfx.pixel_x[1] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0040_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold137 (.A(\gfx.pixel_x[8] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold138 (.A(\music.melody_pos[3] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0008_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold140 (.A(\gfx.pixel_y[7] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0003_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold142 (.A(\music.note_pos[6] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold143 (.A(\gfx.pixel_x[2] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold144 (.A(\music.note_pos[4] ),
    .X(net248));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_4 FILLER_2_133 ();
 sg13g2_fill_2 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_145 ();
 sg13g2_decap_8 FILLER_2_152 ();
 sg13g2_decap_4 FILLER_2_175 ();
 sg13g2_fill_1 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_fill_2 FILLER_2_215 ();
 sg13g2_fill_1 FILLER_2_217 ();
 sg13g2_fill_2 FILLER_2_222 ();
 sg13g2_fill_1 FILLER_2_224 ();
 sg13g2_decap_4 FILLER_2_241 ();
 sg13g2_fill_2 FILLER_2_245 ();
 sg13g2_fill_2 FILLER_2_259 ();
 sg13g2_decap_4 FILLER_2_272 ();
 sg13g2_fill_1 FILLER_2_276 ();
 sg13g2_decap_4 FILLER_2_282 ();
 sg13g2_fill_2 FILLER_2_291 ();
 sg13g2_fill_1 FILLER_2_293 ();
 sg13g2_decap_8 FILLER_2_297 ();
 sg13g2_decap_8 FILLER_2_304 ();
 sg13g2_decap_8 FILLER_2_311 ();
 sg13g2_decap_8 FILLER_2_318 ();
 sg13g2_decap_8 FILLER_2_325 ();
 sg13g2_decap_8 FILLER_2_332 ();
 sg13g2_decap_8 FILLER_2_339 ();
 sg13g2_fill_2 FILLER_2_346 ();
 sg13g2_fill_1 FILLER_2_348 ();
 sg13g2_decap_8 FILLER_2_353 ();
 sg13g2_decap_8 FILLER_2_360 ();
 sg13g2_decap_8 FILLER_2_367 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_4 FILLER_3_126 ();
 sg13g2_fill_1 FILLER_3_136 ();
 sg13g2_decap_4 FILLER_3_151 ();
 sg13g2_fill_2 FILLER_3_200 ();
 sg13g2_fill_2 FILLER_3_222 ();
 sg13g2_fill_1 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_246 ();
 sg13g2_fill_1 FILLER_3_253 ();
 sg13g2_fill_2 FILLER_3_271 ();
 sg13g2_fill_2 FILLER_3_292 ();
 sg13g2_fill_1 FILLER_3_306 ();
 sg13g2_decap_4 FILLER_3_324 ();
 sg13g2_fill_2 FILLER_3_328 ();
 sg13g2_fill_2 FILLER_3_340 ();
 sg13g2_fill_1 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_4 FILLER_4_112 ();
 sg13g2_fill_2 FILLER_4_132 ();
 sg13g2_decap_4 FILLER_4_154 ();
 sg13g2_fill_1 FILLER_4_163 ();
 sg13g2_decap_4 FILLER_4_173 ();
 sg13g2_fill_1 FILLER_4_177 ();
 sg13g2_fill_2 FILLER_4_202 ();
 sg13g2_fill_1 FILLER_4_204 ();
 sg13g2_fill_2 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_fill_1 FILLER_4_224 ();
 sg13g2_fill_1 FILLER_4_246 ();
 sg13g2_decap_4 FILLER_4_255 ();
 sg13g2_fill_1 FILLER_4_259 ();
 sg13g2_decap_4 FILLER_4_275 ();
 sg13g2_fill_2 FILLER_4_279 ();
 sg13g2_decap_4 FILLER_4_301 ();
 sg13g2_fill_1 FILLER_4_305 ();
 sg13g2_fill_1 FILLER_4_315 ();
 sg13g2_fill_1 FILLER_4_344 ();
 sg13g2_fill_2 FILLER_4_351 ();
 sg13g2_fill_1 FILLER_4_353 ();
 sg13g2_fill_2 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_2 FILLER_5_130 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_decap_4 FILLER_5_163 ();
 sg13g2_fill_2 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_184 ();
 sg13g2_fill_1 FILLER_5_198 ();
 sg13g2_fill_2 FILLER_5_207 ();
 sg13g2_decap_4 FILLER_5_245 ();
 sg13g2_fill_2 FILLER_5_249 ();
 sg13g2_fill_2 FILLER_5_256 ();
 sg13g2_fill_2 FILLER_5_266 ();
 sg13g2_fill_1 FILLER_5_268 ();
 sg13g2_fill_2 FILLER_5_302 ();
 sg13g2_fill_1 FILLER_5_304 ();
 sg13g2_decap_4 FILLER_5_328 ();
 sg13g2_decap_4 FILLER_5_341 ();
 sg13g2_fill_2 FILLER_5_345 ();
 sg13g2_fill_2 FILLER_5_351 ();
 sg13g2_fill_1 FILLER_5_353 ();
 sg13g2_fill_2 FILLER_5_370 ();
 sg13g2_fill_2 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_4 FILLER_5_403 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_4 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_134 ();
 sg13g2_fill_1 FILLER_6_136 ();
 sg13g2_fill_2 FILLER_6_166 ();
 sg13g2_fill_1 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_192 ();
 sg13g2_decap_4 FILLER_6_199 ();
 sg13g2_fill_2 FILLER_6_208 ();
 sg13g2_fill_1 FILLER_6_210 ();
 sg13g2_fill_2 FILLER_6_221 ();
 sg13g2_fill_2 FILLER_6_228 ();
 sg13g2_fill_2 FILLER_6_234 ();
 sg13g2_fill_1 FILLER_6_236 ();
 sg13g2_fill_2 FILLER_6_242 ();
 sg13g2_fill_1 FILLER_6_257 ();
 sg13g2_decap_4 FILLER_6_275 ();
 sg13g2_fill_2 FILLER_6_279 ();
 sg13g2_decap_4 FILLER_6_288 ();
 sg13g2_fill_1 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_fill_1 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_4 FILLER_6_356 ();
 sg13g2_fill_1 FILLER_6_360 ();
 sg13g2_decap_4 FILLER_6_375 ();
 sg13g2_fill_1 FILLER_6_379 ();
 sg13g2_fill_1 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_4 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_123 ();
 sg13g2_fill_1 FILLER_7_147 ();
 sg13g2_fill_2 FILLER_7_153 ();
 sg13g2_fill_2 FILLER_7_170 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_decap_4 FILLER_7_189 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_fill_2 FILLER_7_235 ();
 sg13g2_decap_4 FILLER_7_246 ();
 sg13g2_fill_1 FILLER_7_250 ();
 sg13g2_decap_4 FILLER_7_256 ();
 sg13g2_fill_2 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_270 ();
 sg13g2_fill_2 FILLER_7_288 ();
 sg13g2_fill_1 FILLER_7_306 ();
 sg13g2_fill_2 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_fill_2 FILLER_7_346 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_4 FILLER_8_112 ();
 sg13g2_fill_1 FILLER_8_132 ();
 sg13g2_fill_2 FILLER_8_141 ();
 sg13g2_fill_2 FILLER_8_164 ();
 sg13g2_fill_1 FILLER_8_166 ();
 sg13g2_decap_8 FILLER_8_180 ();
 sg13g2_fill_2 FILLER_8_187 ();
 sg13g2_fill_2 FILLER_8_204 ();
 sg13g2_fill_1 FILLER_8_206 ();
 sg13g2_fill_2 FILLER_8_212 ();
 sg13g2_fill_1 FILLER_8_214 ();
 sg13g2_fill_2 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_269 ();
 sg13g2_fill_2 FILLER_8_276 ();
 sg13g2_fill_1 FILLER_8_278 ();
 sg13g2_fill_1 FILLER_8_300 ();
 sg13g2_fill_2 FILLER_8_305 ();
 sg13g2_decap_4 FILLER_8_320 ();
 sg13g2_fill_2 FILLER_8_324 ();
 sg13g2_fill_1 FILLER_8_331 ();
 sg13g2_fill_1 FILLER_8_358 ();
 sg13g2_fill_2 FILLER_8_380 ();
 sg13g2_fill_1 FILLER_8_394 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_112 ();
 sg13g2_fill_1 FILLER_9_114 ();
 sg13g2_fill_2 FILLER_9_124 ();
 sg13g2_fill_1 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_148 ();
 sg13g2_fill_2 FILLER_9_155 ();
 sg13g2_fill_1 FILLER_9_157 ();
 sg13g2_decap_8 FILLER_9_176 ();
 sg13g2_fill_2 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_185 ();
 sg13g2_decap_4 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_234 ();
 sg13g2_fill_2 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_257 ();
 sg13g2_fill_1 FILLER_9_259 ();
 sg13g2_decap_4 FILLER_9_273 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_decap_4 FILLER_9_289 ();
 sg13g2_fill_1 FILLER_9_293 ();
 sg13g2_fill_1 FILLER_9_299 ();
 sg13g2_fill_1 FILLER_9_306 ();
 sg13g2_fill_2 FILLER_9_313 ();
 sg13g2_fill_2 FILLER_9_328 ();
 sg13g2_fill_2 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_367 ();
 sg13g2_decap_4 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_378 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_fill_2 FILLER_10_136 ();
 sg13g2_fill_1 FILLER_10_138 ();
 sg13g2_fill_1 FILLER_10_150 ();
 sg13g2_fill_2 FILLER_10_174 ();
 sg13g2_decap_4 FILLER_10_198 ();
 sg13g2_fill_2 FILLER_10_202 ();
 sg13g2_decap_4 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_fill_1 FILLER_10_231 ();
 sg13g2_fill_2 FILLER_10_236 ();
 sg13g2_fill_2 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_4 FILLER_10_256 ();
 sg13g2_fill_2 FILLER_10_272 ();
 sg13g2_fill_1 FILLER_10_274 ();
 sg13g2_fill_1 FILLER_10_289 ();
 sg13g2_decap_4 FILLER_10_318 ();
 sg13g2_fill_1 FILLER_10_322 ();
 sg13g2_fill_2 FILLER_10_327 ();
 sg13g2_decap_4 FILLER_10_340 ();
 sg13g2_fill_2 FILLER_10_344 ();
 sg13g2_fill_2 FILLER_10_350 ();
 sg13g2_fill_1 FILLER_10_352 ();
 sg13g2_decap_4 FILLER_10_357 ();
 sg13g2_fill_1 FILLER_10_361 ();
 sg13g2_fill_2 FILLER_10_380 ();
 sg13g2_fill_1 FILLER_10_382 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_4 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_38 ();
 sg13g2_fill_1 FILLER_11_45 ();
 sg13g2_fill_2 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_54 ();
 sg13g2_decap_8 FILLER_11_61 ();
 sg13g2_fill_1 FILLER_11_68 ();
 sg13g2_fill_1 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_92 ();
 sg13g2_decap_8 FILLER_11_99 ();
 sg13g2_decap_4 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_110 ();
 sg13g2_fill_1 FILLER_11_131 ();
 sg13g2_fill_2 FILLER_11_144 ();
 sg13g2_fill_1 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_1 FILLER_11_164 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_186 ();
 sg13g2_fill_2 FILLER_11_193 ();
 sg13g2_fill_1 FILLER_11_224 ();
 sg13g2_fill_1 FILLER_11_269 ();
 sg13g2_decap_4 FILLER_11_286 ();
 sg13g2_decap_8 FILLER_11_306 ();
 sg13g2_decap_4 FILLER_11_313 ();
 sg13g2_fill_1 FILLER_11_317 ();
 sg13g2_fill_2 FILLER_11_345 ();
 sg13g2_fill_2 FILLER_11_353 ();
 sg13g2_decap_4 FILLER_11_384 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_9 ();
 sg13g2_decap_4 FILLER_12_106 ();
 sg13g2_fill_2 FILLER_12_110 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_fill_2 FILLER_12_152 ();
 sg13g2_fill_1 FILLER_12_205 ();
 sg13g2_fill_2 FILLER_12_226 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_4 FILLER_12_259 ();
 sg13g2_fill_1 FILLER_12_263 ();
 sg13g2_fill_2 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_fill_2 FILLER_12_328 ();
 sg13g2_fill_1 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_341 ();
 sg13g2_fill_1 FILLER_12_343 ();
 sg13g2_fill_2 FILLER_12_354 ();
 sg13g2_fill_1 FILLER_12_356 ();
 sg13g2_fill_2 FILLER_12_380 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_fill_2 FILLER_13_25 ();
 sg13g2_fill_1 FILLER_13_27 ();
 sg13g2_fill_1 FILLER_13_45 ();
 sg13g2_fill_1 FILLER_13_85 ();
 sg13g2_fill_2 FILLER_13_144 ();
 sg13g2_fill_1 FILLER_13_146 ();
 sg13g2_decap_8 FILLER_13_176 ();
 sg13g2_decap_4 FILLER_13_183 ();
 sg13g2_fill_1 FILLER_13_187 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_fill_2 FILLER_13_209 ();
 sg13g2_fill_1 FILLER_13_211 ();
 sg13g2_fill_2 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_233 ();
 sg13g2_fill_2 FILLER_13_240 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_fill_2 FILLER_13_254 ();
 sg13g2_fill_2 FILLER_13_270 ();
 sg13g2_fill_1 FILLER_13_272 ();
 sg13g2_fill_2 FILLER_13_283 ();
 sg13g2_fill_1 FILLER_13_285 ();
 sg13g2_fill_2 FILLER_13_306 ();
 sg13g2_fill_1 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_343 ();
 sg13g2_fill_1 FILLER_13_360 ();
 sg13g2_decap_4 FILLER_13_381 ();
 sg13g2_fill_1 FILLER_13_385 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_27 ();
 sg13g2_fill_1 FILLER_14_34 ();
 sg13g2_fill_2 FILLER_14_62 ();
 sg13g2_fill_2 FILLER_14_68 ();
 sg13g2_decap_8 FILLER_14_111 ();
 sg13g2_fill_2 FILLER_14_118 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_decap_8 FILLER_14_130 ();
 sg13g2_fill_2 FILLER_14_137 ();
 sg13g2_fill_1 FILLER_14_139 ();
 sg13g2_fill_1 FILLER_14_145 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_175 ();
 sg13g2_decap_4 FILLER_14_203 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_decap_4 FILLER_14_253 ();
 sg13g2_fill_1 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_263 ();
 sg13g2_fill_1 FILLER_14_265 ();
 sg13g2_fill_2 FILLER_14_289 ();
 sg13g2_fill_1 FILLER_14_291 ();
 sg13g2_decap_4 FILLER_14_323 ();
 sg13g2_decap_4 FILLER_14_343 ();
 sg13g2_fill_1 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_364 ();
 sg13g2_fill_1 FILLER_14_397 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_fill_2 FILLER_15_15 ();
 sg13g2_fill_1 FILLER_15_17 ();
 sg13g2_fill_1 FILLER_15_27 ();
 sg13g2_fill_2 FILLER_15_51 ();
 sg13g2_fill_2 FILLER_15_100 ();
 sg13g2_fill_1 FILLER_15_102 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_155 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_178 ();
 sg13g2_decap_4 FILLER_15_188 ();
 sg13g2_fill_2 FILLER_15_204 ();
 sg13g2_fill_1 FILLER_15_206 ();
 sg13g2_fill_1 FILLER_15_220 ();
 sg13g2_fill_2 FILLER_15_230 ();
 sg13g2_fill_1 FILLER_15_237 ();
 sg13g2_decap_4 FILLER_15_251 ();
 sg13g2_fill_2 FILLER_15_288 ();
 sg13g2_decap_4 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_313 ();
 sg13g2_fill_2 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_fill_1 FILLER_15_369 ();
 sg13g2_decap_4 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_fill_1 FILLER_16_33 ();
 sg13g2_fill_2 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_103 ();
 sg13g2_fill_2 FILLER_16_116 ();
 sg13g2_fill_1 FILLER_16_118 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_decap_4 FILLER_16_130 ();
 sg13g2_fill_1 FILLER_16_134 ();
 sg13g2_fill_2 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_153 ();
 sg13g2_decap_4 FILLER_16_178 ();
 sg13g2_decap_4 FILLER_16_202 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_decap_4 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_fill_2 FILLER_16_279 ();
 sg13g2_fill_2 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_fill_2 FILLER_16_345 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_fill_2 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_fill_1 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_10 ();
 sg13g2_fill_2 FILLER_17_16 ();
 sg13g2_fill_2 FILLER_17_78 ();
 sg13g2_fill_1 FILLER_17_80 ();
 sg13g2_fill_1 FILLER_17_99 ();
 sg13g2_fill_2 FILLER_17_141 ();
 sg13g2_fill_1 FILLER_17_143 ();
 sg13g2_fill_2 FILLER_17_159 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_decap_4 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_190 ();
 sg13g2_decap_4 FILLER_17_197 ();
 sg13g2_fill_2 FILLER_17_201 ();
 sg13g2_decap_4 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_211 ();
 sg13g2_fill_2 FILLER_17_221 ();
 sg13g2_decap_4 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_282 ();
 sg13g2_fill_1 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_299 ();
 sg13g2_decap_4 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_decap_4 FILLER_17_353 ();
 sg13g2_fill_1 FILLER_17_357 ();
 sg13g2_decap_4 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_4 FILLER_17_384 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_67 ();
 sg13g2_fill_1 FILLER_18_124 ();
 sg13g2_decap_8 FILLER_18_138 ();
 sg13g2_decap_8 FILLER_18_145 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_decap_8 FILLER_18_180 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_209 ();
 sg13g2_fill_1 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_280 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_fill_1 FILLER_18_306 ();
 sg13g2_decap_4 FILLER_18_342 ();
 sg13g2_fill_2 FILLER_18_351 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_fill_2 FILLER_19_45 ();
 sg13g2_fill_1 FILLER_19_89 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_decap_4 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_169 ();
 sg13g2_decap_4 FILLER_19_183 ();
 sg13g2_decap_4 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_211 ();
 sg13g2_decap_4 FILLER_19_218 ();
 sg13g2_fill_2 FILLER_19_222 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_2 FILLER_19_241 ();
 sg13g2_decap_4 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_decap_4 FILLER_19_281 ();
 sg13g2_fill_2 FILLER_19_290 ();
 sg13g2_decap_4 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_304 ();
 sg13g2_decap_4 FILLER_19_313 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_decap_4 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_353 ();
 sg13g2_fill_1 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_4 FILLER_19_372 ();
 sg13g2_fill_2 FILLER_19_376 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_fill_2 FILLER_20_19 ();
 sg13g2_fill_2 FILLER_20_29 ();
 sg13g2_fill_1 FILLER_20_36 ();
 sg13g2_fill_2 FILLER_20_51 ();
 sg13g2_fill_2 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_decap_4 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_decap_4 FILLER_20_260 ();
 sg13g2_decap_4 FILLER_20_288 ();
 sg13g2_decap_8 FILLER_20_302 ();
 sg13g2_fill_2 FILLER_20_309 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_fill_2 FILLER_20_320 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_decap_4 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_359 ();
 sg13g2_decap_4 FILLER_20_375 ();
 sg13g2_fill_1 FILLER_20_383 ();
 sg13g2_fill_2 FILLER_20_389 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_21_34 ();
 sg13g2_fill_1 FILLER_21_40 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_131 ();
 sg13g2_fill_2 FILLER_21_146 ();
 sg13g2_decap_4 FILLER_21_161 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_4 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_fill_2 FILLER_21_277 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_314 ();
 sg13g2_decap_8 FILLER_21_321 ();
 sg13g2_fill_1 FILLER_21_328 ();
 sg13g2_decap_4 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_fill_2 FILLER_21_381 ();
 sg13g2_fill_1 FILLER_21_383 ();
 sg13g2_fill_2 FILLER_21_390 ();
 sg13g2_fill_1 FILLER_21_392 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_fill_2 FILLER_22_40 ();
 sg13g2_fill_2 FILLER_22_51 ();
 sg13g2_fill_1 FILLER_22_80 ();
 sg13g2_fill_1 FILLER_22_94 ();
 sg13g2_fill_1 FILLER_22_124 ();
 sg13g2_fill_2 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_141 ();
 sg13g2_decap_4 FILLER_22_176 ();
 sg13g2_decap_4 FILLER_22_188 ();
 sg13g2_fill_2 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_fill_1 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_decap_4 FILLER_22_234 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_fill_2 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_256 ();
 sg13g2_fill_2 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_4 FILLER_22_287 ();
 sg13g2_decap_4 FILLER_22_295 ();
 sg13g2_decap_4 FILLER_22_310 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_2 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_173 ();
 sg13g2_decap_8 FILLER_23_180 ();
 sg13g2_decap_4 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_200 ();
 sg13g2_fill_2 FILLER_23_205 ();
 sg13g2_fill_2 FILLER_23_229 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_decap_4 FILLER_23_332 ();
 sg13g2_fill_1 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_364 ();
 sg13g2_fill_1 FILLER_24_67 ();
 sg13g2_fill_1 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_100 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_147 ();
 sg13g2_fill_1 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_176 ();
 sg13g2_fill_2 FILLER_24_205 ();
 sg13g2_decap_4 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_264 ();
 sg13g2_decap_4 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_279 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_decap_4 FILLER_24_293 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_314 ();
 sg13g2_fill_2 FILLER_24_323 ();
 sg13g2_fill_1 FILLER_24_334 ();
 sg13g2_fill_2 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_379 ();
 sg13g2_fill_1 FILLER_24_385 ();
 sg13g2_fill_1 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_fill_2 FILLER_25_241 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_fill_2 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_fill_1 FILLER_25_376 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_388 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_decap_8 FILLER_26_250 ();
 sg13g2_decap_8 FILLER_26_257 ();
 sg13g2_fill_1 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_286 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_308 ();
 sg13g2_decap_4 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_27_38 ();
 sg13g2_fill_1 FILLER_27_115 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_190 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_fill_2 FILLER_27_241 ();
 sg13g2_fill_1 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_fill_2 FILLER_27_384 ();
 sg13g2_fill_1 FILLER_27_386 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_fill_1 FILLER_28_198 ();
 sg13g2_decap_8 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_259 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_fill_2 FILLER_28_361 ();
 sg13g2_fill_1 FILLER_28_363 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_29_34 ();
 sg13g2_fill_2 FILLER_29_90 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_359 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_fill_1 FILLER_29_386 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_27 ();
 sg13g2_fill_2 FILLER_30_38 ();
 sg13g2_fill_2 FILLER_30_64 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_2 FILLER_30_209 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_276 ();
 sg13g2_fill_1 FILLER_30_341 ();
 sg13g2_decap_4 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_71 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_fill_2 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_128 ();
 sg13g2_fill_2 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_342 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_354 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_fill_1 FILLER_31_370 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_fill_2 FILLER_31_383 ();
 sg13g2_fill_1 FILLER_31_385 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_fill_1 FILLER_32_23 ();
 sg13g2_fill_1 FILLER_32_54 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_fill_1 FILLER_32_332 ();
 sg13g2_fill_1 FILLER_32_381 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_27 ();
 sg13g2_fill_1 FILLER_33_76 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_291 ();
 sg13g2_fill_1 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_fill_1 FILLER_35_90 ();
 sg13g2_fill_1 FILLER_35_99 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_2 FILLER_36_44 ();
 sg13g2_fill_1 FILLER_36_97 ();
 sg13g2_fill_2 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_1 FILLER_36_274 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_362 ();
 sg13g2_fill_1 FILLER_36_378 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_81 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_357 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_178 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net104;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
endmodule

module tt_um_rejunity_ternary_dot (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire \i_w_buf[0].A ;
 wire \i_w_buf[100].A ;
 wire \i_w_buf[101].A ;
 wire \i_w_buf[102].A ;
 wire \i_w_buf[103].A ;
 wire \i_w_buf[104].A ;
 wire \i_w_buf[105].A ;
 wire \i_w_buf[106].A ;
 wire \i_w_buf[107].A ;
 wire \i_w_buf[108].A ;
 wire \i_w_buf[109].A ;
 wire \i_w_buf[10].A ;
 wire \i_w_buf[110].A ;
 wire \i_w_buf[111].A ;
 wire \i_w_buf[112].A ;
 wire \i_w_buf[113].A ;
 wire \i_w_buf[114].A ;
 wire \i_w_buf[115].A ;
 wire \i_w_buf[116].A ;
 wire \i_w_buf[117].A ;
 wire \i_w_buf[118].A ;
 wire \i_w_buf[119].A ;
 wire \i_w_buf[11].A ;
 wire \i_w_buf[120].A ;
 wire \i_w_buf[121].A ;
 wire \i_w_buf[122].A ;
 wire \i_w_buf[123].A ;
 wire \i_w_buf[124].A ;
 wire \i_w_buf[125].A ;
 wire \i_w_buf[126].A ;
 wire \i_w_buf[127].A ;
 wire \i_w_buf[128].A ;
 wire \i_w_buf[129].A ;
 wire \i_w_buf[12].A ;
 wire \i_w_buf[130].A ;
 wire \i_w_buf[131].A ;
 wire \i_w_buf[132].A ;
 wire \i_w_buf[133].A ;
 wire \i_w_buf[134].A ;
 wire \i_w_buf[135].A ;
 wire \i_w_buf[136].A ;
 wire \i_w_buf[137].A ;
 wire \i_w_buf[138].A ;
 wire \i_w_buf[139].A ;
 wire \i_w_buf[13].A ;
 wire \i_w_buf[140].A ;
 wire \i_w_buf[141].A ;
 wire \i_w_buf[142].A ;
 wire \i_w_buf[143].A ;
 wire \i_w_buf[144].A ;
 wire \i_w_buf[145].A ;
 wire \i_w_buf[146].A ;
 wire \i_w_buf[147].A ;
 wire \i_w_buf[148].A ;
 wire \i_w_buf[149].A ;
 wire \i_w_buf[14].A ;
 wire \i_w_buf[150].A ;
 wire \i_w_buf[151].A ;
 wire \i_w_buf[152].A ;
 wire \i_w_buf[153].A ;
 wire \i_w_buf[154].A ;
 wire \i_w_buf[155].A ;
 wire \i_w_buf[156].A ;
 wire \i_w_buf[157].A ;
 wire \i_w_buf[158].A ;
 wire \i_w_buf[159].A ;
 wire \i_w_buf[15].A ;
 wire \i_w_buf[160].A ;
 wire \i_w_buf[161].A ;
 wire \i_w_buf[162].A ;
 wire \i_w_buf[163].A ;
 wire \i_w_buf[164].A ;
 wire \i_w_buf[165].A ;
 wire \i_w_buf[166].A ;
 wire \i_w_buf[167].A ;
 wire \i_w_buf[168].A ;
 wire \i_w_buf[169].A ;
 wire \i_w_buf[16].A ;
 wire \i_w_buf[170].A ;
 wire \i_w_buf[171].A ;
 wire \i_w_buf[172].A ;
 wire \i_w_buf[173].A ;
 wire \i_w_buf[174].A ;
 wire \i_w_buf[175].A ;
 wire \i_w_buf[176].A ;
 wire \i_w_buf[177].A ;
 wire \i_w_buf[178].A ;
 wire \i_w_buf[179].A ;
 wire \i_w_buf[17].A ;
 wire \i_w_buf[180].A ;
 wire \i_w_buf[181].A ;
 wire \i_w_buf[182].A ;
 wire \i_w_buf[183].A ;
 wire \i_w_buf[184].A ;
 wire \i_w_buf[185].A ;
 wire \i_w_buf[186].A ;
 wire \i_w_buf[187].A ;
 wire \i_w_buf[188].A ;
 wire \i_w_buf[189].A ;
 wire \i_w_buf[18].A ;
 wire \i_w_buf[190].A ;
 wire \i_w_buf[191].A ;
 wire \i_w_buf[192].A ;
 wire \i_w_buf[193].A ;
 wire \i_w_buf[194].A ;
 wire \i_w_buf[195].A ;
 wire \i_w_buf[196].A ;
 wire \i_w_buf[197].A ;
 wire \i_w_buf[198].A ;
 wire \i_w_buf[199].A ;
 wire \i_w_buf[19].A ;
 wire \i_w_buf[1].A ;
 wire \i_w_buf[200].A ;
 wire \i_w_buf[201].A ;
 wire \i_w_buf[202].A ;
 wire \i_w_buf[203].A ;
 wire \i_w_buf[204].A ;
 wire \i_w_buf[205].A ;
 wire \i_w_buf[206].A ;
 wire \i_w_buf[207].A ;
 wire \i_w_buf[208].A ;
 wire \i_w_buf[209].A ;
 wire \i_w_buf[20].A ;
 wire \i_w_buf[210].A ;
 wire \i_w_buf[211].A ;
 wire \i_w_buf[212].A ;
 wire \i_w_buf[213].A ;
 wire \i_w_buf[214].A ;
 wire \i_w_buf[215].A ;
 wire \i_w_buf[216].A ;
 wire \i_w_buf[217].A ;
 wire \i_w_buf[218].A ;
 wire \i_w_buf[219].A ;
 wire \i_w_buf[21].A ;
 wire \i_w_buf[220].A ;
 wire \i_w_buf[221].A ;
 wire \i_w_buf[222].A ;
 wire \i_w_buf[223].A ;
 wire \i_w_buf[224].A ;
 wire \i_w_buf[225].A ;
 wire \i_w_buf[226].A ;
 wire \i_w_buf[227].A ;
 wire \i_w_buf[228].A ;
 wire \i_w_buf[229].A ;
 wire \i_w_buf[22].A ;
 wire \i_w_buf[230].A ;
 wire \i_w_buf[231].A ;
 wire \i_w_buf[232].A ;
 wire \i_w_buf[233].A ;
 wire \i_w_buf[234].A ;
 wire \i_w_buf[235].A ;
 wire \i_w_buf[236].A ;
 wire \i_w_buf[237].A ;
 wire \i_w_buf[238].A ;
 wire \i_w_buf[239].A ;
 wire \i_w_buf[23].A ;
 wire \i_w_buf[240].A ;
 wire \i_w_buf[241].A ;
 wire \i_w_buf[242].A ;
 wire \i_w_buf[243].A ;
 wire \i_w_buf[244].A ;
 wire \i_w_buf[245].A ;
 wire \i_w_buf[246].A ;
 wire \i_w_buf[247].A ;
 wire \i_w_buf[248].A ;
 wire \i_w_buf[249].A ;
 wire \i_w_buf[24].A ;
 wire \i_w_buf[250].A ;
 wire \i_w_buf[251].A ;
 wire \i_w_buf[252].A ;
 wire \i_w_buf[253].A ;
 wire \i_w_buf[254].A ;
 wire \i_w_buf[255].A ;
 wire \i_w_buf[25].A ;
 wire \i_w_buf[26].A ;
 wire \i_w_buf[27].A ;
 wire \i_w_buf[28].A ;
 wire \i_w_buf[29].A ;
 wire \i_w_buf[2].A ;
 wire \i_w_buf[30].A ;
 wire \i_w_buf[31].A ;
 wire \i_w_buf[32].A ;
 wire \i_w_buf[33].A ;
 wire \i_w_buf[34].A ;
 wire \i_w_buf[35].A ;
 wire \i_w_buf[36].A ;
 wire \i_w_buf[37].A ;
 wire \i_w_buf[38].A ;
 wire \i_w_buf[39].A ;
 wire \i_w_buf[3].A ;
 wire \i_w_buf[40].A ;
 wire \i_w_buf[41].A ;
 wire \i_w_buf[42].A ;
 wire \i_w_buf[43].A ;
 wire \i_w_buf[44].A ;
 wire \i_w_buf[45].A ;
 wire \i_w_buf[46].A ;
 wire \i_w_buf[47].A ;
 wire \i_w_buf[48].A ;
 wire \i_w_buf[49].A ;
 wire \i_w_buf[4].A ;
 wire \i_w_buf[50].A ;
 wire \i_w_buf[51].A ;
 wire \i_w_buf[52].A ;
 wire \i_w_buf[53].A ;
 wire \i_w_buf[54].A ;
 wire \i_w_buf[55].A ;
 wire \i_w_buf[56].A ;
 wire \i_w_buf[57].A ;
 wire \i_w_buf[58].A ;
 wire \i_w_buf[59].A ;
 wire \i_w_buf[5].A ;
 wire \i_w_buf[60].A ;
 wire \i_w_buf[61].A ;
 wire \i_w_buf[62].A ;
 wire \i_w_buf[63].A ;
 wire \i_w_buf[64].A ;
 wire \i_w_buf[65].A ;
 wire \i_w_buf[66].A ;
 wire \i_w_buf[67].A ;
 wire \i_w_buf[68].A ;
 wire \i_w_buf[69].A ;
 wire \i_w_buf[6].A ;
 wire \i_w_buf[70].A ;
 wire \i_w_buf[71].A ;
 wire \i_w_buf[72].A ;
 wire \i_w_buf[73].A ;
 wire \i_w_buf[74].A ;
 wire \i_w_buf[75].A ;
 wire \i_w_buf[76].A ;
 wire \i_w_buf[77].A ;
 wire \i_w_buf[78].A ;
 wire \i_w_buf[79].A ;
 wire \i_w_buf[7].A ;
 wire \i_w_buf[80].A ;
 wire \i_w_buf[81].A ;
 wire \i_w_buf[82].A ;
 wire \i_w_buf[83].A ;
 wire \i_w_buf[84].A ;
 wire \i_w_buf[85].A ;
 wire \i_w_buf[86].A ;
 wire \i_w_buf[87].A ;
 wire \i_w_buf[88].A ;
 wire \i_w_buf[89].A ;
 wire \i_w_buf[8].A ;
 wire \i_w_buf[90].A ;
 wire \i_w_buf[91].A ;
 wire \i_w_buf[92].A ;
 wire \i_w_buf[93].A ;
 wire \i_w_buf[94].A ;
 wire \i_w_buf[95].A ;
 wire \i_w_buf[96].A ;
 wire \i_w_buf[97].A ;
 wire \i_w_buf[98].A ;
 wire \i_w_buf[99].A ;
 wire \i_w_buf[9].A ;
 wire net7;
 wire net8;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire clknet_leaf_0_clk;
 wire net9;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;

 sg13g2_inv_2 _2100_ (.Y(_0862_),
    .A(net101));
 sg13g2_inv_8 _2101_ (.Y(_0863_),
    .A(net96));
 sg13g2_inv_8 _2102_ (.Y(_0864_),
    .A(net103));
 sg13g2_inv_2 _2103_ (.Y(_0865_),
    .A(net91));
 sg13g2_inv_2 _2104_ (.Y(_0866_),
    .A(net106));
 sg13g2_inv_2 _2105_ (.Y(_0867_),
    .A(net93));
 sg13g2_inv_1 _2106_ (.Y(_0868_),
    .A(\i_w_buf[125].A ));
 sg13g2_inv_1 _2107_ (.Y(_0869_),
    .A(net89));
 sg13g2_inv_2 _2108_ (.Y(_0870_),
    .A(net98));
 sg13g2_inv_1 _2109_ (.Y(_0871_),
    .A(\i_w_buf[7].A ));
 sg13g2_inv_1 _2110_ (.Y(_0872_),
    .A(\i_w_buf[159].A ));
 sg13g2_inv_1 _2111_ (.Y(_0873_),
    .A(\i_w_buf[11].A ));
 sg13g2_inv_1 _2112_ (.Y(_0874_),
    .A(\i_w_buf[15].A ));
 sg13g2_inv_1 _2113_ (.Y(_0875_),
    .A(\i_w_buf[27].A ));
 sg13g2_inv_1 _2114_ (.Y(_0876_),
    .A(\i_w_buf[29].A ));
 sg13g2_inv_1 _2115_ (.Y(_0877_),
    .A(\i_w_buf[35].A ));
 sg13g2_inv_1 _2116_ (.Y(_0878_),
    .A(\i_w_buf[37].A ));
 sg13g2_inv_1 _2117_ (.Y(_0879_),
    .A(\i_w_buf[53].A ));
 sg13g2_inv_1 _2118_ (.Y(_0880_),
    .A(\i_w_buf[139].A ));
 sg13g2_inv_1 _2119_ (.Y(_0881_),
    .A(\i_w_buf[57].A ));
 sg13g2_inv_1 _2120_ (.Y(_0882_),
    .A(\i_w_buf[89].A ));
 sg13g2_inv_1 _2121_ (.Y(_0883_),
    .A(\i_w_buf[71].A ));
 sg13g2_inv_1 _2122_ (.Y(_0884_),
    .A(\i_w_buf[75].A ));
 sg13g2_inv_1 _2123_ (.Y(_0885_),
    .A(\i_w_buf[111].A ));
 sg13g2_inv_1 _2124_ (.Y(_0886_),
    .A(\i_w_buf[129].A ));
 sg13g2_inv_1 _2125_ (.Y(_0887_),
    .A(\i_w_buf[9].A ));
 sg13g2_inv_1 _2126_ (.Y(_0888_),
    .A(\i_w_buf[93].A ));
 sg13g2_inv_1 _2127_ (.Y(_0889_),
    .A(\i_w_buf[107].A ));
 sg13g2_inv_1 _2128_ (.Y(_0890_),
    .A(\i_w_buf[143].A ));
 sg13g2_inv_1 _2129_ (.Y(_0891_),
    .A(\i_w_buf[161].A ));
 sg13g2_inv_1 _2130_ (.Y(_0892_),
    .A(\i_w_buf[147].A ));
 sg13g2_inv_1 _2131_ (.Y(_0893_),
    .A(\i_w_buf[165].A ));
 sg13g2_inv_1 _2132_ (.Y(_0894_),
    .A(\i_w_buf[173].A ));
 sg13g2_inv_1 _2133_ (.Y(_0895_),
    .A(\i_w_buf[177].A ));
 sg13g2_nand3b_1 _2134_ (.B(\i_w_buf[81].A ),
    .C(net106),
    .Y(_0896_),
    .A_N(\i_w_buf[80].A ));
 sg13g2_nand3b_1 _2135_ (.B(\i_w_buf[69].A ),
    .C(net100),
    .Y(_0897_),
    .A_N(\i_w_buf[68].A ));
 sg13g2_nor2b_1 _2136_ (.A(\i_w_buf[2].A ),
    .B_N(net105),
    .Y(_0898_));
 sg13g2_nand2_1 _2137_ (.Y(_0899_),
    .A(\i_w_buf[3].A ),
    .B(_0898_));
 sg13g2_nor2b_1 _2138_ (.A(\i_w_buf[136].A ),
    .B_N(net96),
    .Y(_0900_));
 sg13g2_nand2_2 _2139_ (.Y(_0901_),
    .A(\i_w_buf[137].A ),
    .B(_0900_));
 sg13g2_nor2b_1 _2140_ (.A(\i_w_buf[34].A ),
    .B_N(net105),
    .Y(_0902_));
 sg13g2_nand2_1 _2141_ (.Y(_0903_),
    .A(\i_w_buf[35].A ),
    .B(_0902_));
 sg13g2_nand3b_1 _2142_ (.B(\i_w_buf[141].A ),
    .C(net92),
    .Y(_0904_),
    .A_N(\i_w_buf[140].A ));
 sg13g2_inv_1 _2143_ (.Y(_0905_),
    .A(_0904_));
 sg13g2_nor2_1 _2144_ (.A(net82),
    .B(\i_w_buf[30].A ),
    .Y(_0906_));
 sg13g2_nand2b_1 _2145_ (.Y(_0907_),
    .B(_0906_),
    .A_N(\i_w_buf[31].A ));
 sg13g2_nor2_1 _2146_ (.A(net87),
    .B(\i_w_buf[12].A ),
    .Y(_0908_));
 sg13g2_nand2b_1 _2147_ (.Y(_0909_),
    .B(net92),
    .A_N(\i_w_buf[12].A ));
 sg13g2_nand2_1 _2148_ (.Y(_0910_),
    .A(\i_w_buf[31].A ),
    .B(_0906_));
 sg13g2_nor2_1 _2149_ (.A(_0865_),
    .B(\i_w_buf[60].A ),
    .Y(_0911_));
 sg13g2_nor3_2 _2150_ (.A(net87),
    .B(\i_w_buf[60].A ),
    .C(\i_w_buf[61].A ),
    .Y(_0912_));
 sg13g2_nor2b_1 _2151_ (.A(\i_w_buf[98].A ),
    .B_N(net104),
    .Y(_0913_));
 sg13g2_nor2b_2 _2152_ (.A(\i_w_buf[99].A ),
    .B_N(_0913_),
    .Y(_0914_));
 sg13g2_nor2b_1 _2153_ (.A(\i_w_buf[156].A ),
    .B_N(net3),
    .Y(_0915_));
 sg13g2_nand2b_1 _2154_ (.Y(_0916_),
    .B(_0915_),
    .A_N(\i_w_buf[157].A ));
 sg13g2_nor2_1 _2155_ (.A(net82),
    .B(\i_w_buf[46].A ),
    .Y(_0917_));
 sg13g2_nand2_2 _2156_ (.Y(_0918_),
    .A(\i_w_buf[47].A ),
    .B(_0917_));
 sg13g2_nor2_1 _2157_ (.A(_0870_),
    .B(\i_w_buf[246].A ),
    .Y(_0919_));
 sg13g2_nor3_1 _2158_ (.A(net80),
    .B(\i_w_buf[246].A ),
    .C(\i_w_buf[247].A ),
    .Y(_0920_));
 sg13g2_nor3_2 _2159_ (.A(net85),
    .B(\i_w_buf[240].A ),
    .C(\i_w_buf[241].A ),
    .Y(_0921_));
 sg13g2_nor2b_1 _2160_ (.A(\i_w_buf[176].A ),
    .B_N(net106),
    .Y(_0922_));
 sg13g2_nand2_1 _2161_ (.Y(_0923_),
    .A(\i_w_buf[177].A ),
    .B(_0922_));
 sg13g2_and2_1 _2162_ (.A(_0921_),
    .B(_0923_),
    .X(_0924_));
 sg13g2_xor2_1 _2163_ (.B(_0923_),
    .A(_0921_),
    .X(_0925_));
 sg13g2_xnor2_1 _2164_ (.Y(_0926_),
    .A(_0920_),
    .B(_0925_));
 sg13g2_nand2b_1 _2165_ (.Y(_0927_),
    .B(_0918_),
    .A_N(_0926_));
 sg13g2_xor2_1 _2166_ (.B(_0926_),
    .A(_0918_),
    .X(_0928_));
 sg13g2_xor2_1 _2167_ (.B(_0928_),
    .A(_0916_),
    .X(_0929_));
 sg13g2_nand2_1 _2168_ (.Y(_0930_),
    .A(_0914_),
    .B(_0929_));
 sg13g2_xnor2_1 _2169_ (.Y(_0931_),
    .A(_0914_),
    .B(_0929_));
 sg13g2_nor2_1 _2170_ (.A(net82),
    .B(\i_w_buf[254].A ),
    .Y(_0932_));
 sg13g2_nor3_1 _2171_ (.A(net82),
    .B(\i_w_buf[254].A ),
    .C(\i_w_buf[255].A ),
    .Y(_0933_));
 sg13g2_nor3_1 _2172_ (.A(_0863_),
    .B(\i_w_buf[248].A ),
    .C(\i_w_buf[249].A ),
    .Y(_0934_));
 sg13g2_nor2b_1 _2173_ (.A(\i_w_buf[164].A ),
    .B_N(net100),
    .Y(_0935_));
 sg13g2_nand2_2 _2174_ (.Y(_0936_),
    .A(\i_w_buf[165].A ),
    .B(_0935_));
 sg13g2_and2_1 _2175_ (.A(_0934_),
    .B(_0936_),
    .X(_0937_));
 sg13g2_xor2_1 _2176_ (.B(_0936_),
    .A(_0934_),
    .X(_0938_));
 sg13g2_xnor2_1 _2177_ (.Y(_0939_),
    .A(_0933_),
    .B(_0938_));
 sg13g2_xor2_1 _2178_ (.B(_0939_),
    .A(_0931_),
    .X(_0940_));
 sg13g2_xnor2_1 _2179_ (.Y(_0941_),
    .A(_0912_),
    .B(_0940_));
 sg13g2_nor2b_1 _2180_ (.A(_0941_),
    .B_N(_0910_),
    .Y(_0942_));
 sg13g2_xor2_1 _2181_ (.B(_0941_),
    .A(_0910_),
    .X(_0943_));
 sg13g2_nor3_1 _2182_ (.A(\i_w_buf[13].A ),
    .B(_0909_),
    .C(_0943_),
    .Y(_0944_));
 sg13g2_o21ai_1 _2183_ (.B1(_0943_),
    .Y(_0945_),
    .A1(\i_w_buf[13].A ),
    .A2(_0909_));
 sg13g2_nand2b_1 _2184_ (.Y(_0946_),
    .B(_0945_),
    .A_N(_0944_));
 sg13g2_nor2_1 _2185_ (.A(_0907_),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_xnor2_1 _2186_ (.Y(_0948_),
    .A(_0907_),
    .B(_0946_));
 sg13g2_xnor2_1 _2187_ (.Y(_0949_),
    .A(_0905_),
    .B(_0948_));
 sg13g2_nand2b_1 _2188_ (.Y(_0950_),
    .B(_0903_),
    .A_N(_0949_));
 sg13g2_xor2_1 _2189_ (.B(_0949_),
    .A(_0903_),
    .X(_0951_));
 sg13g2_nor2b_1 _2190_ (.A(_0951_),
    .B_N(_0901_),
    .Y(_0952_));
 sg13g2_xor2_1 _2191_ (.B(_0951_),
    .A(_0901_),
    .X(_0953_));
 sg13g2_nor2b_1 _2192_ (.A(_0953_),
    .B_N(_0899_),
    .Y(_0954_));
 sg13g2_xor2_1 _2193_ (.B(_0953_),
    .A(_0899_),
    .X(_0955_));
 sg13g2_nand3b_1 _2194_ (.B(\i_w_buf[131].A ),
    .C(net104),
    .Y(_0956_),
    .A_N(\i_w_buf[130].A ));
 sg13g2_nand2b_1 _2195_ (.Y(_0957_),
    .B(net2),
    .A_N(\i_w_buf[8].A ));
 sg13g2_nor2_1 _2196_ (.A(_0887_),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_nand3b_1 _2197_ (.B(\i_w_buf[33].A ),
    .C(net106),
    .Y(_0959_),
    .A_N(\i_w_buf[32].A ));
 sg13g2_nand2b_1 _2198_ (.Y(_0960_),
    .B(net102),
    .A_N(\i_w_buf[4].A ));
 sg13g2_nor2_1 _2199_ (.A(\i_w_buf[5].A ),
    .B(_0960_),
    .Y(_0961_));
 sg13g2_nor3_2 _2200_ (.A(net86),
    .B(\i_w_buf[16].A ),
    .C(\i_w_buf[17].A ),
    .Y(_0962_));
 sg13g2_nand3b_1 _2201_ (.B(\i_w_buf[117].A ),
    .C(net101),
    .Y(_0963_),
    .A_N(\i_w_buf[116].A ));
 sg13g2_nor3_2 _2202_ (.A(net83),
    .B(\i_w_buf[138].A ),
    .C(_0880_),
    .Y(_0964_));
 sg13g2_nor3_2 _2203_ (.A(net87),
    .B(\i_w_buf[44].A ),
    .C(\i_w_buf[45].A ),
    .Y(_0965_));
 sg13g2_or3_2 _2204_ (.A(net85),
    .B(\i_w_buf[112].A ),
    .C(\i_w_buf[113].A ),
    .X(_0966_));
 sg13g2_nand3b_1 _2205_ (.B(\i_w_buf[189].A ),
    .C(net91),
    .Y(_0967_),
    .A_N(\i_w_buf[188].A ));
 sg13g2_nor2_2 _2206_ (.A(_0865_),
    .B(\i_w_buf[172].A ),
    .Y(_0968_));
 sg13g2_nand2b_1 _2207_ (.Y(_0969_),
    .B(net93),
    .A_N(\i_w_buf[170].A ));
 sg13g2_nand3b_1 _2208_ (.B(\i_w_buf[171].A ),
    .C(net93),
    .Y(_0970_),
    .A_N(\i_w_buf[170].A ));
 sg13g2_xnor2_1 _2209_ (.Y(_0971_),
    .A(_0968_),
    .B(_0970_));
 sg13g2_xor2_1 _2210_ (.B(_0970_),
    .A(_0968_),
    .X(_0972_));
 sg13g2_nor3_2 _2211_ (.A(_0864_),
    .B(\i_w_buf[178].A ),
    .C(\i_w_buf[179].A ),
    .Y(_0973_));
 sg13g2_nor2b_1 _2212_ (.A(\i_w_buf[168].A ),
    .B_N(net97),
    .Y(_0974_));
 sg13g2_nor2b_1 _2213_ (.A(\i_w_buf[169].A ),
    .B_N(_0974_),
    .Y(_0975_));
 sg13g2_nand3b_1 _2214_ (.B(\i_w_buf[179].A ),
    .C(net105),
    .Y(_0976_),
    .A_N(\i_w_buf[178].A ));
 sg13g2_nand3_1 _2215_ (.B(_0935_),
    .C(_0976_),
    .A(_0893_),
    .Y(_0977_));
 sg13g2_a21o_1 _2216_ (.A2(_0935_),
    .A1(_0893_),
    .B1(_0976_),
    .X(_0978_));
 sg13g2_nand3_1 _2217_ (.B(_0977_),
    .C(_0978_),
    .A(_0975_),
    .Y(_0979_));
 sg13g2_a21o_1 _2218_ (.A2(_0978_),
    .A1(_0977_),
    .B1(_0975_),
    .X(_0980_));
 sg13g2_and3_1 _2219_ (.X(_0981_),
    .A(_0973_),
    .B(_0979_),
    .C(_0980_));
 sg13g2_nand3_1 _2220_ (.B(_0979_),
    .C(_0980_),
    .A(_0973_),
    .Y(_0982_));
 sg13g2_a21oi_1 _2221_ (.A1(_0979_),
    .A2(_0980_),
    .Y(_0983_),
    .B1(_0973_));
 sg13g2_a21o_1 _2222_ (.A2(_0980_),
    .A1(_0979_),
    .B1(_0973_),
    .X(_0984_));
 sg13g2_nor3_1 _2223_ (.A(_0972_),
    .B(_0981_),
    .C(_0983_),
    .Y(_0985_));
 sg13g2_nand3_1 _2224_ (.B(_0982_),
    .C(_0984_),
    .A(_0971_),
    .Y(_0986_));
 sg13g2_a21oi_1 _2225_ (.A1(_0982_),
    .A2(_0984_),
    .Y(_0987_),
    .B1(_0971_));
 sg13g2_o21ai_1 _2226_ (.B1(_0972_),
    .Y(_0988_),
    .A1(_0981_),
    .A2(_0983_));
 sg13g2_nand3_1 _2227_ (.B(_0986_),
    .C(_0988_),
    .A(_0967_),
    .Y(_0989_));
 sg13g2_a21oi_1 _2228_ (.A1(_0986_),
    .A2(_0988_),
    .Y(_0990_),
    .B1(_0967_));
 sg13g2_nor3_1 _2229_ (.A(_0967_),
    .B(_0985_),
    .C(_0987_),
    .Y(_0991_));
 sg13g2_o21ai_1 _2230_ (.B1(_0967_),
    .Y(_0992_),
    .A1(_0985_),
    .A2(_0987_));
 sg13g2_nor2b_1 _2231_ (.A(_0991_),
    .B_N(_0992_),
    .Y(_0993_));
 sg13g2_xnor2_1 _2232_ (.Y(_0994_),
    .A(_0966_),
    .B(_0993_));
 sg13g2_nor3_2 _2233_ (.A(_0863_),
    .B(\i_w_buf[72].A ),
    .C(\i_w_buf[73].A ),
    .Y(_0995_));
 sg13g2_nor2b_1 _2234_ (.A(\i_w_buf[180].A ),
    .B_N(net100),
    .Y(_0996_));
 sg13g2_nand2b_1 _2235_ (.Y(_0997_),
    .B(_0996_),
    .A_N(\i_w_buf[181].A ));
 sg13g2_nor2b_1 _2236_ (.A(\i_w_buf[92].A ),
    .B_N(net92),
    .Y(_0998_));
 sg13g2_nand2_2 _2237_ (.Y(_0999_),
    .A(\i_w_buf[93].A ),
    .B(_0998_));
 sg13g2_and2_1 _2238_ (.A(\i_w_buf[181].A ),
    .B(_0996_),
    .X(_1000_));
 sg13g2_nor2b_1 _2239_ (.A(\i_w_buf[158].A ),
    .B_N(net90),
    .Y(_1001_));
 sg13g2_nor2b_2 _2240_ (.A(\i_w_buf[160].A ),
    .B_N(net106),
    .Y(_1002_));
 sg13g2_and4_2 _2241_ (.A(_0872_),
    .B(_0891_),
    .C(_1001_),
    .D(_1002_),
    .X(_1003_));
 sg13g2_a22oi_1 _2242_ (.Y(_1004_),
    .B1(_1002_),
    .B2(_0891_),
    .A2(_1001_),
    .A1(_0872_));
 sg13g2_or3_1 _2243_ (.A(_1000_),
    .B(_1003_),
    .C(_1004_),
    .X(_1005_));
 sg13g2_o21ai_1 _2244_ (.B1(_1000_),
    .Y(_1006_),
    .A1(_1003_),
    .A2(_1004_));
 sg13g2_nand3_1 _2245_ (.B(_1005_),
    .C(_1006_),
    .A(_0999_),
    .Y(_1007_));
 sg13g2_a21oi_1 _2246_ (.A1(_1005_),
    .A2(_1006_),
    .Y(_1008_),
    .B1(_0999_));
 sg13g2_a21o_1 _2247_ (.A2(_1006_),
    .A1(_1005_),
    .B1(_0999_),
    .X(_1009_));
 sg13g2_nand2_1 _2248_ (.Y(_1010_),
    .A(_1007_),
    .B(_1009_));
 sg13g2_xnor2_1 _2249_ (.Y(_1011_),
    .A(_0997_),
    .B(_1010_));
 sg13g2_nor3_2 _2250_ (.A(net88),
    .B(\i_w_buf[116].A ),
    .C(\i_w_buf[117].A ),
    .Y(_1012_));
 sg13g2_nand3b_1 _2251_ (.B(\i_w_buf[199].A ),
    .C(net98),
    .Y(_1013_),
    .A_N(\i_w_buf[198].A ));
 sg13g2_nand3b_1 _2252_ (.B(\i_w_buf[203].A ),
    .C(net93),
    .Y(_1014_),
    .A_N(\i_w_buf[202].A ));
 sg13g2_nor3_2 _2253_ (.A(net84),
    .B(\i_w_buf[154].A ),
    .C(\i_w_buf[155].A ),
    .Y(_1015_));
 sg13g2_nand2_1 _2254_ (.Y(_1016_),
    .A(_1014_),
    .B(_1015_));
 sg13g2_xnor2_1 _2255_ (.Y(_1017_),
    .A(_1014_),
    .B(_1015_));
 sg13g2_nand2b_1 _2256_ (.Y(_1018_),
    .B(_1013_),
    .A_N(_1017_));
 sg13g2_xor2_1 _2257_ (.B(_1017_),
    .A(_1013_),
    .X(_1019_));
 sg13g2_nor2_1 _2258_ (.A(_0863_),
    .B(\i_w_buf[184].A ),
    .Y(_1020_));
 sg13g2_nor3_2 _2259_ (.A(_0863_),
    .B(\i_w_buf[184].A ),
    .C(\i_w_buf[185].A ),
    .Y(_1021_));
 sg13g2_nor2b_1 _2260_ (.A(\i_w_buf[150].A ),
    .B_N(net99),
    .Y(_1022_));
 sg13g2_nor2b_1 _2261_ (.A(\i_w_buf[151].A ),
    .B_N(_1022_),
    .Y(_1023_));
 sg13g2_nor2b_2 _2262_ (.A(\i_w_buf[146].A ),
    .B_N(net103),
    .Y(_1024_));
 sg13g2_nand3b_1 _2263_ (.B(\i_w_buf[205].A ),
    .C(net91),
    .Y(_1025_),
    .A_N(\i_w_buf[204].A ));
 sg13g2_nand3_1 _2264_ (.B(_1024_),
    .C(_1025_),
    .A(_0892_),
    .Y(_1026_));
 sg13g2_a21o_1 _2265_ (.A2(_1024_),
    .A1(_0892_),
    .B1(_1025_),
    .X(_1027_));
 sg13g2_nand3_1 _2266_ (.B(_1026_),
    .C(_1027_),
    .A(_1023_),
    .Y(_1028_));
 sg13g2_a21o_1 _2267_ (.A2(_1027_),
    .A1(_1026_),
    .B1(_1023_),
    .X(_1029_));
 sg13g2_and3_1 _2268_ (.X(_1030_),
    .A(_1021_),
    .B(_1028_),
    .C(_1029_));
 sg13g2_nand3_1 _2269_ (.B(_1028_),
    .C(_1029_),
    .A(_1021_),
    .Y(_1031_));
 sg13g2_a21oi_1 _2270_ (.A1(_1028_),
    .A2(_1029_),
    .Y(_1032_),
    .B1(_1021_));
 sg13g2_or3_1 _2271_ (.A(_1019_),
    .B(_1030_),
    .C(_1032_),
    .X(_1033_));
 sg13g2_o21ai_1 _2272_ (.B1(_1019_),
    .Y(_1034_),
    .A1(_1030_),
    .A2(_1032_));
 sg13g2_and3_1 _2273_ (.X(_1035_),
    .A(_1012_),
    .B(_1033_),
    .C(_1034_));
 sg13g2_nand3_1 _2274_ (.B(_1033_),
    .C(_1034_),
    .A(_1012_),
    .Y(_1036_));
 sg13g2_a21oi_1 _2275_ (.A1(_1033_),
    .A2(_1034_),
    .Y(_1037_),
    .B1(_1012_));
 sg13g2_nor2_1 _2276_ (.A(_1035_),
    .B(_1037_),
    .Y(_1038_));
 sg13g2_xnor2_1 _2277_ (.Y(_1039_),
    .A(_1011_),
    .B(_1038_));
 sg13g2_nand2_1 _2278_ (.Y(_1040_),
    .A(_0995_),
    .B(_1039_));
 sg13g2_xnor2_1 _2279_ (.Y(_1041_),
    .A(_0995_),
    .B(_1039_));
 sg13g2_xor2_1 _2280_ (.B(_1041_),
    .A(_0994_),
    .X(_1042_));
 sg13g2_nand2_1 _2281_ (.Y(_1043_),
    .A(_0965_),
    .B(_1042_));
 sg13g2_xnor2_1 _2282_ (.Y(_1044_),
    .A(_0965_),
    .B(_1042_));
 sg13g2_xnor2_1 _2283_ (.Y(_1045_),
    .A(_0964_),
    .B(_1044_));
 sg13g2_nor2b_1 _2284_ (.A(_1045_),
    .B_N(_0963_),
    .Y(_1046_));
 sg13g2_nand2b_1 _2285_ (.Y(_1047_),
    .B(_1045_),
    .A_N(_0963_));
 sg13g2_xnor2_1 _2286_ (.Y(_1048_),
    .A(_0963_),
    .B(_1045_));
 sg13g2_xnor2_1 _2287_ (.Y(_1049_),
    .A(_0962_),
    .B(_1048_));
 sg13g2_nor3_1 _2288_ (.A(\i_w_buf[5].A ),
    .B(_0960_),
    .C(_1049_),
    .Y(_1050_));
 sg13g2_xor2_1 _2289_ (.B(_1049_),
    .A(_0961_),
    .X(_1051_));
 sg13g2_nor3_2 _2290_ (.A(net86),
    .B(\i_w_buf[32].A ),
    .C(\i_w_buf[33].A ),
    .Y(_1052_));
 sg13g2_nand2_2 _2291_ (.Y(_1053_),
    .A(\i_w_buf[147].A ),
    .B(_1024_));
 sg13g2_nor2_1 _2292_ (.A(net81),
    .B(\i_w_buf[238].A ),
    .Y(_1054_));
 sg13g2_nand2_1 _2293_ (.Y(_1055_),
    .A(\i_w_buf[239].A ),
    .B(_1054_));
 sg13g2_nand2b_1 _2294_ (.Y(_1056_),
    .B(net1),
    .A_N(\i_w_buf[64].A ));
 sg13g2_nor2_1 _2295_ (.A(\i_w_buf[65].A ),
    .B(_1056_),
    .Y(_1057_));
 sg13g2_nor3_1 _2296_ (.A(net88),
    .B(\i_w_buf[100].A ),
    .C(\i_w_buf[101].A ),
    .Y(_1058_));
 sg13g2_nor2_1 _2297_ (.A(net82),
    .B(\i_w_buf[174].A ),
    .Y(_1059_));
 sg13g2_nand2_2 _2298_ (.Y(_1060_),
    .A(\i_w_buf[175].A ),
    .B(_1059_));
 sg13g2_nand2b_1 _2299_ (.Y(_1061_),
    .B(_1054_),
    .A_N(\i_w_buf[239].A ));
 sg13g2_nand3b_1 _2300_ (.B(\i_w_buf[201].A ),
    .C(net96),
    .Y(_1062_),
    .A_N(\i_w_buf[200].A ));
 sg13g2_nor3_2 _2301_ (.A(net87),
    .B(\i_w_buf[236].A ),
    .C(\i_w_buf[237].A ),
    .Y(_1063_));
 sg13g2_nand2_1 _2302_ (.Y(_1064_),
    .A(_1062_),
    .B(_1063_));
 sg13g2_xnor2_1 _2303_ (.Y(_1065_),
    .A(_1062_),
    .B(_1063_));
 sg13g2_xnor2_1 _2304_ (.Y(_1066_),
    .A(_1061_),
    .B(_1065_));
 sg13g2_nor2_2 _2305_ (.A(net80),
    .B(\i_w_buf[54].A ),
    .Y(_1067_));
 sg13g2_nand2_2 _2306_ (.Y(_1068_),
    .A(\i_w_buf[55].A ),
    .B(_1067_));
 sg13g2_nor2_1 _2307_ (.A(net80),
    .B(\i_w_buf[230].A ),
    .Y(_1069_));
 sg13g2_nand2b_1 _2308_ (.Y(_1070_),
    .B(_1069_),
    .A_N(\i_w_buf[231].A ));
 sg13g2_nor2_1 _2309_ (.A(net85),
    .B(\i_w_buf[224].A ),
    .Y(_1071_));
 sg13g2_nand2_1 _2310_ (.Y(_1072_),
    .A(\i_w_buf[225].A ),
    .B(_1071_));
 sg13g2_nor3_1 _2311_ (.A(net88),
    .B(\i_w_buf[228].A ),
    .C(\i_w_buf[229].A ),
    .Y(_1073_));
 sg13g2_nand2_1 _2312_ (.Y(_1074_),
    .A(_1072_),
    .B(_1073_));
 sg13g2_xnor2_1 _2313_ (.Y(_1075_),
    .A(_1072_),
    .B(_1073_));
 sg13g2_xor2_1 _2314_ (.B(_1075_),
    .A(_1070_),
    .X(_1076_));
 sg13g2_nand2_1 _2315_ (.Y(_1077_),
    .A(_1068_),
    .B(_1076_));
 sg13g2_xnor2_1 _2316_ (.Y(_1078_),
    .A(_1068_),
    .B(_1076_));
 sg13g2_xor2_1 _2317_ (.B(_1078_),
    .A(_1066_),
    .X(_1079_));
 sg13g2_xnor2_1 _2318_ (.Y(_1080_),
    .A(_1060_),
    .B(_1079_));
 sg13g2_nor4_1 _2319_ (.A(net88),
    .B(\i_w_buf[100].A ),
    .C(\i_w_buf[101].A ),
    .D(_1080_),
    .Y(_1081_));
 sg13g2_xor2_1 _2320_ (.B(_1080_),
    .A(_1058_),
    .X(_1082_));
 sg13g2_nor3_1 _2321_ (.A(\i_w_buf[65].A ),
    .B(_1056_),
    .C(_1082_),
    .Y(_1083_));
 sg13g2_xor2_1 _2322_ (.B(_1082_),
    .A(_1057_),
    .X(_1084_));
 sg13g2_nand2b_1 _2323_ (.Y(_1085_),
    .B(_1055_),
    .A_N(_1084_));
 sg13g2_xor2_1 _2324_ (.B(_1084_),
    .A(_1055_),
    .X(_1086_));
 sg13g2_nor2b_1 _2325_ (.A(_1086_),
    .B_N(_1053_),
    .Y(_1087_));
 sg13g2_nand2b_1 _2326_ (.Y(_1088_),
    .B(_1086_),
    .A_N(_1053_));
 sg13g2_nor2b_1 _2327_ (.A(_1087_),
    .B_N(_1088_),
    .Y(_1089_));
 sg13g2_xnor2_1 _2328_ (.Y(_1090_),
    .A(_1052_),
    .B(_1089_));
 sg13g2_nand2_1 _2329_ (.Y(_1091_),
    .A(\i_w_buf[185].A ),
    .B(_1020_));
 sg13g2_nand2b_1 _2330_ (.Y(_1092_),
    .B(net103),
    .A_N(\i_w_buf[162].A ));
 sg13g2_nand3b_1 _2331_ (.B(\i_w_buf[59].A ),
    .C(net93),
    .Y(_1093_),
    .A_N(\i_w_buf[58].A ));
 sg13g2_nand2b_1 _2332_ (.Y(_1094_),
    .B(net89),
    .A_N(\i_w_buf[222].A ));
 sg13g2_nor2_1 _2333_ (.A(\i_w_buf[223].A ),
    .B(_1094_),
    .Y(_1095_));
 sg13g2_nor3_2 _2334_ (.A(_0863_),
    .B(\i_w_buf[216].A ),
    .C(\i_w_buf[217].A ),
    .Y(_1096_));
 sg13g2_nor3_2 _2335_ (.A(net87),
    .B(\i_w_buf[220].A ),
    .C(\i_w_buf[221].A ),
    .Y(_1097_));
 sg13g2_xnor2_1 _2336_ (.Y(_1098_),
    .A(_1096_),
    .B(_1097_));
 sg13g2_nor3_1 _2337_ (.A(\i_w_buf[223].A ),
    .B(_1094_),
    .C(_1098_),
    .Y(_1099_));
 sg13g2_xor2_1 _2338_ (.B(_1098_),
    .A(_1095_),
    .X(_1100_));
 sg13g2_nor2b_1 _2339_ (.A(_1100_),
    .B_N(_1093_),
    .Y(_1101_));
 sg13g2_xor2_1 _2340_ (.B(_1100_),
    .A(_1093_),
    .X(_1102_));
 sg13g2_nor3_1 _2341_ (.A(\i_w_buf[163].A ),
    .B(_1092_),
    .C(_1102_),
    .Y(_1103_));
 sg13g2_o21ai_1 _2342_ (.B1(_1102_),
    .Y(_1104_),
    .A1(\i_w_buf[163].A ),
    .A2(_1092_));
 sg13g2_nand2b_1 _2343_ (.Y(_1105_),
    .B(_1104_),
    .A_N(_1103_));
 sg13g2_nor2b_1 _2344_ (.A(\i_w_buf[104].A ),
    .B_N(net96),
    .Y(_1106_));
 sg13g2_nor2b_2 _2345_ (.A(\i_w_buf[105].A ),
    .B_N(_1106_),
    .Y(_1107_));
 sg13g2_nor2_1 _2346_ (.A(net80),
    .B(\i_w_buf[214].A ),
    .Y(_1108_));
 sg13g2_nand2b_1 _2347_ (.Y(_1109_),
    .B(net98),
    .A_N(\i_w_buf[214].A ));
 sg13g2_nor3_1 _2348_ (.A(net85),
    .B(\i_w_buf[208].A ),
    .C(\i_w_buf[209].A ),
    .Y(_1110_));
 sg13g2_nand3b_1 _2349_ (.B(\i_w_buf[19].A ),
    .C(net104),
    .Y(_1111_),
    .A_N(\i_w_buf[18].A ));
 sg13g2_xnor2_1 _2350_ (.Y(_1112_),
    .A(_1110_),
    .B(_1111_));
 sg13g2_nor3_1 _2351_ (.A(\i_w_buf[215].A ),
    .B(_1109_),
    .C(_1112_),
    .Y(_1113_));
 sg13g2_o21ai_1 _2352_ (.B1(_1112_),
    .Y(_1114_),
    .A1(\i_w_buf[215].A ),
    .A2(_1109_));
 sg13g2_nand2b_1 _2353_ (.Y(_1115_),
    .B(_1114_),
    .A_N(_1113_));
 sg13g2_nand2b_1 _2354_ (.Y(_1116_),
    .B(net98),
    .A_N(\i_w_buf[166].A ));
 sg13g2_nor2_1 _2355_ (.A(\i_w_buf[167].A ),
    .B(_1116_),
    .Y(_1117_));
 sg13g2_nor2_1 _2356_ (.A(net81),
    .B(\i_w_buf[206].A ),
    .Y(_1118_));
 sg13g2_nor3_2 _2357_ (.A(net81),
    .B(\i_w_buf[206].A ),
    .C(\i_w_buf[207].A ),
    .Y(_1119_));
 sg13g2_nor3_1 _2358_ (.A(_0863_),
    .B(\i_w_buf[200].A ),
    .C(\i_w_buf[201].A ),
    .Y(_1120_));
 sg13g2_nor2b_1 _2359_ (.A(\i_w_buf[24].A ),
    .B_N(net97),
    .Y(_1121_));
 sg13g2_nand2_2 _2360_ (.Y(_1122_),
    .A(\i_w_buf[25].A ),
    .B(_1121_));
 sg13g2_and2_1 _2361_ (.A(_1120_),
    .B(_1122_),
    .X(_1123_));
 sg13g2_xor2_1 _2362_ (.B(_1122_),
    .A(_1120_),
    .X(_1124_));
 sg13g2_xnor2_1 _2363_ (.Y(_1125_),
    .A(_1119_),
    .B(_1124_));
 sg13g2_or3_1 _2364_ (.A(\i_w_buf[167].A ),
    .B(_1116_),
    .C(_1125_),
    .X(_1126_));
 sg13g2_xor2_1 _2365_ (.B(_1125_),
    .A(_1117_),
    .X(_1127_));
 sg13g2_xor2_1 _2366_ (.B(_1127_),
    .A(_1115_),
    .X(_1128_));
 sg13g2_nand2_1 _2367_ (.Y(_1129_),
    .A(_1107_),
    .B(_1128_));
 sg13g2_xnor2_1 _2368_ (.Y(_1130_),
    .A(_1107_),
    .B(_1128_));
 sg13g2_xor2_1 _2369_ (.B(_1130_),
    .A(_1105_),
    .X(_1131_));
 sg13g2_inv_1 _2370_ (.Y(_1132_),
    .A(_1131_));
 sg13g2_nand2_1 _2371_ (.Y(_1133_),
    .A(\i_w_buf[247].A ),
    .B(_0919_));
 sg13g2_nor2b_1 _2372_ (.A(\i_w_buf[182].A ),
    .B_N(net99),
    .Y(_1134_));
 sg13g2_and2_1 _2373_ (.A(\i_w_buf[183].A ),
    .B(_1134_),
    .X(_1135_));
 sg13g2_nand2b_2 _2374_ (.Y(_1136_),
    .B(net91),
    .A_N(\i_w_buf[108].A ));
 sg13g2_nor2_1 _2375_ (.A(\i_w_buf[109].A ),
    .B(_1136_),
    .Y(_1137_));
 sg13g2_nand2_1 _2376_ (.Y(_1138_),
    .A(\i_w_buf[61].A ),
    .B(_0911_));
 sg13g2_nor2_1 _2377_ (.A(\i_w_buf[171].A ),
    .B(_0969_),
    .Y(_1139_));
 sg13g2_nor3_1 _2378_ (.A(net80),
    .B(\i_w_buf[198].A ),
    .C(\i_w_buf[199].A ),
    .Y(_1140_));
 sg13g2_nor2b_1 _2379_ (.A(\i_w_buf[194].A ),
    .B_N(net103),
    .Y(_1141_));
 sg13g2_nor2b_1 _2380_ (.A(\i_w_buf[195].A ),
    .B_N(_1141_),
    .Y(_1142_));
 sg13g2_nor2b_1 _2381_ (.A(\i_w_buf[120].A ),
    .B_N(net97),
    .Y(_1143_));
 sg13g2_nand2_2 _2382_ (.Y(_1144_),
    .A(\i_w_buf[121].A ),
    .B(_1143_));
 sg13g2_and2_1 _2383_ (.A(_1142_),
    .B(_1144_),
    .X(_1145_));
 sg13g2_xor2_1 _2384_ (.B(_1144_),
    .A(_1142_),
    .X(_1146_));
 sg13g2_xnor2_1 _2385_ (.Y(_1147_),
    .A(_1140_),
    .B(_1146_));
 sg13g2_nor3_1 _2386_ (.A(\i_w_buf[171].A ),
    .B(_0969_),
    .C(_1147_),
    .Y(_1148_));
 sg13g2_xor2_1 _2387_ (.B(_1147_),
    .A(_1139_),
    .X(_1149_));
 sg13g2_nor2b_1 _2388_ (.A(_1149_),
    .B_N(_1138_),
    .Y(_1150_));
 sg13g2_xor2_1 _2389_ (.B(_1149_),
    .A(_1138_),
    .X(_1151_));
 sg13g2_or3_1 _2390_ (.A(\i_w_buf[109].A ),
    .B(_1136_),
    .C(_1151_),
    .X(_1152_));
 sg13g2_xor2_1 _2391_ (.B(_1151_),
    .A(_1137_),
    .X(_1153_));
 sg13g2_xnor2_1 _2392_ (.Y(_1154_),
    .A(_1135_),
    .B(_1153_));
 sg13g2_nand2b_1 _2393_ (.Y(_1155_),
    .B(_1133_),
    .A_N(_1154_));
 sg13g2_xor2_1 _2394_ (.B(_1154_),
    .A(_1133_),
    .X(_1156_));
 sg13g2_xnor2_1 _2395_ (.Y(_1157_),
    .A(_1132_),
    .B(_1156_));
 sg13g2_nand2b_1 _2396_ (.Y(_1158_),
    .B(net99),
    .A_N(\i_w_buf[38].A ));
 sg13g2_nor2_1 _2397_ (.A(\i_w_buf[39].A ),
    .B(_1158_),
    .Y(_1159_));
 sg13g2_nor3_2 _2398_ (.A(_0862_),
    .B(\i_w_buf[68].A ),
    .C(\i_w_buf[69].A ),
    .Y(_1160_));
 sg13g2_nor2_1 _2399_ (.A(net84),
    .B(\i_w_buf[250].A ),
    .Y(_1161_));
 sg13g2_nand2b_1 _2400_ (.Y(_1162_),
    .B(net95),
    .A_N(\i_w_buf[250].A ));
 sg13g2_nor2b_2 _2401_ (.A(\i_w_buf[142].A ),
    .B_N(net89),
    .Y(_1163_));
 sg13g2_nand2_2 _2402_ (.Y(_1164_),
    .A(\i_w_buf[143].A ),
    .B(_1163_));
 sg13g2_nand2_1 _2403_ (.Y(_1165_),
    .A(\i_w_buf[151].A ),
    .B(_1022_));
 sg13g2_nor3_2 _2404_ (.A(net81),
    .B(\i_w_buf[190].A ),
    .C(\i_w_buf[191].A ),
    .Y(_1166_));
 sg13g2_xnor2_1 _2405_ (.Y(_1167_),
    .A(_1165_),
    .B(_1166_));
 sg13g2_nor2b_1 _2406_ (.A(_1167_),
    .B_N(_1164_),
    .Y(_1168_));
 sg13g2_xor2_1 _2407_ (.B(_1167_),
    .A(_1164_),
    .X(_1169_));
 sg13g2_nor2b_1 _2408_ (.A(\i_w_buf[78].A ),
    .B_N(net90),
    .Y(_1170_));
 sg13g2_nand2_1 _2409_ (.Y(_1171_),
    .A(\i_w_buf[79].A ),
    .B(_1170_));
 sg13g2_nor2_1 _2410_ (.A(net84),
    .B(\i_w_buf[186].A ),
    .Y(_1172_));
 sg13g2_nor3_1 _2411_ (.A(net84),
    .B(\i_w_buf[186].A ),
    .C(\i_w_buf[187].A ),
    .Y(_1173_));
 sg13g2_nor2b_1 _2412_ (.A(\i_w_buf[183].A ),
    .B_N(_1134_),
    .Y(_1174_));
 sg13g2_nand3b_1 _2413_ (.B(\i_w_buf[155].A ),
    .C(net95),
    .Y(_1175_),
    .A_N(\i_w_buf[154].A ));
 sg13g2_and2_1 _2414_ (.A(_1174_),
    .B(_1175_),
    .X(_1176_));
 sg13g2_xor2_1 _2415_ (.B(_1175_),
    .A(_1174_),
    .X(_1177_));
 sg13g2_xnor2_1 _2416_ (.Y(_1178_),
    .A(_1173_),
    .B(_1177_));
 sg13g2_nand2b_1 _2417_ (.Y(_1179_),
    .B(_1171_),
    .A_N(_1178_));
 sg13g2_xor2_1 _2418_ (.B(_1178_),
    .A(_1171_),
    .X(_1180_));
 sg13g2_xnor2_1 _2419_ (.Y(_1181_),
    .A(_1169_),
    .B(_1180_));
 sg13g2_nand2_1 _2420_ (.Y(_1182_),
    .A(\i_w_buf[187].A ),
    .B(_1172_));
 sg13g2_nand2b_1 _2421_ (.Y(_1183_),
    .B(_1059_),
    .A_N(\i_w_buf[175].A ));
 sg13g2_nand3b_1 _2422_ (.B(\i_w_buf[87].A ),
    .C(net99),
    .Y(_1184_),
    .A_N(\i_w_buf[86].A ));
 sg13g2_nand2_1 _2423_ (.Y(_1185_),
    .A(\i_w_buf[157].A ),
    .B(_0915_));
 sg13g2_nand3b_1 _2424_ (.B(\i_w_buf[167].A ),
    .C(net99),
    .Y(_1186_),
    .A_N(\i_w_buf[166].A ));
 sg13g2_nand3_1 _2425_ (.B(_0922_),
    .C(_1186_),
    .A(_0895_),
    .Y(_1187_));
 sg13g2_a21o_1 _2426_ (.A2(_0922_),
    .A1(_0895_),
    .B1(_1186_),
    .X(_1188_));
 sg13g2_nand3_1 _2427_ (.B(_1187_),
    .C(_1188_),
    .A(_1185_),
    .Y(_1189_));
 sg13g2_a21o_1 _2428_ (.A2(_1188_),
    .A1(_1187_),
    .B1(_1185_),
    .X(_1190_));
 sg13g2_nand2_1 _2429_ (.Y(_1191_),
    .A(_1189_),
    .B(_1190_));
 sg13g2_nand3_1 _2430_ (.B(_1189_),
    .C(_1190_),
    .A(_1184_),
    .Y(_1192_));
 sg13g2_a21oi_1 _2431_ (.A1(_1189_),
    .A2(_1190_),
    .Y(_1193_),
    .B1(_1184_));
 sg13g2_xnor2_1 _2432_ (.Y(_1194_),
    .A(_1184_),
    .B(_1191_));
 sg13g2_xnor2_1 _2433_ (.Y(_1195_),
    .A(_1183_),
    .B(_1194_));
 sg13g2_nand2_1 _2434_ (.Y(_1196_),
    .A(_1182_),
    .B(_1195_));
 sg13g2_xnor2_1 _2435_ (.Y(_1197_),
    .A(_1182_),
    .B(_1195_));
 sg13g2_xnor2_1 _2436_ (.Y(_1198_),
    .A(_1181_),
    .B(_1197_));
 sg13g2_a21oi_1 _2437_ (.A1(\i_w_buf[251].A ),
    .A2(_1161_),
    .Y(_1199_),
    .B1(_1198_));
 sg13g2_nand3_1 _2438_ (.B(_1161_),
    .C(_1198_),
    .A(\i_w_buf[251].A ),
    .Y(_1200_));
 sg13g2_nand2b_1 _2439_ (.Y(_1201_),
    .B(_1200_),
    .A_N(_1199_));
 sg13g2_xor2_1 _2440_ (.B(_1201_),
    .A(_1160_),
    .X(_1202_));
 sg13g2_or3_1 _2441_ (.A(\i_w_buf[39].A ),
    .B(_1158_),
    .C(_1202_),
    .X(_1203_));
 sg13g2_xor2_1 _2442_ (.B(_1202_),
    .A(_1159_),
    .X(_1204_));
 sg13g2_xor2_1 _2443_ (.B(_1204_),
    .A(_1157_),
    .X(_1205_));
 sg13g2_nand2_1 _2444_ (.Y(_1206_),
    .A(_1091_),
    .B(_1205_));
 sg13g2_xnor2_1 _2445_ (.Y(_1207_),
    .A(_1091_),
    .B(_1205_));
 sg13g2_xor2_1 _2446_ (.B(_1207_),
    .A(_1090_),
    .X(_1208_));
 sg13g2_nand2b_1 _2447_ (.Y(_1209_),
    .B(_1208_),
    .A_N(_1051_));
 sg13g2_xnor2_1 _2448_ (.Y(_1210_),
    .A(_1051_),
    .B(_1208_));
 sg13g2_nand2_1 _2449_ (.Y(_1211_),
    .A(_0959_),
    .B(_1210_));
 sg13g2_xnor2_1 _2450_ (.Y(_1212_),
    .A(_0959_),
    .B(_1210_));
 sg13g2_xnor2_1 _2451_ (.Y(_1213_),
    .A(_0958_),
    .B(_1212_));
 sg13g2_nand2_2 _2452_ (.Y(_1214_),
    .A(\i_w_buf[161].A ),
    .B(_1002_));
 sg13g2_nor2b_1 _2453_ (.A(\i_w_buf[74].A ),
    .B_N(net95),
    .Y(_1215_));
 sg13g2_nand2_2 _2454_ (.Y(_1216_),
    .A(\i_w_buf[75].A ),
    .B(_1215_));
 sg13g2_nor2_1 _2455_ (.A(\i_w_buf[9].A ),
    .B(_0957_),
    .Y(_1217_));
 sg13g2_nand2b_1 _2456_ (.Y(_1218_),
    .B(net92),
    .A_N(\i_w_buf[252].A ));
 sg13g2_nand3b_1 _2457_ (.B(\i_w_buf[253].A ),
    .C(net3),
    .Y(_1219_),
    .A_N(\i_w_buf[252].A ));
 sg13g2_inv_1 _2458_ (.Y(_1220_),
    .A(_1219_));
 sg13g2_nor3_2 _2459_ (.A(_0865_),
    .B(\i_w_buf[76].A ),
    .C(\i_w_buf[77].A ),
    .Y(_1221_));
 sg13g2_nand2_1 _2460_ (.Y(_1222_),
    .A(\i_w_buf[207].A ),
    .B(_1118_));
 sg13g2_inv_1 _2461_ (.Y(_1223_),
    .A(_1222_));
 sg13g2_and2_1 _2462_ (.A(\i_w_buf[215].A ),
    .B(_1108_),
    .X(_1224_));
 sg13g2_nand2_1 _2463_ (.Y(_1225_),
    .A(\i_w_buf[215].A ),
    .B(_1108_));
 sg13g2_nand3b_1 _2464_ (.B(\i_w_buf[103].A ),
    .C(net98),
    .Y(_1226_),
    .A_N(\i_w_buf[102].A ));
 sg13g2_nor3_2 _2465_ (.A(net87),
    .B(\i_w_buf[188].A ),
    .C(\i_w_buf[189].A ),
    .Y(_1227_));
 sg13g2_nor2b_1 _2466_ (.A(\i_w_buf[210].A ),
    .B_N(net103),
    .Y(_1228_));
 sg13g2_nand2_1 _2467_ (.Y(_1229_),
    .A(\i_w_buf[211].A ),
    .B(_1228_));
 sg13g2_nand3b_1 _2468_ (.B(\i_w_buf[213].A ),
    .C(net101),
    .Y(_1230_),
    .A_N(\i_w_buf[212].A ));
 sg13g2_nand3_1 _2469_ (.B(_1163_),
    .C(_1230_),
    .A(_0890_),
    .Y(_1231_));
 sg13g2_a21o_1 _2470_ (.A2(_1163_),
    .A1(_0890_),
    .B1(_1230_),
    .X(_1232_));
 sg13g2_nand3_1 _2471_ (.B(_1231_),
    .C(_1232_),
    .A(_1229_),
    .Y(_1233_));
 sg13g2_a21o_1 _2472_ (.A2(_1232_),
    .A1(_1231_),
    .B1(_1229_),
    .X(_1234_));
 sg13g2_nand3_1 _2473_ (.B(_1233_),
    .C(_1234_),
    .A(_1227_),
    .Y(_1235_));
 sg13g2_a21o_1 _2474_ (.A2(_1234_),
    .A1(_1233_),
    .B1(_1227_),
    .X(_1236_));
 sg13g2_and3_1 _2475_ (.X(_1237_),
    .A(_1226_),
    .B(_1235_),
    .C(_1236_));
 sg13g2_nand3_1 _2476_ (.B(_1235_),
    .C(_1236_),
    .A(_1226_),
    .Y(_1238_));
 sg13g2_a21oi_1 _2477_ (.A1(_1235_),
    .A2(_1236_),
    .Y(_1239_),
    .B1(_1226_));
 sg13g2_a21o_1 _2478_ (.A2(_1236_),
    .A1(_1235_),
    .B1(_1226_),
    .X(_1240_));
 sg13g2_nor3_2 _2479_ (.A(_1224_),
    .B(_1237_),
    .C(_1239_),
    .Y(_1241_));
 sg13g2_nand3_1 _2480_ (.B(_1238_),
    .C(_1240_),
    .A(_1225_),
    .Y(_1242_));
 sg13g2_a21oi_1 _2481_ (.A1(_1238_),
    .A2(_1240_),
    .Y(_1243_),
    .B1(_1225_));
 sg13g2_o21ai_1 _2482_ (.B1(_1224_),
    .Y(_1244_),
    .A1(_1237_),
    .A2(_1239_));
 sg13g2_nor3_1 _2483_ (.A(_1223_),
    .B(_1241_),
    .C(_1243_),
    .Y(_1245_));
 sg13g2_nand3_1 _2484_ (.B(_1242_),
    .C(_1244_),
    .A(_1222_),
    .Y(_1246_));
 sg13g2_a21oi_1 _2485_ (.A1(_1242_),
    .A2(_1244_),
    .Y(_1247_),
    .B1(_1222_));
 sg13g2_o21ai_1 _2486_ (.B1(_1223_),
    .Y(_1248_),
    .A1(_1241_),
    .A2(_1243_));
 sg13g2_nand3_1 _2487_ (.B(_1246_),
    .C(_1248_),
    .A(_1221_),
    .Y(_1249_));
 sg13g2_a21oi_1 _2488_ (.A1(_1246_),
    .A2(_1248_),
    .Y(_1250_),
    .B1(_1221_));
 sg13g2_nor3_1 _2489_ (.A(_1221_),
    .B(_1245_),
    .C(_1247_),
    .Y(_1251_));
 sg13g2_o21ai_1 _2490_ (.B1(_1221_),
    .Y(_1252_),
    .A1(_1245_),
    .A2(_1247_));
 sg13g2_nand2b_1 _2491_ (.Y(_1253_),
    .B(_1252_),
    .A_N(_1251_));
 sg13g2_xnor2_1 _2492_ (.Y(_1254_),
    .A(_1219_),
    .B(_1253_));
 sg13g2_nor3_1 _2493_ (.A(net81),
    .B(\i_w_buf[46].A ),
    .C(\i_w_buf[47].A ),
    .Y(_1255_));
 sg13g2_nand2b_1 _2494_ (.Y(_1256_),
    .B(_0917_),
    .A_N(\i_w_buf[47].A ));
 sg13g2_nor2b_1 _2495_ (.A(\i_w_buf[62].A ),
    .B_N(net89),
    .Y(_1257_));
 sg13g2_nand2_2 _2496_ (.Y(_1258_),
    .A(\i_w_buf[63].A ),
    .B(_1257_));
 sg13g2_nor2_1 _2497_ (.A(net83),
    .B(\i_w_buf[218].A ),
    .Y(_1259_));
 sg13g2_and2_1 _2498_ (.A(\i_w_buf[219].A ),
    .B(_1259_),
    .X(_1260_));
 sg13g2_nand2_1 _2499_ (.Y(_1261_),
    .A(\i_w_buf[219].A ),
    .B(_1259_));
 sg13g2_nor2_1 _2500_ (.A(net81),
    .B(\i_w_buf[126].A ),
    .Y(_1262_));
 sg13g2_nor3_2 _2501_ (.A(net81),
    .B(\i_w_buf[126].A ),
    .C(\i_w_buf[127].A ),
    .Y(_1263_));
 sg13g2_nor2b_1 _2502_ (.A(\i_w_buf[121].A ),
    .B_N(_1143_),
    .Y(_1264_));
 sg13g2_inv_1 _2503_ (.Y(_1265_),
    .A(_1264_));
 sg13g2_nand3b_1 _2504_ (.B(\i_w_buf[23].A ),
    .C(net98),
    .Y(_1266_),
    .A_N(\i_w_buf[22].A ));
 sg13g2_nor2b_1 _2505_ (.A(\i_w_buf[118].A ),
    .B_N(net98),
    .Y(_1267_));
 sg13g2_nor2b_1 _2506_ (.A(\i_w_buf[119].A ),
    .B_N(_1267_),
    .Y(_1268_));
 sg13g2_nand2_1 _2507_ (.Y(_1269_),
    .A(_1266_),
    .B(_1268_));
 sg13g2_xnor2_1 _2508_ (.Y(_1270_),
    .A(_1266_),
    .B(_1268_));
 sg13g2_xnor2_1 _2509_ (.Y(_1271_),
    .A(_1265_),
    .B(_1270_));
 sg13g2_nor2_1 _2510_ (.A(net88),
    .B(\i_w_buf[196].A ),
    .Y(_1272_));
 sg13g2_nor3_2 _2511_ (.A(net88),
    .B(\i_w_buf[196].A ),
    .C(\i_w_buf[197].A ),
    .Y(_1273_));
 sg13g2_nor2b_1 _2512_ (.A(\i_w_buf[114].A ),
    .B_N(net103),
    .Y(_1274_));
 sg13g2_nor2b_1 _2513_ (.A(\i_w_buf[115].A ),
    .B_N(_1274_),
    .Y(_1275_));
 sg13g2_nor2b_2 _2514_ (.A(\i_w_buf[110].A ),
    .B_N(net89),
    .Y(_1276_));
 sg13g2_nor2b_1 _2515_ (.A(\i_w_buf[26].A ),
    .B_N(net94),
    .Y(_1277_));
 sg13g2_nand3b_1 _2516_ (.B(\i_w_buf[27].A ),
    .C(net94),
    .Y(_1278_),
    .A_N(\i_w_buf[26].A ));
 sg13g2_nand3_1 _2517_ (.B(_1276_),
    .C(_1278_),
    .A(_0885_),
    .Y(_1279_));
 sg13g2_a21o_1 _2518_ (.A2(_1276_),
    .A1(_0885_),
    .B1(_1278_),
    .X(_1280_));
 sg13g2_nand3_1 _2519_ (.B(_1279_),
    .C(_1280_),
    .A(_1275_),
    .Y(_1281_));
 sg13g2_a21o_1 _2520_ (.A2(_1280_),
    .A1(_1279_),
    .B1(_1275_),
    .X(_1282_));
 sg13g2_and3_1 _2521_ (.X(_1283_),
    .A(_1273_),
    .B(_1281_),
    .C(_1282_));
 sg13g2_a21oi_1 _2522_ (.A1(_1281_),
    .A2(_1282_),
    .Y(_1284_),
    .B1(_1273_));
 sg13g2_or3_1 _2523_ (.A(_1271_),
    .B(_1283_),
    .C(_1284_),
    .X(_1285_));
 sg13g2_o21ai_1 _2524_ (.B1(_1271_),
    .Y(_1286_),
    .A1(_1283_),
    .A2(_1284_));
 sg13g2_nand3_1 _2525_ (.B(_1285_),
    .C(_1286_),
    .A(_1263_),
    .Y(_1287_));
 sg13g2_a21oi_1 _2526_ (.A1(_1285_),
    .A2(_1286_),
    .Y(_1288_),
    .B1(_1263_));
 sg13g2_a21o_1 _2527_ (.A2(_1286_),
    .A1(_1285_),
    .B1(_1263_),
    .X(_1289_));
 sg13g2_nand3_1 _2528_ (.B(_1287_),
    .C(_1289_),
    .A(_1261_),
    .Y(_1290_));
 sg13g2_a21o_1 _2529_ (.A2(_1289_),
    .A1(_1287_),
    .B1(_1261_),
    .X(_1291_));
 sg13g2_nand3_1 _2530_ (.B(_1290_),
    .C(_1291_),
    .A(_1258_),
    .Y(_1292_));
 sg13g2_a21oi_1 _2531_ (.A1(_1290_),
    .A2(_1291_),
    .Y(_1293_),
    .B1(_1258_));
 sg13g2_a21o_1 _2532_ (.A2(_1291_),
    .A1(_1290_),
    .B1(_1258_),
    .X(_1294_));
 sg13g2_nand3b_1 _2533_ (.B(\i_w_buf[217].A ),
    .C(net96),
    .Y(_1295_),
    .A_N(\i_w_buf[216].A ));
 sg13g2_inv_1 _2534_ (.Y(_1296_),
    .A(_1295_));
 sg13g2_nand3b_1 _2535_ (.B(\i_w_buf[227].A ),
    .C(net103),
    .Y(_1297_),
    .A_N(\i_w_buf[226].A ));
 sg13g2_nor2b_2 _2536_ (.A(\i_w_buf[137].A ),
    .B_N(_0900_),
    .Y(_1298_));
 sg13g2_nand2_1 _2537_ (.Y(_1299_),
    .A(_1297_),
    .B(_1298_));
 sg13g2_xnor2_1 _2538_ (.Y(_1300_),
    .A(_1297_),
    .B(_1298_));
 sg13g2_xnor2_1 _2539_ (.Y(_1301_),
    .A(_1296_),
    .B(_1300_));
 sg13g2_nor2b_1 _2540_ (.A(\i_w_buf[106].A ),
    .B_N(net93),
    .Y(_1302_));
 sg13g2_nand2_1 _2541_ (.Y(_1303_),
    .A(\i_w_buf[107].A ),
    .B(_1302_));
 sg13g2_nor2b_1 _2542_ (.A(\i_w_buf[132].A ),
    .B_N(net101),
    .Y(_1304_));
 sg13g2_nor2b_1 _2543_ (.A(\i_w_buf[133].A ),
    .B_N(_1304_),
    .Y(_1305_));
 sg13g2_nor2b_2 _2544_ (.A(\i_w_buf[128].A ),
    .B_N(net107),
    .Y(_1306_));
 sg13g2_nand3b_1 _2545_ (.B(\i_w_buf[229].A ),
    .C(net101),
    .Y(_1307_),
    .A_N(\i_w_buf[228].A ));
 sg13g2_nand3_1 _2546_ (.B(_1306_),
    .C(_1307_),
    .A(_0886_),
    .Y(_1308_));
 sg13g2_a21o_1 _2547_ (.A2(_1306_),
    .A1(_0886_),
    .B1(_1307_),
    .X(_1309_));
 sg13g2_nand3_1 _2548_ (.B(_1308_),
    .C(_1309_),
    .A(_1305_),
    .Y(_1310_));
 sg13g2_a21o_1 _2549_ (.A2(_1309_),
    .A1(_1308_),
    .B1(_1305_),
    .X(_1311_));
 sg13g2_nand2_1 _2550_ (.Y(_1312_),
    .A(_1310_),
    .B(_1311_));
 sg13g2_nand3_1 _2551_ (.B(_1310_),
    .C(_1311_),
    .A(_1303_),
    .Y(_1313_));
 sg13g2_a21oi_1 _2552_ (.A1(_1310_),
    .A2(_1311_),
    .Y(_1314_),
    .B1(_1303_));
 sg13g2_xor2_1 _2553_ (.B(_1312_),
    .A(_1303_),
    .X(_1315_));
 sg13g2_xnor2_1 _2554_ (.Y(_1316_),
    .A(_1301_),
    .B(_1315_));
 sg13g2_nor3_2 _2555_ (.A(net83),
    .B(\i_w_buf[122].A ),
    .C(\i_w_buf[123].A ),
    .Y(_1317_));
 sg13g2_nor3_2 _2556_ (.A(net85),
    .B(\i_w_buf[192].A ),
    .C(\i_w_buf[193].A ),
    .Y(_1318_));
 sg13g2_nand3b_1 _2557_ (.B(\i_w_buf[109].A ),
    .C(net91),
    .Y(_1319_),
    .A_N(\i_w_buf[108].A ));
 sg13g2_nor2b_1 _2558_ (.A(\i_w_buf[232].A ),
    .B_N(net97),
    .Y(_1320_));
 sg13g2_nand2_1 _2559_ (.Y(_1321_),
    .A(\i_w_buf[233].A ),
    .B(_1320_));
 sg13g2_nand3b_1 _2560_ (.B(\i_w_buf[241].A ),
    .C(net107),
    .Y(_1322_),
    .A_N(\i_w_buf[240].A ));
 sg13g2_nor2b_1 _2561_ (.A(\i_w_buf[124].A ),
    .B_N(net91),
    .Y(_1323_));
 sg13g2_nand3_1 _2562_ (.B(_1322_),
    .C(_1323_),
    .A(_0868_),
    .Y(_1324_));
 sg13g2_a21o_1 _2563_ (.A2(_1323_),
    .A1(_0868_),
    .B1(_1322_),
    .X(_1325_));
 sg13g2_nand3_1 _2564_ (.B(_1324_),
    .C(_1325_),
    .A(_1321_),
    .Y(_1326_));
 sg13g2_a21o_1 _2565_ (.A2(_1325_),
    .A1(_1324_),
    .B1(_1321_),
    .X(_1327_));
 sg13g2_and3_1 _2566_ (.X(_1328_),
    .A(_1319_),
    .B(_1326_),
    .C(_1327_));
 sg13g2_nand3_1 _2567_ (.B(_1326_),
    .C(_1327_),
    .A(_1319_),
    .Y(_1329_));
 sg13g2_a21o_1 _2568_ (.A2(_1327_),
    .A1(_1326_),
    .B1(_1319_),
    .X(_1330_));
 sg13g2_nand3_1 _2569_ (.B(_1329_),
    .C(_1330_),
    .A(_1318_),
    .Y(_1331_));
 sg13g2_a21o_1 _2570_ (.A2(_1330_),
    .A1(_1329_),
    .B1(_1318_),
    .X(_1332_));
 sg13g2_nand2_1 _2571_ (.Y(_1333_),
    .A(_1331_),
    .B(_1332_));
 sg13g2_nand3_1 _2572_ (.B(_1331_),
    .C(_1332_),
    .A(_1317_),
    .Y(_1334_));
 sg13g2_a21oi_1 _2573_ (.A1(_1331_),
    .A2(_1332_),
    .Y(_1335_),
    .B1(_1317_));
 sg13g2_xor2_1 _2574_ (.B(_1333_),
    .A(_1317_),
    .X(_1336_));
 sg13g2_xor2_1 _2575_ (.B(_1336_),
    .A(_1316_),
    .X(_1337_));
 sg13g2_xnor2_1 _2576_ (.Y(_1338_),
    .A(_1316_),
    .B(_1336_));
 sg13g2_nand3_1 _2577_ (.B(_1294_),
    .C(_1337_),
    .A(_1292_),
    .Y(_1339_));
 sg13g2_a21o_1 _2578_ (.A2(_1294_),
    .A1(_1292_),
    .B1(_1337_),
    .X(_1340_));
 sg13g2_nand3_1 _2579_ (.B(_1339_),
    .C(_1340_),
    .A(_1255_),
    .Y(_1341_));
 sg13g2_a21oi_1 _2580_ (.A1(_1339_),
    .A2(_1340_),
    .Y(_1342_),
    .B1(_1255_));
 sg13g2_a21oi_1 _2581_ (.A1(_1339_),
    .A2(_1340_),
    .Y(_1343_),
    .B1(_1256_));
 sg13g2_nand3_1 _2582_ (.B(_1339_),
    .C(_1340_),
    .A(_1256_),
    .Y(_1344_));
 sg13g2_nor2b_1 _2583_ (.A(_1343_),
    .B_N(_1344_),
    .Y(_1345_));
 sg13g2_xnor2_1 _2584_ (.Y(_1346_),
    .A(_1254_),
    .B(_1345_));
 sg13g2_nor2_1 _2585_ (.A(net84),
    .B(\i_w_buf[10].A ),
    .Y(_1347_));
 sg13g2_nand2_2 _2586_ (.Y(_1348_),
    .A(\i_w_buf[11].A ),
    .B(_1347_));
 sg13g2_nand2_2 _2587_ (.Y(_1349_),
    .A(\i_w_buf[255].A ),
    .B(_0932_));
 sg13g2_inv_1 _2588_ (.Y(_1350_),
    .A(_1349_));
 sg13g2_nor3_1 _2589_ (.A(_0864_),
    .B(\i_w_buf[50].A ),
    .C(\i_w_buf[51].A ),
    .Y(_1351_));
 sg13g2_nand3b_1 _2590_ (.B(\i_w_buf[95].A ),
    .C(net89),
    .Y(_1352_),
    .A_N(\i_w_buf[94].A ));
 sg13g2_nor2b_1 _2591_ (.A(\i_w_buf[82].A ),
    .B_N(net105),
    .Y(_1353_));
 sg13g2_nor2b_2 _2592_ (.A(\i_w_buf[83].A ),
    .B_N(_1353_),
    .Y(_1354_));
 sg13g2_nand2_1 _2593_ (.Y(_1355_),
    .A(\i_w_buf[115].A ),
    .B(_1274_));
 sg13g2_inv_1 _2594_ (.Y(_1356_),
    .A(_1355_));
 sg13g2_nor3_2 _2595_ (.A(net83),
    .B(\i_w_buf[202].A ),
    .C(\i_w_buf[203].A ),
    .Y(_1357_));
 sg13g2_nor2b_1 _2596_ (.A(\i_w_buf[28].A ),
    .B_N(net92),
    .Y(_1358_));
 sg13g2_nand2_2 _2597_ (.Y(_1359_),
    .A(\i_w_buf[29].A ),
    .B(_1358_));
 sg13g2_nand3b_1 _2598_ (.B(\i_w_buf[39].A ),
    .C(net99),
    .Y(_1360_),
    .A_N(\i_w_buf[38].A ));
 sg13g2_nand3_1 _2599_ (.B(_1302_),
    .C(_1360_),
    .A(_0889_),
    .Y(_1361_));
 sg13g2_a21o_1 _2600_ (.A2(_1302_),
    .A1(_0889_),
    .B1(_1360_),
    .X(_1362_));
 sg13g2_nand3_1 _2601_ (.B(_1361_),
    .C(_1362_),
    .A(_1359_),
    .Y(_1363_));
 sg13g2_a21o_1 _2602_ (.A2(_1362_),
    .A1(_1361_),
    .B1(_1359_),
    .X(_1364_));
 sg13g2_and3_1 _2603_ (.X(_1365_),
    .A(_1357_),
    .B(_1363_),
    .C(_1364_));
 sg13g2_nand3_1 _2604_ (.B(_1363_),
    .C(_1364_),
    .A(_1357_),
    .Y(_1366_));
 sg13g2_a21oi_1 _2605_ (.A1(_1363_),
    .A2(_1364_),
    .Y(_1367_),
    .B1(_1357_));
 sg13g2_nor2_1 _2606_ (.A(_1365_),
    .B(_1367_),
    .Y(_1368_));
 sg13g2_xnor2_1 _2607_ (.Y(_1369_),
    .A(_1355_),
    .B(_1368_));
 sg13g2_nand3b_1 _2608_ (.B(\i_w_buf[221].A ),
    .C(net91),
    .Y(_1370_),
    .A_N(\i_w_buf[220].A ));
 sg13g2_nor3_2 _2609_ (.A(net80),
    .B(\i_w_buf[102].A ),
    .C(\i_w_buf[103].A ),
    .Y(_1371_));
 sg13g2_nand3b_1 _2610_ (.B(\i_w_buf[45].A ),
    .C(net92),
    .Y(_1372_),
    .A_N(\i_w_buf[44].A ));
 sg13g2_nand3b_1 _2611_ (.B(\i_w_buf[43].A ),
    .C(net93),
    .Y(_1373_),
    .A_N(\i_w_buf[42].A ));
 sg13g2_and2_1 _2612_ (.A(_1372_),
    .B(_1373_),
    .X(_1374_));
 sg13g2_xor2_1 _2613_ (.B(_1373_),
    .A(_1372_),
    .X(_1375_));
 sg13g2_xnor2_1 _2614_ (.Y(_1376_),
    .A(_1371_),
    .B(_1375_));
 sg13g2_nor3_2 _2615_ (.A(net87),
    .B(\i_w_buf[204].A ),
    .C(\i_w_buf[205].A ),
    .Y(_1377_));
 sg13g2_nor2b_1 _2616_ (.A(\i_w_buf[96].A ),
    .B_N(net107),
    .Y(_1378_));
 sg13g2_nor2b_1 _2617_ (.A(\i_w_buf[97].A ),
    .B_N(_1378_),
    .Y(_1379_));
 sg13g2_nand3b_1 _2618_ (.B(\i_w_buf[51].A ),
    .C(net104),
    .Y(_1380_),
    .A_N(\i_w_buf[50].A ));
 sg13g2_nand3_1 _2619_ (.B(_0998_),
    .C(_1380_),
    .A(_0888_),
    .Y(_1381_));
 sg13g2_a21o_1 _2620_ (.A2(_0998_),
    .A1(_0888_),
    .B1(_1380_),
    .X(_1382_));
 sg13g2_nand3_1 _2621_ (.B(_1381_),
    .C(_1382_),
    .A(_1379_),
    .Y(_1383_));
 sg13g2_a21o_1 _2622_ (.A2(_1382_),
    .A1(_1381_),
    .B1(_1379_),
    .X(_1384_));
 sg13g2_and3_1 _2623_ (.X(_1385_),
    .A(_1377_),
    .B(_1383_),
    .C(_1384_));
 sg13g2_nand3_1 _2624_ (.B(_1383_),
    .C(_1384_),
    .A(_1377_),
    .Y(_1386_));
 sg13g2_a21oi_1 _2625_ (.A1(_1383_),
    .A2(_1384_),
    .Y(_1387_),
    .B1(_1377_));
 sg13g2_or3_1 _2626_ (.A(_1376_),
    .B(_1385_),
    .C(_1387_),
    .X(_1388_));
 sg13g2_o21ai_1 _2627_ (.B1(_1376_),
    .Y(_1389_),
    .A1(_1385_),
    .A2(_1387_));
 sg13g2_and3_1 _2628_ (.X(_1390_),
    .A(_1370_),
    .B(_1388_),
    .C(_1389_));
 sg13g2_a21oi_1 _2629_ (.A1(_1388_),
    .A2(_1389_),
    .Y(_1391_),
    .B1(_1370_));
 sg13g2_or3_1 _2630_ (.A(_1369_),
    .B(_1390_),
    .C(_1391_),
    .X(_1392_));
 sg13g2_o21ai_1 _2631_ (.B1(_1369_),
    .Y(_1393_),
    .A1(_1390_),
    .A2(_1391_));
 sg13g2_nand3_1 _2632_ (.B(_1392_),
    .C(_1393_),
    .A(_1354_),
    .Y(_1394_));
 sg13g2_a21o_1 _2633_ (.A2(_1393_),
    .A1(_1392_),
    .B1(_1354_),
    .X(_1395_));
 sg13g2_nand3_1 _2634_ (.B(_1394_),
    .C(_1395_),
    .A(_1352_),
    .Y(_1396_));
 sg13g2_a21o_1 _2635_ (.A2(_1395_),
    .A1(_1394_),
    .B1(_1352_),
    .X(_1397_));
 sg13g2_and3_1 _2636_ (.X(_1398_),
    .A(_1351_),
    .B(_1396_),
    .C(_1397_));
 sg13g2_nand3_1 _2637_ (.B(_1396_),
    .C(_1397_),
    .A(_1351_),
    .Y(_1399_));
 sg13g2_a21oi_1 _2638_ (.A1(_1396_),
    .A2(_1397_),
    .Y(_1400_),
    .B1(_1351_));
 sg13g2_nor3_1 _2639_ (.A(_1350_),
    .B(_1398_),
    .C(_1400_),
    .Y(_1401_));
 sg13g2_o21ai_1 _2640_ (.B1(_1350_),
    .Y(_1402_),
    .A1(_1398_),
    .A2(_1400_));
 sg13g2_nor2b_2 _2641_ (.A(_1401_),
    .B_N(_1402_),
    .Y(_1403_));
 sg13g2_nand2_1 _2642_ (.Y(_1404_),
    .A(_1348_),
    .B(_1403_));
 sg13g2_xnor2_1 _2643_ (.Y(_1405_),
    .A(_1348_),
    .B(_1403_));
 sg13g2_xnor2_1 _2644_ (.Y(_1406_),
    .A(_1346_),
    .B(_1405_));
 sg13g2_nor3_1 _2645_ (.A(\i_w_buf[9].A ),
    .B(_0957_),
    .C(_1406_),
    .Y(_1407_));
 sg13g2_xnor2_1 _2646_ (.Y(_1408_),
    .A(_1217_),
    .B(_1406_));
 sg13g2_xnor2_1 _2647_ (.Y(_1409_),
    .A(_1216_),
    .B(_1408_));
 sg13g2_nand2_2 _2648_ (.Y(_1410_),
    .A(\i_w_buf[129].A ),
    .B(_1306_));
 sg13g2_nor3_2 _2649_ (.A(net80),
    .B(\i_w_buf[22].A ),
    .C(\i_w_buf[23].A ),
    .Y(_1411_));
 sg13g2_nand2b_1 _2650_ (.Y(_1412_),
    .B(_1121_),
    .A_N(\i_w_buf[25].A ));
 sg13g2_nor3_2 _2651_ (.A(_0864_),
    .B(\i_w_buf[130].A ),
    .C(\i_w_buf[131].A ),
    .Y(_1413_));
 sg13g2_and2_1 _2652_ (.A(\i_w_buf[231].A ),
    .B(_1069_),
    .X(_1414_));
 sg13g2_nor2b_1 _2653_ (.A(\i_w_buf[20].A ),
    .B_N(net101),
    .Y(_1415_));
 sg13g2_nand2_2 _2654_ (.Y(_1416_),
    .A(\i_w_buf[21].A ),
    .B(_1415_));
 sg13g2_nor2b_1 _2655_ (.A(\i_w_buf[211].A ),
    .B_N(_1228_),
    .Y(_1417_));
 sg13g2_nor2b_2 _2656_ (.A(\i_w_buf[52].A ),
    .B_N(net101),
    .Y(_1418_));
 sg13g2_nand2_2 _2657_ (.Y(_1419_),
    .A(\i_w_buf[53].A ),
    .B(_1418_));
 sg13g2_nor2b_1 _2658_ (.A(\i_w_buf[56].A ),
    .B_N(net96),
    .Y(_1420_));
 sg13g2_nand3b_1 _2659_ (.B(\i_w_buf[57].A ),
    .C(net96),
    .Y(_1421_),
    .A_N(\i_w_buf[56].A ));
 sg13g2_nor2b_2 _2660_ (.A(\i_w_buf[88].A ),
    .B_N(net96),
    .Y(_1422_));
 sg13g2_nand3_1 _2661_ (.B(_1421_),
    .C(_1422_),
    .A(_0882_),
    .Y(_1423_));
 sg13g2_a21o_1 _2662_ (.A2(_1422_),
    .A1(_0882_),
    .B1(_1421_),
    .X(_1424_));
 sg13g2_nand3_1 _2663_ (.B(_1423_),
    .C(_1424_),
    .A(_1419_),
    .Y(_1425_));
 sg13g2_a21o_1 _2664_ (.A2(_1424_),
    .A1(_1423_),
    .B1(_1419_),
    .X(_1426_));
 sg13g2_nand3_1 _2665_ (.B(_1425_),
    .C(_1426_),
    .A(_1417_),
    .Y(_1427_));
 sg13g2_a21o_1 _2666_ (.A2(_1426_),
    .A1(_1425_),
    .B1(_1417_),
    .X(_1428_));
 sg13g2_and3_1 _2667_ (.X(_1429_),
    .A(_1416_),
    .B(_1427_),
    .C(_1428_));
 sg13g2_nand3_1 _2668_ (.B(_1427_),
    .C(_1428_),
    .A(_1416_),
    .Y(_1430_));
 sg13g2_a21oi_1 _2669_ (.A1(_1427_),
    .A2(_1428_),
    .Y(_1431_),
    .B1(_1416_));
 sg13g2_nor3_1 _2670_ (.A(_1414_),
    .B(_1429_),
    .C(_1431_),
    .Y(_1432_));
 sg13g2_o21ai_1 _2671_ (.B1(_1414_),
    .Y(_1433_),
    .A1(_1429_),
    .A2(_1431_));
 sg13g2_nor2b_1 _2672_ (.A(_1432_),
    .B_N(_1433_),
    .Y(_1434_));
 sg13g2_xnor2_1 _2673_ (.Y(_1435_),
    .A(_1413_),
    .B(_1434_));
 sg13g2_and2_1 _2674_ (.A(\i_w_buf[111].A ),
    .B(_1276_),
    .X(_1436_));
 sg13g2_nand2_1 _2675_ (.Y(_1437_),
    .A(\i_w_buf[111].A ),
    .B(_1276_));
 sg13g2_nor2b_1 _2676_ (.A(\i_w_buf[134].A ),
    .B_N(net98),
    .Y(_1438_));
 sg13g2_nor2b_1 _2677_ (.A(\i_w_buf[135].A ),
    .B_N(_1438_),
    .Y(_1439_));
 sg13g2_and2_1 _2678_ (.A(\i_w_buf[13].A ),
    .B(_0908_),
    .X(_1440_));
 sg13g2_nand2_1 _2679_ (.Y(_1441_),
    .A(\i_w_buf[13].A ),
    .B(_0908_));
 sg13g2_nor3_2 _2680_ (.A(net83),
    .B(\i_w_buf[218].A ),
    .C(\i_w_buf[219].A ),
    .Y(_1442_));
 sg13g2_nand2_1 _2681_ (.Y(_1443_),
    .A(\i_w_buf[83].A ),
    .B(_1353_));
 sg13g2_nand3b_1 _2682_ (.B(\i_w_buf[85].A ),
    .C(net100),
    .Y(_1444_),
    .A_N(\i_w_buf[84].A ));
 sg13g2_nor2b_2 _2683_ (.A(\i_w_buf[70].A ),
    .B_N(net99),
    .Y(_1445_));
 sg13g2_nand3_1 _2684_ (.B(_1444_),
    .C(_1445_),
    .A(_0883_),
    .Y(_1446_));
 sg13g2_a21o_1 _2685_ (.A2(_1445_),
    .A1(_0883_),
    .B1(_1444_),
    .X(_1447_));
 sg13g2_nand3_1 _2686_ (.B(_1446_),
    .C(_1447_),
    .A(_1443_),
    .Y(_1448_));
 sg13g2_a21o_1 _2687_ (.A2(_1447_),
    .A1(_1446_),
    .B1(_1443_),
    .X(_1449_));
 sg13g2_nand3_1 _2688_ (.B(_1448_),
    .C(_1449_),
    .A(_1442_),
    .Y(_1450_));
 sg13g2_a21oi_1 _2689_ (.A1(_1448_),
    .A2(_1449_),
    .Y(_1451_),
    .B1(_1442_));
 sg13g2_a21o_1 _2690_ (.A2(_1449_),
    .A1(_1448_),
    .B1(_1442_),
    .X(_1452_));
 sg13g2_nand3_1 _2691_ (.B(_1450_),
    .C(_1452_),
    .A(_1441_),
    .Y(_1453_));
 sg13g2_a21o_1 _2692_ (.A2(_1452_),
    .A1(_1450_),
    .B1(_1441_),
    .X(_1454_));
 sg13g2_nand3_1 _2693_ (.B(_1453_),
    .C(_1454_),
    .A(_1439_),
    .Y(_1455_));
 sg13g2_a21oi_1 _2694_ (.A1(_1453_),
    .A2(_1454_),
    .Y(_1456_),
    .B1(_1439_));
 sg13g2_a21o_1 _2695_ (.A2(_1454_),
    .A1(_1453_),
    .B1(_1439_),
    .X(_1457_));
 sg13g2_nor3_1 _2696_ (.A(net88),
    .B(\i_w_buf[84].A ),
    .C(\i_w_buf[85].A ),
    .Y(_1458_));
 sg13g2_nor3_1 _2697_ (.A(net86),
    .B(\i_w_buf[80].A ),
    .C(\i_w_buf[81].A ),
    .Y(_1459_));
 sg13g2_nand2_1 _2698_ (.Y(_1460_),
    .A(\i_w_buf[71].A ),
    .B(_1445_));
 sg13g2_and2_1 _2699_ (.A(_1459_),
    .B(_1460_),
    .X(_1461_));
 sg13g2_xor2_1 _2700_ (.B(_1460_),
    .A(_1459_),
    .X(_1462_));
 sg13g2_xnor2_1 _2701_ (.Y(_1463_),
    .A(_1458_),
    .B(_1462_));
 sg13g2_nor3_2 _2702_ (.A(net88),
    .B(\i_w_buf[212].A ),
    .C(\i_w_buf[213].A ),
    .Y(_1464_));
 sg13g2_nor2b_1 _2703_ (.A(\i_w_buf[79].A ),
    .B_N(_1170_),
    .Y(_1465_));
 sg13g2_nand3b_1 _2704_ (.B(\i_w_buf[77].A ),
    .C(net92),
    .Y(_1466_),
    .A_N(\i_w_buf[76].A ));
 sg13g2_nand3_1 _2705_ (.B(_1215_),
    .C(_1466_),
    .A(_0884_),
    .Y(_1467_));
 sg13g2_a21o_1 _2706_ (.A2(_1215_),
    .A1(_0884_),
    .B1(_1466_),
    .X(_1468_));
 sg13g2_nand3_1 _2707_ (.B(_1467_),
    .C(_1468_),
    .A(_1465_),
    .Y(_1469_));
 sg13g2_a21o_2 _2708_ (.A2(_1468_),
    .A1(_1467_),
    .B1(_1465_),
    .X(_1470_));
 sg13g2_nand2_1 _2709_ (.Y(_1471_),
    .A(_1469_),
    .B(_1470_));
 sg13g2_nand3_1 _2710_ (.B(_1469_),
    .C(_1470_),
    .A(_1464_),
    .Y(_1472_));
 sg13g2_xor2_1 _2711_ (.B(_1471_),
    .A(_1464_),
    .X(_1473_));
 sg13g2_xor2_1 _2712_ (.B(_1473_),
    .A(_1463_),
    .X(_1474_));
 sg13g2_xnor2_1 _2713_ (.Y(_1475_),
    .A(_1463_),
    .B(_1473_));
 sg13g2_nand3_1 _2714_ (.B(_1457_),
    .C(_1474_),
    .A(_1455_),
    .Y(_1476_));
 sg13g2_a21o_2 _2715_ (.A2(_1457_),
    .A1(_1455_),
    .B1(_1474_),
    .X(_1477_));
 sg13g2_nand3_1 _2716_ (.B(_1476_),
    .C(_1477_),
    .A(_1437_),
    .Y(_1478_));
 sg13g2_a21oi_1 _2717_ (.A1(_1476_),
    .A2(_1477_),
    .Y(_1479_),
    .B1(_1437_));
 sg13g2_a21oi_1 _2718_ (.A1(_1476_),
    .A2(_1477_),
    .Y(_1480_),
    .B1(_1436_));
 sg13g2_nand3_1 _2719_ (.B(_1476_),
    .C(_1477_),
    .A(_1436_),
    .Y(_1481_));
 sg13g2_nor2b_1 _2720_ (.A(_1480_),
    .B_N(_1481_),
    .Y(_1482_));
 sg13g2_xnor2_1 _2721_ (.Y(_1483_),
    .A(_1435_),
    .B(_1482_));
 sg13g2_and2_1 _2722_ (.A(\i_w_buf[127].A ),
    .B(_1262_),
    .X(_1484_));
 sg13g2_nand2_1 _2723_ (.Y(_1485_),
    .A(\i_w_buf[127].A ),
    .B(_1262_));
 sg13g2_nor3_1 _2724_ (.A(net80),
    .B(\i_w_buf[86].A ),
    .C(\i_w_buf[87].A ),
    .Y(_1486_));
 sg13g2_nand2_2 _2725_ (.Y(_1487_),
    .A(\i_w_buf[119].A ),
    .B(_1267_));
 sg13g2_nand3b_1 _2726_ (.B(\i_w_buf[235].A ),
    .C(net94),
    .Y(_1488_),
    .A_N(\i_w_buf[234].A ));
 sg13g2_nor3_1 _2727_ (.A(net83),
    .B(\i_w_buf[138].A ),
    .C(\i_w_buf[139].A ),
    .Y(_1489_));
 sg13g2_nor2b_1 _2728_ (.A(\i_w_buf[66].A ),
    .B_N(net105),
    .Y(_1490_));
 sg13g2_nor2b_2 _2729_ (.A(\i_w_buf[67].A ),
    .B_N(_1490_),
    .Y(_1491_));
 sg13g2_nor2b_1 _2730_ (.A(\i_w_buf[63].A ),
    .B_N(_1257_),
    .Y(_1492_));
 sg13g2_nand2_2 _2731_ (.Y(_1493_),
    .A(\i_w_buf[89].A ),
    .B(_1422_));
 sg13g2_and2_1 _2732_ (.A(_1492_),
    .B(_1493_),
    .X(_1494_));
 sg13g2_xor2_1 _2733_ (.B(_1493_),
    .A(_1492_),
    .X(_1495_));
 sg13g2_xnor2_1 _2734_ (.Y(_1496_),
    .A(_1491_),
    .B(_1495_));
 sg13g2_nor2b_2 _2735_ (.A(\i_w_buf[6].A ),
    .B_N(net99),
    .Y(_1497_));
 sg13g2_nand2_2 _2736_ (.Y(_1498_),
    .A(\i_w_buf[7].A ),
    .B(_1497_));
 sg13g2_nand2_1 _2737_ (.Y(_1499_),
    .A(\i_w_buf[99].A ),
    .B(_0913_));
 sg13g2_nand3b_1 _2738_ (.B(\i_w_buf[101].A ),
    .C(net101),
    .Y(_1500_),
    .A_N(\i_w_buf[100].A ));
 sg13g2_nand3_1 _2739_ (.B(_1420_),
    .C(_1500_),
    .A(_0881_),
    .Y(_1501_));
 sg13g2_a21o_1 _2740_ (.A2(_1420_),
    .A1(_0881_),
    .B1(_1500_),
    .X(_1502_));
 sg13g2_nand3_1 _2741_ (.B(_1501_),
    .C(_1502_),
    .A(_1499_),
    .Y(_1503_));
 sg13g2_a21o_1 _2742_ (.A2(_1502_),
    .A1(_1501_),
    .B1(_1499_),
    .X(_1504_));
 sg13g2_and3_1 _2743_ (.X(_1505_),
    .A(_1498_),
    .B(_1503_),
    .C(_1504_));
 sg13g2_a21oi_1 _2744_ (.A1(_1503_),
    .A2(_1504_),
    .Y(_1506_),
    .B1(_1498_));
 sg13g2_or3_1 _2745_ (.A(_1496_),
    .B(_1505_),
    .C(_1506_),
    .X(_1507_));
 sg13g2_o21ai_1 _2746_ (.B1(_1496_),
    .Y(_1508_),
    .A1(_1505_),
    .A2(_1506_));
 sg13g2_nand3_1 _2747_ (.B(_1507_),
    .C(_1508_),
    .A(_1489_),
    .Y(_1509_));
 sg13g2_a21o_1 _2748_ (.A2(_1508_),
    .A1(_1507_),
    .B1(_1489_),
    .X(_1510_));
 sg13g2_nand3_1 _2749_ (.B(_1509_),
    .C(_1510_),
    .A(_1488_),
    .Y(_1511_));
 sg13g2_a21o_1 _2750_ (.A2(_1510_),
    .A1(_1509_),
    .B1(_1488_),
    .X(_1512_));
 sg13g2_and3_1 _2751_ (.X(_1513_),
    .A(_1487_),
    .B(_1511_),
    .C(_1512_));
 sg13g2_nand3_1 _2752_ (.B(_1511_),
    .C(_1512_),
    .A(_1487_),
    .Y(_1514_));
 sg13g2_a21o_1 _2753_ (.A2(_1512_),
    .A1(_1511_),
    .B1(_1487_),
    .X(_1515_));
 sg13g2_nand3_1 _2754_ (.B(_1514_),
    .C(_1515_),
    .A(_1486_),
    .Y(_1516_));
 sg13g2_a21o_1 _2755_ (.A2(_1515_),
    .A1(_1514_),
    .B1(_1486_),
    .X(_1517_));
 sg13g2_nand3_1 _2756_ (.B(_1516_),
    .C(_1517_),
    .A(_1485_),
    .Y(_1518_));
 sg13g2_a21oi_1 _2757_ (.A1(_1516_),
    .A2(_1517_),
    .Y(_1519_),
    .B1(_1485_));
 sg13g2_a21o_1 _2758_ (.A2(_1517_),
    .A1(_1516_),
    .B1(_1484_),
    .X(_1520_));
 sg13g2_nand3_1 _2759_ (.B(_1516_),
    .C(_1517_),
    .A(_1484_),
    .Y(_1521_));
 sg13g2_a21oi_1 _2760_ (.A1(_1520_),
    .A2(_1521_),
    .Y(_1522_),
    .B1(_1483_));
 sg13g2_and3_1 _2761_ (.X(_1523_),
    .A(_1483_),
    .B(_1520_),
    .C(_1521_));
 sg13g2_nor3_1 _2762_ (.A(_1412_),
    .B(_1522_),
    .C(_1523_),
    .Y(_1524_));
 sg13g2_o21ai_1 _2763_ (.B1(_1412_),
    .Y(_1525_),
    .A1(_1522_),
    .A2(_1523_));
 sg13g2_nor2b_1 _2764_ (.A(_1524_),
    .B_N(_1525_),
    .Y(_1526_));
 sg13g2_xnor2_1 _2765_ (.Y(_1527_),
    .A(_1411_),
    .B(_1526_));
 sg13g2_nor2b_1 _2766_ (.A(\i_w_buf[14].A ),
    .B_N(net90),
    .Y(_1528_));
 sg13g2_nand2_1 _2767_ (.Y(_1529_),
    .A(\i_w_buf[15].A ),
    .B(_1528_));
 sg13g2_nand2b_2 _2768_ (.Y(_1530_),
    .B(_1067_),
    .A_N(\i_w_buf[55].A ));
 sg13g2_nand3b_1 _2769_ (.B(\i_w_buf[191].A ),
    .C(net89),
    .Y(_1531_),
    .A_N(\i_w_buf[190].A ));
 sg13g2_nor2b_1 _2770_ (.A(\i_w_buf[90].A ),
    .B_N(net93),
    .Y(_1532_));
 sg13g2_nor2b_1 _2771_ (.A(\i_w_buf[91].A ),
    .B_N(_1532_),
    .Y(_1533_));
 sg13g2_nor2_1 _2772_ (.A(_0864_),
    .B(\i_w_buf[242].A ),
    .Y(_1534_));
 sg13g2_nand2_2 _2773_ (.Y(_1535_),
    .A(\i_w_buf[243].A ),
    .B(_1534_));
 sg13g2_nor3_2 _2774_ (.A(net85),
    .B(\i_w_buf[144].A ),
    .C(\i_w_buf[145].A ),
    .Y(_1536_));
 sg13g2_nand2b_1 _2775_ (.Y(_1537_),
    .B(_1320_),
    .A_N(\i_w_buf[233].A ));
 sg13g2_inv_2 _2776_ (.Y(_1538_),
    .A(_1537_));
 sg13g2_nor3_1 _2777_ (.A(net83),
    .B(\i_w_buf[234].A ),
    .C(\i_w_buf[235].A ),
    .Y(_1539_));
 sg13g2_nor2b_1 _2778_ (.A(\i_w_buf[148].A ),
    .B_N(net100),
    .Y(_1540_));
 sg13g2_and2_2 _2779_ (.A(\i_w_buf[149].A ),
    .B(_1540_),
    .X(_1541_));
 sg13g2_and4_1 _2780_ (.A(_0875_),
    .B(_0876_),
    .C(_1277_),
    .D(_1358_),
    .X(_1542_));
 sg13g2_a22oi_1 _2781_ (.Y(_1543_),
    .B1(_1358_),
    .B2(_0876_),
    .A2(_1277_),
    .A1(_0875_));
 sg13g2_or3_1 _2782_ (.A(_1541_),
    .B(_1542_),
    .C(_1543_),
    .X(_1544_));
 sg13g2_o21ai_1 _2783_ (.B1(_1541_),
    .Y(_1545_),
    .A1(_1542_),
    .A2(_1543_));
 sg13g2_nand3_1 _2784_ (.B(_1544_),
    .C(_1545_),
    .A(_1539_),
    .Y(_1546_));
 sg13g2_a21o_1 _2785_ (.A2(_1545_),
    .A1(_1544_),
    .B1(_1539_),
    .X(_1547_));
 sg13g2_nand3_1 _2786_ (.B(_1546_),
    .C(_1547_),
    .A(_1538_),
    .Y(_1548_));
 sg13g2_a21o_1 _2787_ (.A2(_1547_),
    .A1(_1546_),
    .B1(_1538_),
    .X(_1549_));
 sg13g2_and3_1 _2788_ (.X(_1550_),
    .A(_1536_),
    .B(_1548_),
    .C(_1549_));
 sg13g2_nand3_1 _2789_ (.B(_1548_),
    .C(_1549_),
    .A(_1536_),
    .Y(_1551_));
 sg13g2_a21o_1 _2790_ (.A2(_1549_),
    .A1(_1548_),
    .B1(_1536_),
    .X(_1552_));
 sg13g2_nand3_1 _2791_ (.B(_1551_),
    .C(_1552_),
    .A(_1535_),
    .Y(_1553_));
 sg13g2_a21o_1 _2792_ (.A2(_1552_),
    .A1(_1551_),
    .B1(_1535_),
    .X(_1554_));
 sg13g2_nand3_1 _2793_ (.B(_1553_),
    .C(_1554_),
    .A(_1533_),
    .Y(_1555_));
 sg13g2_a21o_1 _2794_ (.A2(_1554_),
    .A1(_1553_),
    .B1(_1533_),
    .X(_1556_));
 sg13g2_nand2b_1 _2795_ (.Y(_1557_),
    .B(_1071_),
    .A_N(\i_w_buf[225].A ));
 sg13g2_nor3_2 _2796_ (.A(_0864_),
    .B(\i_w_buf[226].A ),
    .C(\i_w_buf[227].A ),
    .Y(_1558_));
 sg13g2_and2_1 _2797_ (.A(\i_w_buf[105].A ),
    .B(_1106_),
    .X(_1559_));
 sg13g2_nand2_1 _2798_ (.Y(_1560_),
    .A(\i_w_buf[105].A ),
    .B(_1106_));
 sg13g2_nand3b_1 _2799_ (.B(\i_w_buf[113].A ),
    .C(net107),
    .Y(_1561_),
    .A_N(\i_w_buf[112].A ));
 sg13g2_and3_1 _2800_ (.X(_1562_),
    .A(_0879_),
    .B(_1418_),
    .C(_1561_));
 sg13g2_nand3_1 _2801_ (.B(_1418_),
    .C(_1561_),
    .A(_0879_),
    .Y(_1563_));
 sg13g2_a21oi_1 _2802_ (.A1(_0879_),
    .A2(_1418_),
    .Y(_1564_),
    .B1(_1561_));
 sg13g2_a21o_1 _2803_ (.A2(_1418_),
    .A1(_0879_),
    .B1(_1561_),
    .X(_1565_));
 sg13g2_nor3_1 _2804_ (.A(_1559_),
    .B(_1562_),
    .C(_1564_),
    .Y(_1566_));
 sg13g2_nand3_1 _2805_ (.B(_1563_),
    .C(_1565_),
    .A(_1560_),
    .Y(_1567_));
 sg13g2_a21oi_1 _2806_ (.A1(_1563_),
    .A2(_1565_),
    .Y(_1568_),
    .B1(_1560_));
 sg13g2_o21ai_1 _2807_ (.B1(_1559_),
    .Y(_1569_),
    .A1(_1562_),
    .A2(_1564_));
 sg13g2_nand3_1 _2808_ (.B(_1567_),
    .C(_1569_),
    .A(_1558_),
    .Y(_1570_));
 sg13g2_a21oi_1 _2809_ (.A1(_1567_),
    .A2(_1569_),
    .Y(_1571_),
    .B1(_1558_));
 sg13g2_nor3_1 _2810_ (.A(_1558_),
    .B(_1566_),
    .C(_1568_),
    .Y(_1572_));
 sg13g2_o21ai_1 _2811_ (.B1(_1558_),
    .Y(_1573_),
    .A1(_1566_),
    .A2(_1568_));
 sg13g2_nor2b_1 _2812_ (.A(_1572_),
    .B_N(_1573_),
    .Y(_1574_));
 sg13g2_xnor2_1 _2813_ (.Y(_1575_),
    .A(_1557_),
    .B(_1574_));
 sg13g2_nor3_1 _2814_ (.A(net87),
    .B(\i_w_buf[140].A ),
    .C(\i_w_buf[141].A ),
    .Y(_1576_));
 sg13g2_nor2_1 _2815_ (.A(net85),
    .B(\i_w_buf[48].A ),
    .Y(_1577_));
 sg13g2_nor3_1 _2816_ (.A(net85),
    .B(\i_w_buf[48].A ),
    .C(\i_w_buf[49].A ),
    .Y(_1578_));
 sg13g2_nor3_1 _2817_ (.A(net84),
    .B(\i_w_buf[42].A ),
    .C(\i_w_buf[43].A ),
    .Y(_1579_));
 sg13g2_nand2_1 _2818_ (.Y(_1580_),
    .A(\i_w_buf[135].A ),
    .B(_1438_));
 sg13g2_and2_1 _2819_ (.A(_1579_),
    .B(_1580_),
    .X(_1581_));
 sg13g2_xor2_1 _2820_ (.B(_1580_),
    .A(_1579_),
    .X(_1582_));
 sg13g2_xnor2_1 _2821_ (.Y(_1583_),
    .A(_1578_),
    .B(_1582_));
 sg13g2_nand3b_1 _2822_ (.B(\i_w_buf[209].A ),
    .C(net107),
    .Y(_1584_),
    .A_N(\i_w_buf[208].A ));
 sg13g2_or3_1 _2823_ (.A(\i_w_buf[40].A ),
    .B(\i_w_buf[41].A ),
    .C(_0863_),
    .X(_1585_));
 sg13g2_nor2b_1 _2824_ (.A(\i_w_buf[36].A ),
    .B_N(net100),
    .Y(_1586_));
 sg13g2_and4_2 _2825_ (.A(_0877_),
    .B(_0878_),
    .C(_0902_),
    .D(_1586_),
    .X(_1587_));
 sg13g2_a22oi_1 _2826_ (.Y(_0000_),
    .B1(_1586_),
    .B2(_0878_),
    .A2(_0902_),
    .A1(_0877_));
 sg13g2_or3_2 _2827_ (.A(_1585_),
    .B(_1587_),
    .C(_0000_),
    .X(_0001_));
 sg13g2_inv_1 _2828_ (.Y(_0002_),
    .A(_0001_));
 sg13g2_o21ai_1 _2829_ (.B1(_1585_),
    .Y(_0003_),
    .A1(_1587_),
    .A2(_0000_));
 sg13g2_and3_1 _2830_ (.X(_0004_),
    .A(_1584_),
    .B(_0001_),
    .C(_0003_));
 sg13g2_nand3_1 _2831_ (.B(_0001_),
    .C(_0003_),
    .A(_1584_),
    .Y(_0005_));
 sg13g2_a21oi_1 _2832_ (.A1(_0001_),
    .A2(_0003_),
    .Y(_0006_),
    .B1(_1584_));
 sg13g2_or3_1 _2833_ (.A(_1583_),
    .B(_0004_),
    .C(_0006_),
    .X(_0007_));
 sg13g2_o21ai_1 _2834_ (.B1(_1583_),
    .Y(_0008_),
    .A1(_0004_),
    .A2(_0006_));
 sg13g2_and3_1 _2835_ (.X(_0009_),
    .A(_1576_),
    .B(_0007_),
    .C(_0008_));
 sg13g2_nand3_1 _2836_ (.B(_0007_),
    .C(_0008_),
    .A(_1576_),
    .Y(_0010_));
 sg13g2_a21oi_1 _2837_ (.A1(_0007_),
    .A2(_0008_),
    .Y(_0011_),
    .B1(_1576_));
 sg13g2_nor2_1 _2838_ (.A(_0009_),
    .B(_0011_),
    .Y(_0012_));
 sg13g2_xnor2_1 _2839_ (.Y(_0013_),
    .A(_1575_),
    .B(_0012_));
 sg13g2_nand3_1 _2840_ (.B(_1556_),
    .C(_0013_),
    .A(_1555_),
    .Y(_0014_));
 sg13g2_a21o_1 _2841_ (.A2(_1556_),
    .A1(_1555_),
    .B1(_0013_),
    .X(_0015_));
 sg13g2_nand3_1 _2842_ (.B(_0014_),
    .C(_0015_),
    .A(_1531_),
    .Y(_0016_));
 sg13g2_a21oi_1 _2843_ (.A1(_0014_),
    .A2(_0015_),
    .Y(_0017_),
    .B1(_1531_));
 sg13g2_a21o_1 _2844_ (.A2(_0015_),
    .A1(_0014_),
    .B1(_1531_),
    .X(_0018_));
 sg13g2_nand2_1 _2845_ (.Y(_0019_),
    .A(_0016_),
    .B(_0018_));
 sg13g2_xnor2_1 _2846_ (.Y(_0020_),
    .A(_1530_),
    .B(_0019_));
 sg13g2_nand3b_1 _2847_ (.B(\i_w_buf[153].A ),
    .C(net2),
    .Y(_0021_),
    .A_N(\i_w_buf[152].A ));
 sg13g2_nand3b_1 _2848_ (.B(\i_w_buf[123].A ),
    .C(net94),
    .Y(_0022_),
    .A_N(\i_w_buf[122].A ));
 sg13g2_inv_1 _2849_ (.Y(_0023_),
    .A(_0022_));
 sg13g2_nor3_2 _2850_ (.A(net81),
    .B(\i_w_buf[94].A ),
    .C(\i_w_buf[95].A ),
    .Y(_0024_));
 sg13g2_nand3b_1 _2851_ (.B(\i_w_buf[163].A ),
    .C(net103),
    .Y(_0025_),
    .A_N(\i_w_buf[162].A ));
 sg13g2_nor3_2 _2852_ (.A(_0864_),
    .B(\i_w_buf[18].A ),
    .C(\i_w_buf[19].A ),
    .Y(_0026_));
 sg13g2_nor2b_2 _2853_ (.A(\i_w_buf[21].A ),
    .B_N(_1415_),
    .Y(_0027_));
 sg13g2_and2_1 _2854_ (.A(_0026_),
    .B(_0027_),
    .X(_0028_));
 sg13g2_or2_1 _2855_ (.X(_0029_),
    .B(_0027_),
    .A(_0026_));
 sg13g2_xor2_1 _2856_ (.B(_0027_),
    .A(_0026_),
    .X(_0030_));
 sg13g2_xnor2_1 _2857_ (.Y(_0031_),
    .A(_0025_),
    .B(_0030_));
 sg13g2_nand2_2 _2858_ (.Y(_0032_),
    .A(\i_w_buf[197].A ),
    .B(_1272_));
 sg13g2_nand2_1 _2859_ (.Y(_0033_),
    .A(\i_w_buf[91].A ),
    .B(_1532_));
 sg13g2_nand3b_1 _2860_ (.B(\i_w_buf[237].A ),
    .C(net91),
    .Y(_0034_),
    .A_N(\i_w_buf[236].A ));
 sg13g2_nand3_1 _2861_ (.B(_1528_),
    .C(_0034_),
    .A(_0874_),
    .Y(_0035_));
 sg13g2_a21o_1 _2862_ (.A2(_1528_),
    .A1(_0874_),
    .B1(_0034_),
    .X(_0036_));
 sg13g2_nand3_1 _2863_ (.B(_0035_),
    .C(_0036_),
    .A(_0033_),
    .Y(_0037_));
 sg13g2_a21o_1 _2864_ (.A2(_0036_),
    .A1(_0035_),
    .B1(_0033_),
    .X(_0038_));
 sg13g2_nand3_1 _2865_ (.B(_0037_),
    .C(_0038_),
    .A(_0032_),
    .Y(_0039_));
 sg13g2_a21oi_1 _2866_ (.A1(_0037_),
    .A2(_0038_),
    .Y(_0040_),
    .B1(_0032_));
 sg13g2_a21o_1 _2867_ (.A2(_0038_),
    .A1(_0037_),
    .B1(_0032_),
    .X(_0041_));
 sg13g2_nand2_1 _2868_ (.Y(_0042_),
    .A(_0039_),
    .B(_0041_));
 sg13g2_xnor2_1 _2869_ (.Y(_0043_),
    .A(_0031_),
    .B(_0042_));
 sg13g2_nand2b_1 _2870_ (.Y(_0044_),
    .B(net102),
    .A_N(\i_w_buf[244].A ));
 sg13g2_nand3b_1 _2871_ (.B(\i_w_buf[245].A ),
    .C(net102),
    .Y(_0045_),
    .A_N(\i_w_buf[244].A ));
 sg13g2_nand2_2 _2872_ (.Y(_0046_),
    .A(\i_w_buf[195].A ),
    .B(_1141_));
 sg13g2_nand2b_1 _2873_ (.Y(_0047_),
    .B(_1534_),
    .A_N(\i_w_buf[243].A ));
 sg13g2_and2_1 _2874_ (.A(_0871_),
    .B(_1497_),
    .X(_0048_));
 sg13g2_nand3b_1 _2875_ (.B(\i_w_buf[159].A ),
    .C(net90),
    .Y(_0049_),
    .A_N(\i_w_buf[158].A ));
 sg13g2_nand3_1 _2876_ (.B(_1497_),
    .C(_0049_),
    .A(_0871_),
    .Y(_0050_));
 sg13g2_a21o_1 _2877_ (.A2(_1497_),
    .A1(_0871_),
    .B1(_0049_),
    .X(_0051_));
 sg13g2_and4_2 _2878_ (.A(_0873_),
    .B(_1347_),
    .C(_0050_),
    .D(_0051_),
    .X(_0052_));
 sg13g2_a22oi_1 _2879_ (.Y(_0053_),
    .B1(_0050_),
    .B2(_0051_),
    .A2(_1347_),
    .A1(_0873_));
 sg13g2_nor3_1 _2880_ (.A(_0047_),
    .B(_0052_),
    .C(_0053_),
    .Y(_0054_));
 sg13g2_or3_1 _2881_ (.A(_0047_),
    .B(_0052_),
    .C(_0053_),
    .X(_0055_));
 sg13g2_o21ai_1 _2882_ (.B1(_0047_),
    .Y(_0056_),
    .A1(_0052_),
    .A2(_0053_));
 sg13g2_nand3_1 _2883_ (.B(_0055_),
    .C(_0056_),
    .A(_0046_),
    .Y(_0057_));
 sg13g2_a21o_1 _2884_ (.A2(_0056_),
    .A1(_0055_),
    .B1(_0046_),
    .X(_0058_));
 sg13g2_and3_1 _2885_ (.X(_0059_),
    .A(_0045_),
    .B(_0057_),
    .C(_0058_));
 sg13g2_a21oi_1 _2886_ (.A1(_0057_),
    .A2(_0058_),
    .Y(_0060_),
    .B1(_0045_));
 sg13g2_or3_1 _2887_ (.A(_0043_),
    .B(_0059_),
    .C(_0060_),
    .X(_0061_));
 sg13g2_o21ai_1 _2888_ (.B1(_0043_),
    .Y(_0062_),
    .A1(_0059_),
    .A2(_0060_));
 sg13g2_nand2_1 _2889_ (.Y(_0063_),
    .A(_0061_),
    .B(_0062_));
 sg13g2_nand3_1 _2890_ (.B(_0061_),
    .C(_0062_),
    .A(_0024_),
    .Y(_0064_));
 sg13g2_a21oi_1 _2891_ (.A1(_0061_),
    .A2(_0062_),
    .Y(_0065_),
    .B1(_0024_));
 sg13g2_xnor2_1 _2892_ (.Y(_0066_),
    .A(_0024_),
    .B(_0063_));
 sg13g2_xnor2_1 _2893_ (.Y(_0067_),
    .A(_0022_),
    .B(_0066_));
 sg13g2_nor3_2 _2894_ (.A(net83),
    .B(\i_w_buf[58].A ),
    .C(\i_w_buf[59].A ),
    .Y(_0068_));
 sg13g2_nor2b_1 _2895_ (.A(\i_w_buf[149].A ),
    .B_N(_1540_),
    .Y(_0069_));
 sg13g2_nand3b_1 _2896_ (.B(\i_w_buf[249].A ),
    .C(net97),
    .Y(_0070_),
    .A_N(\i_w_buf[248].A ));
 sg13g2_nand3b_1 _2897_ (.B(\i_w_buf[223].A ),
    .C(net89),
    .Y(_0071_),
    .A_N(\i_w_buf[222].A ));
 sg13g2_nor3_2 _2898_ (.A(net86),
    .B(\i_w_buf[0].A ),
    .C(\i_w_buf[1].A ),
    .Y(_0072_));
 sg13g2_nor2b_2 _2899_ (.A(\i_w_buf[3].A ),
    .B_N(_0898_),
    .Y(_0073_));
 sg13g2_and2_1 _2900_ (.A(_0072_),
    .B(_0073_),
    .X(_0074_));
 sg13g2_or2_1 _2901_ (.X(_0075_),
    .B(_0073_),
    .A(_0072_));
 sg13g2_xor2_1 _2902_ (.B(_0073_),
    .A(_0072_),
    .X(_0076_));
 sg13g2_xnor2_1 _2903_ (.Y(_0077_),
    .A(_0071_),
    .B(_0076_));
 sg13g2_nor2_1 _2904_ (.A(\i_w_buf[245].A ),
    .B(_0044_),
    .Y(_0078_));
 sg13g2_nand3b_1 _2905_ (.B(\i_w_buf[1].A ),
    .C(net106),
    .Y(_0079_),
    .A_N(\i_w_buf[0].A ));
 sg13g2_nand3b_1 _2906_ (.B(\i_w_buf[17].A ),
    .C(net106),
    .Y(_0080_),
    .A_N(\i_w_buf[16].A ));
 sg13g2_nand3b_1 _2907_ (.B(\i_w_buf[65].A ),
    .C(net106),
    .Y(_0081_),
    .A_N(\i_w_buf[64].A ));
 sg13g2_and2_1 _2908_ (.A(_0080_),
    .B(_0081_),
    .X(_0082_));
 sg13g2_xor2_1 _2909_ (.B(_0081_),
    .A(_0080_),
    .X(_0083_));
 sg13g2_xnor2_1 _2910_ (.Y(_0084_),
    .A(_0079_),
    .B(_0083_));
 sg13g2_or3_1 _2911_ (.A(\i_w_buf[245].A ),
    .B(_0044_),
    .C(_0084_),
    .X(_0085_));
 sg13g2_xor2_1 _2912_ (.B(_0084_),
    .A(_0078_),
    .X(_0086_));
 sg13g2_xor2_1 _2913_ (.B(_0086_),
    .A(_0077_),
    .X(_0087_));
 sg13g2_and2_1 _2914_ (.A(_0070_),
    .B(_0087_),
    .X(_0088_));
 sg13g2_xor2_1 _2915_ (.B(_0087_),
    .A(_0070_),
    .X(_0089_));
 sg13g2_xnor2_1 _2916_ (.Y(_0090_),
    .A(_0069_),
    .B(_0089_));
 sg13g2_nand2_2 _2917_ (.Y(_0091_),
    .A(\i_w_buf[125].A ),
    .B(_1323_));
 sg13g2_nand2_2 _2918_ (.Y(_0092_),
    .A(\i_w_buf[169].A ),
    .B(_0974_));
 sg13g2_nor2_1 _2919_ (.A(\i_w_buf[251].A ),
    .B(_1162_),
    .Y(_0093_));
 sg13g2_nand3b_1 _2920_ (.B(\i_w_buf[5].A ),
    .C(net100),
    .Y(_0094_),
    .A_N(\i_w_buf[4].A ));
 sg13g2_nand3b_1 _2921_ (.B(\i_w_buf[145].A ),
    .C(net107),
    .Y(_0095_),
    .A_N(\i_w_buf[144].A ));
 sg13g2_nand3b_1 _2922_ (.B(\i_w_buf[193].A ),
    .C(net107),
    .Y(_0096_),
    .A_N(\i_w_buf[192].A ));
 sg13g2_and2_1 _2923_ (.A(_0095_),
    .B(_0096_),
    .X(_0097_));
 sg13g2_xor2_1 _2924_ (.B(_0096_),
    .A(_0095_),
    .X(_0098_));
 sg13g2_xnor2_1 _2925_ (.Y(_0099_),
    .A(_0094_),
    .B(_0098_));
 sg13g2_nor3_1 _2926_ (.A(\i_w_buf[251].A ),
    .B(_1162_),
    .C(_0099_),
    .Y(_0100_));
 sg13g2_xnor2_1 _2927_ (.Y(_0101_),
    .A(_0093_),
    .B(_0099_));
 sg13g2_xnor2_1 _2928_ (.Y(_0102_),
    .A(_0092_),
    .B(_0101_));
 sg13g2_nor3_2 _2929_ (.A(_0863_),
    .B(\i_w_buf[152].A ),
    .C(\i_w_buf[153].A ),
    .Y(_0103_));
 sg13g2_nand2_2 _2930_ (.Y(_0104_),
    .A(\i_w_buf[133].A ),
    .B(_1304_));
 sg13g2_nand3b_1 _2931_ (.B(\i_w_buf[73].A ),
    .C(net97),
    .Y(_0105_),
    .A_N(\i_w_buf[72].A ));
 sg13g2_nand2_2 _2932_ (.Y(_0106_),
    .A(\i_w_buf[97].A ),
    .B(_1378_));
 sg13g2_and2_1 _2933_ (.A(_0105_),
    .B(_0106_),
    .X(_0107_));
 sg13g2_xor2_1 _2934_ (.B(_0106_),
    .A(_0105_),
    .X(_0108_));
 sg13g2_xnor2_1 _2935_ (.Y(_0109_),
    .A(_0104_),
    .B(_0108_));
 sg13g2_nor2_1 _2936_ (.A(\i_w_buf[253].A ),
    .B(_1218_),
    .Y(_0110_));
 sg13g2_nand2_1 _2937_ (.Y(_0111_),
    .A(\i_w_buf[67].A ),
    .B(_1490_));
 sg13g2_nand3b_1 _2938_ (.B(\i_w_buf[37].A ),
    .C(net100),
    .Y(_0112_),
    .A_N(\i_w_buf[36].A ));
 sg13g2_nand3b_1 _2939_ (.B(\i_w_buf[41].A ),
    .C(net97),
    .Y(_0113_),
    .A_N(\i_w_buf[40].A ));
 sg13g2_and2_1 _2940_ (.A(_0112_),
    .B(_0113_),
    .X(_0114_));
 sg13g2_xor2_1 _2941_ (.B(_0113_),
    .A(_0112_),
    .X(_0115_));
 sg13g2_xnor2_1 _2942_ (.Y(_0116_),
    .A(_0111_),
    .B(_0115_));
 sg13g2_or3_1 _2943_ (.A(\i_w_buf[253].A ),
    .B(_1218_),
    .C(_0116_),
    .X(_0117_));
 sg13g2_xor2_1 _2944_ (.B(_0116_),
    .A(_0110_),
    .X(_0118_));
 sg13g2_xor2_1 _2945_ (.B(_0118_),
    .A(_0109_),
    .X(_0119_));
 sg13g2_nand2_1 _2946_ (.Y(_0120_),
    .A(_0103_),
    .B(_0119_));
 sg13g2_xnor2_1 _2947_ (.Y(_0121_),
    .A(_0103_),
    .B(_0119_));
 sg13g2_xor2_1 _2948_ (.B(_0121_),
    .A(_0102_),
    .X(_0122_));
 sg13g2_nand2_1 _2949_ (.Y(_0123_),
    .A(_0091_),
    .B(_0122_));
 sg13g2_xnor2_1 _2950_ (.Y(_0124_),
    .A(_0091_),
    .B(_0122_));
 sg13g2_xor2_1 _2951_ (.B(_0124_),
    .A(_0090_),
    .X(_0125_));
 sg13g2_nand2_1 _2952_ (.Y(_0126_),
    .A(_0068_),
    .B(_0125_));
 sg13g2_xnor2_1 _2953_ (.Y(_0127_),
    .A(_0068_),
    .B(_0125_));
 sg13g2_xor2_1 _2954_ (.B(_0127_),
    .A(_0067_),
    .X(_0128_));
 sg13g2_nand2_1 _2955_ (.Y(_0129_),
    .A(_0021_),
    .B(_0128_));
 sg13g2_xnor2_1 _2956_ (.Y(_0130_),
    .A(_0021_),
    .B(_0128_));
 sg13g2_xor2_1 _2957_ (.B(_0130_),
    .A(_0020_),
    .X(_0131_));
 sg13g2_nand2_1 _2958_ (.Y(_0132_),
    .A(_1529_),
    .B(_0131_));
 sg13g2_xnor2_1 _2959_ (.Y(_0133_),
    .A(_1529_),
    .B(_0131_));
 sg13g2_xor2_1 _2960_ (.B(_0133_),
    .A(_1527_),
    .X(_0134_));
 sg13g2_nand2_1 _2961_ (.Y(_0135_),
    .A(_1410_),
    .B(_0134_));
 sg13g2_xnor2_1 _2962_ (.Y(_0136_),
    .A(_1410_),
    .B(_0134_));
 sg13g2_xor2_1 _2963_ (.B(_0136_),
    .A(_1409_),
    .X(_0137_));
 sg13g2_nand2_1 _2964_ (.Y(_0138_),
    .A(_1214_),
    .B(_0137_));
 sg13g2_xnor2_1 _2965_ (.Y(_0139_),
    .A(_1214_),
    .B(_0137_));
 sg13g2_xor2_1 _2966_ (.B(_0139_),
    .A(_1213_),
    .X(_0140_));
 sg13g2_nand2_1 _2967_ (.Y(_0141_),
    .A(_0956_),
    .B(_0140_));
 sg13g2_xnor2_1 _2968_ (.Y(_0142_),
    .A(_0956_),
    .B(_0140_));
 sg13g2_xor2_1 _2969_ (.B(_0142_),
    .A(_0955_),
    .X(_0143_));
 sg13g2_and2_1 _2970_ (.A(_0897_),
    .B(_0143_),
    .X(_0144_));
 sg13g2_xor2_1 _2971_ (.B(_0143_),
    .A(_0897_),
    .X(_0145_));
 sg13g2_xnor2_1 _2972_ (.Y(_0146_),
    .A(_0896_),
    .B(_0145_));
 sg13g2_nand2_2 _2973_ (.Y(_0147_),
    .A(\i_w_buf[49].A ),
    .B(_1577_));
 sg13g2_nor2b_1 _2974_ (.A(_0146_),
    .B_N(_0147_),
    .Y(_0148_));
 sg13g2_xnor2_1 _2975_ (.Y(uo_out[0]),
    .A(_0146_),
    .B(_0147_));
 sg13g2_a21oi_1 _2976_ (.A1(_0896_),
    .A2(_0145_),
    .Y(_0149_),
    .B1(_0144_));
 sg13g2_nor2_1 _2977_ (.A(_0952_),
    .B(_0954_),
    .Y(_0150_));
 sg13g2_o21ai_1 _2978_ (.B1(_0141_),
    .Y(_0151_),
    .A1(_0955_),
    .A2(_0142_));
 sg13g2_o21ai_1 _2979_ (.B1(_0950_),
    .Y(_0152_),
    .A1(_0905_),
    .A2(_0948_));
 sg13g2_o21ai_1 _2980_ (.B1(_1211_),
    .Y(_0153_),
    .A1(_0958_),
    .A2(_1212_));
 sg13g2_or2_1 _2981_ (.X(_0154_),
    .B(_0947_),
    .A(_0944_));
 sg13g2_inv_1 _2982_ (.Y(_0155_),
    .A(_0154_));
 sg13g2_o21ai_1 _2983_ (.B1(_1206_),
    .Y(_0156_),
    .A1(_1090_),
    .A2(_1207_));
 sg13g2_a21o_1 _2984_ (.A2(_0940_),
    .A1(_0912_),
    .B1(_0942_),
    .X(_0157_));
 sg13g2_a21oi_1 _2985_ (.A1(_1052_),
    .A2(_1088_),
    .Y(_0158_),
    .B1(_1087_));
 sg13g2_a21o_1 _2986_ (.A2(_0938_),
    .A1(_0933_),
    .B1(_0937_),
    .X(_0159_));
 sg13g2_inv_1 _2987_ (.Y(_0160_),
    .A(_0159_));
 sg13g2_o21ai_1 _2988_ (.B1(_0930_),
    .Y(_0161_),
    .A1(_0931_),
    .A2(_0939_));
 sg13g2_o21ai_1 _2989_ (.B1(_0927_),
    .Y(_0162_),
    .A1(_0916_),
    .A2(_0928_));
 sg13g2_inv_1 _2990_ (.Y(_0163_),
    .A(_0162_));
 sg13g2_o21ai_1 _2991_ (.B1(_1064_),
    .Y(_0164_),
    .A1(_1061_),
    .A2(_1065_));
 sg13g2_a21o_1 _2992_ (.A2(_0925_),
    .A1(_0920_),
    .B1(_0924_),
    .X(_0165_));
 sg13g2_nor2_2 _2993_ (.A(_0164_),
    .B(_0165_),
    .Y(_0166_));
 sg13g2_xor2_1 _2994_ (.B(_0165_),
    .A(_0164_),
    .X(_0167_));
 sg13g2_xnor2_1 _2995_ (.Y(_0168_),
    .A(_0162_),
    .B(_0167_));
 sg13g2_nand2_1 _2996_ (.Y(_0169_),
    .A(_0161_),
    .B(_0168_));
 sg13g2_xnor2_1 _2997_ (.Y(_0170_),
    .A(_0161_),
    .B(_0168_));
 sg13g2_xnor2_1 _2998_ (.Y(_0171_),
    .A(_0160_),
    .B(_0170_));
 sg13g2_nor2_1 _2999_ (.A(_0158_),
    .B(_0171_),
    .Y(_0172_));
 sg13g2_xor2_1 _3000_ (.B(_0171_),
    .A(_0158_),
    .X(_0173_));
 sg13g2_xnor2_1 _3001_ (.Y(_0174_),
    .A(_0157_),
    .B(_0173_));
 sg13g2_nand2b_1 _3002_ (.Y(_0175_),
    .B(_0156_),
    .A_N(_0174_));
 sg13g2_xor2_1 _3003_ (.B(_0174_),
    .A(_0156_),
    .X(_0176_));
 sg13g2_xnor2_1 _3004_ (.Y(_0177_),
    .A(_0155_),
    .B(_0176_));
 sg13g2_nand2b_1 _3005_ (.Y(_0178_),
    .B(_0153_),
    .A_N(_0177_));
 sg13g2_xor2_1 _3006_ (.B(_0177_),
    .A(_0153_),
    .X(_0179_));
 sg13g2_nand2b_1 _3007_ (.Y(_0180_),
    .B(_0152_),
    .A_N(_0179_));
 sg13g2_xor2_1 _3008_ (.B(_0179_),
    .A(_0152_),
    .X(_0181_));
 sg13g2_o21ai_1 _3009_ (.B1(_0138_),
    .Y(_0182_),
    .A1(_1213_),
    .A2(_0139_));
 sg13g2_nand2b_1 _3010_ (.Y(_0183_),
    .B(_1209_),
    .A_N(_1050_));
 sg13g2_a21oi_2 _3011_ (.B1(_1407_),
    .Y(_0184_),
    .A2(_1408_),
    .A1(_1216_));
 sg13g2_nand2b_2 _3012_ (.Y(_0185_),
    .B(_1085_),
    .A_N(_1083_));
 sg13g2_inv_1 _3013_ (.Y(_0186_),
    .A(_0185_));
 sg13g2_o21ai_1 _3014_ (.B1(_1155_),
    .Y(_0187_),
    .A1(_1132_),
    .A2(_1156_));
 sg13g2_a21o_1 _3015_ (.A2(_1079_),
    .A1(_1060_),
    .B1(_1081_),
    .X(_0188_));
 sg13g2_o21ai_1 _3016_ (.B1(_1129_),
    .Y(_0189_),
    .A1(_1105_),
    .A2(_1130_));
 sg13g2_inv_1 _3017_ (.Y(_0190_),
    .A(_0189_));
 sg13g2_o21ai_1 _3018_ (.B1(_1077_),
    .Y(_0191_),
    .A1(_1066_),
    .A2(_1078_));
 sg13g2_o21ai_1 _3019_ (.B1(_1074_),
    .Y(_0192_),
    .A1(_1070_),
    .A2(_1075_));
 sg13g2_o21ai_1 _3020_ (.B1(_0192_),
    .Y(_0193_),
    .A1(_1101_),
    .A2(_1103_));
 sg13g2_inv_1 _3021_ (.Y(_0194_),
    .A(_0193_));
 sg13g2_or3_1 _3022_ (.A(_1101_),
    .B(_1103_),
    .C(_0192_),
    .X(_0195_));
 sg13g2_and2_1 _3023_ (.A(_0193_),
    .B(_0195_),
    .X(_0196_));
 sg13g2_xnor2_1 _3024_ (.Y(_0197_),
    .A(_0191_),
    .B(_0196_));
 sg13g2_xnor2_1 _3025_ (.Y(_0198_),
    .A(_0190_),
    .B(_0197_));
 sg13g2_nand2b_1 _3026_ (.Y(_0199_),
    .B(_0188_),
    .A_N(_0198_));
 sg13g2_xor2_1 _3027_ (.B(_0198_),
    .A(_0188_),
    .X(_0200_));
 sg13g2_nand2b_1 _3028_ (.Y(_0201_),
    .B(_0187_),
    .A_N(_0200_));
 sg13g2_xor2_1 _3029_ (.B(_0200_),
    .A(_0187_),
    .X(_0202_));
 sg13g2_xor2_1 _3030_ (.B(_0202_),
    .A(_0185_),
    .X(_0203_));
 sg13g2_o21ai_1 _3031_ (.B1(_1203_),
    .Y(_0204_),
    .A1(_1157_),
    .A2(_1204_));
 sg13g2_a21o_1 _3032_ (.A2(_1124_),
    .A1(_1119_),
    .B1(_1123_),
    .X(_0205_));
 sg13g2_o21ai_1 _3033_ (.B1(_1126_),
    .Y(_0206_),
    .A1(_1115_),
    .A2(_1127_));
 sg13g2_nand2_1 _3034_ (.Y(_0207_),
    .A(_0205_),
    .B(_0206_));
 sg13g2_nor2_1 _3035_ (.A(_0205_),
    .B(_0206_),
    .Y(_0208_));
 sg13g2_xor2_1 _3036_ (.B(_0206_),
    .A(_0205_),
    .X(_0209_));
 sg13g2_a21oi_1 _3037_ (.A1(_1110_),
    .A2(_1111_),
    .Y(_0210_),
    .B1(_1113_));
 sg13g2_a21oi_2 _3038_ (.B1(_1099_),
    .Y(_0211_),
    .A2(_1097_),
    .A1(_1096_));
 sg13g2_and2_1 _3039_ (.A(_0210_),
    .B(_0211_),
    .X(_0212_));
 sg13g2_xnor2_1 _3040_ (.Y(_0213_),
    .A(_0210_),
    .B(_0211_));
 sg13g2_nand2_1 _3041_ (.Y(_0214_),
    .A(_0209_),
    .B(_0213_));
 sg13g2_xor2_1 _3042_ (.B(_0213_),
    .A(_0209_),
    .X(_0215_));
 sg13g2_o21ai_1 _3043_ (.B1(_1152_),
    .Y(_0216_),
    .A1(_1135_),
    .A2(_1153_));
 sg13g2_or2_2 _3044_ (.X(_0217_),
    .B(_1150_),
    .A(_1148_));
 sg13g2_o21ai_1 _3045_ (.B1(_1179_),
    .Y(_0218_),
    .A1(_1169_),
    .A2(_1180_));
 sg13g2_a21o_1 _3046_ (.A2(_1166_),
    .A1(_1165_),
    .B1(_1168_),
    .X(_0219_));
 sg13g2_a21o_2 _3047_ (.A2(_1146_),
    .A1(_1140_),
    .B1(_1145_),
    .X(_0220_));
 sg13g2_nor2_1 _3048_ (.A(_0219_),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_xor2_1 _3049_ (.B(_0220_),
    .A(_0219_),
    .X(_0222_));
 sg13g2_inv_1 _3050_ (.Y(_0223_),
    .A(_0222_));
 sg13g2_xnor2_1 _3051_ (.Y(_0224_),
    .A(_0218_),
    .B(_0222_));
 sg13g2_and2_1 _3052_ (.A(_0217_),
    .B(_0224_),
    .X(_0225_));
 sg13g2_xnor2_1 _3053_ (.Y(_0226_),
    .A(_0217_),
    .B(_0224_));
 sg13g2_nor2b_1 _3054_ (.A(_0226_),
    .B_N(_0216_),
    .Y(_0227_));
 sg13g2_xor2_1 _3055_ (.B(_0226_),
    .A(_0216_),
    .X(_0228_));
 sg13g2_inv_1 _3056_ (.Y(_0229_),
    .A(_0228_));
 sg13g2_xor2_1 _3057_ (.B(_0228_),
    .A(_0215_),
    .X(_0230_));
 sg13g2_a21o_1 _3058_ (.A2(_1200_),
    .A1(_1160_),
    .B1(_1199_),
    .X(_0231_));
 sg13g2_o21ai_1 _3059_ (.B1(_1196_),
    .Y(_0232_),
    .A1(_1181_),
    .A2(_1197_));
 sg13g2_o21ai_1 _3060_ (.B1(_0989_),
    .Y(_0233_),
    .A1(_0966_),
    .A2(_0990_));
 sg13g2_a21o_1 _3061_ (.A2(_1177_),
    .A1(_1173_),
    .B1(_1176_),
    .X(_0234_));
 sg13g2_o21ai_1 _3062_ (.B1(_1192_),
    .Y(_0235_),
    .A1(_1183_),
    .A2(_1193_));
 sg13g2_mux2_2 _3063_ (.A0(_0970_),
    .A1(_0894_),
    .S(_0968_),
    .X(_0236_));
 sg13g2_nand2_1 _3064_ (.Y(_0237_),
    .A(_1187_),
    .B(_1189_));
 sg13g2_or2_1 _3065_ (.X(_0238_),
    .B(_0237_),
    .A(_0236_));
 sg13g2_xnor2_1 _3066_ (.Y(_0239_),
    .A(_0236_),
    .B(_0237_));
 sg13g2_and2_1 _3067_ (.A(_0235_),
    .B(_0239_),
    .X(_0240_));
 sg13g2_xor2_1 _3068_ (.B(_0239_),
    .A(_0235_),
    .X(_0241_));
 sg13g2_xnor2_1 _3069_ (.Y(_0242_),
    .A(_0234_),
    .B(_0241_));
 sg13g2_nor2b_1 _3070_ (.A(_0242_),
    .B_N(_0233_),
    .Y(_0243_));
 sg13g2_xnor2_1 _3071_ (.Y(_0244_),
    .A(_0233_),
    .B(_0242_));
 sg13g2_xnor2_1 _3072_ (.Y(_0245_),
    .A(_0232_),
    .B(_0244_));
 sg13g2_inv_1 _3073_ (.Y(_0246_),
    .A(_0245_));
 sg13g2_nand2_1 _3074_ (.Y(_0247_),
    .A(_0231_),
    .B(_0246_));
 sg13g2_xnor2_1 _3075_ (.Y(_0248_),
    .A(_0231_),
    .B(_0246_));
 sg13g2_xor2_1 _3076_ (.B(_0248_),
    .A(_0230_),
    .X(_0249_));
 sg13g2_nand2_1 _3077_ (.Y(_0250_),
    .A(_0204_),
    .B(_0249_));
 sg13g2_xnor2_1 _3078_ (.Y(_0251_),
    .A(_0204_),
    .B(_0249_));
 sg13g2_xor2_1 _3079_ (.B(_0251_),
    .A(_0203_),
    .X(_0252_));
 sg13g2_a21oi_2 _3080_ (.B1(_1046_),
    .Y(_0253_),
    .A2(_1047_),
    .A1(_0962_));
 sg13g2_o21ai_1 _3081_ (.B1(_1043_),
    .Y(_0254_),
    .A1(_0964_),
    .A2(_1044_));
 sg13g2_o21ai_1 _3082_ (.B1(_1341_),
    .Y(_0255_),
    .A1(_1254_),
    .A2(_1342_));
 sg13g2_o21ai_1 _3083_ (.B1(_1040_),
    .Y(_0256_),
    .A1(_0994_),
    .A2(_1041_));
 sg13g2_o21ai_1 _3084_ (.B1(_1249_),
    .Y(_0257_),
    .A1(_1220_),
    .A2(_1250_));
 sg13g2_nand2_1 _3085_ (.Y(_0258_),
    .A(_0982_),
    .B(_0986_));
 sg13g2_o21ai_1 _3086_ (.B1(_1007_),
    .Y(_0259_),
    .A1(_0997_),
    .A2(_1008_));
 sg13g2_nand2_1 _3087_ (.Y(_0260_),
    .A(_0977_),
    .B(_0979_));
 sg13g2_and2_1 _3088_ (.A(_0259_),
    .B(_0260_),
    .X(_0261_));
 sg13g2_xor2_1 _3089_ (.B(_0260_),
    .A(_0259_),
    .X(_0262_));
 sg13g2_xnor2_1 _3090_ (.Y(_0263_),
    .A(_0258_),
    .B(_0262_));
 sg13g2_o21ai_1 _3091_ (.B1(_1036_),
    .Y(_0264_),
    .A1(_1011_),
    .A2(_1037_));
 sg13g2_nand2_2 _3092_ (.Y(_0265_),
    .A(_1026_),
    .B(_1028_));
 sg13g2_o21ai_1 _3093_ (.B1(_1031_),
    .Y(_0266_),
    .A1(_1019_),
    .A2(_1032_));
 sg13g2_nand2_1 _3094_ (.Y(_0267_),
    .A(_0265_),
    .B(_0266_));
 sg13g2_xor2_1 _3095_ (.B(_0266_),
    .A(_0265_),
    .X(_0268_));
 sg13g2_nor2b_1 _3096_ (.A(_1003_),
    .B_N(_1005_),
    .Y(_0269_));
 sg13g2_and3_1 _3097_ (.X(_0270_),
    .A(_1016_),
    .B(_1018_),
    .C(_0269_));
 sg13g2_inv_1 _3098_ (.Y(_0271_),
    .A(_0270_));
 sg13g2_a21oi_1 _3099_ (.A1(_1016_),
    .A2(_1018_),
    .Y(_0272_),
    .B1(_0269_));
 sg13g2_or2_1 _3100_ (.X(_0273_),
    .B(_0272_),
    .A(_0270_));
 sg13g2_nand2_1 _3101_ (.Y(_0274_),
    .A(_0268_),
    .B(_0273_));
 sg13g2_xor2_1 _3102_ (.B(_0273_),
    .A(_0268_),
    .X(_0275_));
 sg13g2_nand2_1 _3103_ (.Y(_0276_),
    .A(_0264_),
    .B(_0275_));
 sg13g2_xnor2_1 _3104_ (.Y(_0277_),
    .A(_0264_),
    .B(_0275_));
 sg13g2_xor2_1 _3105_ (.B(_0277_),
    .A(_0263_),
    .X(_0278_));
 sg13g2_and2_1 _3106_ (.A(_0257_),
    .B(_0278_),
    .X(_0279_));
 sg13g2_xor2_1 _3107_ (.B(_0278_),
    .A(_0257_),
    .X(_0280_));
 sg13g2_xnor2_1 _3108_ (.Y(_0281_),
    .A(_0256_),
    .B(_0280_));
 sg13g2_nor2b_1 _3109_ (.A(_0281_),
    .B_N(_0255_),
    .Y(_0282_));
 sg13g2_xnor2_1 _3110_ (.Y(_0283_),
    .A(_0255_),
    .B(_0281_));
 sg13g2_xnor2_1 _3111_ (.Y(_0284_),
    .A(_0254_),
    .B(_0283_));
 sg13g2_nor2_1 _3112_ (.A(_0253_),
    .B(_0284_),
    .Y(_0285_));
 sg13g2_nand2_1 _3113_ (.Y(_0286_),
    .A(_0253_),
    .B(_0284_));
 sg13g2_xor2_1 _3114_ (.B(_0284_),
    .A(_0253_),
    .X(_0287_));
 sg13g2_xnor2_1 _3115_ (.Y(_0288_),
    .A(_0252_),
    .B(_0287_));
 sg13g2_nor2_1 _3116_ (.A(_0184_),
    .B(_0288_),
    .Y(_0289_));
 sg13g2_nand2_1 _3117_ (.Y(_0290_),
    .A(_0184_),
    .B(_0288_));
 sg13g2_xor2_1 _3118_ (.B(_0288_),
    .A(_0184_),
    .X(_0291_));
 sg13g2_xnor2_1 _3119_ (.Y(_0292_),
    .A(_0183_),
    .B(_0291_));
 sg13g2_o21ai_1 _3120_ (.B1(_0135_),
    .Y(_0293_),
    .A1(_1409_),
    .A2(_0136_));
 sg13g2_o21ai_1 _3121_ (.B1(_1404_),
    .Y(_0294_),
    .A1(_1346_),
    .A2(_1405_));
 sg13g2_a21o_2 _3122_ (.A2(_1525_),
    .A1(_1411_),
    .B1(_1524_),
    .X(_0295_));
 sg13g2_nor2_1 _3123_ (.A(_1241_),
    .B(_1245_),
    .Y(_0296_));
 sg13g2_o21ai_1 _3124_ (.B1(_1334_),
    .Y(_0297_),
    .A1(_1316_),
    .A2(_1335_));
 sg13g2_nand2_1 _3125_ (.Y(_0298_),
    .A(_1235_),
    .B(_1238_));
 sg13g2_o21ai_1 _3126_ (.B1(_1313_),
    .Y(_0299_),
    .A1(_1301_),
    .A2(_1314_));
 sg13g2_o21ai_1 _3127_ (.B1(_1299_),
    .Y(_0300_),
    .A1(_1296_),
    .A2(_1300_));
 sg13g2_nand2_1 _3128_ (.Y(_0301_),
    .A(_1231_),
    .B(_1233_));
 sg13g2_nor2_1 _3129_ (.A(_0300_),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_xor2_1 _3130_ (.B(_0301_),
    .A(_0300_),
    .X(_0303_));
 sg13g2_inv_1 _3131_ (.Y(_0304_),
    .A(_0303_));
 sg13g2_and2_1 _3132_ (.A(_0299_),
    .B(_0304_),
    .X(_0305_));
 sg13g2_xnor2_1 _3133_ (.Y(_0306_),
    .A(_0299_),
    .B(_0303_));
 sg13g2_xnor2_1 _3134_ (.Y(_0307_),
    .A(_0298_),
    .B(_0306_));
 sg13g2_nand2b_1 _3135_ (.Y(_0308_),
    .B(_0297_),
    .A_N(_0307_));
 sg13g2_xor2_1 _3136_ (.B(_0307_),
    .A(_0297_),
    .X(_0309_));
 sg13g2_xnor2_1 _3137_ (.Y(_0310_),
    .A(_0296_),
    .B(_0309_));
 sg13g2_o21ai_1 _3138_ (.B1(_1292_),
    .Y(_0311_),
    .A1(_1293_),
    .A2(_1338_));
 sg13g2_nand2_1 _3139_ (.Y(_0312_),
    .A(_1308_),
    .B(_1310_));
 sg13g2_a21oi_1 _3140_ (.A1(_1318_),
    .A2(_1330_),
    .Y(_0313_),
    .B1(_1328_));
 sg13g2_o21ai_1 _3141_ (.B1(_1269_),
    .Y(_0314_),
    .A1(_1265_),
    .A2(_1270_));
 sg13g2_nand2_1 _3142_ (.Y(_0315_),
    .A(_1324_),
    .B(_1326_));
 sg13g2_nor2_2 _3143_ (.A(_0314_),
    .B(_0315_),
    .Y(_0316_));
 sg13g2_xor2_1 _3144_ (.B(_0315_),
    .A(_0314_),
    .X(_0317_));
 sg13g2_nor2_1 _3145_ (.A(_0313_),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_xor2_1 _3146_ (.B(_0317_),
    .A(_0313_),
    .X(_0319_));
 sg13g2_xnor2_1 _3147_ (.Y(_0320_),
    .A(_0312_),
    .B(_0319_));
 sg13g2_o21ai_1 _3148_ (.B1(_1287_),
    .Y(_0321_),
    .A1(_1260_),
    .A2(_1288_));
 sg13g2_nand2b_1 _3149_ (.Y(_0322_),
    .B(_1285_),
    .A_N(_1283_));
 sg13g2_o21ai_1 _3150_ (.B1(_1366_),
    .Y(_0323_),
    .A1(_1356_),
    .A2(_1367_));
 sg13g2_nand2_1 _3151_ (.Y(_0324_),
    .A(_1279_),
    .B(_1281_));
 sg13g2_and2_1 _3152_ (.A(_0323_),
    .B(_0324_),
    .X(_0325_));
 sg13g2_xor2_1 _3153_ (.B(_0324_),
    .A(_0323_),
    .X(_0326_));
 sg13g2_xor2_1 _3154_ (.B(_0326_),
    .A(_0322_),
    .X(_0327_));
 sg13g2_nand2_1 _3155_ (.Y(_0328_),
    .A(_0321_),
    .B(_0327_));
 sg13g2_xnor2_1 _3156_ (.Y(_0329_),
    .A(_0321_),
    .B(_0327_));
 sg13g2_xor2_1 _3157_ (.B(_0329_),
    .A(_0320_),
    .X(_0330_));
 sg13g2_nand2_1 _3158_ (.Y(_0331_),
    .A(_0311_),
    .B(_0330_));
 sg13g2_xnor2_1 _3159_ (.Y(_0332_),
    .A(_0311_),
    .B(_0330_));
 sg13g2_xor2_1 _3160_ (.B(_0332_),
    .A(_0310_),
    .X(_0333_));
 sg13g2_o21ai_1 _3161_ (.B1(_1399_),
    .Y(_0334_),
    .A1(_1350_),
    .A2(_1400_));
 sg13g2_nand2_1 _3162_ (.Y(_0335_),
    .A(_1394_),
    .B(_1396_));
 sg13g2_o21ai_1 _3163_ (.B1(_1478_),
    .Y(_0336_),
    .A1(_1435_),
    .A2(_1479_));
 sg13g2_nand2b_1 _3164_ (.Y(_0337_),
    .B(_1392_),
    .A_N(_1390_));
 sg13g2_a21oi_1 _3165_ (.A1(_1413_),
    .A2(_1433_),
    .Y(_0338_),
    .B1(_1432_));
 sg13g2_nand2_1 _3166_ (.Y(_0339_),
    .A(_1381_),
    .B(_1383_));
 sg13g2_o21ai_1 _3167_ (.B1(_1386_),
    .Y(_0340_),
    .A1(_1376_),
    .A2(_1387_));
 sg13g2_xor2_1 _3168_ (.B(_0340_),
    .A(_0339_),
    .X(_0341_));
 sg13g2_a21o_1 _3169_ (.A2(_1375_),
    .A1(_1371_),
    .B1(_1374_),
    .X(_0342_));
 sg13g2_nand2_1 _3170_ (.Y(_0343_),
    .A(_1361_),
    .B(_1363_));
 sg13g2_nor2_1 _3171_ (.A(_0342_),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_xnor2_1 _3172_ (.Y(_0345_),
    .A(_0342_),
    .B(_0343_));
 sg13g2_and2_1 _3173_ (.A(_0341_),
    .B(_0345_),
    .X(_0346_));
 sg13g2_xor2_1 _3174_ (.B(_0345_),
    .A(_0341_),
    .X(_0347_));
 sg13g2_nor2b_1 _3175_ (.A(_0338_),
    .B_N(_0347_),
    .Y(_0348_));
 sg13g2_xnor2_1 _3176_ (.Y(_0349_),
    .A(_0338_),
    .B(_0347_));
 sg13g2_xnor2_1 _3177_ (.Y(_0350_),
    .A(_0337_),
    .B(_0349_));
 sg13g2_nor2b_1 _3178_ (.A(_0350_),
    .B_N(_0336_),
    .Y(_0351_));
 sg13g2_xnor2_1 _3179_ (.Y(_0352_),
    .A(_0336_),
    .B(_0350_));
 sg13g2_xnor2_1 _3180_ (.Y(_0353_),
    .A(_0335_),
    .B(_0352_));
 sg13g2_nor2b_1 _3181_ (.A(_0353_),
    .B_N(_0334_),
    .Y(_0354_));
 sg13g2_xnor2_1 _3182_ (.Y(_0355_),
    .A(_0334_),
    .B(_0353_));
 sg13g2_xnor2_1 _3183_ (.Y(_0356_),
    .A(_0333_),
    .B(_0355_));
 sg13g2_nor2b_1 _3184_ (.A(_0356_),
    .B_N(_0295_),
    .Y(_0357_));
 sg13g2_xnor2_1 _3185_ (.Y(_0358_),
    .A(_0295_),
    .B(_0356_));
 sg13g2_xnor2_1 _3186_ (.Y(_0359_),
    .A(_0294_),
    .B(_0358_));
 sg13g2_o21ai_1 _3187_ (.B1(_0132_),
    .Y(_0360_),
    .A1(_1527_),
    .A2(_0133_));
 sg13g2_o21ai_1 _3188_ (.B1(_1518_),
    .Y(_0361_),
    .A1(_1483_),
    .A2(_1519_));
 sg13g2_o21ai_1 _3189_ (.B1(_0016_),
    .Y(_0362_),
    .A1(_1530_),
    .A2(_0017_));
 sg13g2_nand2_2 _3190_ (.Y(_0363_),
    .A(_1427_),
    .B(_1430_));
 sg13g2_o21ai_1 _3191_ (.B1(_1472_),
    .Y(_0364_),
    .A1(_1463_),
    .A2(_1473_));
 sg13g2_a21o_1 _3192_ (.A2(_1462_),
    .A1(_1458_),
    .B1(_1461_),
    .X(_0365_));
 sg13g2_nand2_2 _3193_ (.Y(_0366_),
    .A(_1423_),
    .B(_1425_));
 sg13g2_nor2_1 _3194_ (.A(_0365_),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_xnor2_1 _3195_ (.Y(_0368_),
    .A(_0365_),
    .B(_0366_));
 sg13g2_and2_1 _3196_ (.A(_0364_),
    .B(_0368_),
    .X(_0369_));
 sg13g2_xor2_1 _3197_ (.B(_0368_),
    .A(_0364_),
    .X(_0370_));
 sg13g2_xnor2_1 _3198_ (.Y(_0371_),
    .A(_0363_),
    .B(_0370_));
 sg13g2_o21ai_1 _3199_ (.B1(_1455_),
    .Y(_0372_),
    .A1(_1456_),
    .A2(_1475_));
 sg13g2_nand2_2 _3200_ (.Y(_0373_),
    .A(_1467_),
    .B(_1469_));
 sg13g2_o21ai_1 _3201_ (.B1(_1450_),
    .Y(_0374_),
    .A1(_1440_),
    .A2(_1451_));
 sg13g2_a21oi_1 _3202_ (.A1(_1491_),
    .A2(_1495_),
    .Y(_0375_),
    .B1(_1494_));
 sg13g2_nand2_1 _3203_ (.Y(_0376_),
    .A(_1446_),
    .B(_1448_));
 sg13g2_and3_1 _3204_ (.X(_0377_),
    .A(_1446_),
    .B(_1448_),
    .C(_0375_));
 sg13g2_xnor2_1 _3205_ (.Y(_0378_),
    .A(_0375_),
    .B(_0376_));
 sg13g2_a21oi_1 _3206_ (.A1(_1450_),
    .A2(_1453_),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_xnor2_1 _3207_ (.Y(_0380_),
    .A(_0374_),
    .B(_0378_));
 sg13g2_xnor2_1 _3208_ (.Y(_0381_),
    .A(_0373_),
    .B(_0380_));
 sg13g2_nand2b_1 _3209_ (.Y(_0382_),
    .B(_0372_),
    .A_N(_0381_));
 sg13g2_xor2_1 _3210_ (.B(_0381_),
    .A(_0372_),
    .X(_0383_));
 sg13g2_xor2_1 _3211_ (.B(_0383_),
    .A(_0371_),
    .X(_0384_));
 sg13g2_inv_1 _3212_ (.Y(_0385_),
    .A(_0384_));
 sg13g2_a21oi_1 _3213_ (.A1(_1486_),
    .A2(_1515_),
    .Y(_0386_),
    .B1(_1513_));
 sg13g2_and2_1 _3214_ (.A(_1509_),
    .B(_1511_),
    .X(_0387_));
 sg13g2_o21ai_1 _3215_ (.B1(_0010_),
    .Y(_0388_),
    .A1(_1575_),
    .A2(_0011_));
 sg13g2_nand2b_1 _3216_ (.Y(_0389_),
    .B(_1507_),
    .A_N(_1505_));
 sg13g2_o21ai_1 _3217_ (.B1(_1570_),
    .Y(_0390_),
    .A1(_1557_),
    .A2(_1571_));
 sg13g2_nand2_1 _3218_ (.Y(_0391_),
    .A(_1501_),
    .B(_1503_));
 sg13g2_and2_1 _3219_ (.A(_0390_),
    .B(_0391_),
    .X(_0392_));
 sg13g2_xor2_1 _3220_ (.B(_0391_),
    .A(_0390_),
    .X(_0393_));
 sg13g2_xnor2_1 _3221_ (.Y(_0394_),
    .A(_0389_),
    .B(_0393_));
 sg13g2_nand2b_1 _3222_ (.Y(_0395_),
    .B(_0388_),
    .A_N(_0394_));
 sg13g2_xor2_1 _3223_ (.B(_0394_),
    .A(_0388_),
    .X(_0396_));
 sg13g2_xnor2_1 _3224_ (.Y(_0397_),
    .A(_0387_),
    .B(_0396_));
 sg13g2_nor2_1 _3225_ (.A(_0386_),
    .B(_0397_),
    .Y(_0398_));
 sg13g2_xnor2_1 _3226_ (.Y(_0399_),
    .A(_0386_),
    .B(_0397_));
 sg13g2_nor2_1 _3227_ (.A(_0385_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_xnor2_1 _3228_ (.Y(_0401_),
    .A(_0385_),
    .B(_0399_));
 sg13g2_nor2b_1 _3229_ (.A(_0401_),
    .B_N(_0362_),
    .Y(_0402_));
 sg13g2_xnor2_1 _3230_ (.Y(_0403_),
    .A(_0362_),
    .B(_0401_));
 sg13g2_xnor2_1 _3231_ (.Y(_0404_),
    .A(_0361_),
    .B(_0403_));
 sg13g2_o21ai_1 _3232_ (.B1(_0129_),
    .Y(_0405_),
    .A1(_0020_),
    .A2(_0130_));
 sg13g2_o21ai_1 _3233_ (.B1(_0126_),
    .Y(_0406_),
    .A1(_0067_),
    .A2(_0127_));
 sg13g2_nand2b_1 _3234_ (.Y(_0407_),
    .B(_0061_),
    .A_N(_0059_));
 sg13g2_a21oi_1 _3235_ (.A1(_0069_),
    .A2(_0089_),
    .Y(_0408_),
    .B1(_0088_));
 sg13g2_nand2_2 _3236_ (.Y(_0409_),
    .A(_0035_),
    .B(_0037_));
 sg13g2_a21o_1 _3237_ (.A2(_0056_),
    .A1(_0046_),
    .B1(_0054_),
    .X(_0410_));
 sg13g2_a21oi_1 _3238_ (.A1(_0071_),
    .A2(_0075_),
    .Y(_0411_),
    .B1(_0074_));
 sg13g2_a21oi_1 _3239_ (.A1(_0048_),
    .A2(_0049_),
    .Y(_0412_),
    .B1(_0052_));
 sg13g2_and2_1 _3240_ (.A(_0411_),
    .B(_0412_),
    .X(_0413_));
 sg13g2_xnor2_1 _3241_ (.Y(_0414_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_and2_1 _3242_ (.A(_0410_),
    .B(_0414_),
    .X(_0415_));
 sg13g2_xor2_1 _3243_ (.B(_0414_),
    .A(_0410_),
    .X(_0416_));
 sg13g2_xnor2_1 _3244_ (.Y(_0417_),
    .A(_0409_),
    .B(_0416_));
 sg13g2_nor2_1 _3245_ (.A(_0408_),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_xor2_1 _3246_ (.B(_0417_),
    .A(_0408_),
    .X(_0419_));
 sg13g2_xnor2_1 _3247_ (.Y(_0420_),
    .A(_0407_),
    .B(_0419_));
 sg13g2_o21ai_1 _3248_ (.B1(_0123_),
    .Y(_0421_),
    .A1(_0090_),
    .A2(_0124_));
 sg13g2_o21ai_1 _3249_ (.B1(_0085_),
    .Y(_0422_),
    .A1(_0077_),
    .A2(_0086_));
 sg13g2_a21oi_2 _3250_ (.B1(_0100_),
    .Y(_0423_),
    .A2(_0101_),
    .A1(_0092_));
 sg13g2_a21o_1 _3251_ (.A2(_0083_),
    .A1(_0079_),
    .B1(_0082_),
    .X(_0424_));
 sg13g2_nor2b_1 _3252_ (.A(_0423_),
    .B_N(_0424_),
    .Y(_0425_));
 sg13g2_xor2_1 _3253_ (.B(_0424_),
    .A(_0423_),
    .X(_0426_));
 sg13g2_nor2b_1 _3254_ (.A(_0426_),
    .B_N(_0422_),
    .Y(_0427_));
 sg13g2_xor2_1 _3255_ (.B(_0426_),
    .A(_0422_),
    .X(_0428_));
 sg13g2_o21ai_1 _3256_ (.B1(_0120_),
    .Y(_0429_),
    .A1(_0102_),
    .A2(_0121_));
 sg13g2_a21oi_2 _3257_ (.B1(_0114_),
    .Y(_0430_),
    .A2(_0115_),
    .A1(_0111_));
 sg13g2_o21ai_1 _3258_ (.B1(_0117_),
    .Y(_0431_),
    .A1(_0109_),
    .A2(_0118_));
 sg13g2_inv_1 _3259_ (.Y(_0432_),
    .A(_0431_));
 sg13g2_xor2_1 _3260_ (.B(_0431_),
    .A(_0430_),
    .X(_0433_));
 sg13g2_a21oi_1 _3261_ (.A1(_0104_),
    .A2(_0108_),
    .Y(_0434_),
    .B1(_0107_));
 sg13g2_a21oi_2 _3262_ (.B1(_0097_),
    .Y(_0435_),
    .A2(_0098_),
    .A1(_0094_));
 sg13g2_nand2_1 _3263_ (.Y(_0436_),
    .A(_0434_),
    .B(_0435_));
 sg13g2_xnor2_1 _3264_ (.Y(_0437_),
    .A(_0434_),
    .B(_0435_));
 sg13g2_nand2b_1 _3265_ (.Y(_0438_),
    .B(_0437_),
    .A_N(_0433_));
 sg13g2_xor2_1 _3266_ (.B(_0437_),
    .A(_0433_),
    .X(_0439_));
 sg13g2_nand2b_1 _3267_ (.Y(_0440_),
    .B(_0429_),
    .A_N(_0439_));
 sg13g2_xor2_1 _3268_ (.B(_0439_),
    .A(_0429_),
    .X(_0441_));
 sg13g2_or2_1 _3269_ (.X(_0442_),
    .B(_0441_),
    .A(_0428_));
 sg13g2_xor2_1 _3270_ (.B(_0441_),
    .A(_0428_),
    .X(_0443_));
 sg13g2_nand2_1 _3271_ (.Y(_0444_),
    .A(_0421_),
    .B(_0443_));
 sg13g2_xnor2_1 _3272_ (.Y(_0445_),
    .A(_0421_),
    .B(_0443_));
 sg13g2_xor2_1 _3273_ (.B(_0445_),
    .A(_0420_),
    .X(_0446_));
 sg13g2_nand2_1 _3274_ (.Y(_0447_),
    .A(_0406_),
    .B(_0446_));
 sg13g2_xnor2_1 _3275_ (.Y(_0448_),
    .A(_0406_),
    .B(_0446_));
 sg13g2_and2_1 _3276_ (.A(_1555_),
    .B(_0014_),
    .X(_0449_));
 sg13g2_o21ai_1 _3277_ (.B1(_0064_),
    .Y(_0450_),
    .A1(_0023_),
    .A2(_0065_));
 sg13g2_nor2_1 _3278_ (.A(_1587_),
    .B(_0002_),
    .Y(_0451_));
 sg13g2_o21ai_1 _3279_ (.B1(_0005_),
    .Y(_0452_),
    .A1(_1583_),
    .A2(_0006_));
 sg13g2_nand2b_1 _3280_ (.Y(_0453_),
    .B(_0452_),
    .A_N(_0451_));
 sg13g2_xor2_1 _3281_ (.B(_0452_),
    .A(_0451_),
    .X(_0454_));
 sg13g2_a21o_1 _3282_ (.A2(_1582_),
    .A1(_1578_),
    .B1(_1581_),
    .X(_0455_));
 sg13g2_nand2_2 _3283_ (.Y(_0456_),
    .A(_1563_),
    .B(_1567_));
 sg13g2_or2_1 _3284_ (.X(_0457_),
    .B(_0456_),
    .A(_0455_));
 sg13g2_xor2_1 _3285_ (.B(_0456_),
    .A(_0455_),
    .X(_0458_));
 sg13g2_xnor2_1 _3286_ (.Y(_0459_),
    .A(_0454_),
    .B(_0458_));
 sg13g2_a21oi_1 _3287_ (.A1(_1535_),
    .A2(_1552_),
    .Y(_0460_),
    .B1(_1550_));
 sg13g2_nand2_1 _3288_ (.Y(_0461_),
    .A(_1546_),
    .B(_1548_));
 sg13g2_o21ai_1 _3289_ (.B1(_0039_),
    .Y(_0462_),
    .A1(_0031_),
    .A2(_0040_));
 sg13g2_a21oi_1 _3290_ (.A1(_0025_),
    .A2(_0029_),
    .Y(_0463_),
    .B1(_0028_));
 sg13g2_nor2b_1 _3291_ (.A(_1542_),
    .B_N(_1544_),
    .Y(_0464_));
 sg13g2_and2_1 _3292_ (.A(_0463_),
    .B(_0464_),
    .X(_0465_));
 sg13g2_xnor2_1 _3293_ (.Y(_0466_),
    .A(_0463_),
    .B(_0464_));
 sg13g2_and2_1 _3294_ (.A(_0462_),
    .B(_0466_),
    .X(_0467_));
 sg13g2_xor2_1 _3295_ (.B(_0466_),
    .A(_0462_),
    .X(_0468_));
 sg13g2_xnor2_1 _3296_ (.Y(_0469_),
    .A(_0461_),
    .B(_0468_));
 sg13g2_or2_1 _3297_ (.X(_0470_),
    .B(_0469_),
    .A(_0460_));
 sg13g2_xnor2_1 _3298_ (.Y(_0471_),
    .A(_0460_),
    .B(_0469_));
 sg13g2_xor2_1 _3299_ (.B(_0471_),
    .A(_0459_),
    .X(_0472_));
 sg13g2_nand2_1 _3300_ (.Y(_0473_),
    .A(_0450_),
    .B(_0472_));
 sg13g2_xnor2_1 _3301_ (.Y(_0474_),
    .A(_0450_),
    .B(_0472_));
 sg13g2_xnor2_1 _3302_ (.Y(_0475_),
    .A(_0449_),
    .B(_0474_));
 sg13g2_xor2_1 _3303_ (.B(_0475_),
    .A(_0448_),
    .X(_0476_));
 sg13g2_nand2_1 _3304_ (.Y(_0477_),
    .A(_0405_),
    .B(_0476_));
 sg13g2_xnor2_1 _3305_ (.Y(_0478_),
    .A(_0405_),
    .B(_0476_));
 sg13g2_xor2_1 _3306_ (.B(_0478_),
    .A(_0404_),
    .X(_0479_));
 sg13g2_nand2_1 _3307_ (.Y(_0480_),
    .A(_0360_),
    .B(_0479_));
 sg13g2_xnor2_1 _3308_ (.Y(_0481_),
    .A(_0360_),
    .B(_0479_));
 sg13g2_xor2_1 _3309_ (.B(_0481_),
    .A(_0359_),
    .X(_0482_));
 sg13g2_nand2_1 _3310_ (.Y(_0483_),
    .A(_0293_),
    .B(_0482_));
 sg13g2_xnor2_1 _3311_ (.Y(_0484_),
    .A(_0293_),
    .B(_0482_));
 sg13g2_xor2_1 _3312_ (.B(_0484_),
    .A(_0292_),
    .X(_0485_));
 sg13g2_nand2_1 _3313_ (.Y(_0486_),
    .A(_0182_),
    .B(_0485_));
 sg13g2_xnor2_1 _3314_ (.Y(_0487_),
    .A(_0182_),
    .B(_0485_));
 sg13g2_xor2_1 _3315_ (.B(_0487_),
    .A(_0181_),
    .X(_0488_));
 sg13g2_nand2_1 _3316_ (.Y(_0489_),
    .A(_0151_),
    .B(_0488_));
 sg13g2_xnor2_1 _3317_ (.Y(_0490_),
    .A(_0151_),
    .B(_0488_));
 sg13g2_xnor2_1 _3318_ (.Y(_0491_),
    .A(_0150_),
    .B(_0490_));
 sg13g2_nor2_1 _3319_ (.A(_0149_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_xor2_1 _3320_ (.B(_0491_),
    .A(_0149_),
    .X(_0493_));
 sg13g2_xor2_1 _3321_ (.B(_0493_),
    .A(_0148_),
    .X(uo_out[1]));
 sg13g2_nand2_1 _3322_ (.Y(_0494_),
    .A(_0178_),
    .B(_0180_));
 sg13g2_inv_1 _3323_ (.Y(_0495_),
    .A(_0494_));
 sg13g2_o21ai_1 _3324_ (.B1(_0486_),
    .Y(_0496_),
    .A1(_0181_),
    .A2(_0487_));
 sg13g2_o21ai_1 _3325_ (.B1(_0175_),
    .Y(_0497_),
    .A1(_0155_),
    .A2(_0176_));
 sg13g2_a21oi_1 _3326_ (.A1(_0183_),
    .A2(_0290_),
    .Y(_0498_),
    .B1(_0289_));
 sg13g2_a21oi_1 _3327_ (.A1(_0157_),
    .A2(_0173_),
    .Y(_0499_),
    .B1(_0172_));
 sg13g2_o21ai_1 _3328_ (.B1(_0250_),
    .Y(_0500_),
    .A1(_0203_),
    .A2(_0251_));
 sg13g2_o21ai_1 _3329_ (.B1(_0169_),
    .Y(_0501_),
    .A1(_0160_),
    .A2(_0170_));
 sg13g2_o21ai_1 _3330_ (.B1(_0201_),
    .Y(_0502_),
    .A1(_0186_),
    .A2(_0202_));
 sg13g2_nor3_2 _3331_ (.A(_0163_),
    .B(_0166_),
    .C(_0167_),
    .Y(_0503_));
 sg13g2_a21oi_1 _3332_ (.A1(_0163_),
    .A2(_0166_),
    .Y(_0504_),
    .B1(_0503_));
 sg13g2_xnor2_1 _3333_ (.Y(_0505_),
    .A(_0502_),
    .B(_0504_));
 sg13g2_nor2b_1 _3334_ (.A(_0505_),
    .B_N(_0501_),
    .Y(_0506_));
 sg13g2_xor2_1 _3335_ (.B(_0505_),
    .A(_0501_),
    .X(_0507_));
 sg13g2_nand2b_1 _3336_ (.Y(_0508_),
    .B(_0500_),
    .A_N(_0507_));
 sg13g2_xor2_1 _3337_ (.B(_0507_),
    .A(_0500_),
    .X(_0509_));
 sg13g2_xor2_1 _3338_ (.B(_0509_),
    .A(_0499_),
    .X(_0510_));
 sg13g2_nor2b_1 _3339_ (.A(_0498_),
    .B_N(_0510_),
    .Y(_0511_));
 sg13g2_xnor2_1 _3340_ (.Y(_0512_),
    .A(_0498_),
    .B(_0510_));
 sg13g2_xnor2_1 _3341_ (.Y(_0513_),
    .A(_0497_),
    .B(_0512_));
 sg13g2_o21ai_1 _3342_ (.B1(_0483_),
    .Y(_0514_),
    .A1(_0292_),
    .A2(_0484_));
 sg13g2_a21oi_1 _3343_ (.A1(_0252_),
    .A2(_0286_),
    .Y(_0515_),
    .B1(_0285_));
 sg13g2_a21oi_2 _3344_ (.B1(_0357_),
    .Y(_0516_),
    .A2(_0358_),
    .A1(_0294_));
 sg13g2_o21ai_1 _3345_ (.B1(_0199_),
    .Y(_0517_),
    .A1(_0190_),
    .A2(_0197_));
 sg13g2_a21oi_1 _3346_ (.A1(_0215_),
    .A2(_0229_),
    .Y(_0518_),
    .B1(_0227_));
 sg13g2_a21oi_1 _3347_ (.A1(_0191_),
    .A2(_0196_),
    .Y(_0519_),
    .B1(_0194_));
 sg13g2_nand2_1 _3348_ (.Y(_0520_),
    .A(_0208_),
    .B(_0212_));
 sg13g2_a21o_1 _3349_ (.A2(_0214_),
    .A1(_0207_),
    .B1(_0212_),
    .X(_0521_));
 sg13g2_nand2_1 _3350_ (.Y(_0522_),
    .A(_0520_),
    .B(_0521_));
 sg13g2_xor2_1 _3351_ (.B(_0522_),
    .A(_0519_),
    .X(_0523_));
 sg13g2_nor2b_1 _3352_ (.A(_0518_),
    .B_N(_0523_),
    .Y(_0524_));
 sg13g2_xnor2_1 _3353_ (.Y(_0525_),
    .A(_0518_),
    .B(_0523_));
 sg13g2_xnor2_1 _3354_ (.Y(_0526_),
    .A(_0517_),
    .B(_0525_));
 sg13g2_o21ai_1 _3355_ (.B1(_0247_),
    .Y(_0527_),
    .A1(_0230_),
    .A2(_0248_));
 sg13g2_a21oi_1 _3356_ (.A1(_0218_),
    .A2(_0223_),
    .Y(_0528_),
    .B1(_0225_));
 sg13g2_nand2_1 _3357_ (.Y(_0529_),
    .A(_0221_),
    .B(_0528_));
 sg13g2_xnor2_1 _3358_ (.Y(_0530_),
    .A(_0221_),
    .B(_0528_));
 sg13g2_a21oi_1 _3359_ (.A1(_0232_),
    .A2(_0244_),
    .Y(_0531_),
    .B1(_0243_));
 sg13g2_a21o_1 _3360_ (.A2(_0241_),
    .A1(_0234_),
    .B1(_0240_),
    .X(_0532_));
 sg13g2_a21oi_2 _3361_ (.B1(_0261_),
    .Y(_0533_),
    .A2(_0262_),
    .A1(_0258_));
 sg13g2_inv_1 _3362_ (.Y(_0534_),
    .A(_0533_));
 sg13g2_xnor2_1 _3363_ (.Y(_0535_),
    .A(_0238_),
    .B(_0533_));
 sg13g2_and2_1 _3364_ (.A(_0532_),
    .B(_0535_),
    .X(_0536_));
 sg13g2_xnor2_1 _3365_ (.Y(_0537_),
    .A(_0532_),
    .B(_0535_));
 sg13g2_xor2_1 _3366_ (.B(_0537_),
    .A(_0531_),
    .X(_0538_));
 sg13g2_nand2_1 _3367_ (.Y(_0539_),
    .A(_0530_),
    .B(_0538_));
 sg13g2_xnor2_1 _3368_ (.Y(_0540_),
    .A(_0530_),
    .B(_0538_));
 sg13g2_nand2b_1 _3369_ (.Y(_0541_),
    .B(_0527_),
    .A_N(_0540_));
 sg13g2_xor2_1 _3370_ (.B(_0540_),
    .A(_0527_),
    .X(_0542_));
 sg13g2_xor2_1 _3371_ (.B(_0542_),
    .A(_0526_),
    .X(_0543_));
 sg13g2_a21oi_1 _3372_ (.A1(_0254_),
    .A2(_0283_),
    .Y(_0544_),
    .B1(_0282_));
 sg13g2_a21oi_1 _3373_ (.A1(_0256_),
    .A2(_0280_),
    .Y(_0545_),
    .B1(_0279_));
 sg13g2_o21ai_1 _3374_ (.B1(_0331_),
    .Y(_0546_),
    .A1(_0310_),
    .A2(_0332_));
 sg13g2_o21ai_1 _3375_ (.B1(_0276_),
    .Y(_0547_),
    .A1(_0263_),
    .A2(_0277_));
 sg13g2_o21ai_1 _3376_ (.B1(_0308_),
    .Y(_0548_),
    .A1(_0296_),
    .A2(_0309_));
 sg13g2_nor3_2 _3377_ (.A(_0265_),
    .B(_0266_),
    .C(_0271_),
    .Y(_0549_));
 sg13g2_a21oi_1 _3378_ (.A1(_0267_),
    .A2(_0274_),
    .Y(_0550_),
    .B1(_0270_));
 sg13g2_nor2_1 _3379_ (.A(_0549_),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_or2_1 _3380_ (.X(_0552_),
    .B(_0550_),
    .A(_0549_));
 sg13g2_and2_1 _3381_ (.A(_0548_),
    .B(_0552_),
    .X(_0553_));
 sg13g2_xnor2_1 _3382_ (.Y(_0554_),
    .A(_0548_),
    .B(_0551_));
 sg13g2_xnor2_1 _3383_ (.Y(_0555_),
    .A(_0547_),
    .B(_0554_));
 sg13g2_nand2b_1 _3384_ (.Y(_0556_),
    .B(_0546_),
    .A_N(_0555_));
 sg13g2_xor2_1 _3385_ (.B(_0555_),
    .A(_0546_),
    .X(_0557_));
 sg13g2_xor2_1 _3386_ (.B(_0557_),
    .A(_0545_),
    .X(_0558_));
 sg13g2_nor2b_1 _3387_ (.A(_0544_),
    .B_N(_0558_),
    .Y(_0559_));
 sg13g2_xnor2_1 _3388_ (.Y(_0560_),
    .A(_0544_),
    .B(_0558_));
 sg13g2_xnor2_1 _3389_ (.Y(_0561_),
    .A(_0543_),
    .B(_0560_));
 sg13g2_nor2_1 _3390_ (.A(_0516_),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_xor2_1 _3391_ (.B(_0561_),
    .A(_0516_),
    .X(_0563_));
 sg13g2_nor2b_1 _3392_ (.A(_0515_),
    .B_N(_0563_),
    .Y(_0564_));
 sg13g2_xor2_1 _3393_ (.B(_0563_),
    .A(_0515_),
    .X(_0565_));
 sg13g2_o21ai_1 _3394_ (.B1(_0480_),
    .Y(_0566_),
    .A1(_0359_),
    .A2(_0481_));
 sg13g2_a21o_2 _3395_ (.A2(_0355_),
    .A1(_0333_),
    .B1(_0354_),
    .X(_0567_));
 sg13g2_a21oi_1 _3396_ (.A1(_0361_),
    .A2(_0403_),
    .Y(_0568_),
    .B1(_0402_));
 sg13g2_a21oi_1 _3397_ (.A1(_0298_),
    .A2(_0306_),
    .Y(_0569_),
    .B1(_0305_));
 sg13g2_a21oi_1 _3398_ (.A1(_0312_),
    .A2(_0319_),
    .Y(_0570_),
    .B1(_0318_));
 sg13g2_nor2_1 _3399_ (.A(_0302_),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_xnor2_1 _3400_ (.Y(_0572_),
    .A(_0302_),
    .B(_0570_));
 sg13g2_nor2_1 _3401_ (.A(_0569_),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_xnor2_1 _3402_ (.Y(_0574_),
    .A(_0569_),
    .B(_0572_));
 sg13g2_o21ai_1 _3403_ (.B1(_0328_),
    .Y(_0575_),
    .A1(_0320_),
    .A2(_0329_));
 sg13g2_a21oi_1 _3404_ (.A1(_0322_),
    .A2(_0326_),
    .Y(_0576_),
    .B1(_0325_));
 sg13g2_or2_1 _3405_ (.X(_0577_),
    .B(_0576_),
    .A(_0344_));
 sg13g2_xnor2_1 _3406_ (.Y(_0578_),
    .A(_0344_),
    .B(_0576_));
 sg13g2_xor2_1 _3407_ (.B(_0578_),
    .A(_0316_),
    .X(_0579_));
 sg13g2_nand2_1 _3408_ (.Y(_0580_),
    .A(_0575_),
    .B(_0579_));
 sg13g2_xnor2_1 _3409_ (.Y(_0581_),
    .A(_0575_),
    .B(_0579_));
 sg13g2_xnor2_1 _3410_ (.Y(_0582_),
    .A(_0574_),
    .B(_0581_));
 sg13g2_a21oi_2 _3411_ (.B1(_0351_),
    .Y(_0583_),
    .A2(_0352_),
    .A1(_0335_));
 sg13g2_a21oi_2 _3412_ (.B1(_0348_),
    .Y(_0584_),
    .A2(_0349_),
    .A1(_0337_));
 sg13g2_o21ai_1 _3413_ (.B1(_0382_),
    .Y(_0585_),
    .A1(_0371_),
    .A2(_0383_));
 sg13g2_a21oi_1 _3414_ (.A1(_0363_),
    .A2(_0370_),
    .Y(_0586_),
    .B1(_0369_));
 sg13g2_inv_1 _3415_ (.Y(_0587_),
    .A(_0586_));
 sg13g2_a21o_2 _3416_ (.A2(_0340_),
    .A1(_0339_),
    .B1(_0346_),
    .X(_0588_));
 sg13g2_nor2_1 _3417_ (.A(_0587_),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_xor2_1 _3418_ (.B(_0588_),
    .A(_0586_),
    .X(_0590_));
 sg13g2_nand2_1 _3419_ (.Y(_0591_),
    .A(_0585_),
    .B(_0590_));
 sg13g2_nor2_1 _3420_ (.A(_0585_),
    .B(_0590_),
    .Y(_0592_));
 sg13g2_xor2_1 _3421_ (.B(_0590_),
    .A(_0585_),
    .X(_0593_));
 sg13g2_xnor2_1 _3422_ (.Y(_0594_),
    .A(_0584_),
    .B(_0593_));
 sg13g2_nand2b_1 _3423_ (.Y(_0595_),
    .B(_0594_),
    .A_N(_0583_));
 sg13g2_xnor2_1 _3424_ (.Y(_0596_),
    .A(_0583_),
    .B(_0594_));
 sg13g2_nand2b_1 _3425_ (.Y(_0597_),
    .B(_0596_),
    .A_N(_0582_));
 sg13g2_xor2_1 _3426_ (.B(_0596_),
    .A(_0582_),
    .X(_0598_));
 sg13g2_nor2_1 _3427_ (.A(_0568_),
    .B(_0598_),
    .Y(_0599_));
 sg13g2_xor2_1 _3428_ (.B(_0598_),
    .A(_0568_),
    .X(_0600_));
 sg13g2_xnor2_1 _3429_ (.Y(_0601_),
    .A(_0567_),
    .B(_0600_));
 sg13g2_o21ai_1 _3430_ (.B1(_0477_),
    .Y(_0602_),
    .A1(_0404_),
    .A2(_0478_));
 sg13g2_nor2_2 _3431_ (.A(_0398_),
    .B(_0400_),
    .Y(_0603_));
 sg13g2_o21ai_1 _3432_ (.B1(_0473_),
    .Y(_0604_),
    .A1(_0449_),
    .A2(_0474_));
 sg13g2_a21oi_1 _3433_ (.A1(_0373_),
    .A2(_0380_),
    .Y(_0605_),
    .B1(_0379_));
 sg13g2_or2_1 _3434_ (.X(_0606_),
    .B(_0605_),
    .A(_0377_));
 sg13g2_xnor2_1 _3435_ (.Y(_0607_),
    .A(_0377_),
    .B(_0605_));
 sg13g2_xor2_1 _3436_ (.B(_0607_),
    .A(_0367_),
    .X(_0608_));
 sg13g2_inv_1 _3437_ (.Y(_0609_),
    .A(_0608_));
 sg13g2_o21ai_1 _3438_ (.B1(_0395_),
    .Y(_0610_),
    .A1(_0387_),
    .A2(_0396_));
 sg13g2_a21o_1 _3439_ (.A2(_0393_),
    .A1(_0389_),
    .B1(_0392_),
    .X(_0611_));
 sg13g2_nor4_1 _3440_ (.A(_1587_),
    .B(_0002_),
    .C(_0452_),
    .D(_0457_),
    .Y(_0612_));
 sg13g2_o21ai_1 _3441_ (.B1(_0453_),
    .Y(_0613_),
    .A1(_0454_),
    .A2(_0458_));
 sg13g2_a21oi_1 _3442_ (.A1(_0457_),
    .A2(_0613_),
    .Y(_0614_),
    .B1(_0612_));
 sg13g2_xor2_1 _3443_ (.B(_0614_),
    .A(_0611_),
    .X(_0615_));
 sg13g2_xnor2_1 _3444_ (.Y(_0616_),
    .A(_0610_),
    .B(_0615_));
 sg13g2_nor2_1 _3445_ (.A(_0609_),
    .B(_0616_),
    .Y(_0617_));
 sg13g2_xnor2_1 _3446_ (.Y(_0618_),
    .A(_0609_),
    .B(_0616_));
 sg13g2_nand2b_1 _3447_ (.Y(_0619_),
    .B(_0604_),
    .A_N(_0618_));
 sg13g2_xor2_1 _3448_ (.B(_0618_),
    .A(_0604_),
    .X(_0620_));
 sg13g2_xor2_1 _3449_ (.B(_0620_),
    .A(_0603_),
    .X(_0621_));
 sg13g2_o21ai_1 _3450_ (.B1(_0447_),
    .Y(_0622_),
    .A1(_0448_),
    .A2(_0475_));
 sg13g2_o21ai_1 _3451_ (.B1(_0470_),
    .Y(_0623_),
    .A1(_0459_),
    .A2(_0471_));
 sg13g2_a21oi_2 _3452_ (.B1(_0418_),
    .Y(_0624_),
    .A2(_0419_),
    .A1(_0407_));
 sg13g2_a21oi_2 _3453_ (.B1(_0467_),
    .Y(_0625_),
    .A2(_0468_),
    .A1(_0461_));
 sg13g2_nand2_2 _3454_ (.Y(_0626_),
    .A(_0465_),
    .B(_0625_));
 sg13g2_xnor2_1 _3455_ (.Y(_0627_),
    .A(_0465_),
    .B(_0625_));
 sg13g2_nor2b_1 _3456_ (.A(_0624_),
    .B_N(_0627_),
    .Y(_0628_));
 sg13g2_xnor2_1 _3457_ (.Y(_0629_),
    .A(_0624_),
    .B(_0627_));
 sg13g2_xnor2_1 _3458_ (.Y(_0630_),
    .A(_0623_),
    .B(_0629_));
 sg13g2_o21ai_1 _3459_ (.B1(_0444_),
    .Y(_0631_),
    .A1(_0420_),
    .A2(_0445_));
 sg13g2_a21oi_1 _3460_ (.A1(_0409_),
    .A2(_0416_),
    .Y(_0632_),
    .B1(_0415_));
 sg13g2_nor2_1 _3461_ (.A(_0425_),
    .B(_0427_),
    .Y(_0633_));
 sg13g2_nor2_1 _3462_ (.A(_0413_),
    .B(_0633_),
    .Y(_0634_));
 sg13g2_xnor2_1 _3463_ (.Y(_0635_),
    .A(_0413_),
    .B(_0633_));
 sg13g2_nor2_1 _3464_ (.A(_0632_),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_xor2_1 _3465_ (.B(_0635_),
    .A(_0632_),
    .X(_0637_));
 sg13g2_o21ai_1 _3466_ (.B1(_0440_),
    .Y(_0638_),
    .A1(_0428_),
    .A2(_0441_));
 sg13g2_and4_1 _3467_ (.A(_0430_),
    .B(_0432_),
    .C(_0434_),
    .D(_0435_),
    .X(_0639_));
 sg13g2_o21ai_1 _3468_ (.B1(_0438_),
    .Y(_0640_),
    .A1(_0430_),
    .A2(_0432_));
 sg13g2_a21oi_1 _3469_ (.A1(_0436_),
    .A2(_0640_),
    .Y(_0641_),
    .B1(_0639_));
 sg13g2_a21oi_1 _3470_ (.A1(_0440_),
    .A2(_0442_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_xnor2_1 _3471_ (.Y(_0643_),
    .A(_0638_),
    .B(_0641_));
 sg13g2_xnor2_1 _3472_ (.Y(_0644_),
    .A(_0637_),
    .B(_0643_));
 sg13g2_nand2b_1 _3473_ (.Y(_0645_),
    .B(_0631_),
    .A_N(_0644_));
 sg13g2_xor2_1 _3474_ (.B(_0644_),
    .A(_0631_),
    .X(_0646_));
 sg13g2_xor2_1 _3475_ (.B(_0646_),
    .A(_0630_),
    .X(_0647_));
 sg13g2_and2_1 _3476_ (.A(_0622_),
    .B(_0647_),
    .X(_0648_));
 sg13g2_or2_1 _3477_ (.X(_0649_),
    .B(_0647_),
    .A(_0622_));
 sg13g2_xnor2_1 _3478_ (.Y(_0650_),
    .A(_0622_),
    .B(_0647_));
 sg13g2_xnor2_1 _3479_ (.Y(_0651_),
    .A(_0621_),
    .B(_0650_));
 sg13g2_nand2_1 _3480_ (.Y(_0652_),
    .A(_0602_),
    .B(_0651_));
 sg13g2_xnor2_1 _3481_ (.Y(_0653_),
    .A(_0602_),
    .B(_0651_));
 sg13g2_xor2_1 _3482_ (.B(_0653_),
    .A(_0601_),
    .X(_0654_));
 sg13g2_nand2_1 _3483_ (.Y(_0655_),
    .A(_0566_),
    .B(_0654_));
 sg13g2_xnor2_1 _3484_ (.Y(_0656_),
    .A(_0566_),
    .B(_0654_));
 sg13g2_xnor2_1 _3485_ (.Y(_0657_),
    .A(_0565_),
    .B(_0656_));
 sg13g2_nand2b_1 _3486_ (.Y(_0658_),
    .B(_0514_),
    .A_N(_0657_));
 sg13g2_xor2_1 _3487_ (.B(_0657_),
    .A(_0514_),
    .X(_0659_));
 sg13g2_xor2_1 _3488_ (.B(_0659_),
    .A(_0513_),
    .X(_0660_));
 sg13g2_nand2_1 _3489_ (.Y(_0661_),
    .A(_0496_),
    .B(_0660_));
 sg13g2_xnor2_1 _3490_ (.Y(_0662_),
    .A(_0496_),
    .B(_0660_));
 sg13g2_xnor2_1 _3491_ (.Y(_0663_),
    .A(_0495_),
    .B(_0662_));
 sg13g2_o21ai_1 _3492_ (.B1(_0489_),
    .Y(_0664_),
    .A1(_0150_),
    .A2(_0490_));
 sg13g2_nand2b_1 _3493_ (.Y(_0665_),
    .B(_0664_),
    .A_N(_0663_));
 sg13g2_xor2_1 _3494_ (.B(_0664_),
    .A(_0663_),
    .X(_0666_));
 sg13g2_a21oi_2 _3495_ (.B1(_0492_),
    .Y(_0667_),
    .A2(_0493_),
    .A1(_0148_));
 sg13g2_xor2_1 _3496_ (.B(_0667_),
    .A(_0666_),
    .X(uo_out[2]));
 sg13g2_o21ai_1 _3497_ (.B1(_0661_),
    .Y(_0668_),
    .A1(_0495_),
    .A2(_0662_));
 sg13g2_a21oi_2 _3498_ (.B1(_0511_),
    .Y(_0669_),
    .A2(_0512_),
    .A1(_0497_));
 sg13g2_o21ai_1 _3499_ (.B1(_0658_),
    .Y(_0670_),
    .A1(_0513_),
    .A2(_0659_));
 sg13g2_o21ai_1 _3500_ (.B1(_0508_),
    .Y(_0671_),
    .A1(_0499_),
    .A2(_0509_));
 sg13g2_nor2_1 _3501_ (.A(_0562_),
    .B(_0564_),
    .Y(_0672_));
 sg13g2_a21oi_1 _3502_ (.A1(_0502_),
    .A2(_0504_),
    .Y(_0673_),
    .B1(_0506_));
 sg13g2_o21ai_1 _3503_ (.B1(_0541_),
    .Y(_0674_),
    .A1(_0526_),
    .A2(_0542_));
 sg13g2_a21oi_2 _3504_ (.B1(_0524_),
    .Y(_0675_),
    .A2(_0525_),
    .A1(_0517_));
 sg13g2_nor2b_1 _3505_ (.A(_0675_),
    .B_N(_0503_),
    .Y(_0676_));
 sg13g2_xnor2_1 _3506_ (.Y(_0677_),
    .A(_0503_),
    .B(_0675_));
 sg13g2_nand2_1 _3507_ (.Y(_0678_),
    .A(_0674_),
    .B(_0677_));
 sg13g2_xnor2_1 _3508_ (.Y(_0679_),
    .A(_0674_),
    .B(_0677_));
 sg13g2_xor2_1 _3509_ (.B(_0679_),
    .A(_0673_),
    .X(_0680_));
 sg13g2_nor2b_1 _3510_ (.A(_0672_),
    .B_N(_0680_),
    .Y(_0681_));
 sg13g2_xnor2_1 _3511_ (.Y(_0682_),
    .A(_0672_),
    .B(_0680_));
 sg13g2_xnor2_1 _3512_ (.Y(_0683_),
    .A(_0671_),
    .B(_0682_));
 sg13g2_o21ai_1 _3513_ (.B1(_0655_),
    .Y(_0684_),
    .A1(_0565_),
    .A2(_0656_));
 sg13g2_a21oi_1 _3514_ (.A1(_0543_),
    .A2(_0560_),
    .Y(_0685_),
    .B1(_0559_));
 sg13g2_a21oi_2 _3515_ (.B1(_0599_),
    .Y(_0686_),
    .A2(_0600_),
    .A1(_0567_));
 sg13g2_a21o_1 _3516_ (.A2(_0534_),
    .A1(_0238_),
    .B1(_0536_),
    .X(_0687_));
 sg13g2_o21ai_1 _3517_ (.B1(_0539_),
    .Y(_0688_),
    .A1(_0531_),
    .A2(_0537_));
 sg13g2_nand2_1 _3518_ (.Y(_0689_),
    .A(_0687_),
    .B(_0688_));
 sg13g2_xnor2_1 _3519_ (.Y(_0690_),
    .A(_0687_),
    .B(_0688_));
 sg13g2_o21ai_1 _3520_ (.B1(_0521_),
    .Y(_0691_),
    .A1(_0519_),
    .A2(_0522_));
 sg13g2_nor2_2 _3521_ (.A(_0529_),
    .B(_0691_),
    .Y(_0692_));
 sg13g2_xor2_1 _3522_ (.B(_0691_),
    .A(_0529_),
    .X(_0693_));
 sg13g2_xnor2_1 _3523_ (.Y(_0694_),
    .A(_0690_),
    .B(_0693_));
 sg13g2_o21ai_1 _3524_ (.B1(_0556_),
    .Y(_0695_),
    .A1(_0545_),
    .A2(_0557_));
 sg13g2_a21oi_1 _3525_ (.A1(_0547_),
    .A2(_0554_),
    .Y(_0696_),
    .B1(_0553_));
 sg13g2_o21ai_1 _3526_ (.B1(_0580_),
    .Y(_0697_),
    .A1(_0574_),
    .A2(_0581_));
 sg13g2_nor2_2 _3527_ (.A(_0571_),
    .B(_0573_),
    .Y(_0698_));
 sg13g2_nand2_1 _3528_ (.Y(_0699_),
    .A(_0549_),
    .B(_0698_));
 sg13g2_xnor2_1 _3529_ (.Y(_0700_),
    .A(_0549_),
    .B(_0698_));
 sg13g2_xor2_1 _3530_ (.B(_0700_),
    .A(_0697_),
    .X(_0701_));
 sg13g2_nor2b_1 _3531_ (.A(_0696_),
    .B_N(_0701_),
    .Y(_0702_));
 sg13g2_xnor2_1 _3532_ (.Y(_0703_),
    .A(_0696_),
    .B(_0701_));
 sg13g2_nand2_1 _3533_ (.Y(_0704_),
    .A(_0695_),
    .B(_0703_));
 sg13g2_xnor2_1 _3534_ (.Y(_0705_),
    .A(_0695_),
    .B(_0703_));
 sg13g2_xor2_1 _3535_ (.B(_0705_),
    .A(_0694_),
    .X(_0706_));
 sg13g2_nor2b_1 _3536_ (.A(_0686_),
    .B_N(_0706_),
    .Y(_0707_));
 sg13g2_xor2_1 _3537_ (.B(_0706_),
    .A(_0686_),
    .X(_0708_));
 sg13g2_nor2_1 _3538_ (.A(_0685_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_xnor2_1 _3539_ (.Y(_0710_),
    .A(_0685_),
    .B(_0708_));
 sg13g2_o21ai_1 _3540_ (.B1(_0652_),
    .Y(_0711_),
    .A1(_0601_),
    .A2(_0653_));
 sg13g2_nand2_2 _3541_ (.Y(_0712_),
    .A(_0595_),
    .B(_0597_));
 sg13g2_o21ai_1 _3542_ (.B1(_0619_),
    .Y(_0713_),
    .A1(_0603_),
    .A2(_0620_));
 sg13g2_o21ai_1 _3543_ (.B1(_0577_),
    .Y(_0714_),
    .A1(_0316_),
    .A2(_0578_));
 sg13g2_o21ai_1 _3544_ (.B1(_0591_),
    .Y(_0715_),
    .A1(_0584_),
    .A2(_0592_));
 sg13g2_o21ai_1 _3545_ (.B1(_0606_),
    .Y(_0716_),
    .A1(_0367_),
    .A2(_0607_));
 sg13g2_nor3_1 _3546_ (.A(_0587_),
    .B(_0588_),
    .C(_0716_),
    .Y(_0717_));
 sg13g2_xor2_1 _3547_ (.B(_0716_),
    .A(_0589_),
    .X(_0718_));
 sg13g2_and2_1 _3548_ (.A(_0715_),
    .B(_0718_),
    .X(_0719_));
 sg13g2_xor2_1 _3549_ (.B(_0718_),
    .A(_0715_),
    .X(_0720_));
 sg13g2_xnor2_1 _3550_ (.Y(_0721_),
    .A(_0714_),
    .B(_0720_));
 sg13g2_nor2b_1 _3551_ (.A(_0721_),
    .B_N(_0713_),
    .Y(_0722_));
 sg13g2_xnor2_1 _3552_ (.Y(_0723_),
    .A(_0713_),
    .B(_0721_));
 sg13g2_xnor2_1 _3553_ (.Y(_0724_),
    .A(_0712_),
    .B(_0723_));
 sg13g2_a21o_1 _3554_ (.A2(_0649_),
    .A1(_0621_),
    .B1(_0648_),
    .X(_0725_));
 sg13g2_a21oi_1 _3555_ (.A1(_0610_),
    .A2(_0615_),
    .Y(_0726_),
    .B1(_0617_));
 sg13g2_a21oi_1 _3556_ (.A1(_0623_),
    .A2(_0629_),
    .Y(_0727_),
    .B1(_0628_));
 sg13g2_a22oi_1 _3557_ (.Y(_0728_),
    .B1(_0614_),
    .B2(_0611_),
    .A2(_0613_),
    .A1(_0457_));
 sg13g2_nor2_1 _3558_ (.A(_0727_),
    .B(_0728_),
    .Y(_0729_));
 sg13g2_xnor2_1 _3559_ (.Y(_0730_),
    .A(_0727_),
    .B(_0728_));
 sg13g2_nor2_1 _3560_ (.A(_0726_),
    .B(_0730_),
    .Y(_0731_));
 sg13g2_xnor2_1 _3561_ (.Y(_0732_),
    .A(_0726_),
    .B(_0730_));
 sg13g2_o21ai_1 _3562_ (.B1(_0645_),
    .Y(_0733_),
    .A1(_0630_),
    .A2(_0646_));
 sg13g2_a21oi_2 _3563_ (.B1(_0642_),
    .Y(_0734_),
    .A2(_0643_),
    .A1(_0637_));
 sg13g2_or2_1 _3564_ (.X(_0735_),
    .B(_0734_),
    .A(_0639_));
 sg13g2_xnor2_1 _3565_ (.Y(_0736_),
    .A(_0639_),
    .B(_0734_));
 sg13g2_nor3_2 _3566_ (.A(_0626_),
    .B(_0634_),
    .C(_0636_),
    .Y(_0737_));
 sg13g2_o21ai_1 _3567_ (.B1(_0626_),
    .Y(_0738_),
    .A1(_0634_),
    .A2(_0636_));
 sg13g2_nor2b_1 _3568_ (.A(_0737_),
    .B_N(_0738_),
    .Y(_0739_));
 sg13g2_xnor2_1 _3569_ (.Y(_0740_),
    .A(_0736_),
    .B(_0739_));
 sg13g2_nand2b_1 _3570_ (.Y(_0741_),
    .B(_0733_),
    .A_N(_0740_));
 sg13g2_xor2_1 _3571_ (.B(_0740_),
    .A(_0733_),
    .X(_0742_));
 sg13g2_xnor2_1 _3572_ (.Y(_0743_),
    .A(_0732_),
    .B(_0742_));
 sg13g2_nand2b_1 _3573_ (.Y(_0744_),
    .B(_0725_),
    .A_N(_0743_));
 sg13g2_xor2_1 _3574_ (.B(_0743_),
    .A(_0725_),
    .X(_0745_));
 sg13g2_xor2_1 _3575_ (.B(_0745_),
    .A(_0724_),
    .X(_0746_));
 sg13g2_nand2_1 _3576_ (.Y(_0747_),
    .A(_0711_),
    .B(_0746_));
 sg13g2_xnor2_1 _3577_ (.Y(_0748_),
    .A(_0711_),
    .B(_0746_));
 sg13g2_xor2_1 _3578_ (.B(_0748_),
    .A(_0710_),
    .X(_0749_));
 sg13g2_nand2_1 _3579_ (.Y(_0750_),
    .A(_0684_),
    .B(_0749_));
 sg13g2_xnor2_1 _3580_ (.Y(_0751_),
    .A(_0684_),
    .B(_0749_));
 sg13g2_xor2_1 _3581_ (.B(_0751_),
    .A(_0683_),
    .X(_0752_));
 sg13g2_nand2_1 _3582_ (.Y(_0753_),
    .A(_0670_),
    .B(_0752_));
 sg13g2_xnor2_1 _3583_ (.Y(_0754_),
    .A(_0670_),
    .B(_0752_));
 sg13g2_xor2_1 _3584_ (.B(_0754_),
    .A(_0669_),
    .X(_0755_));
 sg13g2_nand2_1 _3585_ (.Y(_0756_),
    .A(_0668_),
    .B(_0755_));
 sg13g2_nor2_1 _3586_ (.A(_0668_),
    .B(_0755_),
    .Y(_0757_));
 sg13g2_xnor2_1 _3587_ (.Y(_0758_),
    .A(_0668_),
    .B(_0755_));
 sg13g2_o21ai_1 _3588_ (.B1(_0665_),
    .Y(_0759_),
    .A1(_0666_),
    .A2(_0667_));
 sg13g2_xnor2_1 _3589_ (.Y(uo_out[3]),
    .A(_0758_),
    .B(_0759_));
 sg13g2_a21oi_2 _3590_ (.B1(_0681_),
    .Y(_0760_),
    .A2(_0682_),
    .A1(_0671_));
 sg13g2_o21ai_1 _3591_ (.B1(_0750_),
    .Y(_0761_),
    .A1(_0683_),
    .A2(_0751_));
 sg13g2_o21ai_1 _3592_ (.B1(_0678_),
    .Y(_0762_),
    .A1(_0673_),
    .A2(_0679_));
 sg13g2_nor2_2 _3593_ (.A(_0707_),
    .B(_0709_),
    .Y(_0763_));
 sg13g2_nor2_1 _3594_ (.A(_0166_),
    .B(_0676_),
    .Y(_0764_));
 sg13g2_o21ai_1 _3595_ (.B1(_0689_),
    .Y(_0765_),
    .A1(_0690_),
    .A2(_0693_));
 sg13g2_nor2_1 _3596_ (.A(_0166_),
    .B(_0692_),
    .Y(_0766_));
 sg13g2_xnor2_1 _3597_ (.Y(_0767_),
    .A(_0166_),
    .B(_0692_));
 sg13g2_nand2b_1 _3598_ (.Y(_0768_),
    .B(_0765_),
    .A_N(_0767_));
 sg13g2_xor2_1 _3599_ (.B(_0767_),
    .A(_0765_),
    .X(_0769_));
 sg13g2_xor2_1 _3600_ (.B(_0769_),
    .A(_0764_),
    .X(_0770_));
 sg13g2_nor2b_1 _3601_ (.A(_0763_),
    .B_N(_0770_),
    .Y(_0771_));
 sg13g2_xnor2_1 _3602_ (.Y(_0772_),
    .A(_0763_),
    .B(_0770_));
 sg13g2_xnor2_1 _3603_ (.Y(_0773_),
    .A(_0762_),
    .B(_0772_));
 sg13g2_o21ai_1 _3604_ (.B1(_0747_),
    .Y(_0774_),
    .A1(_0710_),
    .A2(_0748_));
 sg13g2_o21ai_1 _3605_ (.B1(_0744_),
    .Y(_0775_),
    .A1(_0724_),
    .A2(_0745_));
 sg13g2_a21oi_1 _3606_ (.A1(_0714_),
    .A2(_0720_),
    .Y(_0776_),
    .B1(_0719_));
 sg13g2_nor2_1 _3607_ (.A(_0729_),
    .B(_0731_),
    .Y(_0777_));
 sg13g2_nor2_1 _3608_ (.A(_0717_),
    .B(_0777_),
    .Y(_0778_));
 sg13g2_xnor2_1 _3609_ (.Y(_0779_),
    .A(_0717_),
    .B(_0777_));
 sg13g2_nor2_1 _3610_ (.A(_0776_),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_xnor2_1 _3611_ (.Y(_0781_),
    .A(_0776_),
    .B(_0779_));
 sg13g2_o21ai_1 _3612_ (.B1(_0741_),
    .Y(_0782_),
    .A1(_0732_),
    .A2(_0742_));
 sg13g2_nand3_1 _3613_ (.B(_0734_),
    .C(_0737_),
    .A(_0639_),
    .Y(_0783_));
 sg13g2_o21ai_1 _3614_ (.B1(_0735_),
    .Y(_0784_),
    .A1(_0736_),
    .A2(_0739_));
 sg13g2_inv_1 _3615_ (.Y(_0785_),
    .A(_0784_));
 sg13g2_o21ai_1 _3616_ (.B1(_0783_),
    .Y(_0786_),
    .A1(_0737_),
    .A2(_0785_));
 sg13g2_nand2_1 _3617_ (.Y(_0787_),
    .A(_0782_),
    .B(_0786_));
 sg13g2_xnor2_1 _3618_ (.Y(_0788_),
    .A(_0782_),
    .B(_0786_));
 sg13g2_xnor2_1 _3619_ (.Y(_0789_),
    .A(_0781_),
    .B(_0788_));
 sg13g2_nand2b_1 _3620_ (.Y(_0790_),
    .B(_0775_),
    .A_N(_0789_));
 sg13g2_xor2_1 _3621_ (.B(_0789_),
    .A(_0775_),
    .X(_0791_));
 sg13g2_o21ai_1 _3622_ (.B1(_0704_),
    .Y(_0792_),
    .A1(_0694_),
    .A2(_0705_));
 sg13g2_a21oi_2 _3623_ (.B1(_0722_),
    .Y(_0793_),
    .A2(_0723_),
    .A1(_0712_));
 sg13g2_a21o_1 _3624_ (.A2(_0700_),
    .A1(_0697_),
    .B1(_0702_),
    .X(_0794_));
 sg13g2_nor2_1 _3625_ (.A(_0699_),
    .B(_0794_),
    .Y(_0795_));
 sg13g2_xor2_1 _3626_ (.B(_0794_),
    .A(_0699_),
    .X(_0796_));
 sg13g2_nor2_1 _3627_ (.A(_0793_),
    .B(_0796_),
    .Y(_0797_));
 sg13g2_nand2_1 _3628_ (.Y(_0798_),
    .A(_0793_),
    .B(_0796_));
 sg13g2_nand2b_1 _3629_ (.Y(_0799_),
    .B(_0798_),
    .A_N(_0797_));
 sg13g2_xor2_1 _3630_ (.B(_0799_),
    .A(_0792_),
    .X(_0800_));
 sg13g2_xor2_1 _3631_ (.B(_0800_),
    .A(_0791_),
    .X(_0801_));
 sg13g2_nand2_1 _3632_ (.Y(_0802_),
    .A(_0774_),
    .B(_0801_));
 sg13g2_xnor2_1 _3633_ (.Y(_0803_),
    .A(_0774_),
    .B(_0801_));
 sg13g2_xor2_1 _3634_ (.B(_0803_),
    .A(_0773_),
    .X(_0804_));
 sg13g2_nand2_1 _3635_ (.Y(_0805_),
    .A(_0761_),
    .B(_0804_));
 sg13g2_xnor2_1 _3636_ (.Y(_0806_),
    .A(_0761_),
    .B(_0804_));
 sg13g2_or2_1 _3637_ (.X(_0807_),
    .B(_0806_),
    .A(_0760_));
 sg13g2_xor2_1 _3638_ (.B(_0806_),
    .A(_0760_),
    .X(_0808_));
 sg13g2_o21ai_1 _3639_ (.B1(_0753_),
    .Y(_0809_),
    .A1(_0669_),
    .A2(_0754_));
 sg13g2_and2_1 _3640_ (.A(_0808_),
    .B(_0809_),
    .X(_0810_));
 sg13g2_xor2_1 _3641_ (.B(_0809_),
    .A(_0808_),
    .X(_0811_));
 sg13g2_or2_1 _3642_ (.X(_0812_),
    .B(_0758_),
    .A(_0666_));
 sg13g2_a21o_1 _3643_ (.A2(_0756_),
    .A1(_0665_),
    .B1(_0757_),
    .X(_0813_));
 sg13g2_o21ai_1 _3644_ (.B1(_0813_),
    .Y(_0814_),
    .A1(_0667_),
    .A2(_0812_));
 sg13g2_xor2_1 _3645_ (.B(_0814_),
    .A(_0811_),
    .X(uo_out[4]));
 sg13g2_a21oi_2 _3646_ (.B1(_0771_),
    .Y(_0815_),
    .A2(_0772_),
    .A1(_0762_));
 sg13g2_o21ai_1 _3647_ (.B1(_0802_),
    .Y(_0816_),
    .A1(_0773_),
    .A2(_0803_));
 sg13g2_o21ai_1 _3648_ (.B1(_0768_),
    .Y(_0817_),
    .A1(_0764_),
    .A2(_0769_));
 sg13g2_a21oi_2 _3649_ (.B1(_0797_),
    .Y(_0818_),
    .A2(_0798_),
    .A1(_0792_));
 sg13g2_nor2_1 _3650_ (.A(_0766_),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_nand2_1 _3651_ (.Y(_0820_),
    .A(_0766_),
    .B(_0818_));
 sg13g2_nor2b_1 _3652_ (.A(_0819_),
    .B_N(_0820_),
    .Y(_0821_));
 sg13g2_xnor2_1 _3653_ (.Y(_0822_),
    .A(_0817_),
    .B(_0821_));
 sg13g2_o21ai_1 _3654_ (.B1(_0790_),
    .Y(_0823_),
    .A1(_0791_),
    .A2(_0800_));
 sg13g2_nor2_2 _3655_ (.A(_0778_),
    .B(_0780_),
    .Y(_0824_));
 sg13g2_and2_2 _3656_ (.A(_0795_),
    .B(_0824_),
    .X(_0825_));
 sg13g2_xnor2_1 _3657_ (.Y(_0826_),
    .A(_0795_),
    .B(_0824_));
 sg13g2_o21ai_1 _3658_ (.B1(_0787_),
    .Y(_0827_),
    .A1(_0781_),
    .A2(_0788_));
 sg13g2_and2_1 _3659_ (.A(_0783_),
    .B(_0827_),
    .X(_0828_));
 sg13g2_xor2_1 _3660_ (.B(_0827_),
    .A(_0783_),
    .X(_0829_));
 sg13g2_xnor2_1 _3661_ (.Y(_0830_),
    .A(_0826_),
    .B(_0829_));
 sg13g2_nand2b_1 _3662_ (.Y(_0831_),
    .B(_0823_),
    .A_N(_0830_));
 sg13g2_xor2_1 _3663_ (.B(_0830_),
    .A(_0823_),
    .X(_0832_));
 sg13g2_xor2_1 _3664_ (.B(_0832_),
    .A(_0822_),
    .X(_0833_));
 sg13g2_nand2_1 _3665_ (.Y(_0834_),
    .A(_0816_),
    .B(_0833_));
 sg13g2_xnor2_1 _3666_ (.Y(_0835_),
    .A(_0816_),
    .B(_0833_));
 sg13g2_xnor2_1 _3667_ (.Y(_0836_),
    .A(_0815_),
    .B(_0835_));
 sg13g2_a21oi_1 _3668_ (.A1(_0805_),
    .A2(_0807_),
    .Y(_0837_),
    .B1(_0836_));
 sg13g2_nand3_1 _3669_ (.B(_0807_),
    .C(_0836_),
    .A(_0805_),
    .Y(_0838_));
 sg13g2_nor2b_1 _3670_ (.A(_0837_),
    .B_N(_0838_),
    .Y(_0839_));
 sg13g2_a21oi_1 _3671_ (.A1(_0811_),
    .A2(_0814_),
    .Y(_0840_),
    .B1(_0810_));
 sg13g2_xnor2_1 _3672_ (.Y(uo_out[5]),
    .A(_0839_),
    .B(_0840_));
 sg13g2_a21oi_1 _3673_ (.A1(_0817_),
    .A2(_0820_),
    .Y(_0841_),
    .B1(_0819_));
 sg13g2_o21ai_1 _3674_ (.B1(_0831_),
    .Y(_0842_),
    .A1(_0822_),
    .A2(_0832_));
 sg13g2_a21oi_2 _3675_ (.B1(_0828_),
    .Y(_0843_),
    .A2(_0829_),
    .A1(_0826_));
 sg13g2_xor2_1 _3676_ (.B(_0825_),
    .A(_0766_),
    .X(_0844_));
 sg13g2_xnor2_1 _3677_ (.Y(_0845_),
    .A(_0843_),
    .B(_0844_));
 sg13g2_xnor2_1 _3678_ (.Y(_0846_),
    .A(_0842_),
    .B(_0845_));
 sg13g2_nor2_1 _3679_ (.A(_0841_),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_xnor2_1 _3680_ (.Y(_0848_),
    .A(_0841_),
    .B(_0846_));
 sg13g2_o21ai_1 _3681_ (.B1(_0834_),
    .Y(_0849_),
    .A1(_0815_),
    .A2(_0835_));
 sg13g2_nor2b_1 _3682_ (.A(_0848_),
    .B_N(_0849_),
    .Y(_0850_));
 sg13g2_xnor2_1 _3683_ (.Y(_0851_),
    .A(_0848_),
    .B(_0849_));
 sg13g2_and2_1 _3684_ (.A(_0811_),
    .B(_0839_),
    .X(_0852_));
 sg13g2_nand2_1 _3685_ (.Y(_0853_),
    .A(_0810_),
    .B(_0838_));
 sg13g2_nand2b_1 _3686_ (.Y(_0854_),
    .B(_0853_),
    .A_N(_0837_));
 sg13g2_a21o_1 _3687_ (.A2(_0852_),
    .A1(_0814_),
    .B1(_0854_),
    .X(_0855_));
 sg13g2_xor2_1 _3688_ (.B(_0855_),
    .A(_0851_),
    .X(uo_out[6]));
 sg13g2_a21oi_1 _3689_ (.A1(_0851_),
    .A2(_0855_),
    .Y(_0856_),
    .B1(_0850_));
 sg13g2_a21oi_1 _3690_ (.A1(_0842_),
    .A2(_0845_),
    .Y(_0857_),
    .B1(_0847_));
 sg13g2_nor4_2 _3691_ (.A(_0166_),
    .B(_0692_),
    .C(_0825_),
    .Y(_0858_),
    .D(_0843_));
 sg13g2_nor2b_1 _3692_ (.A(_0857_),
    .B_N(_0858_),
    .Y(_0859_));
 sg13g2_xnor2_1 _3693_ (.Y(_0860_),
    .A(_0857_),
    .B(_0858_));
 sg13g2_xnor2_1 _3694_ (.Y(uo_out[7]),
    .A(_0856_),
    .B(_0860_));
 sg13g2_and2_1 _3695_ (.A(_0851_),
    .B(_0860_),
    .X(_0861_));
 sg13g2_a221oi_1 _3696_ (.B2(_0855_),
    .C1(_0859_),
    .B1(_0861_),
    .A1(_0850_),
    .Y(uio_out[7]),
    .A2(_0860_));
 sg13g2_dfrbp_1 _3697_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net11),
    .D(net4),
    .Q_N(_1589_),
    .Q(\i_w_buf[0].A ));
 sg13g2_dfrbp_1 _3698_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net12),
    .D(net5),
    .Q_N(_1590_),
    .Q(\i_w_buf[1].A ));
 sg13g2_dfrbp_1 _3699_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net13),
    .D(net438),
    .Q_N(_1591_),
    .Q(\i_w_buf[2].A ));
 sg13g2_dfrbp_1 _3700_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net14),
    .D(net473),
    .Q_N(_1592_),
    .Q(\i_w_buf[3].A ));
 sg13g2_dfrbp_1 _3701_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net15),
    .D(net325),
    .Q_N(_1593_),
    .Q(\i_w_buf[4].A ));
 sg13g2_dfrbp_1 _3702_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net16),
    .D(net448),
    .Q_N(_1594_),
    .Q(\i_w_buf[5].A ));
 sg13g2_dfrbp_1 _3703_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net17),
    .D(net359),
    .Q_N(_1595_),
    .Q(\i_w_buf[6].A ));
 sg13g2_dfrbp_1 _3704_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net18),
    .D(net446),
    .Q_N(_1596_),
    .Q(\i_w_buf[7].A ));
 sg13g2_dfrbp_1 _3705_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net19),
    .D(net417),
    .Q_N(_1597_),
    .Q(\i_w_buf[8].A ));
 sg13g2_dfrbp_1 _3706_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net20),
    .D(net509),
    .Q_N(_1598_),
    .Q(\i_w_buf[9].A ));
 sg13g2_dfrbp_1 _3707_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net21),
    .D(net319),
    .Q_N(_1599_),
    .Q(\i_w_buf[10].A ));
 sg13g2_dfrbp_1 _3708_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net22),
    .D(net402),
    .Q_N(_1600_),
    .Q(\i_w_buf[11].A ));
 sg13g2_dfrbp_1 _3709_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net23),
    .D(net302),
    .Q_N(_1601_),
    .Q(\i_w_buf[12].A ));
 sg13g2_dfrbp_1 _3710_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net24),
    .D(net463),
    .Q_N(_1602_),
    .Q(\i_w_buf[13].A ));
 sg13g2_dfrbp_1 _3711_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net25),
    .D(net539),
    .Q_N(_1603_),
    .Q(\i_w_buf[14].A ));
 sg13g2_dfrbp_1 _3712_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net26),
    .D(net551),
    .Q_N(_1604_),
    .Q(\i_w_buf[15].A ));
 sg13g2_dfrbp_1 _3713_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net27),
    .D(net316),
    .Q_N(_1605_),
    .Q(\i_w_buf[16].A ));
 sg13g2_dfrbp_1 _3714_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net28),
    .D(net334),
    .Q_N(_1606_),
    .Q(\i_w_buf[17].A ));
 sg13g2_dfrbp_1 _3715_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net29),
    .D(net385),
    .Q_N(_1607_),
    .Q(\i_w_buf[18].A ));
 sg13g2_dfrbp_1 _3716_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net30),
    .D(net435),
    .Q_N(_1608_),
    .Q(\i_w_buf[19].A ));
 sg13g2_dfrbp_1 _3717_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net31),
    .D(net545),
    .Q_N(_1609_),
    .Q(\i_w_buf[20].A ));
 sg13g2_dfrbp_1 _3718_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net32),
    .D(net512),
    .Q_N(_1610_),
    .Q(\i_w_buf[21].A ));
 sg13g2_dfrbp_1 _3719_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net33),
    .D(net313),
    .Q_N(_1611_),
    .Q(\i_w_buf[22].A ));
 sg13g2_dfrbp_1 _3720_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net34),
    .D(net503),
    .Q_N(_1612_),
    .Q(\i_w_buf[23].A ));
 sg13g2_dfrbp_1 _3721_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net35),
    .D(net335),
    .Q_N(_1613_),
    .Q(\i_w_buf[24].A ));
 sg13g2_dfrbp_1 _3722_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net36),
    .D(net437),
    .Q_N(_1614_),
    .Q(\i_w_buf[25].A ));
 sg13g2_dfrbp_1 _3723_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net37),
    .D(net372),
    .Q_N(_1615_),
    .Q(\i_w_buf[26].A ));
 sg13g2_dfrbp_1 _3724_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net38),
    .D(net368),
    .Q_N(_1616_),
    .Q(\i_w_buf[27].A ));
 sg13g2_dfrbp_1 _3725_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net39),
    .D(net386),
    .Q_N(_1617_),
    .Q(\i_w_buf[28].A ));
 sg13g2_dfrbp_1 _3726_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net40),
    .D(net413),
    .Q_N(_1618_),
    .Q(\i_w_buf[29].A ));
 sg13g2_dfrbp_1 _3727_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net41),
    .D(net500),
    .Q_N(_1619_),
    .Q(\i_w_buf[30].A ));
 sg13g2_dfrbp_1 _3728_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net42),
    .D(net525),
    .Q_N(_1620_),
    .Q(\i_w_buf[31].A ));
 sg13g2_dfrbp_1 _3729_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net43),
    .D(net351),
    .Q_N(_1621_),
    .Q(\i_w_buf[32].A ));
 sg13g2_dfrbp_1 _3730_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net44),
    .D(net462),
    .Q_N(_1622_),
    .Q(\i_w_buf[33].A ));
 sg13g2_dfrbp_1 _3731_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net45),
    .D(net471),
    .Q_N(_1623_),
    .Q(\i_w_buf[34].A ));
 sg13g2_dfrbp_1 _3732_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net46),
    .D(net429),
    .Q_N(_1624_),
    .Q(\i_w_buf[35].A ));
 sg13g2_dfrbp_1 _3733_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net47),
    .D(net332),
    .Q_N(_1625_),
    .Q(\i_w_buf[36].A ));
 sg13g2_dfrbp_1 _3734_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net48),
    .D(net384),
    .Q_N(_1626_),
    .Q(\i_w_buf[37].A ));
 sg13g2_dfrbp_1 _3735_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net49),
    .D(net514),
    .Q_N(_1627_),
    .Q(\i_w_buf[38].A ));
 sg13g2_dfrbp_1 _3736_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net50),
    .D(net534),
    .Q_N(_1628_),
    .Q(\i_w_buf[39].A ));
 sg13g2_dfrbp_1 _3737_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net51),
    .D(net329),
    .Q_N(_1629_),
    .Q(\i_w_buf[40].A ));
 sg13g2_dfrbp_1 _3738_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net52),
    .D(net461),
    .Q_N(_1630_),
    .Q(\i_w_buf[41].A ));
 sg13g2_dfrbp_1 _3739_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net53),
    .D(net541),
    .Q_N(_1631_),
    .Q(\i_w_buf[42].A ));
 sg13g2_dfrbp_1 _3740_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net54),
    .D(net544),
    .Q_N(_1632_),
    .Q(\i_w_buf[43].A ));
 sg13g2_dfrbp_1 _3741_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net55),
    .D(net381),
    .Q_N(_1633_),
    .Q(\i_w_buf[44].A ));
 sg13g2_dfrbp_1 _3742_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net56),
    .D(net409),
    .Q_N(_1634_),
    .Q(\i_w_buf[45].A ));
 sg13g2_dfrbp_1 _3743_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net57),
    .D(net479),
    .Q_N(_1635_),
    .Q(\i_w_buf[46].A ));
 sg13g2_dfrbp_1 _3744_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net58),
    .D(net445),
    .Q_N(_1636_),
    .Q(\i_w_buf[47].A ));
 sg13g2_dfrbp_1 _3745_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net59),
    .D(net374),
    .Q_N(_1637_),
    .Q(\i_w_buf[48].A ));
 sg13g2_dfrbp_1 _3746_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net60),
    .D(net455),
    .Q_N(_1638_),
    .Q(\i_w_buf[49].A ));
 sg13g2_dfrbp_1 _3747_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net61),
    .D(net538),
    .Q_N(_1639_),
    .Q(\i_w_buf[50].A ));
 sg13g2_dfrbp_1 _3748_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net62),
    .D(net441),
    .Q_N(_1640_),
    .Q(\i_w_buf[51].A ));
 sg13g2_dfrbp_1 _3749_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net63),
    .D(net442),
    .Q_N(_1641_),
    .Q(\i_w_buf[52].A ));
 sg13g2_dfrbp_1 _3750_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net64),
    .D(net533),
    .Q_N(_1642_),
    .Q(\i_w_buf[53].A ));
 sg13g2_dfrbp_1 _3751_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net65),
    .D(net345),
    .Q_N(_1643_),
    .Q(\i_w_buf[54].A ));
 sg13g2_dfrbp_1 _3752_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net66),
    .D(net347),
    .Q_N(_1644_),
    .Q(\i_w_buf[55].A ));
 sg13g2_dfrbp_1 _3753_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net67),
    .D(net449),
    .Q_N(_1645_),
    .Q(\i_w_buf[56].A ));
 sg13g2_dfrbp_1 _3754_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net68),
    .D(net491),
    .Q_N(_1646_),
    .Q(\i_w_buf[57].A ));
 sg13g2_dfrbp_1 _3755_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net69),
    .D(net364),
    .Q_N(_1647_),
    .Q(\i_w_buf[58].A ));
 sg13g2_dfrbp_1 _3756_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net70),
    .D(net458),
    .Q_N(_1648_),
    .Q(\i_w_buf[59].A ));
 sg13g2_dfrbp_1 _3757_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net71),
    .D(net492),
    .Q_N(_1649_),
    .Q(\i_w_buf[60].A ));
 sg13g2_dfrbp_1 _3758_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net72),
    .D(net481),
    .Q_N(_1650_),
    .Q(\i_w_buf[61].A ));
 sg13g2_dfrbp_1 _3759_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net73),
    .D(net444),
    .Q_N(_1651_),
    .Q(\i_w_buf[62].A ));
 sg13g2_dfrbp_1 _3760_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net74),
    .D(net460),
    .Q_N(_1652_),
    .Q(\i_w_buf[63].A ));
 sg13g2_dfrbp_1 _3761_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net75),
    .D(net308),
    .Q_N(_1653_),
    .Q(\i_w_buf[64].A ));
 sg13g2_dfrbp_1 _3762_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net76),
    .D(net376),
    .Q_N(_1654_),
    .Q(\i_w_buf[65].A ));
 sg13g2_dfrbp_1 _3763_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net77),
    .D(net548),
    .Q_N(_1655_),
    .Q(\i_w_buf[66].A ));
 sg13g2_dfrbp_1 _3764_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net78),
    .D(net546),
    .Q_N(_1656_),
    .Q(\i_w_buf[67].A ));
 sg13g2_dfrbp_1 _3765_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net79),
    .D(net337),
    .Q_N(_1657_),
    .Q(\i_w_buf[68].A ));
 sg13g2_dfrbp_1 _3766_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net108),
    .D(net552),
    .Q_N(_1658_),
    .Q(\i_w_buf[69].A ));
 sg13g2_dfrbp_1 _3767_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net109),
    .D(net497),
    .Q_N(_1659_),
    .Q(\i_w_buf[70].A ));
 sg13g2_dfrbp_1 _3768_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net110),
    .D(net299),
    .Q_N(_1660_),
    .Q(\i_w_buf[71].A ));
 sg13g2_dfrbp_1 _3769_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net111),
    .D(net474),
    .Q_N(_1661_),
    .Q(\i_w_buf[72].A ));
 sg13g2_dfrbp_1 _3770_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net112),
    .D(net485),
    .Q_N(_1662_),
    .Q(\i_w_buf[73].A ));
 sg13g2_dfrbp_1 _3771_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net113),
    .D(net516),
    .Q_N(_1663_),
    .Q(\i_w_buf[74].A ));
 sg13g2_dfrbp_1 _3772_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net114),
    .D(net505),
    .Q_N(_1664_),
    .Q(\i_w_buf[75].A ));
 sg13g2_dfrbp_1 _3773_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net115),
    .D(net380),
    .Q_N(_1665_),
    .Q(\i_w_buf[76].A ));
 sg13g2_dfrbp_1 _3774_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net116),
    .D(net432),
    .Q_N(_1666_),
    .Q(\i_w_buf[77].A ));
 sg13g2_dfrbp_1 _3775_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net117),
    .D(net542),
    .Q_N(_1667_),
    .Q(\i_w_buf[78].A ));
 sg13g2_dfrbp_1 _3776_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net118),
    .D(net532),
    .Q_N(_1668_),
    .Q(\i_w_buf[79].A ));
 sg13g2_dfrbp_1 _3777_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net119),
    .D(net331),
    .Q_N(_1669_),
    .Q(\i_w_buf[80].A ));
 sg13g2_dfrbp_1 _3778_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net120),
    .D(net377),
    .Q_N(_1670_),
    .Q(\i_w_buf[81].A ));
 sg13g2_dfrbp_1 _3779_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net121),
    .D(net482),
    .Q_N(_1671_),
    .Q(\i_w_buf[82].A ));
 sg13g2_dfrbp_1 _3780_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net122),
    .D(net452),
    .Q_N(_1672_),
    .Q(\i_w_buf[83].A ));
 sg13g2_dfrbp_1 _3781_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net123),
    .D(net312),
    .Q_N(_1673_),
    .Q(\i_w_buf[84].A ));
 sg13g2_dfrbp_1 _3782_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net124),
    .D(net416),
    .Q_N(_1674_),
    .Q(\i_w_buf[85].A ));
 sg13g2_dfrbp_1 _3783_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net125),
    .D(net401),
    .Q_N(_1675_),
    .Q(\i_w_buf[86].A ));
 sg13g2_dfrbp_1 _3784_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net126),
    .D(net427),
    .Q_N(_1676_),
    .Q(\i_w_buf[87].A ));
 sg13g2_dfrbp_1 _3785_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net127),
    .D(net499),
    .Q_N(_1677_),
    .Q(\i_w_buf[88].A ));
 sg13g2_dfrbp_1 _3786_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net128),
    .D(net522),
    .Q_N(_1678_),
    .Q(\i_w_buf[89].A ));
 sg13g2_dfrbp_1 _3787_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net129),
    .D(net333),
    .Q_N(_1679_),
    .Q(\i_w_buf[90].A ));
 sg13g2_dfrbp_1 _3788_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net130),
    .D(net483),
    .Q_N(_1680_),
    .Q(\i_w_buf[91].A ));
 sg13g2_dfrbp_1 _3789_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net131),
    .D(net511),
    .Q_N(_1681_),
    .Q(\i_w_buf[92].A ));
 sg13g2_dfrbp_1 _3790_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net132),
    .D(net484),
    .Q_N(_1682_),
    .Q(\i_w_buf[93].A ));
 sg13g2_dfrbp_1 _3791_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net133),
    .D(net301),
    .Q_N(_1683_),
    .Q(\i_w_buf[94].A ));
 sg13g2_dfrbp_1 _3792_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net134),
    .D(net470),
    .Q_N(_1684_),
    .Q(\i_w_buf[95].A ));
 sg13g2_dfrbp_1 _3793_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net135),
    .D(net493),
    .Q_N(_1685_),
    .Q(\i_w_buf[96].A ));
 sg13g2_dfrbp_1 _3794_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net136),
    .D(net355),
    .Q_N(_1686_),
    .Q(\i_w_buf[97].A ));
 sg13g2_dfrbp_1 _3795_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net137),
    .D(net305),
    .Q_N(_1687_),
    .Q(\i_w_buf[98].A ));
 sg13g2_dfrbp_1 _3796_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net138),
    .D(net447),
    .Q_N(_1688_),
    .Q(\i_w_buf[99].A ));
 sg13g2_dfrbp_1 _3797_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net139),
    .D(net344),
    .Q_N(_1689_),
    .Q(\i_w_buf[100].A ));
 sg13g2_dfrbp_1 _3798_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net140),
    .D(net450),
    .Q_N(_1690_),
    .Q(\i_w_buf[101].A ));
 sg13g2_dfrbp_1 _3799_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net141),
    .D(net550),
    .Q_N(_1691_),
    .Q(\i_w_buf[102].A ));
 sg13g2_dfrbp_1 _3800_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net142),
    .D(net549),
    .Q_N(_1692_),
    .Q(\i_w_buf[103].A ));
 sg13g2_dfrbp_1 _3801_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net143),
    .D(net487),
    .Q_N(_1693_),
    .Q(\i_w_buf[104].A ));
 sg13g2_dfrbp_1 _3802_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net144),
    .D(net498),
    .Q_N(_1694_),
    .Q(\i_w_buf[105].A ));
 sg13g2_dfrbp_1 _3803_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net145),
    .D(net309),
    .Q_N(_1695_),
    .Q(\i_w_buf[106].A ));
 sg13g2_dfrbp_1 _3804_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net146),
    .D(net378),
    .Q_N(_1696_),
    .Q(\i_w_buf[107].A ));
 sg13g2_dfrbp_1 _3805_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net147),
    .D(net324),
    .Q_N(_1697_),
    .Q(\i_w_buf[108].A ));
 sg13g2_dfrbp_1 _3806_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net148),
    .D(net440),
    .Q_N(_1698_),
    .Q(\i_w_buf[109].A ));
 sg13g2_dfrbp_1 _3807_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net149),
    .D(net453),
    .Q_N(_1699_),
    .Q(\i_w_buf[110].A ));
 sg13g2_dfrbp_1 _3808_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net150),
    .D(net547),
    .Q_N(_1700_),
    .Q(\i_w_buf[111].A ));
 sg13g2_dfrbp_1 _3809_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net151),
    .D(net502),
    .Q_N(_1701_),
    .Q(\i_w_buf[112].A ));
 sg13g2_dfrbp_1 _3810_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net152),
    .D(net530),
    .Q_N(_1702_),
    .Q(\i_w_buf[113].A ));
 sg13g2_dfrbp_1 _3811_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net153),
    .D(net354),
    .Q_N(_1703_),
    .Q(\i_w_buf[114].A ));
 sg13g2_dfrbp_1 _3812_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net154),
    .D(net340),
    .Q_N(_1704_),
    .Q(\i_w_buf[115].A ));
 sg13g2_dfrbp_1 _3813_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net155),
    .D(net348),
    .Q_N(_1705_),
    .Q(\i_w_buf[116].A ));
 sg13g2_dfrbp_1 _3814_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net156),
    .D(net395),
    .Q_N(_1706_),
    .Q(\i_w_buf[117].A ));
 sg13g2_dfrbp_1 _3815_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net157),
    .D(net400),
    .Q_N(_1707_),
    .Q(\i_w_buf[118].A ));
 sg13g2_dfrbp_1 _3816_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net158),
    .D(net397),
    .Q_N(_1708_),
    .Q(\i_w_buf[119].A ));
 sg13g2_dfrbp_1 _3817_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net159),
    .D(net391),
    .Q_N(_1709_),
    .Q(\i_w_buf[120].A ));
 sg13g2_dfrbp_1 _3818_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net160),
    .D(net504),
    .Q_N(_1710_),
    .Q(\i_w_buf[121].A ));
 sg13g2_dfrbp_1 _3819_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net161),
    .D(net320),
    .Q_N(_1711_),
    .Q(\i_w_buf[122].A ));
 sg13g2_dfrbp_1 _3820_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net162),
    .D(net404),
    .Q_N(_1712_),
    .Q(\i_w_buf[123].A ));
 sg13g2_dfrbp_1 _3821_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net163),
    .D(net508),
    .Q_N(_1713_),
    .Q(\i_w_buf[124].A ));
 sg13g2_dfrbp_1 _3822_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net164),
    .D(net513),
    .Q_N(_1714_),
    .Q(\i_w_buf[125].A ));
 sg13g2_dfrbp_1 _3823_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net165),
    .D(net420),
    .Q_N(_1715_),
    .Q(\i_w_buf[126].A ));
 sg13g2_dfrbp_1 _3824_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net166),
    .D(net507),
    .Q_N(_1716_),
    .Q(\i_w_buf[127].A ));
 sg13g2_dfrbp_1 _3825_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net167),
    .D(net528),
    .Q_N(_1717_),
    .Q(\i_w_buf[128].A ));
 sg13g2_dfrbp_1 _3826_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net168),
    .D(net535),
    .Q_N(_1718_),
    .Q(\i_w_buf[129].A ));
 sg13g2_dfrbp_1 _3827_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net169),
    .D(net352),
    .Q_N(_1719_),
    .Q(\i_w_buf[130].A ));
 sg13g2_dfrbp_1 _3828_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net170),
    .D(net421),
    .Q_N(_1720_),
    .Q(\i_w_buf[131].A ));
 sg13g2_dfrbp_1 _3829_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net171),
    .D(net478),
    .Q_N(_1721_),
    .Q(\i_w_buf[132].A ));
 sg13g2_dfrbp_1 _3830_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net172),
    .D(net469),
    .Q_N(_1722_),
    .Q(\i_w_buf[133].A ));
 sg13g2_dfrbp_1 _3831_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net173),
    .D(net306),
    .Q_N(_1723_),
    .Q(\i_w_buf[134].A ));
 sg13g2_dfrbp_1 _3832_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net174),
    .D(net424),
    .Q_N(_1724_),
    .Q(\i_w_buf[135].A ));
 sg13g2_dfrbp_1 _3833_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net175),
    .D(net520),
    .Q_N(_1725_),
    .Q(\i_w_buf[136].A ));
 sg13g2_dfrbp_1 _3834_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net176),
    .D(net529),
    .Q_N(_1726_),
    .Q(\i_w_buf[137].A ));
 sg13g2_dfrbp_1 _3835_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net177),
    .D(net303),
    .Q_N(_1727_),
    .Q(\i_w_buf[138].A ));
 sg13g2_dfrbp_1 _3836_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net178),
    .D(net439),
    .Q_N(_1728_),
    .Q(\i_w_buf[139].A ));
 sg13g2_dfrbp_1 _3837_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net179),
    .D(net490),
    .Q_N(_1729_),
    .Q(\i_w_buf[140].A ));
 sg13g2_dfrbp_1 _3838_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net180),
    .D(net363),
    .Q_N(_1730_),
    .Q(\i_w_buf[141].A ));
 sg13g2_dfrbp_1 _3839_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net181),
    .D(net468),
    .Q_N(_1731_),
    .Q(\i_w_buf[142].A ));
 sg13g2_dfrbp_1 _3840_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net182),
    .D(net488),
    .Q_N(_1732_),
    .Q(\i_w_buf[143].A ));
 sg13g2_dfrbp_1 _3841_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net183),
    .D(net370),
    .Q_N(_1733_),
    .Q(\i_w_buf[144].A ));
 sg13g2_dfrbp_1 _3842_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net184),
    .D(net521),
    .Q_N(_1734_),
    .Q(\i_w_buf[145].A ));
 sg13g2_dfrbp_1 _3843_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net185),
    .D(net361),
    .Q_N(_1735_),
    .Q(\i_w_buf[146].A ));
 sg13g2_dfrbp_1 _3844_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net186),
    .D(net362),
    .Q_N(_1736_),
    .Q(\i_w_buf[147].A ));
 sg13g2_dfrbp_1 _3845_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net187),
    .D(net367),
    .Q_N(_1737_),
    .Q(\i_w_buf[148].A ));
 sg13g2_dfrbp_1 _3846_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net188),
    .D(net480),
    .Q_N(_1738_),
    .Q(\i_w_buf[149].A ));
 sg13g2_dfrbp_1 _3847_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net189),
    .D(net410),
    .Q_N(_1739_),
    .Q(\i_w_buf[150].A ));
 sg13g2_dfrbp_1 _3848_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net190),
    .D(net477),
    .Q_N(_1740_),
    .Q(\i_w_buf[151].A ));
 sg13g2_dfrbp_1 _3849_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net191),
    .D(net486),
    .Q_N(_1741_),
    .Q(\i_w_buf[152].A ));
 sg13g2_dfrbp_1 _3850_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net192),
    .D(net523),
    .Q_N(_1742_),
    .Q(\i_w_buf[153].A ));
 sg13g2_dfrbp_1 _3851_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net193),
    .D(net518),
    .Q_N(_1743_),
    .Q(\i_w_buf[154].A ));
 sg13g2_dfrbp_1 _3852_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net194),
    .D(net433),
    .Q_N(_1744_),
    .Q(\i_w_buf[155].A ));
 sg13g2_dfrbp_1 _3853_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net195),
    .D(net406),
    .Q_N(_1745_),
    .Q(\i_w_buf[156].A ));
 sg13g2_dfrbp_1 _3854_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net196),
    .D(net506),
    .Q_N(_1746_),
    .Q(\i_w_buf[157].A ));
 sg13g2_dfrbp_1 _3855_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net197),
    .D(net451),
    .Q_N(_1747_),
    .Q(\i_w_buf[158].A ));
 sg13g2_dfrbp_1 _3856_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net198),
    .D(net466),
    .Q_N(_1748_),
    .Q(\i_w_buf[159].A ));
 sg13g2_dfrbp_1 _3857_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net199),
    .D(net373),
    .Q_N(_1749_),
    .Q(\i_w_buf[160].A ));
 sg13g2_dfrbp_1 _3858_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net200),
    .D(net357),
    .Q_N(_1750_),
    .Q(\i_w_buf[161].A ));
 sg13g2_dfrbp_1 _3859_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net201),
    .D(net343),
    .Q_N(_1751_),
    .Q(\i_w_buf[162].A ));
 sg13g2_dfrbp_1 _3860_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net202),
    .D(net387),
    .Q_N(_1752_),
    .Q(\i_w_buf[163].A ));
 sg13g2_dfrbp_1 _3861_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net203),
    .D(net537),
    .Q_N(_1753_),
    .Q(\i_w_buf[164].A ));
 sg13g2_dfrbp_1 _3862_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net204),
    .D(net543),
    .Q_N(_1754_),
    .Q(\i_w_buf[165].A ));
 sg13g2_dfrbp_1 _3863_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net205),
    .D(net311),
    .Q_N(_1755_),
    .Q(\i_w_buf[166].A ));
 sg13g2_dfrbp_1 _3864_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net206),
    .D(net393),
    .Q_N(_1756_),
    .Q(\i_w_buf[167].A ));
 sg13g2_dfrbp_1 _3865_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net207),
    .D(net495),
    .Q_N(_1757_),
    .Q(\i_w_buf[168].A ));
 sg13g2_dfrbp_1 _3866_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net208),
    .D(net524),
    .Q_N(_1758_),
    .Q(\i_w_buf[169].A ));
 sg13g2_dfrbp_1 _3867_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net209),
    .D(net317),
    .Q_N(_1759_),
    .Q(\i_w_buf[170].A ));
 sg13g2_dfrbp_1 _3868_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net210),
    .D(net392),
    .Q_N(_1760_),
    .Q(\i_w_buf[171].A ));
 sg13g2_dfrbp_1 _3869_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net211),
    .D(net338),
    .Q_N(_1761_),
    .Q(\i_w_buf[172].A ));
 sg13g2_dfrbp_1 _3870_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net212),
    .D(net412),
    .Q_N(_1762_),
    .Q(\i_w_buf[173].A ));
 sg13g2_dfrbp_1 _3871_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net213),
    .D(net328),
    .Q_N(_1763_),
    .Q(\i_w_buf[174].A ));
 sg13g2_dfrbp_1 _3872_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net214),
    .D(net315),
    .Q_N(_1764_),
    .Q(\i_w_buf[175].A ));
 sg13g2_dfrbp_1 _3873_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net215),
    .D(net369),
    .Q_N(_1765_),
    .Q(\i_w_buf[176].A ));
 sg13g2_dfrbp_1 _3874_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net216),
    .D(net422),
    .Q_N(_1766_),
    .Q(\i_w_buf[177].A ));
 sg13g2_dfrbp_1 _3875_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net217),
    .D(net326),
    .Q_N(_1767_),
    .Q(\i_w_buf[178].A ));
 sg13g2_dfrbp_1 _3876_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net218),
    .D(net353),
    .Q_N(_1768_),
    .Q(\i_w_buf[179].A ));
 sg13g2_dfrbp_1 _3877_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net219),
    .D(net430),
    .Q_N(_1769_),
    .Q(\i_w_buf[180].A ));
 sg13g2_dfrbp_1 _3878_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net220),
    .D(net457),
    .Q_N(_1770_),
    .Q(\i_w_buf[181].A ));
 sg13g2_dfrbp_1 _3879_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net221),
    .D(net431),
    .Q_N(_1771_),
    .Q(\i_w_buf[182].A ));
 sg13g2_dfrbp_1 _3880_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net222),
    .D(net476),
    .Q_N(_1772_),
    .Q(\i_w_buf[183].A ));
 sg13g2_dfrbp_1 _3881_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net223),
    .D(net323),
    .Q_N(_1773_),
    .Q(\i_w_buf[184].A ));
 sg13g2_dfrbp_1 _3882_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net224),
    .D(net307),
    .Q_N(_1774_),
    .Q(\i_w_buf[185].A ));
 sg13g2_dfrbp_1 _3883_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net225),
    .D(net327),
    .Q_N(_1775_),
    .Q(\i_w_buf[186].A ));
 sg13g2_dfrbp_1 _3884_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net226),
    .D(net405),
    .Q_N(_1776_),
    .Q(\i_w_buf[187].A ));
 sg13g2_dfrbp_1 _3885_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net227),
    .D(net531),
    .Q_N(_1777_),
    .Q(\i_w_buf[188].A ));
 sg13g2_dfrbp_1 _3886_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net228),
    .D(net526),
    .Q_N(_1778_),
    .Q(\i_w_buf[189].A ));
 sg13g2_dfrbp_1 _3887_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net229),
    .D(net434),
    .Q_N(_1779_),
    .Q(\i_w_buf[190].A ));
 sg13g2_dfrbp_1 _3888_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net230),
    .D(net425),
    .Q_N(_1780_),
    .Q(\i_w_buf[191].A ));
 sg13g2_dfrbp_1 _3889_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net231),
    .D(net389),
    .Q_N(_1781_),
    .Q(\i_w_buf[192].A ));
 sg13g2_dfrbp_1 _3890_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net232),
    .D(net365),
    .Q_N(_1782_),
    .Q(\i_w_buf[193].A ));
 sg13g2_dfrbp_1 _3891_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net233),
    .D(net475),
    .Q_N(_1783_),
    .Q(\i_w_buf[194].A ));
 sg13g2_dfrbp_1 _3892_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net234),
    .D(net472),
    .Q_N(_1784_),
    .Q(\i_w_buf[195].A ));
 sg13g2_dfrbp_1 _3893_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net235),
    .D(net310),
    .Q_N(_1785_),
    .Q(\i_w_buf[196].A ));
 sg13g2_dfrbp_1 _3894_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net236),
    .D(net396),
    .Q_N(_1786_),
    .Q(\i_w_buf[197].A ));
 sg13g2_dfrbp_1 _3895_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net237),
    .D(net467),
    .Q_N(_1787_),
    .Q(\i_w_buf[198].A ));
 sg13g2_dfrbp_1 _3896_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net238),
    .D(net494),
    .Q_N(_1788_),
    .Q(\i_w_buf[199].A ));
 sg13g2_dfrbp_1 _3897_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net239),
    .D(net390),
    .Q_N(_1789_),
    .Q(\i_w_buf[200].A ));
 sg13g2_dfrbp_1 _3898_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net240),
    .D(net366),
    .Q_N(_1790_),
    .Q(\i_w_buf[201].A ));
 sg13g2_dfrbp_1 _3899_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net241),
    .D(net336),
    .Q_N(_1791_),
    .Q(\i_w_buf[202].A ));
 sg13g2_dfrbp_1 _3900_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net242),
    .D(net356),
    .Q_N(_1792_),
    .Q(\i_w_buf[203].A ));
 sg13g2_dfrbp_1 _3901_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net243),
    .D(net383),
    .Q_N(_1793_),
    .Q(\i_w_buf[204].A ));
 sg13g2_dfrbp_1 _3902_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net244),
    .D(net407),
    .Q_N(_1794_),
    .Q(\i_w_buf[205].A ));
 sg13g2_dfrbp_1 _3903_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net245),
    .D(net403),
    .Q_N(_1795_),
    .Q(\i_w_buf[206].A ));
 sg13g2_dfrbp_1 _3904_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net246),
    .D(net379),
    .Q_N(_1796_),
    .Q(\i_w_buf[207].A ));
 sg13g2_dfrbp_1 _3905_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net247),
    .D(net443),
    .Q_N(_1797_),
    .Q(\i_w_buf[208].A ));
 sg13g2_dfrbp_1 _3906_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net248),
    .D(net394),
    .Q_N(_1798_),
    .Q(\i_w_buf[209].A ));
 sg13g2_dfrbp_1 _3907_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net249),
    .D(net375),
    .Q_N(_1799_),
    .Q(\i_w_buf[210].A ));
 sg13g2_dfrbp_1 _3908_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net250),
    .D(net388),
    .Q_N(_1800_),
    .Q(\i_w_buf[211].A ));
 sg13g2_dfrbp_1 _3909_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net251),
    .D(net318),
    .Q_N(_1801_),
    .Q(\i_w_buf[212].A ));
 sg13g2_dfrbp_1 _3910_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net252),
    .D(net342),
    .Q_N(_1802_),
    .Q(\i_w_buf[213].A ));
 sg13g2_dfrbp_1 _3911_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net253),
    .D(net426),
    .Q_N(_1803_),
    .Q(\i_w_buf[214].A ));
 sg13g2_dfrbp_1 _3912_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net254),
    .D(net418),
    .Q_N(_1804_),
    .Q(\i_w_buf[215].A ));
 sg13g2_dfrbp_1 _3913_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net255),
    .D(net501),
    .Q_N(_1805_),
    .Q(\i_w_buf[216].A ));
 sg13g2_dfrbp_1 _3914_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net256),
    .D(net489),
    .Q_N(_1806_),
    .Q(\i_w_buf[217].A ));
 sg13g2_dfrbp_1 _3915_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net257),
    .D(net414),
    .Q_N(_1807_),
    .Q(\i_w_buf[218].A ));
 sg13g2_dfrbp_1 _3916_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net258),
    .D(net415),
    .Q_N(_1808_),
    .Q(\i_w_buf[219].A ));
 sg13g2_dfrbp_1 _3917_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net259),
    .D(net519),
    .Q_N(_1809_),
    .Q(\i_w_buf[220].A ));
 sg13g2_dfrbp_1 _3918_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net260),
    .D(net540),
    .Q_N(_1810_),
    .Q(\i_w_buf[221].A ));
 sg13g2_dfrbp_1 _3919_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net261),
    .D(net456),
    .Q_N(_1811_),
    .Q(\i_w_buf[222].A ));
 sg13g2_dfrbp_1 _3920_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net262),
    .D(net382),
    .Q_N(_1812_),
    .Q(\i_w_buf[223].A ));
 sg13g2_dfrbp_1 _3921_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net263),
    .D(net436),
    .Q_N(_1813_),
    .Q(\i_w_buf[224].A ));
 sg13g2_dfrbp_1 _3922_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net264),
    .D(net465),
    .Q_N(_1814_),
    .Q(\i_w_buf[225].A ));
 sg13g2_dfrbp_1 _3923_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net265),
    .D(net300),
    .Q_N(_1815_),
    .Q(\i_w_buf[226].A ));
 sg13g2_dfrbp_1 _3924_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net266),
    .D(net321),
    .Q_N(_1816_),
    .Q(\i_w_buf[227].A ));
 sg13g2_dfrbp_1 _3925_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net267),
    .D(net398),
    .Q_N(_1817_),
    .Q(\i_w_buf[228].A ));
 sg13g2_dfrbp_1 _3926_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net268),
    .D(net411),
    .Q_N(_1818_),
    .Q(\i_w_buf[229].A ));
 sg13g2_dfrbp_1 _3927_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net269),
    .D(net371),
    .Q_N(_1819_),
    .Q(\i_w_buf[230].A ));
 sg13g2_dfrbp_1 _3928_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net270),
    .D(net330),
    .Q_N(_1820_),
    .Q(\i_w_buf[231].A ));
 sg13g2_dfrbp_1 _3929_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net271),
    .D(net322),
    .Q_N(_1821_),
    .Q(\i_w_buf[232].A ));
 sg13g2_dfrbp_1 _3930_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net272),
    .D(net339),
    .Q_N(_1822_),
    .Q(\i_w_buf[233].A ));
 sg13g2_dfrbp_1 _3931_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net273),
    .D(net304),
    .Q_N(_1823_),
    .Q(\i_w_buf[234].A ));
 sg13g2_dfrbp_1 _3932_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net274),
    .D(net346),
    .Q_N(_1824_),
    .Q(\i_w_buf[235].A ));
 sg13g2_dfrbp_1 _3933_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net275),
    .D(net515),
    .Q_N(_1825_),
    .Q(\i_w_buf[236].A ));
 sg13g2_dfrbp_1 _3934_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net276),
    .D(net510),
    .Q_N(_1826_),
    .Q(\i_w_buf[237].A ));
 sg13g2_dfrbp_1 _3935_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net277),
    .D(net349),
    .Q_N(_1827_),
    .Q(\i_w_buf[238].A ));
 sg13g2_dfrbp_1 _3936_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net278),
    .D(net360),
    .Q_N(_1828_),
    .Q(\i_w_buf[239].A ));
 sg13g2_dfrbp_1 _3937_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net279),
    .D(net419),
    .Q_N(_1829_),
    .Q(\i_w_buf[240].A ));
 sg13g2_dfrbp_1 _3938_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net280),
    .D(net496),
    .Q_N(_1830_),
    .Q(\i_w_buf[241].A ));
 sg13g2_dfrbp_1 _3939_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net281),
    .D(net536),
    .Q_N(_1831_),
    .Q(\i_w_buf[242].A ));
 sg13g2_dfrbp_1 _3940_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net282),
    .D(net527),
    .Q_N(_1832_),
    .Q(\i_w_buf[243].A ));
 sg13g2_dfrbp_1 _3941_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net283),
    .D(net314),
    .Q_N(_1833_),
    .Q(\i_w_buf[244].A ));
 sg13g2_dfrbp_1 _3942_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net284),
    .D(net341),
    .Q_N(_1834_),
    .Q(\i_w_buf[245].A ));
 sg13g2_dfrbp_1 _3943_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net285),
    .D(net358),
    .Q_N(_1835_),
    .Q(\i_w_buf[246].A ));
 sg13g2_dfrbp_1 _3944_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net286),
    .D(net464),
    .Q_N(_1836_),
    .Q(\i_w_buf[247].A ));
 sg13g2_dfrbp_1 _3945_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net287),
    .D(net423),
    .Q_N(_1837_),
    .Q(\i_w_buf[248].A ));
 sg13g2_dfrbp_1 _3946_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net288),
    .D(net459),
    .Q_N(_1838_),
    .Q(\i_w_buf[249].A ));
 sg13g2_dfrbp_1 _3947_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net289),
    .D(net408),
    .Q_N(_1839_),
    .Q(\i_w_buf[250].A ));
 sg13g2_dfrbp_1 _3948_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net290),
    .D(net350),
    .Q_N(_1840_),
    .Q(\i_w_buf[251].A ));
 sg13g2_dfrbp_1 _3949_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net291),
    .D(net399),
    .Q_N(_1841_),
    .Q(\i_w_buf[252].A ));
 sg13g2_dfrbp_1 _3950_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net292),
    .D(net517),
    .Q_N(_1842_),
    .Q(\i_w_buf[253].A ));
 sg13g2_dfrbp_1 _3951_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net9),
    .D(net428),
    .Q_N(_1843_),
    .Q(\i_w_buf[254].A ));
 sg13g2_dfrbp_1 _3952_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net10),
    .D(net454),
    .Q_N(_1588_),
    .Q(\i_w_buf[255].A ));
 sg13g2_tiehi _3952__10 (.L_HI(net10));
 sg13g2_tiehi _3697__11 (.L_HI(net11));
 sg13g2_tiehi _3698__12 (.L_HI(net12));
 sg13g2_tiehi _3699__13 (.L_HI(net13));
 sg13g2_tiehi _3700__14 (.L_HI(net14));
 sg13g2_tiehi _3701__15 (.L_HI(net15));
 sg13g2_tiehi _3702__16 (.L_HI(net16));
 sg13g2_tiehi _3703__17 (.L_HI(net17));
 sg13g2_tiehi _3704__18 (.L_HI(net18));
 sg13g2_tiehi _3705__19 (.L_HI(net19));
 sg13g2_tiehi _3706__20 (.L_HI(net20));
 sg13g2_tiehi _3707__21 (.L_HI(net21));
 sg13g2_tiehi _3708__22 (.L_HI(net22));
 sg13g2_tiehi _3709__23 (.L_HI(net23));
 sg13g2_tiehi _3710__24 (.L_HI(net24));
 sg13g2_tiehi _3711__25 (.L_HI(net25));
 sg13g2_tiehi _3712__26 (.L_HI(net26));
 sg13g2_tiehi _3713__27 (.L_HI(net27));
 sg13g2_tiehi _3714__28 (.L_HI(net28));
 sg13g2_tiehi _3715__29 (.L_HI(net29));
 sg13g2_tiehi _3716__30 (.L_HI(net30));
 sg13g2_tiehi _3717__31 (.L_HI(net31));
 sg13g2_tiehi _3718__32 (.L_HI(net32));
 sg13g2_tiehi _3719__33 (.L_HI(net33));
 sg13g2_tiehi _3720__34 (.L_HI(net34));
 sg13g2_tiehi _3721__35 (.L_HI(net35));
 sg13g2_tiehi _3722__36 (.L_HI(net36));
 sg13g2_tiehi _3723__37 (.L_HI(net37));
 sg13g2_tiehi _3724__38 (.L_HI(net38));
 sg13g2_tiehi _3725__39 (.L_HI(net39));
 sg13g2_tiehi _3726__40 (.L_HI(net40));
 sg13g2_tiehi _3727__41 (.L_HI(net41));
 sg13g2_tiehi _3728__42 (.L_HI(net42));
 sg13g2_tiehi _3729__43 (.L_HI(net43));
 sg13g2_tiehi _3730__44 (.L_HI(net44));
 sg13g2_tiehi _3731__45 (.L_HI(net45));
 sg13g2_tiehi _3732__46 (.L_HI(net46));
 sg13g2_tiehi _3733__47 (.L_HI(net47));
 sg13g2_tiehi _3734__48 (.L_HI(net48));
 sg13g2_tiehi _3735__49 (.L_HI(net49));
 sg13g2_tiehi _3736__50 (.L_HI(net50));
 sg13g2_tiehi _3737__51 (.L_HI(net51));
 sg13g2_tiehi _3738__52 (.L_HI(net52));
 sg13g2_tiehi _3739__53 (.L_HI(net53));
 sg13g2_tiehi _3740__54 (.L_HI(net54));
 sg13g2_tiehi _3741__55 (.L_HI(net55));
 sg13g2_tiehi _3742__56 (.L_HI(net56));
 sg13g2_tiehi _3743__57 (.L_HI(net57));
 sg13g2_tiehi _3744__58 (.L_HI(net58));
 sg13g2_tiehi _3745__59 (.L_HI(net59));
 sg13g2_tiehi _3746__60 (.L_HI(net60));
 sg13g2_tiehi _3747__61 (.L_HI(net61));
 sg13g2_tiehi _3748__62 (.L_HI(net62));
 sg13g2_tiehi _3749__63 (.L_HI(net63));
 sg13g2_tiehi _3750__64 (.L_HI(net64));
 sg13g2_tiehi _3751__65 (.L_HI(net65));
 sg13g2_tiehi _3752__66 (.L_HI(net66));
 sg13g2_tiehi _3753__67 (.L_HI(net67));
 sg13g2_tiehi _3754__68 (.L_HI(net68));
 sg13g2_tiehi _3755__69 (.L_HI(net69));
 sg13g2_tiehi _3756__70 (.L_HI(net70));
 sg13g2_tiehi _3757__71 (.L_HI(net71));
 sg13g2_tiehi _3758__72 (.L_HI(net72));
 sg13g2_tiehi _3759__73 (.L_HI(net73));
 sg13g2_tiehi _3760__74 (.L_HI(net74));
 sg13g2_tiehi _3761__75 (.L_HI(net75));
 sg13g2_tiehi _3762__76 (.L_HI(net76));
 sg13g2_tiehi _3763__77 (.L_HI(net77));
 sg13g2_tiehi _3764__78 (.L_HI(net78));
 sg13g2_tiehi _3765__79 (.L_HI(net79));
 sg13g2_tiehi _3766__80 (.L_HI(net108));
 sg13g2_tiehi _3767__81 (.L_HI(net109));
 sg13g2_tiehi _3768__82 (.L_HI(net110));
 sg13g2_tiehi _3769__83 (.L_HI(net111));
 sg13g2_tiehi _3770__84 (.L_HI(net112));
 sg13g2_tiehi _3771__85 (.L_HI(net113));
 sg13g2_tiehi _3772__86 (.L_HI(net114));
 sg13g2_tiehi _3773__87 (.L_HI(net115));
 sg13g2_tiehi _3774__88 (.L_HI(net116));
 sg13g2_tiehi _3775__89 (.L_HI(net117));
 sg13g2_tiehi _3776__90 (.L_HI(net118));
 sg13g2_tiehi _3777__91 (.L_HI(net119));
 sg13g2_tiehi _3778__92 (.L_HI(net120));
 sg13g2_tiehi _3779__93 (.L_HI(net121));
 sg13g2_tiehi _3780__94 (.L_HI(net122));
 sg13g2_tiehi _3781__95 (.L_HI(net123));
 sg13g2_tiehi _3782__96 (.L_HI(net124));
 sg13g2_tiehi _3783__97 (.L_HI(net125));
 sg13g2_tiehi _3784__98 (.L_HI(net126));
 sg13g2_tiehi _3785__99 (.L_HI(net127));
 sg13g2_tiehi _3786__100 (.L_HI(net128));
 sg13g2_tiehi _3787__101 (.L_HI(net129));
 sg13g2_tiehi _3788__102 (.L_HI(net130));
 sg13g2_tiehi _3789__103 (.L_HI(net131));
 sg13g2_tiehi _3790__104 (.L_HI(net132));
 sg13g2_tiehi _3791__105 (.L_HI(net133));
 sg13g2_tiehi _3792__106 (.L_HI(net134));
 sg13g2_tiehi _3793__107 (.L_HI(net135));
 sg13g2_tiehi _3794__108 (.L_HI(net136));
 sg13g2_tiehi _3795__109 (.L_HI(net137));
 sg13g2_tiehi _3796__110 (.L_HI(net138));
 sg13g2_tiehi _3797__111 (.L_HI(net139));
 sg13g2_tiehi _3798__112 (.L_HI(net140));
 sg13g2_tiehi _3799__113 (.L_HI(net141));
 sg13g2_tiehi _3800__114 (.L_HI(net142));
 sg13g2_tiehi _3801__115 (.L_HI(net143));
 sg13g2_tiehi _3802__116 (.L_HI(net144));
 sg13g2_tiehi _3803__117 (.L_HI(net145));
 sg13g2_tiehi _3804__118 (.L_HI(net146));
 sg13g2_tiehi _3805__119 (.L_HI(net147));
 sg13g2_tiehi _3806__120 (.L_HI(net148));
 sg13g2_tiehi _3807__121 (.L_HI(net149));
 sg13g2_tiehi _3808__122 (.L_HI(net150));
 sg13g2_tiehi _3809__123 (.L_HI(net151));
 sg13g2_tiehi _3810__124 (.L_HI(net152));
 sg13g2_tiehi _3811__125 (.L_HI(net153));
 sg13g2_tiehi _3812__126 (.L_HI(net154));
 sg13g2_tiehi _3813__127 (.L_HI(net155));
 sg13g2_tiehi _3814__128 (.L_HI(net156));
 sg13g2_tiehi _3815__129 (.L_HI(net157));
 sg13g2_tiehi _3816__130 (.L_HI(net158));
 sg13g2_tiehi _3817__131 (.L_HI(net159));
 sg13g2_tiehi _3818__132 (.L_HI(net160));
 sg13g2_tiehi _3819__133 (.L_HI(net161));
 sg13g2_tiehi _3820__134 (.L_HI(net162));
 sg13g2_tiehi _3821__135 (.L_HI(net163));
 sg13g2_tiehi _3822__136 (.L_HI(net164));
 sg13g2_tiehi _3823__137 (.L_HI(net165));
 sg13g2_tiehi _3824__138 (.L_HI(net166));
 sg13g2_tiehi _3825__139 (.L_HI(net167));
 sg13g2_tiehi _3826__140 (.L_HI(net168));
 sg13g2_tiehi _3827__141 (.L_HI(net169));
 sg13g2_tiehi _3828__142 (.L_HI(net170));
 sg13g2_tiehi _3829__143 (.L_HI(net171));
 sg13g2_tiehi _3830__144 (.L_HI(net172));
 sg13g2_tiehi _3831__145 (.L_HI(net173));
 sg13g2_tiehi _3832__146 (.L_HI(net174));
 sg13g2_tiehi _3833__147 (.L_HI(net175));
 sg13g2_tiehi _3834__148 (.L_HI(net176));
 sg13g2_tiehi _3835__149 (.L_HI(net177));
 sg13g2_tiehi _3836__150 (.L_HI(net178));
 sg13g2_tiehi _3837__151 (.L_HI(net179));
 sg13g2_tiehi _3838__152 (.L_HI(net180));
 sg13g2_tiehi _3839__153 (.L_HI(net181));
 sg13g2_tiehi _3840__154 (.L_HI(net182));
 sg13g2_tiehi _3841__155 (.L_HI(net183));
 sg13g2_tiehi _3842__156 (.L_HI(net184));
 sg13g2_tiehi _3843__157 (.L_HI(net185));
 sg13g2_tiehi _3844__158 (.L_HI(net186));
 sg13g2_tiehi _3845__159 (.L_HI(net187));
 sg13g2_tiehi _3846__160 (.L_HI(net188));
 sg13g2_tiehi _3847__161 (.L_HI(net189));
 sg13g2_tiehi _3848__162 (.L_HI(net190));
 sg13g2_tiehi _3849__163 (.L_HI(net191));
 sg13g2_tiehi _3850__164 (.L_HI(net192));
 sg13g2_tiehi _3851__165 (.L_HI(net193));
 sg13g2_tiehi _3852__166 (.L_HI(net194));
 sg13g2_tiehi _3853__167 (.L_HI(net195));
 sg13g2_tiehi _3854__168 (.L_HI(net196));
 sg13g2_tiehi _3855__169 (.L_HI(net197));
 sg13g2_tiehi _3856__170 (.L_HI(net198));
 sg13g2_tiehi _3857__171 (.L_HI(net199));
 sg13g2_tiehi _3858__172 (.L_HI(net200));
 sg13g2_tiehi _3859__173 (.L_HI(net201));
 sg13g2_tiehi _3860__174 (.L_HI(net202));
 sg13g2_tiehi _3861__175 (.L_HI(net203));
 sg13g2_tiehi _3862__176 (.L_HI(net204));
 sg13g2_tiehi _3863__177 (.L_HI(net205));
 sg13g2_tiehi _3864__178 (.L_HI(net206));
 sg13g2_tiehi _3865__179 (.L_HI(net207));
 sg13g2_tiehi _3866__180 (.L_HI(net208));
 sg13g2_tiehi _3867__181 (.L_HI(net209));
 sg13g2_tiehi _3868__182 (.L_HI(net210));
 sg13g2_tiehi _3869__183 (.L_HI(net211));
 sg13g2_tiehi _3870__184 (.L_HI(net212));
 sg13g2_tiehi _3871__185 (.L_HI(net213));
 sg13g2_tiehi _3872__186 (.L_HI(net214));
 sg13g2_tiehi _3873__187 (.L_HI(net215));
 sg13g2_tiehi _3874__188 (.L_HI(net216));
 sg13g2_tiehi _3875__189 (.L_HI(net217));
 sg13g2_tiehi _3876__190 (.L_HI(net218));
 sg13g2_tiehi _3877__191 (.L_HI(net219));
 sg13g2_tiehi _3878__192 (.L_HI(net220));
 sg13g2_tiehi _3879__193 (.L_HI(net221));
 sg13g2_tiehi _3880__194 (.L_HI(net222));
 sg13g2_tiehi _3881__195 (.L_HI(net223));
 sg13g2_tiehi _3882__196 (.L_HI(net224));
 sg13g2_tiehi _3883__197 (.L_HI(net225));
 sg13g2_tiehi _3884__198 (.L_HI(net226));
 sg13g2_tiehi _3885__199 (.L_HI(net227));
 sg13g2_tiehi _3886__200 (.L_HI(net228));
 sg13g2_tiehi _3887__201 (.L_HI(net229));
 sg13g2_tiehi _3888__202 (.L_HI(net230));
 sg13g2_tiehi _3889__203 (.L_HI(net231));
 sg13g2_tiehi _3890__204 (.L_HI(net232));
 sg13g2_tiehi _3891__205 (.L_HI(net233));
 sg13g2_tiehi _3892__206 (.L_HI(net234));
 sg13g2_tiehi _3893__207 (.L_HI(net235));
 sg13g2_tiehi _3894__208 (.L_HI(net236));
 sg13g2_tiehi _3895__209 (.L_HI(net237));
 sg13g2_tiehi _3896__210 (.L_HI(net238));
 sg13g2_tiehi _3897__211 (.L_HI(net239));
 sg13g2_tiehi _3898__212 (.L_HI(net240));
 sg13g2_tiehi _3899__213 (.L_HI(net241));
 sg13g2_tiehi _3900__214 (.L_HI(net242));
 sg13g2_tiehi _3901__215 (.L_HI(net243));
 sg13g2_tiehi _3902__216 (.L_HI(net244));
 sg13g2_tiehi _3903__217 (.L_HI(net245));
 sg13g2_tiehi _3904__218 (.L_HI(net246));
 sg13g2_tiehi _3905__219 (.L_HI(net247));
 sg13g2_tiehi _3906__220 (.L_HI(net248));
 sg13g2_tiehi _3907__221 (.L_HI(net249));
 sg13g2_tiehi _3908__222 (.L_HI(net250));
 sg13g2_tiehi _3909__223 (.L_HI(net251));
 sg13g2_tiehi _3910__224 (.L_HI(net252));
 sg13g2_tiehi _3911__225 (.L_HI(net253));
 sg13g2_tiehi _3912__226 (.L_HI(net254));
 sg13g2_tiehi _3913__227 (.L_HI(net255));
 sg13g2_tiehi _3914__228 (.L_HI(net256));
 sg13g2_tiehi _3915__229 (.L_HI(net257));
 sg13g2_tiehi _3916__230 (.L_HI(net258));
 sg13g2_tiehi _3917__231 (.L_HI(net259));
 sg13g2_tiehi _3918__232 (.L_HI(net260));
 sg13g2_tiehi _3919__233 (.L_HI(net261));
 sg13g2_tiehi _3920__234 (.L_HI(net262));
 sg13g2_tiehi _3921__235 (.L_HI(net263));
 sg13g2_tiehi _3922__236 (.L_HI(net264));
 sg13g2_tiehi _3923__237 (.L_HI(net265));
 sg13g2_tiehi _3924__238 (.L_HI(net266));
 sg13g2_tiehi _3925__239 (.L_HI(net267));
 sg13g2_tiehi _3926__240 (.L_HI(net268));
 sg13g2_tiehi _3927__241 (.L_HI(net269));
 sg13g2_tiehi _3928__242 (.L_HI(net270));
 sg13g2_tiehi _3929__243 (.L_HI(net271));
 sg13g2_tiehi _3930__244 (.L_HI(net272));
 sg13g2_tiehi _3931__245 (.L_HI(net273));
 sg13g2_tiehi _3932__246 (.L_HI(net274));
 sg13g2_tiehi _3933__247 (.L_HI(net275));
 sg13g2_tiehi _3934__248 (.L_HI(net276));
 sg13g2_tiehi _3935__249 (.L_HI(net277));
 sg13g2_tiehi _3936__250 (.L_HI(net278));
 sg13g2_tiehi _3937__251 (.L_HI(net279));
 sg13g2_tiehi _3938__252 (.L_HI(net280));
 sg13g2_tiehi _3939__253 (.L_HI(net281));
 sg13g2_tiehi _3940__254 (.L_HI(net282));
 sg13g2_tiehi _3941__255 (.L_HI(net283));
 sg13g2_tiehi _3942__256 (.L_HI(net284));
 sg13g2_tiehi _3943__257 (.L_HI(net285));
 sg13g2_tiehi _3944__258 (.L_HI(net286));
 sg13g2_tiehi _3945__259 (.L_HI(net287));
 sg13g2_tiehi _3946__260 (.L_HI(net288));
 sg13g2_tiehi _3947__261 (.L_HI(net289));
 sg13g2_tiehi _3948__262 (.L_HI(net290));
 sg13g2_tiehi _3949__263 (.L_HI(net291));
 sg13g2_tiehi _3950__264 (.L_HI(net292));
 sg13g2_tiehi tt_um_rejunity_ternary_dot_265 (.L_HI(net293));
 sg13g2_tiehi tt_um_rejunity_ternary_dot_266 (.L_HI(net294));
 sg13g2_tiehi tt_um_rejunity_ternary_dot_267 (.L_HI(net295));
 sg13g2_tiehi tt_um_rejunity_ternary_dot_268 (.L_HI(net296));
 sg13g2_tiehi tt_um_rejunity_ternary_dot_269 (.L_HI(net297));
 sg13g2_tiehi tt_um_rejunity_ternary_dot_270 (.L_HI(net298));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_rejunity_ternary_dot_7 (.L_LO(net7));
 sg13g2_tielo tt_um_rejunity_ternary_dot_8 (.L_LO(net8));
 sg13g2_tiehi _3951__9 (.L_HI(net9));
 sg13g2_buf_1 _4218_ (.A(uio_out[7]),
    .X(uio_out[1]));
 sg13g2_buf_1 _4219_ (.A(uio_out[7]),
    .X(uio_out[2]));
 sg13g2_buf_1 _4220_ (.A(uio_out[7]),
    .X(uio_out[3]));
 sg13g2_buf_1 _4221_ (.A(uio_out[7]),
    .X(uio_out[4]));
 sg13g2_buf_1 _4222_ (.A(uio_out[7]),
    .X(uio_out[5]));
 sg13g2_buf_1 _4223_ (.A(uio_out[7]),
    .X(uio_out[6]));
 sg13g2_buf_8 fanout80 (.A(_0870_),
    .X(net80));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(net82));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_0869_));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_0867_));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(_0867_));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_0866_));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(_0866_));
 sg13g2_buf_8 fanout87 (.A(_0865_),
    .X(net87));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(_0862_));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(ui_in[7]));
 sg13g2_buf_2 fanout90 (.A(ui_in[7]),
    .X(net90));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(net92));
 sg13g2_buf_8 fanout92 (.A(net3),
    .X(net92));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(net95));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(ui_in[5]));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(net97));
 sg13g2_buf_8 fanout97 (.A(net2),
    .X(net97));
 sg13g2_buf_8 fanout98 (.A(ui_in[3]),
    .X(net98));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(ui_in[3]));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(net102));
 sg13g2_buf_8 fanout101 (.A(ui_in[2]),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(ui_in[2]),
    .X(net102));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net105));
 sg13g2_buf_2 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_8 fanout105 (.A(ui_in[1]),
    .X(net105));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(net107));
 sg13g2_buf_8 fanout107 (.A(net1),
    .X(net107));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ui_in[0]));
 sg13g2_buf_2 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[0]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[1]),
    .X(net5));
 sg13g2_tielo tt_um_rejunity_ternary_dot_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_leaf_36_clk));
 sg13g2_inv_8 clkload3 (.A(clknet_leaf_37_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_32_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_31_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_23_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_26_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_5_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_13_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_21_clk));
 sg13g2_inv_8 clkload13 (.A(clknet_leaf_22_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_19_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\i_w_buf[69].A ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold2 (.A(\i_w_buf[224].A ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold3 (.A(\i_w_buf[92].A ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold4 (.A(\i_w_buf[10].A ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i_w_buf[136].A ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_w_buf[232].A ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_w_buf[96].A ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_w_buf[132].A ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_w_buf[183].A ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_w_buf[62].A ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_w_buf[104].A ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_w_buf[194].A ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_w_buf[164].A ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_w_buf[82].A ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_w_buf[20].A ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_w_buf[242].A ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_w_buf[173].A ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_w_buf[14].A ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_w_buf[168].A ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_w_buf[210].A ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_w_buf[8].A ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_w_buf[120].A ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i_w_buf[225].A ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_w_buf[230].A ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_w_buf[182].A ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_w_buf[106].A ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i_w_buf[2].A ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_w_buf[176].A ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i_w_buf[184].A ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_w_buf[172].A ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_w_buf[38].A ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_w_buf[229].A ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold33 (.A(\i_w_buf[78].A ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_w_buf[34].A ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_w_buf[88].A ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_w_buf[15].A ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold37 (.A(\i_w_buf[22].A ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_w_buf[200].A ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_w_buf[66].A ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_w_buf[170].A ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_w_buf[231].A ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_w_buf[113].A ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold43 (.A(\i_w_buf[243].A ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_w_buf[211].A ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold45 (.A(\i_w_buf[160].A ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_w_buf[98].A ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold47 (.A(\i_w_buf[52].A ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_w_buf[233].A ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_w_buf[53].A ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_w_buf[114].A ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold51 (.A(\i_w_buf[236].A ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_w_buf[249].A ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_w_buf[30].A ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_w_buf[128].A ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_w_buf[177].A ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_w_buf[112].A ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold57 (.A(\i_w_buf[95].A ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_w_buf[201].A ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_w_buf[159].A ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_w_buf[244].A ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold61 (.A(\i_w_buf[4].A ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_w_buf[237].A ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_w_buf[144].A ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold64 (.A(\i_w_buf[145].A ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_w_buf[139].A ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_w_buf[56].A ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold67 (.A(\i_w_buf[191].A ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_w_buf[199].A ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold69 (.A(\i_w_buf[146].A ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_w_buf[25].A ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold71 (.A(\i_w_buf[174].A ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_w_buf[142].A ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold73 (.A(\i_w_buf[228].A ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_w_buf[24].A ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_w_buf[158].A ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_w_buf[46].A ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold77 (.A(\i_w_buf[208].A ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_w_buf[63].A ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold79 (.A(\i_w_buf[79].A ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_w_buf[105].A ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_w_buf[205].A ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_w_buf[74].A ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold83 (.A(\i_w_buf[42].A ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_w_buf[221].A ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold85 (.A(\i_w_buf[202].A ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_w_buf[35].A ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_w_buf[16].A ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_w_buf[26].A ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_w_buf[161].A ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold90 (.A(\i_w_buf[209].A ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_w_buf[190].A ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold92 (.A(\i_w_buf[198].A ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_w_buf[118].A ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold94 (.A(\i_w_buf[169].A ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_w_buf[165].A ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_w_buf[207].A ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_w_buf[115].A ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_w_buf[195].A ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_w_buf[117].A ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold100 (.A(\i_w_buf[226].A ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_w_buf[250].A ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold102 (.A(\i_w_buf[116].A ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_w_buf[84].A ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold104 (.A(\i_w_buf[9].A ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold105 (.A(\i_w_buf[204].A ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_w_buf[121].A ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold107 (.A(\i_w_buf[185].A ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_w_buf[154].A ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_w_buf[203].A ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_w_buf[248].A ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_w_buf[43].A ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_w_buf[148].A ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_w_buf[227].A ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_w_buf[171].A ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold115 (.A(\i_w_buf[27].A ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_w_buf[216].A ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold117 (.A(\i_w_buf[217].A ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_w_buf[83].A ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_w_buf[6].A ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_w_buf[213].A ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold121 (.A(\i_w_buf[238].A ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_w_buf[124].A ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_w_buf[129].A ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_w_buf[175].A ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_w_buf[246].A ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_w_buf[133].A ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_w_buf[189].A ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_w_buf[212].A ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_w_buf[85].A ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_w_buf[252].A ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_w_buf[33].A ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_w_buf[178].A ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_w_buf[180].A ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_w_buf[75].A ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_w_buf[153].A ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold136 (.A(\i_w_buf[188].A ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold137 (.A(\i_w_buf[17].A ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_w_buf[222].A ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_w_buf[23].A ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_w_buf[0].A ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_w_buf[137].A ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold142 (.A(\i_w_buf[107].A ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_w_buf[49].A ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_w_buf[50].A ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_w_buf[206].A ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_w_buf[60].A ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_w_buf[45].A ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_w_buf[5].A ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_w_buf[97].A ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold150 (.A(\i_w_buf[3].A ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_w_buf[54].A ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold152 (.A(\i_w_buf[99].A ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_w_buf[156].A ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_w_buf[81].A ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_w_buf[108].A ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_w_buf[253].A ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_w_buf[47].A ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_w_buf[220].A ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_w_buf[179].A ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_w_buf[57].A ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_w_buf[247].A ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_w_buf[61].A ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_w_buf[39].A ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_w_buf[31].A ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_w_buf[11].A ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_w_buf[245].A ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_w_buf[223].A ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_w_buf[157].A ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_w_buf[196].A ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_w_buf[140].A ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_w_buf[131].A ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold172 (.A(\i_w_buf[93].A ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_w_buf[32].A ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_w_buf[193].A ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_w_buf[1].A ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_w_buf[70].A ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_w_buf[192].A ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_w_buf[181].A ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_w_buf[149].A ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold180 (.A(\i_w_buf[130].A ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_w_buf[44].A ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_w_buf[147].A ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_w_buf[59].A ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold184 (.A(\i_w_buf[80].A ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_w_buf[89].A ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_w_buf[91].A ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_w_buf[71].A ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_w_buf[150].A ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold189 (.A(\i_w_buf[102].A ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold190 (.A(\i_w_buf[141].A ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_w_buf[215].A ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_w_buf[138].A ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold193 (.A(\i_w_buf[55].A ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_w_buf[58].A ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_w_buf[94].A ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold196 (.A(\i_w_buf[197].A ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold197 (.A(\i_w_buf[166].A ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold198 (.A(\i_w_buf[239].A ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_w_buf[68].A ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_w_buf[103].A ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold201 (.A(\i_w_buf[86].A ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold202 (.A(\i_w_buf[28].A ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold203 (.A(\i_w_buf[214].A ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_w_buf[110].A ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold205 (.A(\i_w_buf[21].A ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_w_buf[119].A ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_w_buf[73].A ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold208 (.A(\i_w_buf[155].A ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold209 (.A(\i_w_buf[125].A ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold210 (.A(\i_w_buf[122].A ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_w_buf[7].A ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold212 (.A(\i_w_buf[235].A ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_w_buf[90].A ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold214 (.A(\i_w_buf[19].A ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_w_buf[123].A ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold216 (.A(\i_w_buf[36].A ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_w_buf[234].A ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold218 (.A(\i_w_buf[72].A ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_w_buf[251].A ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_w_buf[152].A ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold221 (.A(\i_w_buf[218].A ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_w_buf[134].A ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_w_buf[143].A ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold224 (.A(\i_w_buf[87].A ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold225 (.A(\i_w_buf[151].A ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold226 (.A(\i_w_buf[167].A ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold227 (.A(\i_w_buf[29].A ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_w_buf[187].A ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold229 (.A(\i_w_buf[241].A ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_w_buf[126].A ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold231 (.A(\i_w_buf[135].A ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_w_buf[111].A ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold233 (.A(\i_w_buf[186].A ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_w_buf[77].A ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_w_buf[51].A ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold236 (.A(\i_w_buf[37].A ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_w_buf[127].A ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_w_buf[240].A ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold239 (.A(\i_w_buf[162].A ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold240 (.A(\i_w_buf[48].A ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold241 (.A(\i_w_buf[12].A ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold242 (.A(\i_w_buf[219].A ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold243 (.A(\i_w_buf[40].A ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_w_buf[76].A ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold245 (.A(\i_w_buf[163].A ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_w_buf[41].A ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold247 (.A(\i_w_buf[18].A ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_w_buf[65].A ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold249 (.A(\i_w_buf[109].A ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_w_buf[64].A ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold251 (.A(\i_w_buf[101].A ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_w_buf[100].A ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold253 (.A(\i_w_buf[13].A ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_w_buf[67].A ),
    .X(net552));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_4 FILLER_0_147 ();
 sg13g2_fill_2 FILLER_0_151 ();
 sg13g2_decap_8 FILLER_0_162 ();
 sg13g2_fill_1 FILLER_0_169 ();
 sg13g2_fill_1 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_fill_2 FILLER_0_245 ();
 sg13g2_fill_1 FILLER_0_247 ();
 sg13g2_decap_4 FILLER_0_261 ();
 sg13g2_fill_1 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_288 ();
 sg13g2_decap_4 FILLER_0_295 ();
 sg13g2_fill_2 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_4 FILLER_0_321 ();
 sg13g2_fill_2 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_fill_2 FILLER_1_182 ();
 sg13g2_fill_2 FILLER_1_218 ();
 sg13g2_fill_1 FILLER_1_220 ();
 sg13g2_fill_2 FILLER_1_312 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_fill_2 FILLER_2_194 ();
 sg13g2_fill_1 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_353 ();
 sg13g2_decap_8 FILLER_2_360 ();
 sg13g2_decap_8 FILLER_2_367 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_4 FILLER_3_133 ();
 sg13g2_fill_2 FILLER_3_172 ();
 sg13g2_fill_1 FILLER_3_174 ();
 sg13g2_fill_2 FILLER_3_201 ();
 sg13g2_fill_2 FILLER_3_242 ();
 sg13g2_fill_1 FILLER_3_244 ();
 sg13g2_fill_1 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_4 FILLER_4_126 ();
 sg13g2_fill_1 FILLER_4_130 ();
 sg13g2_fill_2 FILLER_4_183 ();
 sg13g2_fill_1 FILLER_4_185 ();
 sg13g2_fill_1 FILLER_4_190 ();
 sg13g2_fill_1 FILLER_4_226 ();
 sg13g2_fill_2 FILLER_4_236 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_fill_2 FILLER_4_279 ();
 sg13g2_fill_1 FILLER_4_281 ();
 sg13g2_fill_2 FILLER_4_317 ();
 sg13g2_fill_1 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_4 FILLER_5_119 ();
 sg13g2_fill_2 FILLER_5_165 ();
 sg13g2_fill_1 FILLER_5_184 ();
 sg13g2_fill_2 FILLER_5_189 ();
 sg13g2_fill_1 FILLER_5_191 ();
 sg13g2_fill_2 FILLER_5_205 ();
 sg13g2_decap_8 FILLER_5_212 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_decap_8 FILLER_5_251 ();
 sg13g2_decap_4 FILLER_5_258 ();
 sg13g2_fill_2 FILLER_5_262 ();
 sg13g2_decap_4 FILLER_5_272 ();
 sg13g2_fill_1 FILLER_5_276 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_4 FILLER_6_112 ();
 sg13g2_fill_2 FILLER_6_116 ();
 sg13g2_fill_1 FILLER_6_126 ();
 sg13g2_fill_2 FILLER_6_146 ();
 sg13g2_fill_1 FILLER_6_187 ();
 sg13g2_decap_4 FILLER_6_196 ();
 sg13g2_fill_2 FILLER_6_200 ();
 sg13g2_fill_1 FILLER_6_210 ();
 sg13g2_decap_4 FILLER_6_218 ();
 sg13g2_fill_2 FILLER_6_246 ();
 sg13g2_fill_2 FILLER_6_255 ();
 sg13g2_fill_1 FILLER_6_257 ();
 sg13g2_decap_4 FILLER_6_267 ();
 sg13g2_fill_1 FILLER_6_271 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_222 ();
 sg13g2_fill_1 FILLER_7_233 ();
 sg13g2_fill_2 FILLER_7_271 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_fill_2 FILLER_7_301 ();
 sg13g2_fill_1 FILLER_7_307 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_4 FILLER_8_105 ();
 sg13g2_fill_2 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_fill_2 FILLER_8_222 ();
 sg13g2_fill_1 FILLER_8_237 ();
 sg13g2_fill_1 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_362 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_4 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_109 ();
 sg13g2_fill_2 FILLER_9_227 ();
 sg13g2_fill_2 FILLER_9_288 ();
 sg13g2_fill_2 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_fill_2 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_104 ();
 sg13g2_fill_1 FILLER_10_106 ();
 sg13g2_fill_2 FILLER_10_142 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_fill_1 FILLER_10_150 ();
 sg13g2_fill_1 FILLER_10_160 ();
 sg13g2_fill_1 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_195 ();
 sg13g2_fill_2 FILLER_10_209 ();
 sg13g2_fill_1 FILLER_10_211 ();
 sg13g2_decap_4 FILLER_10_217 ();
 sg13g2_fill_2 FILLER_10_235 ();
 sg13g2_fill_1 FILLER_10_268 ();
 sg13g2_fill_2 FILLER_10_295 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_4 FILLER_11_91 ();
 sg13g2_fill_2 FILLER_11_95 ();
 sg13g2_fill_1 FILLER_11_127 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_fill_1 FILLER_11_187 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_fill_1 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_4 FILLER_11_231 ();
 sg13g2_fill_2 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_251 ();
 sg13g2_decap_4 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_262 ();
 sg13g2_fill_2 FILLER_11_268 ();
 sg13g2_fill_2 FILLER_11_287 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_2 FILLER_11_351 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_4 FILLER_12_98 ();
 sg13g2_fill_1 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_4 FILLER_12_171 ();
 sg13g2_fill_1 FILLER_12_175 ();
 sg13g2_fill_2 FILLER_12_185 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_12_192 ();
 sg13g2_decap_4 FILLER_12_199 ();
 sg13g2_fill_2 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_209 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_decap_4 FILLER_12_223 ();
 sg13g2_fill_2 FILLER_12_227 ();
 sg13g2_fill_1 FILLER_12_251 ();
 sg13g2_fill_2 FILLER_12_261 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_fill_1 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_fill_1 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_234 ();
 sg13g2_fill_1 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_84 ();
 sg13g2_fill_1 FILLER_14_155 ();
 sg13g2_decap_4 FILLER_14_184 ();
 sg13g2_fill_2 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_229 ();
 sg13g2_fill_2 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_fill_2 FILLER_15_119 ();
 sg13g2_decap_4 FILLER_15_130 ();
 sg13g2_fill_2 FILLER_15_134 ();
 sg13g2_fill_1 FILLER_15_150 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_171 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_fill_1 FILLER_15_224 ();
 sg13g2_fill_2 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_278 ();
 sg13g2_fill_1 FILLER_15_285 ();
 sg13g2_decap_8 FILLER_15_292 ();
 sg13g2_fill_2 FILLER_15_304 ();
 sg13g2_fill_2 FILLER_15_324 ();
 sg13g2_fill_2 FILLER_15_331 ();
 sg13g2_decap_4 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_84 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_146 ();
 sg13g2_decap_8 FILLER_16_162 ();
 sg13g2_decap_8 FILLER_16_169 ();
 sg13g2_fill_1 FILLER_16_176 ();
 sg13g2_decap_4 FILLER_16_196 ();
 sg13g2_fill_2 FILLER_16_211 ();
 sg13g2_fill_1 FILLER_16_213 ();
 sg13g2_decap_8 FILLER_16_218 ();
 sg13g2_decap_4 FILLER_16_225 ();
 sg13g2_fill_2 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_fill_2 FILLER_16_248 ();
 sg13g2_fill_1 FILLER_16_250 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_4 FILLER_16_346 ();
 sg13g2_fill_2 FILLER_16_350 ();
 sg13g2_fill_1 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_4 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_fill_2 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_fill_1 FILLER_17_137 ();
 sg13g2_decap_8 FILLER_17_150 ();
 sg13g2_fill_2 FILLER_17_157 ();
 sg13g2_fill_1 FILLER_17_159 ();
 sg13g2_decap_8 FILLER_17_167 ();
 sg13g2_decap_8 FILLER_17_199 ();
 sg13g2_decap_4 FILLER_17_206 ();
 sg13g2_fill_2 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_decap_4 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_decap_4 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_323 ();
 sg13g2_fill_1 FILLER_17_325 ();
 sg13g2_fill_1 FILLER_17_335 ();
 sg13g2_fill_2 FILLER_17_345 ();
 sg13g2_fill_2 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_84 ();
 sg13g2_decap_4 FILLER_18_99 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_8 FILLER_18_142 ();
 sg13g2_decap_4 FILLER_18_149 ();
 sg13g2_decap_8 FILLER_18_195 ();
 sg13g2_decap_4 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_227 ();
 sg13g2_fill_1 FILLER_18_234 ();
 sg13g2_fill_2 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_299 ();
 sg13g2_decap_4 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_127 ();
 sg13g2_decap_4 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_237 ();
 sg13g2_fill_2 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_289 ();
 sg13g2_decap_4 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_97 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_159 ();
 sg13g2_fill_1 FILLER_20_161 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_fill_1 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_274 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_317 ();
 sg13g2_fill_1 FILLER_20_335 ();
 sg13g2_fill_1 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_118 ();
 sg13g2_decap_4 FILLER_21_155 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_fill_2 FILLER_21_169 ();
 sg13g2_fill_1 FILLER_21_177 ();
 sg13g2_decap_4 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_230 ();
 sg13g2_decap_8 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_fill_2 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_295 ();
 sg13g2_fill_1 FILLER_21_297 ();
 sg13g2_fill_2 FILLER_21_324 ();
 sg13g2_fill_2 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_21_347 ();
 sg13g2_decap_4 FILLER_21_383 ();
 sg13g2_fill_1 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_4 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_60 ();
 sg13g2_fill_2 FILLER_22_87 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_decap_4 FILLER_22_164 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_fill_2 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_212 ();
 sg13g2_decap_4 FILLER_22_219 ();
 sg13g2_decap_4 FILLER_22_258 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_decap_4 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_75 ();
 sg13g2_decap_8 FILLER_23_82 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_102 ();
 sg13g2_fill_2 FILLER_23_133 ();
 sg13g2_fill_2 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_156 ();
 sg13g2_fill_1 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_decap_4 FILLER_23_186 ();
 sg13g2_fill_1 FILLER_23_190 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_decap_8 FILLER_23_216 ();
 sg13g2_fill_2 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_225 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_decap_4 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_fill_1 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_4 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_decap_8 FILLER_24_219 ();
 sg13g2_decap_4 FILLER_24_226 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_fill_2 FILLER_24_263 ();
 sg13g2_fill_1 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_279 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_114 ();
 sg13g2_decap_8 FILLER_25_124 ();
 sg13g2_decap_8 FILLER_25_131 ();
 sg13g2_decap_8 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_250 ();
 sg13g2_decap_8 FILLER_25_257 ();
 sg13g2_decap_4 FILLER_25_264 ();
 sg13g2_decap_4 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_fill_2 FILLER_25_321 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_fill_2 FILLER_25_390 ();
 sg13g2_fill_1 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_decap_8 FILLER_26_146 ();
 sg13g2_decap_4 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_171 ();
 sg13g2_decap_4 FILLER_26_178 ();
 sg13g2_fill_1 FILLER_26_182 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_decap_8 FILLER_26_230 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_4 FILLER_26_266 ();
 sg13g2_fill_2 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_fill_2 FILLER_26_281 ();
 sg13g2_fill_1 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_310 ();
 sg13g2_decap_4 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_4 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_decap_8 FILLER_27_148 ();
 sg13g2_decap_8 FILLER_27_155 ();
 sg13g2_decap_8 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_172 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_196 ();
 sg13g2_fill_2 FILLER_27_212 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_84 ();
 sg13g2_decap_4 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_4 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_decap_4 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_318 ();
 sg13g2_fill_2 FILLER_28_331 ();
 sg13g2_fill_1 FILLER_28_333 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_fill_1 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_4 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_100 ();
 sg13g2_fill_1 FILLER_29_102 ();
 sg13g2_fill_2 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_148 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_281 ();
 sg13g2_fill_2 FILLER_29_288 ();
 sg13g2_decap_8 FILLER_29_295 ();
 sg13g2_decap_4 FILLER_29_302 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_decap_4 FILLER_29_338 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_138 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_decap_4 FILLER_30_197 ();
 sg13g2_fill_2 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_decap_4 FILLER_30_283 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_297 ();
 sg13g2_fill_1 FILLER_30_299 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_fill_2 FILLER_30_351 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_4 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_97 ();
 sg13g2_decap_4 FILLER_31_104 ();
 sg13g2_fill_2 FILLER_31_108 ();
 sg13g2_fill_1 FILLER_31_149 ();
 sg13g2_fill_2 FILLER_31_155 ();
 sg13g2_decap_8 FILLER_31_193 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_fill_2 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_decap_4 FILLER_31_241 ();
 sg13g2_decap_8 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_256 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_decap_8 FILLER_31_269 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_decap_8 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_decap_8 FILLER_31_321 ();
 sg13g2_decap_8 FILLER_31_328 ();
 sg13g2_decap_4 FILLER_31_335 ();
 sg13g2_fill_1 FILLER_31_339 ();
 sg13g2_fill_2 FILLER_31_345 ();
 sg13g2_fill_2 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_4 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_decap_4 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_decap_4 FILLER_32_139 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_88 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_145 ();
 sg13g2_decap_8 FILLER_33_152 ();
 sg13g2_decap_8 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_166 ();
 sg13g2_decap_8 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_decap_4 FILLER_33_189 ();
 sg13g2_fill_1 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_217 ();
 sg13g2_fill_2 FILLER_33_228 ();
 sg13g2_decap_4 FILLER_33_256 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_348 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_69 ();
 sg13g2_decap_4 FILLER_34_74 ();
 sg13g2_decap_8 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_fill_2 FILLER_34_118 ();
 sg13g2_fill_2 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_155 ();
 sg13g2_decap_4 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_decap_4 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_308 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_330 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_4 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_decap_8 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_decap_4 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_272 ();
 sg13g2_fill_1 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_283 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_294 ();
 sg13g2_decap_4 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_318 ();
 sg13g2_fill_2 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_357 ();
 sg13g2_fill_2 FILLER_35_362 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_1 FILLER_36_181 ();
 sg13g2_fill_2 FILLER_36_212 ();
 sg13g2_decap_8 FILLER_36_218 ();
 sg13g2_decap_4 FILLER_36_225 ();
 sg13g2_fill_1 FILLER_36_229 ();
 sg13g2_fill_2 FILLER_36_238 ();
 sg13g2_fill_1 FILLER_36_240 ();
 sg13g2_decap_4 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_decap_4 FILLER_36_258 ();
 sg13g2_fill_1 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_293 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_316 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_349 ();
 sg13g2_decap_8 FILLER_36_356 ();
 sg13g2_decap_4 FILLER_36_368 ();
 sg13g2_fill_1 FILLER_36_372 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_4 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_decap_4 FILLER_37_105 ();
 sg13g2_fill_2 FILLER_37_142 ();
 sg13g2_fill_2 FILLER_37_162 ();
 sg13g2_fill_1 FILLER_37_164 ();
 sg13g2_decap_8 FILLER_37_185 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_decap_8 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_213 ();
 sg13g2_decap_4 FILLER_37_220 ();
 sg13g2_decap_4 FILLER_37_229 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_decap_4 FILLER_37_313 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_4 FILLER_37_329 ();
 sg13g2_fill_1 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_fill_2 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_373 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_4 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_53 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_4 FILLER_38_207 ();
 sg13g2_fill_2 FILLER_38_211 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_decap_8 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_decap_8 FILLER_38_297 ();
 sg13g2_fill_2 FILLER_38_304 ();
 sg13g2_fill_1 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_339 ();
 sg13g2_fill_1 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_fill_1 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_73 ();
 sg13g2_fill_2 FILLER_39_80 ();
 sg13g2_fill_1 FILLER_39_82 ();
 sg13g2_decap_8 FILLER_39_87 ();
 sg13g2_decap_8 FILLER_39_94 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_fill_1 FILLER_39_103 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_fill_2 FILLER_39_162 ();
 sg13g2_fill_1 FILLER_39_164 ();
 sg13g2_fill_2 FILLER_39_172 ();
 sg13g2_decap_4 FILLER_39_178 ();
 sg13g2_decap_8 FILLER_39_213 ();
 sg13g2_fill_1 FILLER_39_225 ();
 sg13g2_fill_2 FILLER_39_233 ();
 sg13g2_fill_1 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_268 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_290 ();
 sg13g2_fill_2 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_370 ();
 sg13g2_decap_8 FILLER_39_377 ();
 sg13g2_decap_8 FILLER_39_388 ();
 sg13g2_decap_8 FILLER_39_395 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_4 FILLER_40_63 ();
 sg13g2_fill_1 FILLER_40_71 ();
 sg13g2_decap_8 FILLER_40_102 ();
 sg13g2_decap_8 FILLER_40_109 ();
 sg13g2_fill_1 FILLER_40_133 ();
 sg13g2_fill_2 FILLER_40_144 ();
 sg13g2_fill_1 FILLER_40_146 ();
 sg13g2_fill_1 FILLER_40_165 ();
 sg13g2_fill_2 FILLER_40_170 ();
 sg13g2_fill_1 FILLER_40_195 ();
 sg13g2_decap_4 FILLER_40_242 ();
 sg13g2_fill_2 FILLER_40_254 ();
 sg13g2_fill_1 FILLER_40_256 ();
 sg13g2_fill_1 FILLER_40_292 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_decap_4 FILLER_40_321 ();
 sg13g2_fill_2 FILLER_40_325 ();
 sg13g2_fill_2 FILLER_40_340 ();
 sg13g2_fill_2 FILLER_40_370 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_49 ();
 sg13g2_fill_1 FILLER_41_51 ();
 sg13g2_fill_1 FILLER_41_130 ();
 sg13g2_fill_1 FILLER_41_187 ();
 sg13g2_fill_1 FILLER_41_192 ();
 sg13g2_decap_4 FILLER_41_219 ();
 sg13g2_fill_2 FILLER_41_239 ();
 sg13g2_fill_1 FILLER_41_241 ();
 sg13g2_decap_8 FILLER_41_263 ();
 sg13g2_fill_2 FILLER_41_291 ();
 sg13g2_fill_1 FILLER_41_293 ();
 sg13g2_fill_2 FILLER_41_318 ();
 sg13g2_fill_1 FILLER_41_320 ();
 sg13g2_fill_1 FILLER_41_326 ();
 sg13g2_decap_8 FILLER_41_331 ();
 sg13g2_fill_2 FILLER_41_338 ();
 sg13g2_fill_1 FILLER_41_340 ();
 sg13g2_fill_2 FILLER_41_392 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_4 FILLER_42_42 ();
 sg13g2_fill_1 FILLER_42_46 ();
 sg13g2_fill_1 FILLER_42_82 ();
 sg13g2_fill_2 FILLER_42_103 ();
 sg13g2_fill_1 FILLER_42_138 ();
 sg13g2_fill_2 FILLER_42_179 ();
 sg13g2_decap_8 FILLER_42_207 ();
 sg13g2_decap_8 FILLER_42_214 ();
 sg13g2_fill_1 FILLER_42_221 ();
 sg13g2_decap_4 FILLER_42_234 ();
 sg13g2_fill_1 FILLER_42_238 ();
 sg13g2_fill_1 FILLER_42_244 ();
 sg13g2_fill_2 FILLER_42_275 ();
 sg13g2_fill_1 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_fill_1 FILLER_42_317 ();
 sg13g2_fill_2 FILLER_42_339 ();
 sg13g2_fill_1 FILLER_42_341 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_fill_1 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_fill_1 FILLER_43_49 ();
 sg13g2_fill_2 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_78 ();
 sg13g2_fill_1 FILLER_43_114 ();
 sg13g2_fill_2 FILLER_43_154 ();
 sg13g2_fill_1 FILLER_43_156 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_174 ();
 sg13g2_fill_1 FILLER_43_183 ();
 sg13g2_decap_8 FILLER_43_197 ();
 sg13g2_decap_8 FILLER_43_204 ();
 sg13g2_decap_8 FILLER_43_211 ();
 sg13g2_decap_8 FILLER_43_218 ();
 sg13g2_decap_8 FILLER_43_236 ();
 sg13g2_fill_1 FILLER_43_243 ();
 sg13g2_fill_2 FILLER_43_275 ();
 sg13g2_fill_1 FILLER_43_277 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_349 ();
 sg13g2_decap_8 FILLER_43_395 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_fill_2 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_58 ();
 sg13g2_fill_2 FILLER_44_93 ();
 sg13g2_fill_1 FILLER_44_95 ();
 sg13g2_fill_2 FILLER_44_109 ();
 sg13g2_fill_1 FILLER_44_115 ();
 sg13g2_decap_4 FILLER_44_124 ();
 sg13g2_fill_2 FILLER_44_154 ();
 sg13g2_fill_1 FILLER_44_156 ();
 sg13g2_fill_1 FILLER_44_164 ();
 sg13g2_decap_8 FILLER_44_172 ();
 sg13g2_decap_4 FILLER_44_179 ();
 sg13g2_fill_2 FILLER_44_188 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_decap_8 FILLER_44_242 ();
 sg13g2_fill_2 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_fill_2 FILLER_44_301 ();
 sg13g2_fill_1 FILLER_44_303 ();
 sg13g2_decap_8 FILLER_44_309 ();
 sg13g2_decap_8 FILLER_44_316 ();
 sg13g2_decap_8 FILLER_44_323 ();
 sg13g2_fill_2 FILLER_44_333 ();
 sg13g2_decap_8 FILLER_44_340 ();
 sg13g2_decap_8 FILLER_44_347 ();
 sg13g2_decap_8 FILLER_44_354 ();
 sg13g2_decap_4 FILLER_44_388 ();
 sg13g2_fill_1 FILLER_44_392 ();
 sg13g2_fill_1 FILLER_44_397 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_4 FILLER_45_49 ();
 sg13g2_fill_1 FILLER_45_53 ();
 sg13g2_decap_8 FILLER_45_121 ();
 sg13g2_decap_8 FILLER_45_128 ();
 sg13g2_decap_4 FILLER_45_135 ();
 sg13g2_fill_2 FILLER_45_139 ();
 sg13g2_fill_1 FILLER_45_193 ();
 sg13g2_fill_2 FILLER_45_207 ();
 sg13g2_fill_1 FILLER_45_209 ();
 sg13g2_decap_8 FILLER_45_250 ();
 sg13g2_decap_8 FILLER_45_257 ();
 sg13g2_decap_8 FILLER_45_268 ();
 sg13g2_decap_4 FILLER_45_275 ();
 sg13g2_fill_2 FILLER_45_279 ();
 sg13g2_decap_4 FILLER_45_290 ();
 sg13g2_fill_1 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_319 ();
 sg13g2_fill_1 FILLER_45_326 ();
 sg13g2_fill_2 FILLER_45_352 ();
 sg13g2_fill_1 FILLER_45_354 ();
 sg13g2_fill_1 FILLER_45_381 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_fill_2 FILLER_46_111 ();
 sg13g2_decap_8 FILLER_46_118 ();
 sg13g2_decap_8 FILLER_46_125 ();
 sg13g2_decap_8 FILLER_46_132 ();
 sg13g2_fill_2 FILLER_46_143 ();
 sg13g2_fill_1 FILLER_46_145 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_fill_2 FILLER_46_175 ();
 sg13g2_fill_1 FILLER_46_177 ();
 sg13g2_decap_4 FILLER_46_182 ();
 sg13g2_decap_4 FILLER_46_202 ();
 sg13g2_fill_1 FILLER_46_230 ();
 sg13g2_decap_4 FILLER_46_260 ();
 sg13g2_fill_1 FILLER_46_264 ();
 sg13g2_decap_4 FILLER_46_278 ();
 sg13g2_fill_1 FILLER_46_282 ();
 sg13g2_fill_1 FILLER_46_300 ();
 sg13g2_decap_8 FILLER_46_330 ();
 sg13g2_fill_1 FILLER_46_337 ();
 sg13g2_decap_4 FILLER_46_343 ();
 sg13g2_fill_1 FILLER_46_347 ();
 sg13g2_fill_2 FILLER_46_360 ();
 sg13g2_fill_1 FILLER_46_362 ();
 sg13g2_fill_2 FILLER_46_398 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_4 FILLER_47_63 ();
 sg13g2_fill_2 FILLER_47_71 ();
 sg13g2_fill_1 FILLER_47_73 ();
 sg13g2_fill_2 FILLER_47_83 ();
 sg13g2_fill_1 FILLER_47_85 ();
 sg13g2_decap_4 FILLER_47_89 ();
 sg13g2_fill_1 FILLER_47_93 ();
 sg13g2_decap_8 FILLER_47_132 ();
 sg13g2_decap_8 FILLER_47_139 ();
 sg13g2_decap_4 FILLER_47_146 ();
 sg13g2_fill_2 FILLER_47_150 ();
 sg13g2_decap_8 FILLER_47_156 ();
 sg13g2_decap_8 FILLER_47_167 ();
 sg13g2_decap_4 FILLER_47_174 ();
 sg13g2_fill_1 FILLER_47_178 ();
 sg13g2_decap_4 FILLER_47_187 ();
 sg13g2_fill_2 FILLER_47_282 ();
 sg13g2_fill_1 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_293 ();
 sg13g2_decap_4 FILLER_47_342 ();
 sg13g2_decap_4 FILLER_47_351 ();
 sg13g2_fill_1 FILLER_47_355 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_51 ();
 sg13g2_decap_4 FILLER_48_78 ();
 sg13g2_decap_4 FILLER_48_126 ();
 sg13g2_fill_2 FILLER_48_130 ();
 sg13g2_fill_1 FILLER_48_137 ();
 sg13g2_fill_1 FILLER_48_172 ();
 sg13g2_fill_2 FILLER_48_178 ();
 sg13g2_fill_1 FILLER_48_180 ();
 sg13g2_fill_1 FILLER_48_185 ();
 sg13g2_decap_8 FILLER_48_195 ();
 sg13g2_fill_2 FILLER_48_202 ();
 sg13g2_fill_1 FILLER_48_204 ();
 sg13g2_decap_4 FILLER_48_221 ();
 sg13g2_fill_2 FILLER_48_234 ();
 sg13g2_fill_1 FILLER_48_244 ();
 sg13g2_fill_2 FILLER_48_249 ();
 sg13g2_fill_2 FILLER_48_260 ();
 sg13g2_fill_1 FILLER_48_262 ();
 sg13g2_fill_1 FILLER_48_316 ();
 sg13g2_fill_2 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_333 ();
 sg13g2_decap_8 FILLER_48_340 ();
 sg13g2_fill_2 FILLER_48_347 ();
 sg13g2_fill_2 FILLER_48_361 ();
 sg13g2_fill_1 FILLER_48_363 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_4 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_46 ();
 sg13g2_fill_1 FILLER_49_82 ();
 sg13g2_fill_1 FILLER_49_114 ();
 sg13g2_fill_2 FILLER_49_175 ();
 sg13g2_fill_2 FILLER_49_185 ();
 sg13g2_decap_4 FILLER_49_206 ();
 sg13g2_fill_2 FILLER_49_210 ();
 sg13g2_fill_1 FILLER_49_221 ();
 sg13g2_fill_2 FILLER_49_227 ();
 sg13g2_decap_8 FILLER_49_240 ();
 sg13g2_decap_4 FILLER_49_247 ();
 sg13g2_fill_1 FILLER_49_251 ();
 sg13g2_decap_4 FILLER_49_271 ();
 sg13g2_fill_2 FILLER_49_275 ();
 sg13g2_fill_1 FILLER_49_302 ();
 sg13g2_fill_1 FILLER_49_310 ();
 sg13g2_fill_2 FILLER_49_321 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_decap_4 FILLER_49_357 ();
 sg13g2_fill_2 FILLER_49_368 ();
 sg13g2_fill_1 FILLER_49_383 ();
 sg13g2_decap_8 FILLER_49_401 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_4 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_150 ();
 sg13g2_fill_1 FILLER_50_173 ();
 sg13g2_fill_1 FILLER_50_198 ();
 sg13g2_decap_8 FILLER_50_226 ();
 sg13g2_decap_4 FILLER_50_233 ();
 sg13g2_fill_2 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_253 ();
 sg13g2_decap_8 FILLER_50_260 ();
 sg13g2_decap_8 FILLER_50_267 ();
 sg13g2_decap_8 FILLER_50_274 ();
 sg13g2_decap_4 FILLER_50_281 ();
 sg13g2_fill_2 FILLER_50_295 ();
 sg13g2_fill_2 FILLER_50_317 ();
 sg13g2_fill_2 FILLER_50_340 ();
 sg13g2_fill_1 FILLER_50_342 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_fill_1 FILLER_51_56 ();
 sg13g2_fill_2 FILLER_51_83 ();
 sg13g2_fill_1 FILLER_51_101 ();
 sg13g2_fill_2 FILLER_51_135 ();
 sg13g2_fill_2 FILLER_51_145 ();
 sg13g2_fill_1 FILLER_51_163 ();
 sg13g2_fill_2 FILLER_51_177 ();
 sg13g2_fill_1 FILLER_51_179 ();
 sg13g2_decap_8 FILLER_51_210 ();
 sg13g2_decap_8 FILLER_51_225 ();
 sg13g2_decap_4 FILLER_51_236 ();
 sg13g2_fill_2 FILLER_51_274 ();
 sg13g2_fill_2 FILLER_51_289 ();
 sg13g2_fill_1 FILLER_51_291 ();
 sg13g2_fill_1 FILLER_51_316 ();
 sg13g2_fill_1 FILLER_51_346 ();
 sg13g2_decap_4 FILLER_51_367 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_fill_1 FILLER_52_63 ();
 sg13g2_fill_2 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_83 ();
 sg13g2_decap_4 FILLER_52_90 ();
 sg13g2_fill_2 FILLER_52_104 ();
 sg13g2_fill_1 FILLER_52_106 ();
 sg13g2_fill_2 FILLER_52_120 ();
 sg13g2_fill_2 FILLER_52_157 ();
 sg13g2_fill_2 FILLER_52_163 ();
 sg13g2_decap_8 FILLER_52_173 ();
 sg13g2_decap_4 FILLER_52_180 ();
 sg13g2_fill_1 FILLER_52_184 ();
 sg13g2_fill_2 FILLER_52_232 ();
 sg13g2_fill_2 FILLER_52_257 ();
 sg13g2_fill_1 FILLER_52_299 ();
 sg13g2_fill_2 FILLER_52_304 ();
 sg13g2_fill_1 FILLER_52_306 ();
 sg13g2_decap_8 FILLER_52_312 ();
 sg13g2_decap_4 FILLER_52_319 ();
 sg13g2_fill_1 FILLER_52_323 ();
 sg13g2_decap_8 FILLER_52_337 ();
 sg13g2_decap_8 FILLER_52_344 ();
 sg13g2_decap_8 FILLER_52_351 ();
 sg13g2_fill_2 FILLER_52_358 ();
 sg13g2_fill_1 FILLER_52_365 ();
 sg13g2_fill_2 FILLER_52_371 ();
 sg13g2_fill_1 FILLER_52_373 ();
 sg13g2_decap_4 FILLER_52_378 ();
 sg13g2_fill_1 FILLER_52_386 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_4 FILLER_53_42 ();
 sg13g2_fill_2 FILLER_53_46 ();
 sg13g2_decap_4 FILLER_53_52 ();
 sg13g2_fill_1 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_83 ();
 sg13g2_fill_1 FILLER_53_90 ();
 sg13g2_fill_2 FILLER_53_95 ();
 sg13g2_fill_2 FILLER_53_102 ();
 sg13g2_decap_4 FILLER_53_117 ();
 sg13g2_fill_1 FILLER_53_136 ();
 sg13g2_fill_1 FILLER_53_151 ();
 sg13g2_fill_1 FILLER_53_156 ();
 sg13g2_decap_8 FILLER_53_163 ();
 sg13g2_decap_8 FILLER_53_170 ();
 sg13g2_decap_8 FILLER_53_177 ();
 sg13g2_fill_2 FILLER_53_184 ();
 sg13g2_decap_4 FILLER_53_194 ();
 sg13g2_fill_1 FILLER_53_198 ();
 sg13g2_fill_1 FILLER_53_226 ();
 sg13g2_fill_1 FILLER_53_308 ();
 sg13g2_fill_2 FILLER_53_327 ();
 sg13g2_fill_1 FILLER_53_334 ();
 sg13g2_fill_2 FILLER_53_340 ();
 sg13g2_fill_1 FILLER_53_342 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_42 ();
 sg13g2_fill_2 FILLER_54_78 ();
 sg13g2_fill_2 FILLER_54_106 ();
 sg13g2_fill_1 FILLER_54_122 ();
 sg13g2_decap_8 FILLER_54_137 ();
 sg13g2_decap_8 FILLER_54_144 ();
 sg13g2_fill_2 FILLER_54_151 ();
 sg13g2_fill_1 FILLER_54_153 ();
 sg13g2_decap_8 FILLER_54_183 ();
 sg13g2_fill_2 FILLER_54_190 ();
 sg13g2_fill_2 FILLER_54_214 ();
 sg13g2_fill_2 FILLER_54_221 ();
 sg13g2_fill_1 FILLER_54_223 ();
 sg13g2_fill_1 FILLER_54_250 ();
 sg13g2_decap_8 FILLER_54_282 ();
 sg13g2_decap_8 FILLER_54_289 ();
 sg13g2_fill_2 FILLER_54_303 ();
 sg13g2_fill_2 FILLER_54_323 ();
 sg13g2_fill_2 FILLER_54_381 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_fill_2 FILLER_55_56 ();
 sg13g2_decap_4 FILLER_55_84 ();
 sg13g2_fill_1 FILLER_55_88 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_fill_1 FILLER_55_112 ();
 sg13g2_fill_2 FILLER_55_138 ();
 sg13g2_fill_1 FILLER_55_140 ();
 sg13g2_decap_4 FILLER_55_150 ();
 sg13g2_fill_1 FILLER_55_154 ();
 sg13g2_decap_4 FILLER_55_191 ();
 sg13g2_fill_1 FILLER_55_195 ();
 sg13g2_fill_1 FILLER_55_220 ();
 sg13g2_fill_1 FILLER_55_230 ();
 sg13g2_fill_1 FILLER_55_239 ();
 sg13g2_decap_8 FILLER_55_271 ();
 sg13g2_fill_2 FILLER_55_283 ();
 sg13g2_fill_1 FILLER_55_293 ();
 sg13g2_fill_2 FILLER_55_316 ();
 sg13g2_fill_2 FILLER_55_334 ();
 sg13g2_fill_1 FILLER_55_336 ();
 sg13g2_fill_2 FILLER_55_347 ();
 sg13g2_decap_4 FILLER_55_388 ();
 sg13g2_fill_2 FILLER_55_392 ();
 sg13g2_fill_2 FILLER_55_398 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_fill_2 FILLER_56_56 ();
 sg13g2_fill_2 FILLER_56_97 ();
 sg13g2_decap_4 FILLER_56_117 ();
 sg13g2_fill_1 FILLER_56_121 ();
 sg13g2_fill_1 FILLER_56_134 ();
 sg13g2_fill_1 FILLER_56_161 ();
 sg13g2_decap_4 FILLER_56_170 ();
 sg13g2_fill_1 FILLER_56_174 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_fill_1 FILLER_56_201 ();
 sg13g2_fill_1 FILLER_56_216 ();
 sg13g2_decap_8 FILLER_56_237 ();
 sg13g2_decap_4 FILLER_56_244 ();
 sg13g2_fill_1 FILLER_56_261 ();
 sg13g2_decap_4 FILLER_56_266 ();
 sg13g2_fill_1 FILLER_56_270 ();
 sg13g2_fill_1 FILLER_56_312 ();
 sg13g2_fill_2 FILLER_56_321 ();
 sg13g2_fill_1 FILLER_56_349 ();
 sg13g2_fill_1 FILLER_56_354 ();
 sg13g2_decap_8 FILLER_56_376 ();
 sg13g2_fill_2 FILLER_56_383 ();
 sg13g2_decap_8 FILLER_56_389 ();
 sg13g2_fill_2 FILLER_56_396 ();
 sg13g2_decap_8 FILLER_56_402 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_4 FILLER_57_63 ();
 sg13g2_decap_4 FILLER_57_71 ();
 sg13g2_decap_4 FILLER_57_88 ();
 sg13g2_decap_8 FILLER_57_121 ();
 sg13g2_fill_2 FILLER_57_151 ();
 sg13g2_fill_1 FILLER_57_153 ();
 sg13g2_decap_4 FILLER_57_180 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_fill_2 FILLER_57_196 ();
 sg13g2_fill_1 FILLER_57_198 ();
 sg13g2_decap_4 FILLER_57_212 ();
 sg13g2_fill_2 FILLER_57_216 ();
 sg13g2_fill_2 FILLER_57_235 ();
 sg13g2_fill_1 FILLER_57_237 ();
 sg13g2_decap_8 FILLER_57_251 ();
 sg13g2_decap_8 FILLER_57_258 ();
 sg13g2_decap_8 FILLER_57_265 ();
 sg13g2_decap_8 FILLER_57_272 ();
 sg13g2_fill_2 FILLER_57_279 ();
 sg13g2_fill_2 FILLER_57_289 ();
 sg13g2_fill_1 FILLER_57_291 ();
 sg13g2_decap_8 FILLER_57_337 ();
 sg13g2_decap_4 FILLER_57_344 ();
 sg13g2_fill_2 FILLER_57_348 ();
 sg13g2_fill_1 FILLER_57_363 ();
 sg13g2_fill_2 FILLER_57_372 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_fill_2 FILLER_58_63 ();
 sg13g2_fill_1 FILLER_58_65 ();
 sg13g2_fill_2 FILLER_58_92 ();
 sg13g2_fill_1 FILLER_58_103 ();
 sg13g2_decap_8 FILLER_58_125 ();
 sg13g2_decap_4 FILLER_58_132 ();
 sg13g2_fill_2 FILLER_58_141 ();
 sg13g2_decap_8 FILLER_58_156 ();
 sg13g2_fill_2 FILLER_58_163 ();
 sg13g2_decap_8 FILLER_58_169 ();
 sg13g2_decap_8 FILLER_58_176 ();
 sg13g2_fill_2 FILLER_58_183 ();
 sg13g2_fill_1 FILLER_58_185 ();
 sg13g2_fill_2 FILLER_58_199 ();
 sg13g2_fill_2 FILLER_58_222 ();
 sg13g2_fill_1 FILLER_58_224 ();
 sg13g2_fill_1 FILLER_58_249 ();
 sg13g2_fill_2 FILLER_58_263 ();
 sg13g2_decap_8 FILLER_58_269 ();
 sg13g2_fill_2 FILLER_58_276 ();
 sg13g2_fill_1 FILLER_58_278 ();
 sg13g2_fill_1 FILLER_58_283 ();
 sg13g2_fill_1 FILLER_58_324 ();
 sg13g2_decap_8 FILLER_58_330 ();
 sg13g2_decap_8 FILLER_58_337 ();
 sg13g2_fill_2 FILLER_58_344 ();
 sg13g2_fill_1 FILLER_58_346 ();
 sg13g2_fill_1 FILLER_58_350 ();
 sg13g2_fill_2 FILLER_58_362 ();
 sg13g2_decap_4 FILLER_58_403 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_81 ();
 sg13g2_fill_2 FILLER_59_88 ();
 sg13g2_fill_1 FILLER_59_90 ();
 sg13g2_fill_2 FILLER_59_116 ();
 sg13g2_fill_2 FILLER_59_139 ();
 sg13g2_fill_2 FILLER_59_149 ();
 sg13g2_decap_4 FILLER_59_169 ();
 sg13g2_fill_2 FILLER_59_173 ();
 sg13g2_fill_1 FILLER_59_201 ();
 sg13g2_decap_4 FILLER_59_211 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_fill_2 FILLER_59_250 ();
 sg13g2_fill_1 FILLER_59_252 ();
 sg13g2_decap_8 FILLER_59_314 ();
 sg13g2_decap_8 FILLER_59_321 ();
 sg13g2_decap_8 FILLER_59_328 ();
 sg13g2_fill_2 FILLER_59_335 ();
 sg13g2_decap_8 FILLER_59_375 ();
 sg13g2_decap_4 FILLER_59_382 ();
 sg13g2_fill_2 FILLER_59_386 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_4 FILLER_60_63 ();
 sg13g2_fill_1 FILLER_60_67 ();
 sg13g2_fill_1 FILLER_60_108 ();
 sg13g2_decap_4 FILLER_60_144 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_fill_1 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_275 ();
 sg13g2_decap_8 FILLER_60_290 ();
 sg13g2_decap_8 FILLER_60_297 ();
 sg13g2_decap_8 FILLER_60_304 ();
 sg13g2_decap_4 FILLER_60_311 ();
 sg13g2_fill_1 FILLER_60_315 ();
 sg13g2_decap_8 FILLER_60_324 ();
 sg13g2_decap_4 FILLER_60_331 ();
 sg13g2_fill_1 FILLER_60_335 ();
 sg13g2_decap_4 FILLER_60_343 ();
 sg13g2_fill_1 FILLER_60_347 ();
 sg13g2_decap_4 FILLER_60_365 ();
 sg13g2_decap_8 FILLER_60_395 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_fill_2 FILLER_61_63 ();
 sg13g2_fill_2 FILLER_61_91 ();
 sg13g2_fill_2 FILLER_61_137 ();
 sg13g2_fill_1 FILLER_61_139 ();
 sg13g2_fill_2 FILLER_61_154 ();
 sg13g2_fill_2 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_189 ();
 sg13g2_decap_4 FILLER_61_221 ();
 sg13g2_fill_1 FILLER_61_233 ();
 sg13g2_fill_2 FILLER_61_246 ();
 sg13g2_decap_4 FILLER_61_297 ();
 sg13g2_fill_1 FILLER_61_301 ();
 sg13g2_decap_4 FILLER_61_322 ();
 sg13g2_fill_2 FILLER_61_326 ();
 sg13g2_fill_2 FILLER_61_336 ();
 sg13g2_fill_2 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_396 ();
 sg13g2_decap_4 FILLER_61_403 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_fill_2 FILLER_62_63 ();
 sg13g2_fill_2 FILLER_62_74 ();
 sg13g2_fill_1 FILLER_62_76 ();
 sg13g2_decap_4 FILLER_62_109 ();
 sg13g2_fill_2 FILLER_62_121 ();
 sg13g2_fill_1 FILLER_62_131 ();
 sg13g2_decap_8 FILLER_62_167 ();
 sg13g2_decap_8 FILLER_62_174 ();
 sg13g2_fill_1 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_194 ();
 sg13g2_decap_4 FILLER_62_216 ();
 sg13g2_fill_2 FILLER_62_220 ();
 sg13g2_decap_4 FILLER_62_235 ();
 sg13g2_fill_2 FILLER_62_239 ();
 sg13g2_fill_2 FILLER_62_262 ();
 sg13g2_fill_1 FILLER_62_264 ();
 sg13g2_decap_8 FILLER_62_277 ();
 sg13g2_decap_8 FILLER_62_284 ();
 sg13g2_decap_8 FILLER_62_291 ();
 sg13g2_decap_4 FILLER_62_298 ();
 sg13g2_fill_1 FILLER_62_302 ();
 sg13g2_fill_2 FILLER_62_313 ();
 sg13g2_fill_2 FILLER_62_349 ();
 sg13g2_decap_4 FILLER_62_404 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_fill_2 FILLER_63_63 ();
 sg13g2_decap_4 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_109 ();
 sg13g2_decap_4 FILLER_63_118 ();
 sg13g2_fill_1 FILLER_63_122 ();
 sg13g2_fill_1 FILLER_63_150 ();
 sg13g2_fill_1 FILLER_63_160 ();
 sg13g2_fill_2 FILLER_63_220 ();
 sg13g2_decap_8 FILLER_63_247 ();
 sg13g2_fill_1 FILLER_63_254 ();
 sg13g2_decap_8 FILLER_63_265 ();
 sg13g2_decap_4 FILLER_63_272 ();
 sg13g2_decap_8 FILLER_63_288 ();
 sg13g2_fill_1 FILLER_63_295 ();
 sg13g2_fill_2 FILLER_63_303 ();
 sg13g2_fill_1 FILLER_63_305 ();
 sg13g2_fill_2 FILLER_63_311 ();
 sg13g2_fill_2 FILLER_63_317 ();
 sg13g2_fill_2 FILLER_63_331 ();
 sg13g2_fill_1 FILLER_63_333 ();
 sg13g2_decap_4 FILLER_63_338 ();
 sg13g2_fill_2 FILLER_63_372 ();
 sg13g2_fill_2 FILLER_63_383 ();
 sg13g2_fill_1 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_395 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_fill_2 FILLER_64_56 ();
 sg13g2_fill_1 FILLER_64_58 ();
 sg13g2_fill_1 FILLER_64_111 ();
 sg13g2_decap_4 FILLER_64_146 ();
 sg13g2_fill_2 FILLER_64_150 ();
 sg13g2_decap_8 FILLER_64_155 ();
 sg13g2_fill_2 FILLER_64_162 ();
 sg13g2_fill_1 FILLER_64_176 ();
 sg13g2_fill_2 FILLER_64_192 ();
 sg13g2_fill_1 FILLER_64_211 ();
 sg13g2_fill_1 FILLER_64_233 ();
 sg13g2_fill_2 FILLER_64_239 ();
 sg13g2_fill_1 FILLER_64_241 ();
 sg13g2_fill_1 FILLER_64_267 ();
 sg13g2_decap_8 FILLER_64_282 ();
 sg13g2_fill_2 FILLER_64_289 ();
 sg13g2_fill_1 FILLER_64_291 ();
 sg13g2_fill_2 FILLER_64_307 ();
 sg13g2_fill_2 FILLER_64_344 ();
 sg13g2_fill_1 FILLER_64_346 ();
 sg13g2_decap_8 FILLER_64_382 ();
 sg13g2_decap_8 FILLER_64_389 ();
 sg13g2_decap_8 FILLER_64_396 ();
 sg13g2_decap_4 FILLER_64_403 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_fill_1 FILLER_65_111 ();
 sg13g2_fill_2 FILLER_65_124 ();
 sg13g2_fill_1 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_148 ();
 sg13g2_decap_8 FILLER_65_155 ();
 sg13g2_decap_8 FILLER_65_162 ();
 sg13g2_decap_4 FILLER_65_169 ();
 sg13g2_fill_1 FILLER_65_173 ();
 sg13g2_fill_2 FILLER_65_181 ();
 sg13g2_fill_1 FILLER_65_183 ();
 sg13g2_fill_2 FILLER_65_192 ();
 sg13g2_fill_1 FILLER_65_220 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_fill_2 FILLER_65_289 ();
 sg13g2_fill_1 FILLER_65_308 ();
 sg13g2_fill_1 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_349 ();
 sg13g2_decap_8 FILLER_65_389 ();
 sg13g2_decap_8 FILLER_65_396 ();
 sg13g2_decap_4 FILLER_65_403 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_fill_2 FILLER_66_84 ();
 sg13g2_fill_1 FILLER_66_92 ();
 sg13g2_fill_1 FILLER_66_102 ();
 sg13g2_fill_1 FILLER_66_116 ();
 sg13g2_fill_2 FILLER_66_129 ();
 sg13g2_fill_1 FILLER_66_131 ();
 sg13g2_fill_2 FILLER_66_140 ();
 sg13g2_fill_1 FILLER_66_142 ();
 sg13g2_fill_2 FILLER_66_178 ();
 sg13g2_decap_4 FILLER_66_195 ();
 sg13g2_decap_8 FILLER_66_211 ();
 sg13g2_fill_1 FILLER_66_218 ();
 sg13g2_fill_1 FILLER_66_231 ();
 sg13g2_decap_4 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_241 ();
 sg13g2_fill_2 FILLER_66_255 ();
 sg13g2_fill_1 FILLER_66_257 ();
 sg13g2_decap_4 FILLER_66_271 ();
 sg13g2_decap_8 FILLER_66_402 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_4 FILLER_67_84 ();
 sg13g2_fill_1 FILLER_67_134 ();
 sg13g2_decap_4 FILLER_67_140 ();
 sg13g2_fill_2 FILLER_67_144 ();
 sg13g2_decap_4 FILLER_67_172 ();
 sg13g2_fill_1 FILLER_67_176 ();
 sg13g2_decap_8 FILLER_67_200 ();
 sg13g2_decap_8 FILLER_67_207 ();
 sg13g2_decap_4 FILLER_67_214 ();
 sg13g2_decap_8 FILLER_67_225 ();
 sg13g2_decap_8 FILLER_67_232 ();
 sg13g2_decap_8 FILLER_67_239 ();
 sg13g2_fill_2 FILLER_67_246 ();
 sg13g2_fill_1 FILLER_67_248 ();
 sg13g2_decap_8 FILLER_67_262 ();
 sg13g2_decap_8 FILLER_67_269 ();
 sg13g2_fill_1 FILLER_67_276 ();
 sg13g2_fill_2 FILLER_67_306 ();
 sg13g2_fill_1 FILLER_67_308 ();
 sg13g2_fill_1 FILLER_67_326 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_fill_2 FILLER_68_77 ();
 sg13g2_fill_1 FILLER_68_79 ();
 sg13g2_decap_8 FILLER_68_106 ();
 sg13g2_decap_4 FILLER_68_113 ();
 sg13g2_decap_8 FILLER_68_121 ();
 sg13g2_fill_2 FILLER_68_128 ();
 sg13g2_fill_1 FILLER_68_130 ();
 sg13g2_fill_1 FILLER_68_134 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_4 FILLER_68_162 ();
 sg13g2_fill_2 FILLER_68_170 ();
 sg13g2_fill_1 FILLER_68_172 ();
 sg13g2_decap_8 FILLER_68_178 ();
 sg13g2_decap_4 FILLER_68_185 ();
 sg13g2_decap_8 FILLER_68_192 ();
 sg13g2_decap_8 FILLER_68_199 ();
 sg13g2_fill_2 FILLER_68_206 ();
 sg13g2_fill_1 FILLER_68_208 ();
 sg13g2_decap_8 FILLER_68_234 ();
 sg13g2_decap_8 FILLER_68_253 ();
 sg13g2_fill_1 FILLER_68_260 ();
 sg13g2_decap_4 FILLER_68_297 ();
 sg13g2_fill_2 FILLER_68_301 ();
 sg13g2_decap_4 FILLER_68_307 ();
 sg13g2_fill_2 FILLER_68_311 ();
 sg13g2_fill_2 FILLER_68_325 ();
 sg13g2_decap_8 FILLER_68_334 ();
 sg13g2_fill_1 FILLER_68_341 ();
 sg13g2_fill_1 FILLER_68_346 ();
 sg13g2_fill_1 FILLER_68_361 ();
 sg13g2_decap_8 FILLER_68_396 ();
 sg13g2_decap_4 FILLER_68_403 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_fill_2 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_4 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_140 ();
 sg13g2_fill_2 FILLER_69_156 ();
 sg13g2_decap_4 FILLER_69_194 ();
 sg13g2_fill_1 FILLER_69_241 ();
 sg13g2_decap_8 FILLER_69_258 ();
 sg13g2_decap_8 FILLER_69_265 ();
 sg13g2_decap_4 FILLER_69_272 ();
 sg13g2_fill_2 FILLER_69_292 ();
 sg13g2_fill_1 FILLER_69_299 ();
 sg13g2_fill_2 FILLER_69_308 ();
 sg13g2_decap_8 FILLER_69_323 ();
 sg13g2_decap_8 FILLER_69_330 ();
 sg13g2_decap_8 FILLER_69_337 ();
 sg13g2_fill_1 FILLER_69_344 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_4 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_fill_2 FILLER_70_95 ();
 sg13g2_fill_1 FILLER_70_101 ();
 sg13g2_fill_1 FILLER_70_111 ();
 sg13g2_fill_2 FILLER_70_206 ();
 sg13g2_fill_1 FILLER_70_208 ();
 sg13g2_fill_1 FILLER_70_213 ();
 sg13g2_decap_4 FILLER_70_220 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_decap_8 FILLER_70_261 ();
 sg13g2_decap_8 FILLER_70_268 ();
 sg13g2_decap_4 FILLER_70_275 ();
 sg13g2_fill_1 FILLER_70_279 ();
 sg13g2_fill_2 FILLER_70_296 ();
 sg13g2_fill_1 FILLER_70_298 ();
 sg13g2_fill_1 FILLER_70_307 ();
 sg13g2_decap_4 FILLER_70_313 ();
 sg13g2_fill_1 FILLER_70_317 ();
 sg13g2_decap_8 FILLER_70_342 ();
 sg13g2_decap_8 FILLER_70_349 ();
 sg13g2_decap_8 FILLER_70_360 ();
 sg13g2_decap_8 FILLER_70_367 ();
 sg13g2_decap_8 FILLER_70_374 ();
 sg13g2_decap_8 FILLER_70_381 ();
 sg13g2_decap_4 FILLER_70_388 ();
 sg13g2_decap_8 FILLER_70_401 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_fill_2 FILLER_71_159 ();
 sg13g2_fill_2 FILLER_71_236 ();
 sg13g2_fill_1 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_247 ();
 sg13g2_fill_2 FILLER_71_254 ();
 sg13g2_decap_4 FILLER_71_281 ();
 sg13g2_decap_4 FILLER_71_290 ();
 sg13g2_fill_2 FILLER_71_294 ();
 sg13g2_fill_1 FILLER_71_304 ();
 sg13g2_decap_4 FILLER_71_321 ();
 sg13g2_fill_2 FILLER_71_325 ();
 sg13g2_decap_8 FILLER_71_354 ();
 sg13g2_fill_2 FILLER_71_361 ();
 sg13g2_decap_8 FILLER_71_367 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_399 ();
 sg13g2_fill_2 FILLER_71_406 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_4 FILLER_72_91 ();
 sg13g2_fill_1 FILLER_72_104 ();
 sg13g2_decap_4 FILLER_72_177 ();
 sg13g2_fill_2 FILLER_72_181 ();
 sg13g2_decap_8 FILLER_72_187 ();
 sg13g2_fill_2 FILLER_72_194 ();
 sg13g2_fill_2 FILLER_72_251 ();
 sg13g2_fill_1 FILLER_72_253 ();
 sg13g2_fill_2 FILLER_72_302 ();
 sg13g2_fill_1 FILLER_72_304 ();
 sg13g2_fill_2 FILLER_72_322 ();
 sg13g2_fill_1 FILLER_72_324 ();
 sg13g2_decap_4 FILLER_72_359 ();
 sg13g2_decap_8 FILLER_72_389 ();
 sg13g2_decap_8 FILLER_72_396 ();
 sg13g2_decap_4 FILLER_72_403 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_fill_2 FILLER_73_98 ();
 sg13g2_fill_1 FILLER_73_100 ();
 sg13g2_fill_2 FILLER_73_170 ();
 sg13g2_fill_2 FILLER_73_198 ();
 sg13g2_fill_2 FILLER_73_209 ();
 sg13g2_fill_2 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_248 ();
 sg13g2_fill_1 FILLER_73_262 ();
 sg13g2_decap_8 FILLER_73_275 ();
 sg13g2_fill_1 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_292 ();
 sg13g2_decap_8 FILLER_73_299 ();
 sg13g2_decap_4 FILLER_73_306 ();
 sg13g2_fill_1 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_391 ();
 sg13g2_decap_8 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_fill_1 FILLER_74_112 ();
 sg13g2_decap_4 FILLER_74_169 ();
 sg13g2_fill_2 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_184 ();
 sg13g2_fill_2 FILLER_74_211 ();
 sg13g2_decap_8 FILLER_74_268 ();
 sg13g2_fill_2 FILLER_74_275 ();
 sg13g2_fill_1 FILLER_74_277 ();
 sg13g2_decap_4 FILLER_74_283 ();
 sg13g2_fill_1 FILLER_74_304 ();
 sg13g2_fill_2 FILLER_74_321 ();
 sg13g2_fill_1 FILLER_74_328 ();
 sg13g2_fill_2 FILLER_74_338 ();
 sg13g2_fill_1 FILLER_74_345 ();
 sg13g2_decap_4 FILLER_74_355 ();
 sg13g2_decap_8 FILLER_74_372 ();
 sg13g2_decap_8 FILLER_74_379 ();
 sg13g2_decap_8 FILLER_74_386 ();
 sg13g2_decap_8 FILLER_74_393 ();
 sg13g2_decap_8 FILLER_74_400 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_fill_2 FILLER_75_119 ();
 sg13g2_fill_1 FILLER_75_121 ();
 sg13g2_decap_8 FILLER_75_157 ();
 sg13g2_decap_4 FILLER_75_164 ();
 sg13g2_fill_1 FILLER_75_168 ();
 sg13g2_decap_4 FILLER_75_216 ();
 sg13g2_fill_2 FILLER_75_220 ();
 sg13g2_decap_4 FILLER_75_230 ();
 sg13g2_fill_1 FILLER_75_234 ();
 sg13g2_fill_2 FILLER_75_260 ();
 sg13g2_fill_1 FILLER_75_262 ();
 sg13g2_fill_2 FILLER_75_275 ();
 sg13g2_fill_1 FILLER_75_277 ();
 sg13g2_fill_2 FILLER_75_287 ();
 sg13g2_fill_2 FILLER_75_336 ();
 sg13g2_fill_1 FILLER_75_338 ();
 sg13g2_fill_2 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_378 ();
 sg13g2_decap_8 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_fill_2 FILLER_75_406 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_fill_2 FILLER_76_191 ();
 sg13g2_decap_8 FILLER_76_223 ();
 sg13g2_decap_8 FILLER_76_230 ();
 sg13g2_decap_4 FILLER_76_237 ();
 sg13g2_fill_1 FILLER_76_241 ();
 sg13g2_decap_8 FILLER_76_255 ();
 sg13g2_fill_2 FILLER_76_262 ();
 sg13g2_fill_2 FILLER_76_312 ();
 sg13g2_fill_1 FILLER_76_327 ();
 sg13g2_fill_2 FILLER_76_354 ();
 sg13g2_fill_1 FILLER_76_360 ();
 sg13g2_decap_8 FILLER_76_370 ();
 sg13g2_decap_8 FILLER_76_377 ();
 sg13g2_decap_8 FILLER_76_384 ();
 sg13g2_decap_8 FILLER_76_391 ();
 sg13g2_decap_8 FILLER_76_398 ();
 sg13g2_decap_4 FILLER_76_405 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_4 FILLER_77_147 ();
 sg13g2_fill_1 FILLER_77_151 ();
 sg13g2_decap_4 FILLER_77_187 ();
 sg13g2_fill_2 FILLER_77_191 ();
 sg13g2_fill_2 FILLER_77_236 ();
 sg13g2_fill_1 FILLER_77_238 ();
 sg13g2_fill_2 FILLER_77_274 ();
 sg13g2_fill_1 FILLER_77_276 ();
 sg13g2_fill_2 FILLER_77_290 ();
 sg13g2_fill_1 FILLER_77_292 ();
 sg13g2_decap_8 FILLER_77_334 ();
 sg13g2_decap_8 FILLER_77_341 ();
 sg13g2_decap_8 FILLER_77_348 ();
 sg13g2_decap_8 FILLER_77_355 ();
 sg13g2_decap_8 FILLER_77_362 ();
 sg13g2_decap_8 FILLER_77_369 ();
 sg13g2_decap_8 FILLER_77_376 ();
 sg13g2_decap_8 FILLER_77_383 ();
 sg13g2_decap_8 FILLER_77_390 ();
 sg13g2_decap_8 FILLER_77_397 ();
 sg13g2_decap_4 FILLER_77_404 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_fill_2 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_156 ();
 sg13g2_decap_4 FILLER_78_161 ();
 sg13g2_fill_2 FILLER_78_165 ();
 sg13g2_fill_2 FILLER_78_175 ();
 sg13g2_fill_1 FILLER_78_177 ();
 sg13g2_decap_8 FILLER_78_239 ();
 sg13g2_fill_1 FILLER_78_246 ();
 sg13g2_fill_1 FILLER_78_268 ();
 sg13g2_fill_2 FILLER_78_292 ();
 sg13g2_fill_2 FILLER_78_322 ();
 sg13g2_fill_1 FILLER_78_324 ();
 sg13g2_decap_8 FILLER_78_351 ();
 sg13g2_decap_8 FILLER_78_358 ();
 sg13g2_decap_8 FILLER_78_365 ();
 sg13g2_decap_8 FILLER_78_372 ();
 sg13g2_decap_8 FILLER_78_379 ();
 sg13g2_decap_8 FILLER_78_386 ();
 sg13g2_decap_8 FILLER_78_393 ();
 sg13g2_decap_8 FILLER_78_400 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_fill_2 FILLER_79_161 ();
 sg13g2_fill_1 FILLER_79_193 ();
 sg13g2_decap_4 FILLER_79_270 ();
 sg13g2_decap_8 FILLER_79_289 ();
 sg13g2_fill_2 FILLER_79_296 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_fill_2 FILLER_79_322 ();
 sg13g2_fill_1 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_8 FILLER_80_123 ();
 sg13g2_decap_8 FILLER_80_130 ();
 sg13g2_decap_8 FILLER_80_137 ();
 sg13g2_decap_8 FILLER_80_144 ();
 sg13g2_decap_8 FILLER_80_151 ();
 sg13g2_decap_8 FILLER_80_158 ();
 sg13g2_decap_8 FILLER_80_165 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_fill_2 FILLER_80_180 ();
 sg13g2_fill_1 FILLER_80_182 ();
 sg13g2_decap_4 FILLER_80_227 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_decap_4 FILLER_80_249 ();
 sg13g2_fill_1 FILLER_80_253 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_decap_4 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_273 ();
 sg13g2_decap_8 FILLER_80_283 ();
 sg13g2_decap_4 FILLER_80_290 ();
 sg13g2_fill_2 FILLER_80_294 ();
 sg13g2_decap_4 FILLER_80_300 ();
 sg13g2_decap_8 FILLER_80_308 ();
 sg13g2_decap_4 FILLER_80_315 ();
 sg13g2_fill_1 FILLER_80_319 ();
 sg13g2_decap_8 FILLER_80_325 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_345 ();
 sg13g2_decap_8 FILLER_80_352 ();
 sg13g2_decap_8 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_366 ();
 sg13g2_decap_8 FILLER_80_376 ();
 sg13g2_decap_8 FILLER_80_383 ();
 sg13g2_decap_8 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_397 ();
 sg13g2_decap_4 FILLER_80_404 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net293;
 assign uio_oe[3] = net294;
 assign uio_oe[4] = net295;
 assign uio_oe[5] = net296;
 assign uio_oe[6] = net297;
 assign uio_oe[7] = net298;
 assign uio_out[0] = net8;
endmodule

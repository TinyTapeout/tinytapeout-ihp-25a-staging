module tt_um_tetrap_triggerer (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire DAT_OUT;
 wire DAT_RDY;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire clknet_0_clk;
 wire \trgg.cnt0.cnt[0] ;
 wire \trgg.cnt0.cnt[10] ;
 wire \trgg.cnt0.cnt[11] ;
 wire \trgg.cnt0.cnt[12] ;
 wire \trgg.cnt0.cnt[13] ;
 wire \trgg.cnt0.cnt[14] ;
 wire \trgg.cnt0.cnt[15] ;
 wire \trgg.cnt0.cnt[16] ;
 wire \trgg.cnt0.cnt[17] ;
 wire \trgg.cnt0.cnt[18] ;
 wire \trgg.cnt0.cnt[19] ;
 wire \trgg.cnt0.cnt[1] ;
 wire \trgg.cnt0.cnt[20] ;
 wire \trgg.cnt0.cnt[21] ;
 wire \trgg.cnt0.cnt[22] ;
 wire \trgg.cnt0.cnt[23] ;
 wire \trgg.cnt0.cnt[2] ;
 wire \trgg.cnt0.cnt[3] ;
 wire \trgg.cnt0.cnt[4] ;
 wire \trgg.cnt0.cnt[5] ;
 wire \trgg.cnt0.cnt[6] ;
 wire \trgg.cnt0.cnt[7] ;
 wire \trgg.cnt0.cnt[8] ;
 wire \trgg.cnt0.cnt[9] ;
 wire \trgg.is_timestamp_popped_from_q ;
 wire \trgg.shft.prev_dat_clk ;
 wire \trgg.shft.prev_ena ;
 wire \trgg.shft.tx_word[0] ;
 wire \trgg.shft.tx_word[10] ;
 wire \trgg.shft.tx_word[11] ;
 wire \trgg.shft.tx_word[12] ;
 wire \trgg.shft.tx_word[13] ;
 wire \trgg.shft.tx_word[14] ;
 wire \trgg.shft.tx_word[15] ;
 wire \trgg.shft.tx_word[16] ;
 wire \trgg.shft.tx_word[17] ;
 wire \trgg.shft.tx_word[18] ;
 wire \trgg.shft.tx_word[19] ;
 wire \trgg.shft.tx_word[1] ;
 wire \trgg.shft.tx_word[20] ;
 wire \trgg.shft.tx_word[21] ;
 wire \trgg.shft.tx_word[22] ;
 wire \trgg.shft.tx_word[2] ;
 wire \trgg.shft.tx_word[3] ;
 wire \trgg.shft.tx_word[4] ;
 wire \trgg.shft.tx_word[5] ;
 wire \trgg.shft.tx_word[6] ;
 wire \trgg.shft.tx_word[7] ;
 wire \trgg.shft.tx_word[8] ;
 wire \trgg.shft.tx_word[9] ;
 wire \trgg.shft.word_to_tx[0] ;
 wire \trgg.shft.word_to_tx[10] ;
 wire \trgg.shft.word_to_tx[11] ;
 wire \trgg.shft.word_to_tx[12] ;
 wire \trgg.shft.word_to_tx[13] ;
 wire \trgg.shft.word_to_tx[14] ;
 wire \trgg.shft.word_to_tx[15] ;
 wire \trgg.shft.word_to_tx[16] ;
 wire \trgg.shft.word_to_tx[17] ;
 wire \trgg.shft.word_to_tx[18] ;
 wire \trgg.shft.word_to_tx[19] ;
 wire \trgg.shft.word_to_tx[1] ;
 wire \trgg.shft.word_to_tx[20] ;
 wire \trgg.shft.word_to_tx[21] ;
 wire \trgg.shft.word_to_tx[22] ;
 wire \trgg.shft.word_to_tx[23] ;
 wire \trgg.shft.word_to_tx[2] ;
 wire \trgg.shft.word_to_tx[3] ;
 wire \trgg.shft.word_to_tx[4] ;
 wire \trgg.shft.word_to_tx[5] ;
 wire \trgg.shft.word_to_tx[6] ;
 wire \trgg.shft.word_to_tx[7] ;
 wire \trgg.shft.word_to_tx[8] ;
 wire \trgg.shft.word_to_tx[9] ;
 wire \trgg.trigg_channel.is_mem_full ;
 wire \trgg.trigg_channel.is_timestamp_present ;
 wire \trgg.trigg_channel.ltch.latched_time[0] ;
 wire \trgg.trigg_channel.ltch.latched_time[10] ;
 wire \trgg.trigg_channel.ltch.latched_time[11] ;
 wire \trgg.trigg_channel.ltch.latched_time[12] ;
 wire \trgg.trigg_channel.ltch.latched_time[13] ;
 wire \trgg.trigg_channel.ltch.latched_time[14] ;
 wire \trgg.trigg_channel.ltch.latched_time[15] ;
 wire \trgg.trigg_channel.ltch.latched_time[16] ;
 wire \trgg.trigg_channel.ltch.latched_time[17] ;
 wire \trgg.trigg_channel.ltch.latched_time[18] ;
 wire \trgg.trigg_channel.ltch.latched_time[19] ;
 wire \trgg.trigg_channel.ltch.latched_time[1] ;
 wire \trgg.trigg_channel.ltch.latched_time[20] ;
 wire \trgg.trigg_channel.ltch.latched_time[21] ;
 wire \trgg.trigg_channel.ltch.latched_time[22] ;
 wire \trgg.trigg_channel.ltch.latched_time[23] ;
 wire \trgg.trigg_channel.ltch.latched_time[2] ;
 wire \trgg.trigg_channel.ltch.latched_time[3] ;
 wire \trgg.trigg_channel.ltch.latched_time[4] ;
 wire \trgg.trigg_channel.ltch.latched_time[5] ;
 wire \trgg.trigg_channel.ltch.latched_time[6] ;
 wire \trgg.trigg_channel.ltch.latched_time[7] ;
 wire \trgg.trigg_channel.ltch.latched_time[8] ;
 wire \trgg.trigg_channel.ltch.latched_time[9] ;
 wire \trgg.trigg_channel.ltch.prev_trigger ;
 wire \trgg.trigg_channel.mem.mem_regs[1][0] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][10] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][11] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][12] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][13] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][14] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][15] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][16] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][17] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][18] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][19] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][1] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][20] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][21] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][22] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][23] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][2] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][3] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][4] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][5] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][6] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][7] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][8] ;
 wire \trgg.trigg_channel.mem.mem_regs[1][9] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][0] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][10] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][11] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][12] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][13] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][14] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][15] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][16] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][17] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][18] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][19] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][1] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][20] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][21] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][22] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][23] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][2] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][3] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][4] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][5] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][6] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][7] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][8] ;
 wire \trgg.trigg_channel.mem.mem_regs[2][9] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][0] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][10] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][11] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][12] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][13] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][14] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][15] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][16] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][17] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][18] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][19] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][1] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][20] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][21] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][22] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][23] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][2] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][3] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][4] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][5] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][6] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][7] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][8] ;
 wire \trgg.trigg_channel.mem.mem_regs[3][9] ;
 wire \trgg.trigg_channel.mem.shift_gen[0].mem.if_will_be_data ;
 wire \trgg.trigg_channel.mem.shift_gen[0].mem.is_in ;
 wire \trgg.trigg_channel.mem.shift_gen[1].mem.if_will_be_data ;
 wire \trgg.trigg_channel.mem.shift_gen[1].mem.is_in ;
 wire \trgg.trigg_channel.mem.shift_gen[2].mem.if_will_be_data ;
 wire \trgg.trigg_channel.mem.shift_gen[3].mem.if_will_be_data ;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;

 sg13g2_inv_1 _0618_ (.Y(_0170_),
    .A(\trgg.shft.prev_dat_clk ));
 sg13g2_inv_1 _0619_ (.Y(_0171_),
    .A(\trgg.shft.tx_word[0] ));
 sg13g2_inv_1 _0620_ (.Y(_0172_),
    .A(net4));
 sg13g2_inv_1 _0621_ (.Y(_0173_),
    .A(net447));
 sg13g2_inv_1 _0622_ (.Y(_0174_),
    .A(net437));
 sg13g2_inv_1 _0623_ (.Y(_0175_),
    .A(net282));
 sg13g2_inv_1 _0624_ (.Y(_0176_),
    .A(net411));
 sg13g2_inv_1 _0625_ (.Y(_0177_),
    .A(net469));
 sg13g2_inv_1 _0626_ (.Y(_0178_),
    .A(net455));
 sg13g2_nand2b_1 _0627_ (.Y(_0179_),
    .B(net3),
    .A_N(net471));
 sg13g2_inv_1 _0628_ (.Y(_0000_),
    .A(net157));
 sg13g2_nor2b_1 _0629_ (.A(net351),
    .B_N(\trgg.trigg_channel.is_mem_full ),
    .Y(_0180_));
 sg13g2_nor2b_1 _0630_ (.A(net366),
    .B_N(net398),
    .Y(_0181_));
 sg13g2_a21o_1 _0631_ (.A2(net351),
    .A1(net366),
    .B1(_0181_),
    .X(\trgg.trigg_channel.mem.shift_gen[3].mem.if_will_be_data ));
 sg13g2_nor2b_1 _0632_ (.A(net370),
    .B_N(net351),
    .Y(_0182_));
 sg13g2_a21o_1 _0633_ (.A2(net351),
    .A1(net370),
    .B1(net352),
    .X(\trgg.trigg_channel.mem.shift_gen[2].mem.if_will_be_data ));
 sg13g2_nor2b_1 _0634_ (.A(DAT_RDY),
    .B_N(\trgg.trigg_channel.mem.shift_gen[0].mem.is_in ),
    .Y(_0183_));
 sg13g2_a21o_1 _0635_ (.A2(net370),
    .A1(net466),
    .B1(_0182_),
    .X(\trgg.trigg_channel.mem.shift_gen[1].mem.if_will_be_data ));
 sg13g2_a21o_1 _0636_ (.A2(net219),
    .A1(DAT_RDY),
    .B1(_0183_),
    .X(\trgg.trigg_channel.mem.shift_gen[0].mem.if_will_be_data ));
 sg13g2_xor2_1 _0637_ (.B(net463),
    .A(net338),
    .X(_0011_));
 sg13g2_nand3_1 _0638_ (.B(\trgg.cnt0.cnt[1] ),
    .C(net257),
    .A(\trgg.cnt0.cnt[0] ),
    .Y(_0184_));
 sg13g2_a21o_1 _0639_ (.A2(net463),
    .A1(net338),
    .B1(net257),
    .X(_0185_));
 sg13g2_and2_1 _0640_ (.A(net258),
    .B(_0185_),
    .X(_0016_));
 sg13g2_nand4_1 _0641_ (.B(\trgg.cnt0.cnt[1] ),
    .C(\trgg.cnt0.cnt[2] ),
    .A(\trgg.cnt0.cnt[0] ),
    .Y(_0186_),
    .D(\trgg.cnt0.cnt[3] ));
 sg13g2_xnor2_1 _0642_ (.Y(_0017_),
    .A(net234),
    .B(net258));
 sg13g2_xnor2_1 _0643_ (.Y(_0018_),
    .A(net447),
    .B(_0186_));
 sg13g2_nor3_2 _0644_ (.A(_0173_),
    .B(_0174_),
    .C(_0186_),
    .Y(_0187_));
 sg13g2_o21ai_1 _0645_ (.B1(_0174_),
    .Y(_0188_),
    .A1(_0173_),
    .A2(_0186_));
 sg13g2_nor2b_1 _0646_ (.A(_0187_),
    .B_N(_0188_),
    .Y(_0019_));
 sg13g2_xor2_1 _0647_ (.B(_0187_),
    .A(net317),
    .X(_0020_));
 sg13g2_nand4_1 _0648_ (.B(net437),
    .C(\trgg.cnt0.cnt[6] ),
    .A(net468),
    .Y(_0189_),
    .D(net345));
 sg13g2_nor2_2 _0649_ (.A(_0186_),
    .B(_0189_),
    .Y(_0190_));
 sg13g2_a21oi_1 _0650_ (.A1(net317),
    .A2(_0187_),
    .Y(_0191_),
    .B1(net345));
 sg13g2_nor2_1 _0651_ (.A(_0190_),
    .B(net346),
    .Y(_0021_));
 sg13g2_xor2_1 _0652_ (.B(_0190_),
    .A(net233),
    .X(_0022_));
 sg13g2_a21oi_1 _0653_ (.A1(net233),
    .A2(_0190_),
    .Y(_0192_),
    .B1(net261));
 sg13g2_nand3_1 _0654_ (.B(net261),
    .C(_0190_),
    .A(net233),
    .Y(_0193_));
 sg13g2_nor2b_1 _0655_ (.A(_0192_),
    .B_N(_0193_),
    .Y(_0023_));
 sg13g2_nand4_1 _0656_ (.B(net261),
    .C(net268),
    .A(net233),
    .Y(_0194_),
    .D(_0190_));
 sg13g2_xnor2_1 _0657_ (.Y(_0001_),
    .A(net268),
    .B(_0193_));
 sg13g2_nand4_1 _0658_ (.B(net261),
    .C(net268),
    .A(net438),
    .Y(_0195_),
    .D(net282));
 sg13g2_nor3_2 _0659_ (.A(_0186_),
    .B(_0189_),
    .C(_0195_),
    .Y(_0196_));
 sg13g2_a21oi_1 _0660_ (.A1(_0175_),
    .A2(_0194_),
    .Y(_0002_),
    .B1(_0196_));
 sg13g2_xor2_1 _0661_ (.B(_0196_),
    .A(net464),
    .X(_0003_));
 sg13g2_a21oi_1 _0662_ (.A1(net464),
    .A2(_0196_),
    .Y(_0197_),
    .B1(net228));
 sg13g2_nand3_1 _0663_ (.B(net228),
    .C(_0196_),
    .A(net464),
    .Y(_0198_));
 sg13g2_nor2b_1 _0664_ (.A(_0197_),
    .B_N(_0198_),
    .Y(_0004_));
 sg13g2_nand4_1 _0665_ (.B(net228),
    .C(net409),
    .A(\trgg.cnt0.cnt[12] ),
    .Y(_0199_),
    .D(_0196_));
 sg13g2_xnor2_1 _0666_ (.Y(_0005_),
    .A(net409),
    .B(_0198_));
 sg13g2_nand4_1 _0667_ (.B(net228),
    .C(net409),
    .A(net464),
    .Y(_0200_),
    .D(net411));
 sg13g2_nor4_2 _0668_ (.A(_0186_),
    .B(_0189_),
    .C(_0195_),
    .Y(_0201_),
    .D(_0200_));
 sg13g2_a21oi_1 _0669_ (.A1(_0176_),
    .A2(_0199_),
    .Y(_0006_),
    .B1(_0201_));
 sg13g2_xor2_1 _0670_ (.B(net149),
    .A(net460),
    .X(_0007_));
 sg13g2_a21oi_1 _0671_ (.A1(\trgg.cnt0.cnt[16] ),
    .A2(net149),
    .Y(_0202_),
    .B1(net457));
 sg13g2_nand3_1 _0672_ (.B(net457),
    .C(net149),
    .A(net460),
    .Y(_0203_));
 sg13g2_nor2b_1 _0673_ (.A(net458),
    .B_N(_0203_),
    .Y(_0008_));
 sg13g2_nand4_1 _0674_ (.B(net457),
    .C(net283),
    .A(net460),
    .Y(_0204_),
    .D(net149));
 sg13g2_xnor2_1 _0675_ (.Y(_0009_),
    .A(net283),
    .B(_0203_));
 sg13g2_and4_2 _0676_ (.A(\trgg.cnt0.cnt[16] ),
    .B(net457),
    .C(net283),
    .D(net469),
    .X(_0205_));
 sg13g2_a22oi_1 _0677_ (.Y(_0010_),
    .B1(_0205_),
    .B2(_0201_),
    .A2(_0204_),
    .A1(_0177_));
 sg13g2_a21oi_1 _0678_ (.A1(net149),
    .A2(_0205_),
    .Y(_0206_),
    .B1(net421));
 sg13g2_nand3_1 _0679_ (.B(net149),
    .C(_0205_),
    .A(net421),
    .Y(_0207_));
 sg13g2_nor2b_1 _0680_ (.A(net422),
    .B_N(_0207_),
    .Y(_0012_));
 sg13g2_and2_1 _0681_ (.A(\trgg.cnt0.cnt[20] ),
    .B(net455),
    .X(_0208_));
 sg13g2_and3_1 _0682_ (.X(_0209_),
    .A(net149),
    .B(_0205_),
    .C(_0208_));
 sg13g2_a21oi_1 _0683_ (.A1(_0178_),
    .A2(_0207_),
    .Y(_0013_),
    .B1(_0209_));
 sg13g2_nand4_1 _0684_ (.B(net149),
    .C(_0205_),
    .A(net225),
    .Y(_0210_),
    .D(_0208_));
 sg13g2_xor2_1 _0685_ (.B(_0209_),
    .A(net225),
    .X(_0014_));
 sg13g2_xnor2_1 _0686_ (.Y(_0015_),
    .A(net237),
    .B(_0210_));
 sg13g2_o21ai_1 _0687_ (.B1(net157),
    .Y(_0211_),
    .A1(_0170_),
    .A2(net2));
 sg13g2_nand2_1 _0688_ (.Y(_0212_),
    .A(net269),
    .B(_0000_));
 sg13g2_o21ai_1 _0689_ (.B1(_0212_),
    .Y(_0120_),
    .A1(_0171_),
    .A2(net147));
 sg13g2_nor2_1 _0690_ (.A(\trgg.shft.tx_word[1] ),
    .B(net148),
    .Y(_0213_));
 sg13g2_nor2_1 _0691_ (.A(\trgg.shft.word_to_tx[1] ),
    .B(net158),
    .Y(_0214_));
 sg13g2_nand3b_1 _0692_ (.B(net157),
    .C(\trgg.shft.prev_dat_clk ),
    .Y(_0215_),
    .A_N(net2));
 sg13g2_nor2_1 _0693_ (.A(net406),
    .B(net143),
    .Y(_0216_));
 sg13g2_nor3_1 _0694_ (.A(_0213_),
    .B(_0214_),
    .C(_0216_),
    .Y(_0121_));
 sg13g2_nor2_1 _0695_ (.A(net419),
    .B(net148),
    .Y(_0217_));
 sg13g2_nor2_1 _0696_ (.A(net439),
    .B(net158),
    .Y(_0218_));
 sg13g2_nor2_1 _0697_ (.A(net443),
    .B(net143),
    .Y(_0219_));
 sg13g2_nor3_1 _0698_ (.A(_0217_),
    .B(_0218_),
    .C(_0219_),
    .Y(_0122_));
 sg13g2_nor2_1 _0699_ (.A(net419),
    .B(net144),
    .Y(_0220_));
 sg13g2_nor2_1 _0700_ (.A(\trgg.shft.tx_word[3] ),
    .B(net147),
    .Y(_0221_));
 sg13g2_nor2_1 _0701_ (.A(\trgg.shft.word_to_tx[3] ),
    .B(net157),
    .Y(_0222_));
 sg13g2_nor3_1 _0702_ (.A(_0220_),
    .B(_0221_),
    .C(_0222_),
    .Y(_0123_));
 sg13g2_nor2_1 _0703_ (.A(net399),
    .B(net146),
    .Y(_0223_));
 sg13g2_nor2_1 _0704_ (.A(net408),
    .B(net156),
    .Y(_0224_));
 sg13g2_nor2_1 _0705_ (.A(net467),
    .B(net143),
    .Y(_0225_));
 sg13g2_nor3_1 _0706_ (.A(_0223_),
    .B(_0224_),
    .C(_0225_),
    .Y(_0124_));
 sg13g2_nor2_1 _0707_ (.A(net399),
    .B(net142),
    .Y(_0226_));
 sg13g2_nor2_1 _0708_ (.A(\trgg.shft.tx_word[5] ),
    .B(net146),
    .Y(_0227_));
 sg13g2_nor2_1 _0709_ (.A(\trgg.shft.word_to_tx[5] ),
    .B(net156),
    .Y(_0228_));
 sg13g2_nor3_1 _0710_ (.A(_0226_),
    .B(_0227_),
    .C(_0228_),
    .Y(_0125_));
 sg13g2_nor2_1 _0711_ (.A(\trgg.shft.tx_word[5] ),
    .B(net142),
    .Y(_0229_));
 sg13g2_nor2_1 _0712_ (.A(\trgg.shft.tx_word[6] ),
    .B(net145),
    .Y(_0230_));
 sg13g2_nor2_1 _0713_ (.A(net333),
    .B(net156),
    .Y(_0231_));
 sg13g2_nor3_1 _0714_ (.A(_0229_),
    .B(_0230_),
    .C(_0231_),
    .Y(_0126_));
 sg13g2_nor2_1 _0715_ (.A(\trgg.shft.tx_word[7] ),
    .B(net146),
    .Y(_0232_));
 sg13g2_nor2_1 _0716_ (.A(net404),
    .B(net155),
    .Y(_0233_));
 sg13g2_nor2_1 _0717_ (.A(\trgg.shft.tx_word[6] ),
    .B(net142),
    .Y(_0234_));
 sg13g2_nor3_1 _0718_ (.A(_0232_),
    .B(_0233_),
    .C(_0234_),
    .Y(_0127_));
 sg13g2_nor2_1 _0719_ (.A(\trgg.shft.tx_word[7] ),
    .B(net141),
    .Y(_0235_));
 sg13g2_nor2_1 _0720_ (.A(\trgg.shft.tx_word[8] ),
    .B(net145),
    .Y(_0236_));
 sg13g2_nor2_1 _0721_ (.A(net388),
    .B(net155),
    .Y(_0237_));
 sg13g2_nor3_1 _0722_ (.A(_0235_),
    .B(_0236_),
    .C(_0237_),
    .Y(_0128_));
 sg13g2_nor2_1 _0723_ (.A(net453),
    .B(net145),
    .Y(_0238_));
 sg13g2_nor2_1 _0724_ (.A(\trgg.shft.word_to_tx[9] ),
    .B(net155),
    .Y(_0239_));
 sg13g2_nor2_1 _0725_ (.A(\trgg.shft.tx_word[8] ),
    .B(net141),
    .Y(_0240_));
 sg13g2_nor3_1 _0726_ (.A(_0238_),
    .B(_0239_),
    .C(_0240_),
    .Y(_0129_));
 sg13g2_nor2_1 _0727_ (.A(\trgg.shft.tx_word[9] ),
    .B(net141),
    .Y(_0241_));
 sg13g2_nor2_1 _0728_ (.A(\trgg.shft.tx_word[10] ),
    .B(net145),
    .Y(_0242_));
 sg13g2_nor2_1 _0729_ (.A(net445),
    .B(net155),
    .Y(_0243_));
 sg13g2_nor3_1 _0730_ (.A(_0241_),
    .B(_0242_),
    .C(_0243_),
    .Y(_0130_));
 sg13g2_nor2_1 _0731_ (.A(\trgg.shft.tx_word[10] ),
    .B(net141),
    .Y(_0244_));
 sg13g2_nor2_1 _0732_ (.A(\trgg.shft.tx_word[11] ),
    .B(net145),
    .Y(_0245_));
 sg13g2_nor2_1 _0733_ (.A(net449),
    .B(net155),
    .Y(_0246_));
 sg13g2_nor3_1 _0734_ (.A(_0244_),
    .B(_0245_),
    .C(_0246_),
    .Y(_0131_));
 sg13g2_nor2_1 _0735_ (.A(net386),
    .B(net145),
    .Y(_0247_));
 sg13g2_nor2_1 _0736_ (.A(\trgg.shft.word_to_tx[12] ),
    .B(net155),
    .Y(_0248_));
 sg13g2_nor2_1 _0737_ (.A(\trgg.shft.tx_word[11] ),
    .B(net141),
    .Y(_0249_));
 sg13g2_nor3_1 _0738_ (.A(_0247_),
    .B(_0248_),
    .C(_0249_),
    .Y(_0132_));
 sg13g2_nor2_1 _0739_ (.A(net386),
    .B(net141),
    .Y(_0250_));
 sg13g2_nor2_1 _0740_ (.A(net384),
    .B(net145),
    .Y(_0251_));
 sg13g2_nor2_1 _0741_ (.A(net417),
    .B(net155),
    .Y(_0252_));
 sg13g2_nor3_1 _0742_ (.A(_0250_),
    .B(_0251_),
    .C(_0252_),
    .Y(_0133_));
 sg13g2_nor2_1 _0743_ (.A(net384),
    .B(net141),
    .Y(_0253_));
 sg13g2_nor2_1 _0744_ (.A(net378),
    .B(net146),
    .Y(_0254_));
 sg13g2_nor2_1 _0745_ (.A(\trgg.shft.word_to_tx[14] ),
    .B(net156),
    .Y(_0255_));
 sg13g2_nor3_1 _0746_ (.A(_0253_),
    .B(_0254_),
    .C(_0255_),
    .Y(_0134_));
 sg13g2_nor2_1 _0747_ (.A(\trgg.shft.tx_word[15] ),
    .B(net145),
    .Y(_0256_));
 sg13g2_nor2_1 _0748_ (.A(\trgg.shft.word_to_tx[15] ),
    .B(net155),
    .Y(_0257_));
 sg13g2_nor2_1 _0749_ (.A(net378),
    .B(net141),
    .Y(_0258_));
 sg13g2_nor3_1 _0750_ (.A(_0256_),
    .B(_0257_),
    .C(_0258_),
    .Y(_0135_));
 sg13g2_nor2_1 _0751_ (.A(\trgg.shft.tx_word[16] ),
    .B(net146),
    .Y(_0259_));
 sg13g2_nor2_1 _0752_ (.A(net336),
    .B(net156),
    .Y(_0260_));
 sg13g2_nor2_1 _0753_ (.A(\trgg.shft.tx_word[15] ),
    .B(net142),
    .Y(_0261_));
 sg13g2_nor3_1 _0754_ (.A(_0259_),
    .B(_0260_),
    .C(_0261_),
    .Y(_0136_));
 sg13g2_nor2_1 _0755_ (.A(\trgg.shft.tx_word[17] ),
    .B(net146),
    .Y(_0262_));
 sg13g2_nor2_1 _0756_ (.A(net326),
    .B(net156),
    .Y(_0263_));
 sg13g2_nor2_1 _0757_ (.A(\trgg.shft.tx_word[16] ),
    .B(net142),
    .Y(_0264_));
 sg13g2_nor3_1 _0758_ (.A(_0262_),
    .B(_0263_),
    .C(_0264_),
    .Y(_0137_));
 sg13g2_nor2_1 _0759_ (.A(net429),
    .B(net147),
    .Y(_0265_));
 sg13g2_nor2_1 _0760_ (.A(net435),
    .B(net157),
    .Y(_0266_));
 sg13g2_nor2_1 _0761_ (.A(\trgg.shft.tx_word[17] ),
    .B(net143),
    .Y(_0267_));
 sg13g2_nor3_1 _0762_ (.A(_0265_),
    .B(_0266_),
    .C(_0267_),
    .Y(_0138_));
 sg13g2_nor2_1 _0763_ (.A(net429),
    .B(net143),
    .Y(_0268_));
 sg13g2_nor2_1 _0764_ (.A(net425),
    .B(net147),
    .Y(_0269_));
 sg13g2_nor2_1 _0765_ (.A(\trgg.shft.word_to_tx[19] ),
    .B(net157),
    .Y(_0270_));
 sg13g2_nor3_1 _0766_ (.A(_0268_),
    .B(_0269_),
    .C(_0270_),
    .Y(_0139_));
 sg13g2_nor2_1 _0767_ (.A(\trgg.shft.tx_word[20] ),
    .B(net147),
    .Y(_0271_));
 sg13g2_nor2_1 _0768_ (.A(\trgg.shft.word_to_tx[20] ),
    .B(net157),
    .Y(_0272_));
 sg13g2_nor2_1 _0769_ (.A(net425),
    .B(net143),
    .Y(_0273_));
 sg13g2_nor3_1 _0770_ (.A(_0271_),
    .B(_0272_),
    .C(_0273_),
    .Y(_0140_));
 sg13g2_nor2_1 _0771_ (.A(\trgg.shft.tx_word[20] ),
    .B(net144),
    .Y(_0274_));
 sg13g2_nor2_1 _0772_ (.A(\trgg.shft.tx_word[21] ),
    .B(net147),
    .Y(_0275_));
 sg13g2_nor2_1 _0773_ (.A(net427),
    .B(net158),
    .Y(_0276_));
 sg13g2_nor3_1 _0774_ (.A(_0274_),
    .B(_0275_),
    .C(_0276_),
    .Y(_0141_));
 sg13g2_nor2_1 _0775_ (.A(\trgg.shft.tx_word[21] ),
    .B(net143),
    .Y(_0277_));
 sg13g2_nor2_1 _0776_ (.A(\trgg.shft.tx_word[22] ),
    .B(net147),
    .Y(_0278_));
 sg13g2_nor2_1 _0777_ (.A(net415),
    .B(net157),
    .Y(_0279_));
 sg13g2_nor3_1 _0778_ (.A(_0277_),
    .B(_0278_),
    .C(_0279_),
    .Y(_0142_));
 sg13g2_nor2_1 _0779_ (.A(DAT_OUT),
    .B(net147),
    .Y(_0280_));
 sg13g2_nor2_1 _0780_ (.A(\trgg.shft.word_to_tx[23] ),
    .B(net158),
    .Y(_0281_));
 sg13g2_nor2_1 _0781_ (.A(net423),
    .B(net143),
    .Y(_0282_));
 sg13g2_nor3_1 _0782_ (.A(_0280_),
    .B(_0281_),
    .C(_0282_),
    .Y(_0143_));
 sg13g2_nand2_1 _0783_ (.Y(_0283_),
    .A(net1),
    .B(_0181_));
 sg13g2_mux2_1 _0784_ (.A0(net319),
    .A1(\trgg.trigg_channel.mem.mem_regs[3][0] ),
    .S(net139),
    .X(_0144_));
 sg13g2_mux2_1 _0785_ (.A0(net264),
    .A1(net290),
    .S(net138),
    .X(_0145_));
 sg13g2_mux2_1 _0786_ (.A0(net279),
    .A1(net300),
    .S(net138),
    .X(_0146_));
 sg13g2_mux2_1 _0787_ (.A0(net229),
    .A1(\trgg.trigg_channel.mem.mem_regs[3][3] ),
    .S(net139),
    .X(_0147_));
 sg13g2_mux2_1 _0788_ (.A0(net339),
    .A1(net354),
    .S(net137),
    .X(_0148_));
 sg13g2_mux2_1 _0789_ (.A0(net274),
    .A1(net293),
    .S(net137),
    .X(_0149_));
 sg13g2_mux2_1 _0790_ (.A0(net277),
    .A1(net297),
    .S(net137),
    .X(_0150_));
 sg13g2_mux2_1 _0791_ (.A0(net252),
    .A1(net276),
    .S(net136),
    .X(_0151_));
 sg13g2_mux2_1 _0792_ (.A0(net221),
    .A1(\trgg.trigg_channel.mem.mem_regs[3][8] ),
    .S(net136),
    .X(_0152_));
 sg13g2_mux2_1 _0793_ (.A0(net223),
    .A1(\trgg.trigg_channel.mem.mem_regs[3][9] ),
    .S(net136),
    .X(_0153_));
 sg13g2_mux2_1 _0794_ (.A0(net243),
    .A1(\trgg.trigg_channel.mem.mem_regs[3][10] ),
    .S(net136),
    .X(_0154_));
 sg13g2_mux2_1 _0795_ (.A0(net231),
    .A1(\trgg.trigg_channel.mem.mem_regs[3][11] ),
    .S(net136),
    .X(_0155_));
 sg13g2_mux2_1 _0796_ (.A0(net241),
    .A1(net254),
    .S(net136),
    .X(_0156_));
 sg13g2_mux2_1 _0797_ (.A0(net226),
    .A1(\trgg.trigg_channel.mem.mem_regs[3][13] ),
    .S(net136),
    .X(_0157_));
 sg13g2_mux2_1 _0798_ (.A0(net245),
    .A1(net284),
    .S(net136),
    .X(_0158_));
 sg13g2_mux2_1 _0799_ (.A0(net262),
    .A1(net358),
    .S(net137),
    .X(_0159_));
 sg13g2_mux2_1 _0800_ (.A0(net239),
    .A1(net247),
    .S(net138),
    .X(_0160_));
 sg13g2_mux2_1 _0801_ (.A0(net255),
    .A1(net273),
    .S(net138),
    .X(_0161_));
 sg13g2_mux2_1 _0802_ (.A0(net271),
    .A1(\trgg.trigg_channel.mem.mem_regs[3][18] ),
    .S(net138),
    .X(_0162_));
 sg13g2_mux2_1 _0803_ (.A0(net235),
    .A1(net325),
    .S(net138),
    .X(_0163_));
 sg13g2_mux2_1 _0804_ (.A0(net250),
    .A1(net267),
    .S(net139),
    .X(_0164_));
 sg13g2_mux2_1 _0805_ (.A0(net259),
    .A1(net359),
    .S(net139),
    .X(_0165_));
 sg13g2_mux2_1 _0806_ (.A0(net248),
    .A1(\trgg.trigg_channel.mem.mem_regs[3][22] ),
    .S(net138),
    .X(_0166_));
 sg13g2_mux2_1 _0807_ (.A0(net266),
    .A1(net285),
    .S(net138),
    .X(_0167_));
 sg13g2_nor3_1 _0808_ (.A(\trgg.trigg_channel.is_timestamp_present ),
    .B(_0172_),
    .C(net280),
    .Y(_0284_));
 sg13g2_a21o_1 _0809_ (.A2(net366),
    .A1(net398),
    .B1(net154),
    .X(_0168_));
 sg13g2_nand2_1 _0810_ (.Y(_0285_),
    .A(net1),
    .B(_0180_));
 sg13g2_mux2_1 _0811_ (.A0(net362),
    .A1(\trgg.trigg_channel.mem.mem_regs[2][0] ),
    .S(net134),
    .X(_0169_));
 sg13g2_mux2_1 _0812_ (.A0(net290),
    .A1(net307),
    .S(net134),
    .X(_0025_));
 sg13g2_mux2_1 _0813_ (.A0(net300),
    .A1(net402),
    .S(net133),
    .X(_0026_));
 sg13g2_mux2_1 _0814_ (.A0(net348),
    .A1(net341),
    .S(net134),
    .X(_0027_));
 sg13g2_mux2_1 _0815_ (.A0(net354),
    .A1(\trgg.trigg_channel.mem.mem_regs[2][4] ),
    .S(net132),
    .X(_0028_));
 sg13g2_mux2_1 _0816_ (.A0(net293),
    .A1(net321),
    .S(net132),
    .X(_0029_));
 sg13g2_mux2_1 _0817_ (.A0(net297),
    .A1(net309),
    .S(net132),
    .X(_0030_));
 sg13g2_mux2_1 _0818_ (.A0(net276),
    .A1(net294),
    .S(net131),
    .X(_0031_));
 sg13g2_mux2_1 _0819_ (.A0(net397),
    .A1(net286),
    .S(net131),
    .X(_0032_));
 sg13g2_mux2_1 _0820_ (.A0(net393),
    .A1(net288),
    .S(net131),
    .X(_0033_));
 sg13g2_mux2_1 _0821_ (.A0(net418),
    .A1(net377),
    .S(net131),
    .X(_0034_));
 sg13g2_mux2_1 _0822_ (.A0(net401),
    .A1(net298),
    .S(net131),
    .X(_0035_));
 sg13g2_mux2_1 _0823_ (.A0(net254),
    .A1(net368),
    .S(net131),
    .X(_0036_));
 sg13g2_mux2_1 _0824_ (.A0(net394),
    .A1(net390),
    .S(net131),
    .X(_0037_));
 sg13g2_mux2_1 _0825_ (.A0(net284),
    .A1(net367),
    .S(net131),
    .X(_0038_));
 sg13g2_mux2_1 _0826_ (.A0(net358),
    .A1(net313),
    .S(net132),
    .X(_0039_));
 sg13g2_mux2_1 _0827_ (.A0(net247),
    .A1(net343),
    .S(net133),
    .X(_0040_));
 sg13g2_mux2_1 _0828_ (.A0(net273),
    .A1(net335),
    .S(net133),
    .X(_0041_));
 sg13g2_mux2_1 _0829_ (.A0(net303),
    .A1(\trgg.trigg_channel.mem.mem_regs[2][18] ),
    .S(net133),
    .X(_0042_));
 sg13g2_mux2_1 _0830_ (.A0(net325),
    .A1(net356),
    .S(net133),
    .X(_0043_));
 sg13g2_mux2_1 _0831_ (.A0(net267),
    .A1(net291),
    .S(net134),
    .X(_0044_));
 sg13g2_mux2_1 _0832_ (.A0(net359),
    .A1(net330),
    .S(net133),
    .X(_0045_));
 sg13g2_mux2_1 _0833_ (.A0(net392),
    .A1(net331),
    .S(net133),
    .X(_0046_));
 sg13g2_mux2_1 _0834_ (.A0(net285),
    .A1(net305),
    .S(net133),
    .X(_0047_));
 sg13g2_nand2_1 _0835_ (.Y(_0286_),
    .A(net1),
    .B(_0182_));
 sg13g2_mux2_1 _0836_ (.A0(net431),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][0] ),
    .S(net129),
    .X(_0048_));
 sg13g2_mux2_1 _0837_ (.A0(net307),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][1] ),
    .S(net129),
    .X(_0049_));
 sg13g2_mux2_1 _0838_ (.A0(net402),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][2] ),
    .S(net129),
    .X(_0050_));
 sg13g2_mux2_1 _0839_ (.A0(net341),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][3] ),
    .S(net128),
    .X(_0051_));
 sg13g2_mux2_1 _0840_ (.A0(\trgg.trigg_channel.mem.mem_regs[2][4] ),
    .A1(net380),
    .S(net128),
    .X(_0052_));
 sg13g2_mux2_1 _0841_ (.A0(net321),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][5] ),
    .S(net127),
    .X(_0053_));
 sg13g2_mux2_1 _0842_ (.A0(net309),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][6] ),
    .S(net127),
    .X(_0054_));
 sg13g2_mux2_1 _0843_ (.A0(net294),
    .A1(net349),
    .S(net127),
    .X(_0055_));
 sg13g2_mux2_1 _0844_ (.A0(net286),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][8] ),
    .S(net126),
    .X(_0056_));
 sg13g2_mux2_1 _0845_ (.A0(net288),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][9] ),
    .S(net126),
    .X(_0057_));
 sg13g2_mux2_1 _0846_ (.A0(net377),
    .A1(net360),
    .S(net126),
    .X(_0058_));
 sg13g2_mux2_1 _0847_ (.A0(net298),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][11] ),
    .S(net126),
    .X(_0059_));
 sg13g2_mux2_1 _0848_ (.A0(net368),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][12] ),
    .S(net126),
    .X(_0060_));
 sg13g2_mux2_1 _0849_ (.A0(net390),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][13] ),
    .S(net126),
    .X(_0061_));
 sg13g2_mux2_1 _0850_ (.A0(net367),
    .A1(net311),
    .S(net126),
    .X(_0062_));
 sg13g2_mux2_1 _0851_ (.A0(net313),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][15] ),
    .S(net127),
    .X(_0063_));
 sg13g2_mux2_1 _0852_ (.A0(net343),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][16] ),
    .S(net126),
    .X(_0064_));
 sg13g2_mux2_1 _0853_ (.A0(net335),
    .A1(net374),
    .S(net128),
    .X(_0065_));
 sg13g2_mux2_1 _0854_ (.A0(net353),
    .A1(net295),
    .S(net128),
    .X(_0066_));
 sg13g2_mux2_1 _0855_ (.A0(net356),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][19] ),
    .S(net128),
    .X(_0067_));
 sg13g2_mux2_1 _0856_ (.A0(net291),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][20] ),
    .S(net129),
    .X(_0068_));
 sg13g2_mux2_1 _0857_ (.A0(net330),
    .A1(net301),
    .S(net128),
    .X(_0069_));
 sg13g2_mux2_1 _0858_ (.A0(net331),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][22] ),
    .S(net128),
    .X(_0070_));
 sg13g2_mux2_1 _0859_ (.A0(net305),
    .A1(\trgg.trigg_channel.mem.mem_regs[1][23] ),
    .S(net128),
    .X(_0071_));
 sg13g2_nand2_1 _0860_ (.Y(_0287_),
    .A(net162),
    .B(_0183_));
 sg13g2_mux2_1 _0861_ (.A0(net444),
    .A1(net269),
    .S(net124),
    .X(_0072_));
 sg13g2_mux2_1 _0862_ (.A0(net461),
    .A1(\trgg.shft.word_to_tx[1] ),
    .S(net124),
    .X(_0073_));
 sg13g2_mux2_1 _0863_ (.A0(\trgg.trigg_channel.mem.mem_regs[1][2] ),
    .A1(net439),
    .S(net124),
    .X(_0074_));
 sg13g2_mux2_1 _0864_ (.A0(net364),
    .A1(\trgg.shft.word_to_tx[3] ),
    .S(net123),
    .X(_0075_));
 sg13g2_mux2_1 _0865_ (.A0(net380),
    .A1(net408),
    .S(net123),
    .X(_0076_));
 sg13g2_mux2_1 _0866_ (.A0(net413),
    .A1(\trgg.shft.word_to_tx[5] ),
    .S(net122),
    .X(_0077_));
 sg13g2_mux2_1 _0867_ (.A0(net328),
    .A1(\trgg.shft.word_to_tx[6] ),
    .S(net122),
    .X(_0078_));
 sg13g2_mux2_1 _0868_ (.A0(net349),
    .A1(\trgg.shft.word_to_tx[7] ),
    .S(net121),
    .X(_0079_));
 sg13g2_mux2_1 _0869_ (.A0(net375),
    .A1(\trgg.shft.word_to_tx[8] ),
    .S(net121),
    .X(_0080_));
 sg13g2_mux2_1 _0870_ (.A0(net433),
    .A1(\trgg.shft.word_to_tx[9] ),
    .S(net121),
    .X(_0081_));
 sg13g2_mux2_1 _0871_ (.A0(net360),
    .A1(\trgg.shft.word_to_tx[10] ),
    .S(net121),
    .X(_0082_));
 sg13g2_mux2_1 _0872_ (.A0(net323),
    .A1(\trgg.shft.word_to_tx[11] ),
    .S(net121),
    .X(_0083_));
 sg13g2_mux2_1 _0873_ (.A0(net382),
    .A1(\trgg.shft.word_to_tx[12] ),
    .S(net121),
    .X(_0084_));
 sg13g2_mux2_1 _0874_ (.A0(net395),
    .A1(\trgg.shft.word_to_tx[13] ),
    .S(net121),
    .X(_0085_));
 sg13g2_mux2_1 _0875_ (.A0(net311),
    .A1(\trgg.shft.word_to_tx[14] ),
    .S(net121),
    .X(_0086_));
 sg13g2_mux2_1 _0876_ (.A0(net315),
    .A1(\trgg.shft.word_to_tx[15] ),
    .S(net122),
    .X(_0087_));
 sg13g2_mux2_1 _0877_ (.A0(net373),
    .A1(net336),
    .S(net122),
    .X(_0088_));
 sg13g2_mux2_1 _0878_ (.A0(net374),
    .A1(net326),
    .S(net123),
    .X(_0089_));
 sg13g2_mux2_1 _0879_ (.A0(net295),
    .A1(\trgg.shft.word_to_tx[18] ),
    .S(net123),
    .X(_0090_));
 sg13g2_mux2_1 _0880_ (.A0(net371),
    .A1(\trgg.shft.word_to_tx[19] ),
    .S(net123),
    .X(_0091_));
 sg13g2_mux2_1 _0881_ (.A0(\trgg.trigg_channel.mem.mem_regs[1][20] ),
    .A1(net451),
    .S(net124),
    .X(_0092_));
 sg13g2_mux2_1 _0882_ (.A0(net301),
    .A1(\trgg.shft.word_to_tx[21] ),
    .S(net123),
    .X(_0093_));
 sg13g2_mux2_1 _0883_ (.A0(net465),
    .A1(net415),
    .S(net123),
    .X(_0094_));
 sg13g2_mux2_1 _0884_ (.A0(net441),
    .A1(\trgg.shft.word_to_tx[23] ),
    .S(net123),
    .X(_0095_));
 sg13g2_mux2_1 _0885_ (.A0(net319),
    .A1(net338),
    .S(net153),
    .X(_0096_));
 sg13g2_mux2_1 _0886_ (.A0(net264),
    .A1(\trgg.cnt0.cnt[1] ),
    .S(net153),
    .X(_0097_));
 sg13g2_mux2_1 _0887_ (.A0(net279),
    .A1(net257),
    .S(net153),
    .X(_0098_));
 sg13g2_mux2_1 _0888_ (.A0(net229),
    .A1(net234),
    .S(net153),
    .X(_0099_));
 sg13g2_nor2_1 _0889_ (.A(net339),
    .B(net151),
    .Y(_0288_));
 sg13g2_a21oi_1 _0890_ (.A1(_0173_),
    .A2(net151),
    .Y(_0100_),
    .B1(_0288_));
 sg13g2_nor2_1 _0891_ (.A(net274),
    .B(net151),
    .Y(_0289_));
 sg13g2_a21oi_1 _0892_ (.A1(_0174_),
    .A2(net151),
    .Y(_0101_),
    .B1(_0289_));
 sg13g2_mux2_1 _0893_ (.A0(net277),
    .A1(\trgg.cnt0.cnt[6] ),
    .S(net151),
    .X(_0102_));
 sg13g2_mux2_1 _0894_ (.A0(net252),
    .A1(\trgg.cnt0.cnt[7] ),
    .S(net154),
    .X(_0103_));
 sg13g2_mux2_1 _0895_ (.A0(net221),
    .A1(net233),
    .S(net150),
    .X(_0104_));
 sg13g2_mux2_1 _0896_ (.A0(net223),
    .A1(net261),
    .S(net150),
    .X(_0105_));
 sg13g2_mux2_1 _0897_ (.A0(net243),
    .A1(net268),
    .S(net150),
    .X(_0106_));
 sg13g2_mux2_1 _0898_ (.A0(net231),
    .A1(net282),
    .S(net150),
    .X(_0107_));
 sg13g2_mux2_1 _0899_ (.A0(net241),
    .A1(\trgg.cnt0.cnt[12] ),
    .S(net150),
    .X(_0108_));
 sg13g2_mux2_1 _0900_ (.A0(net226),
    .A1(net228),
    .S(net150),
    .X(_0109_));
 sg13g2_mux2_1 _0901_ (.A0(net245),
    .A1(\trgg.cnt0.cnt[14] ),
    .S(net150),
    .X(_0110_));
 sg13g2_nor2_1 _0902_ (.A(net262),
    .B(net151),
    .Y(_0290_));
 sg13g2_a21oi_1 _0903_ (.A1(_0176_),
    .A2(net150),
    .Y(_0111_),
    .B1(_0290_));
 sg13g2_mux2_1 _0904_ (.A0(net239),
    .A1(\trgg.cnt0.cnt[16] ),
    .S(net151),
    .X(_0112_));
 sg13g2_mux2_1 _0905_ (.A0(net255),
    .A1(\trgg.cnt0.cnt[17] ),
    .S(net152),
    .X(_0113_));
 sg13g2_mux2_1 _0906_ (.A0(net271),
    .A1(net283),
    .S(net152),
    .X(_0114_));
 sg13g2_nor2_1 _0907_ (.A(net235),
    .B(net152),
    .Y(_0291_));
 sg13g2_a21oi_1 _0908_ (.A1(_0177_),
    .A2(net152),
    .Y(_0115_),
    .B1(_0291_));
 sg13g2_mux2_1 _0909_ (.A0(net250),
    .A1(\trgg.cnt0.cnt[20] ),
    .S(net152),
    .X(_0116_));
 sg13g2_nor2_1 _0910_ (.A(net259),
    .B(net152),
    .Y(_0292_));
 sg13g2_a21oi_1 _0911_ (.A1(_0178_),
    .A2(net152),
    .Y(_0117_),
    .B1(_0292_));
 sg13g2_mux2_1 _0912_ (.A0(net248),
    .A1(net225),
    .S(net152),
    .X(_0118_));
 sg13g2_mux2_1 _0913_ (.A0(net266),
    .A1(net237),
    .S(net153),
    .X(_0119_));
 sg13g2_dfrbp_1 _0914_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net74),
    .D(net270),
    .Q_N(_0438_),
    .Q(\trgg.shft.tx_word[0] ));
 sg13g2_dfrbp_1 _0915_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net68),
    .D(net407),
    .Q_N(_0437_),
    .Q(\trgg.shft.tx_word[1] ));
 sg13g2_dfrbp_1 _0916_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net67),
    .D(_0122_),
    .Q_N(_0436_),
    .Q(\trgg.shft.tx_word[2] ));
 sg13g2_dfrbp_1 _0917_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net66),
    .D(net420),
    .Q_N(_0435_),
    .Q(\trgg.shft.tx_word[3] ));
 sg13g2_dfrbp_1 _0918_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net65),
    .D(_0124_),
    .Q_N(_0434_),
    .Q(\trgg.shft.tx_word[4] ));
 sg13g2_dfrbp_1 _0919_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net64),
    .D(net400),
    .Q_N(_0433_),
    .Q(\trgg.shft.tx_word[5] ));
 sg13g2_dfrbp_1 _0920_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net63),
    .D(net334),
    .Q_N(_0432_),
    .Q(\trgg.shft.tx_word[6] ));
 sg13g2_dfrbp_1 _0921_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net62),
    .D(net405),
    .Q_N(_0431_),
    .Q(\trgg.shft.tx_word[7] ));
 sg13g2_dfrbp_1 _0922_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net61),
    .D(net389),
    .Q_N(_0430_),
    .Q(\trgg.shft.tx_word[8] ));
 sg13g2_dfrbp_1 _0923_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net60),
    .D(net454),
    .Q_N(_0429_),
    .Q(\trgg.shft.tx_word[9] ));
 sg13g2_dfrbp_1 _0924_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net59),
    .D(net446),
    .Q_N(_0428_),
    .Q(\trgg.shft.tx_word[10] ));
 sg13g2_dfrbp_1 _0925_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net58),
    .D(net450),
    .Q_N(_0427_),
    .Q(\trgg.shft.tx_word[11] ));
 sg13g2_dfrbp_1 _0926_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net57),
    .D(net387),
    .Q_N(_0426_),
    .Q(\trgg.shft.tx_word[12] ));
 sg13g2_dfrbp_1 _0927_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net56),
    .D(_0133_),
    .Q_N(_0425_),
    .Q(\trgg.shft.tx_word[13] ));
 sg13g2_dfrbp_1 _0928_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net55),
    .D(net385),
    .Q_N(_0424_),
    .Q(\trgg.shft.tx_word[14] ));
 sg13g2_dfrbp_1 _0929_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net54),
    .D(net379),
    .Q_N(_0423_),
    .Q(\trgg.shft.tx_word[15] ));
 sg13g2_dfrbp_1 _0930_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net53),
    .D(net337),
    .Q_N(_0422_),
    .Q(\trgg.shft.tx_word[16] ));
 sg13g2_dfrbp_1 _0931_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net52),
    .D(net327),
    .Q_N(_0421_),
    .Q(\trgg.shft.tx_word[17] ));
 sg13g2_dfrbp_1 _0932_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net51),
    .D(net436),
    .Q_N(_0420_),
    .Q(\trgg.shft.tx_word[18] ));
 sg13g2_dfrbp_1 _0933_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net50),
    .D(net430),
    .Q_N(_0419_),
    .Q(\trgg.shft.tx_word[19] ));
 sg13g2_dfrbp_1 _0934_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net49),
    .D(net426),
    .Q_N(_0418_),
    .Q(\trgg.shft.tx_word[20] ));
 sg13g2_dfrbp_1 _0935_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net48),
    .D(net428),
    .Q_N(_0417_),
    .Q(\trgg.shft.tx_word[21] ));
 sg13g2_dfrbp_1 _0936_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net47),
    .D(net416),
    .Q_N(_0416_),
    .Q(\trgg.shft.tx_word[22] ));
 sg13g2_dfrbp_1 _0937_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net46),
    .D(net424),
    .Q_N(_0415_),
    .Q(DAT_OUT));
 sg13g2_dfrbp_1 _0938_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net45),
    .D(net320),
    .Q_N(_0414_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][0] ));
 sg13g2_dfrbp_1 _0939_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net44),
    .D(_0145_),
    .Q_N(_0413_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][1] ));
 sg13g2_dfrbp_1 _0940_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net43),
    .D(_0146_),
    .Q_N(_0412_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][2] ));
 sg13g2_dfrbp_1 _0941_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net42),
    .D(net230),
    .Q_N(_0411_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][3] ));
 sg13g2_dfrbp_1 _0942_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net41),
    .D(_0148_),
    .Q_N(_0410_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][4] ));
 sg13g2_dfrbp_1 _0943_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net40),
    .D(_0149_),
    .Q_N(_0409_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][5] ));
 sg13g2_dfrbp_1 _0944_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net39),
    .D(_0150_),
    .Q_N(_0408_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][6] ));
 sg13g2_dfrbp_1 _0945_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net38),
    .D(_0151_),
    .Q_N(_0407_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][7] ));
 sg13g2_dfrbp_1 _0946_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net37),
    .D(net222),
    .Q_N(_0406_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][8] ));
 sg13g2_dfrbp_1 _0947_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net36),
    .D(net224),
    .Q_N(_0405_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][9] ));
 sg13g2_dfrbp_1 _0948_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net35),
    .D(net244),
    .Q_N(_0404_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][10] ));
 sg13g2_dfrbp_1 _0949_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net34),
    .D(net232),
    .Q_N(_0403_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][11] ));
 sg13g2_dfrbp_1 _0950_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net33),
    .D(_0156_),
    .Q_N(_0402_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][12] ));
 sg13g2_dfrbp_1 _0951_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net32),
    .D(net227),
    .Q_N(_0401_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][13] ));
 sg13g2_dfrbp_1 _0952_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net31),
    .D(_0158_),
    .Q_N(_0400_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][14] ));
 sg13g2_dfrbp_1 _0953_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net30),
    .D(_0159_),
    .Q_N(_0399_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][15] ));
 sg13g2_dfrbp_1 _0954_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net29),
    .D(_0160_),
    .Q_N(_0398_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][16] ));
 sg13g2_dfrbp_1 _0955_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net28),
    .D(_0161_),
    .Q_N(_0397_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][17] ));
 sg13g2_dfrbp_1 _0956_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net27),
    .D(net272),
    .Q_N(_0396_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][18] ));
 sg13g2_dfrbp_1 _0957_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net215),
    .D(_0163_),
    .Q_N(_0395_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][19] ));
 sg13g2_dfrbp_1 _0958_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net214),
    .D(_0164_),
    .Q_N(_0394_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][20] ));
 sg13g2_dfrbp_1 _0959_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net213),
    .D(_0165_),
    .Q_N(_0393_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][21] ));
 sg13g2_dfrbp_1 _0960_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net212),
    .D(net249),
    .Q_N(_0392_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][22] ));
 sg13g2_dfrbp_1 _0961_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net75),
    .D(_0167_),
    .Q_N(_0439_),
    .Q(\trgg.trigg_channel.mem.mem_regs[3][23] ));
 sg13g2_dfrbp_1 _0962_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net76),
    .D(_0000_),
    .Q_N(_0024_),
    .Q(\trgg.is_timestamp_popped_from_q ));
 sg13g2_dfrbp_1 _0963_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net77),
    .D(net3),
    .Q_N(_0440_),
    .Q(\trgg.shft.prev_ena ));
 sg13g2_dfrbp_1 _0964_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net102),
    .D(net2),
    .Q_N(_0441_),
    .Q(\trgg.shft.prev_dat_clk ));
 sg13g2_dfrbp_1 _0965_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net211),
    .D(net4),
    .Q_N(_0391_),
    .Q(\trgg.trigg_channel.ltch.prev_trigger ));
 sg13g2_dfrbp_1 _0966_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net210),
    .D(_0168_),
    .Q_N(_0390_),
    .Q(\trgg.trigg_channel.is_timestamp_present ));
 sg13g2_dfrbp_1 _0967_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net209),
    .D(net363),
    .Q_N(_0389_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][0] ));
 sg13g2_dfrbp_1 _0968_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net208),
    .D(_0025_),
    .Q_N(_0388_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][1] ));
 sg13g2_dfrbp_1 _0969_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net207),
    .D(_0026_),
    .Q_N(_0387_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][2] ));
 sg13g2_dfrbp_1 _0970_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net206),
    .D(_0027_),
    .Q_N(_0386_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][3] ));
 sg13g2_dfrbp_1 _0971_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net205),
    .D(net355),
    .Q_N(_0385_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][4] ));
 sg13g2_dfrbp_1 _0972_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net204),
    .D(_0029_),
    .Q_N(_0384_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][5] ));
 sg13g2_dfrbp_1 _0973_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net203),
    .D(_0030_),
    .Q_N(_0383_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][6] ));
 sg13g2_dfrbp_1 _0974_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net202),
    .D(_0031_),
    .Q_N(_0382_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][7] ));
 sg13g2_dfrbp_1 _0975_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net201),
    .D(_0032_),
    .Q_N(_0381_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][8] ));
 sg13g2_dfrbp_1 _0976_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net200),
    .D(_0033_),
    .Q_N(_0380_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][9] ));
 sg13g2_dfrbp_1 _0977_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net199),
    .D(_0034_),
    .Q_N(_0379_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][10] ));
 sg13g2_dfrbp_1 _0978_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net198),
    .D(_0035_),
    .Q_N(_0378_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][11] ));
 sg13g2_dfrbp_1 _0979_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net197),
    .D(_0036_),
    .Q_N(_0377_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][12] ));
 sg13g2_dfrbp_1 _0980_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net196),
    .D(_0037_),
    .Q_N(_0376_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][13] ));
 sg13g2_dfrbp_1 _0981_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net195),
    .D(_0038_),
    .Q_N(_0375_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][14] ));
 sg13g2_dfrbp_1 _0982_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net194),
    .D(_0039_),
    .Q_N(_0374_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][15] ));
 sg13g2_dfrbp_1 _0983_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net193),
    .D(_0040_),
    .Q_N(_0373_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][16] ));
 sg13g2_dfrbp_1 _0984_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net191),
    .D(_0041_),
    .Q_N(_0372_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][17] ));
 sg13g2_dfrbp_1 _0985_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net190),
    .D(net304),
    .Q_N(_0371_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][18] ));
 sg13g2_dfrbp_1 _0986_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net189),
    .D(_0043_),
    .Q_N(_0370_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][19] ));
 sg13g2_dfrbp_1 _0987_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net188),
    .D(_0044_),
    .Q_N(_0369_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][20] ));
 sg13g2_dfrbp_1 _0988_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net187),
    .D(_0045_),
    .Q_N(_0368_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][21] ));
 sg13g2_dfrbp_1 _0989_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net186),
    .D(_0046_),
    .Q_N(_0367_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][22] ));
 sg13g2_dfrbp_1 _0990_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net168),
    .D(_0047_),
    .Q_N(_0442_),
    .Q(\trgg.trigg_channel.mem.mem_regs[2][23] ));
 sg13g2_dfrbp_1 _0991_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net162),
    .D(\trgg.trigg_channel.mem.shift_gen[3].mem.if_will_be_data ),
    .Q_N(_0366_),
    .Q(\trgg.trigg_channel.is_mem_full ));
 sg13g2_dfrbp_1 _0992_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net185),
    .D(net432),
    .Q_N(_0365_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][0] ));
 sg13g2_dfrbp_1 _0993_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net184),
    .D(net308),
    .Q_N(_0364_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][1] ));
 sg13g2_dfrbp_1 _0994_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net183),
    .D(net403),
    .Q_N(_0363_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][2] ));
 sg13g2_dfrbp_1 _0995_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net182),
    .D(net342),
    .Q_N(_0362_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][3] ));
 sg13g2_dfrbp_1 _0996_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net181),
    .D(net381),
    .Q_N(_0361_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][4] ));
 sg13g2_dfrbp_1 _0997_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net180),
    .D(net322),
    .Q_N(_0360_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][5] ));
 sg13g2_dfrbp_1 _0998_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net179),
    .D(net310),
    .Q_N(_0359_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][6] ));
 sg13g2_dfrbp_1 _0999_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net178),
    .D(_0055_),
    .Q_N(_0358_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][7] ));
 sg13g2_dfrbp_1 _1000_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net177),
    .D(net287),
    .Q_N(_0357_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][8] ));
 sg13g2_dfrbp_1 _1001_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net176),
    .D(net289),
    .Q_N(_0356_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][9] ));
 sg13g2_dfrbp_1 _1002_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net175),
    .D(_0058_),
    .Q_N(_0355_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][10] ));
 sg13g2_dfrbp_1 _1003_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net174),
    .D(net299),
    .Q_N(_0354_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][11] ));
 sg13g2_dfrbp_1 _1004_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net173),
    .D(net369),
    .Q_N(_0353_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][12] ));
 sg13g2_dfrbp_1 _1005_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net172),
    .D(net391),
    .Q_N(_0352_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][13] ));
 sg13g2_dfrbp_1 _1006_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net171),
    .D(_0062_),
    .Q_N(_0351_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][14] ));
 sg13g2_dfrbp_1 _1007_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net170),
    .D(net314),
    .Q_N(_0350_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][15] ));
 sg13g2_dfrbp_1 _1008_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net169),
    .D(net344),
    .Q_N(_0349_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][16] ));
 sg13g2_dfrbp_1 _1009_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net167),
    .D(_0065_),
    .Q_N(_0348_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][17] ));
 sg13g2_dfrbp_1 _1010_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net166),
    .D(_0066_),
    .Q_N(_0347_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][18] ));
 sg13g2_dfrbp_1 _1011_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net165),
    .D(net357),
    .Q_N(_0346_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][19] ));
 sg13g2_dfrbp_1 _1012_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net164),
    .D(net292),
    .Q_N(_0345_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][20] ));
 sg13g2_dfrbp_1 _1013_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net163),
    .D(_0069_),
    .Q_N(_0344_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][21] ));
 sg13g2_dfrbp_1 _1014_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net120),
    .D(net332),
    .Q_N(_0343_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][22] ));
 sg13g2_dfrbp_1 _1015_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net192),
    .D(net306),
    .Q_N(_0443_),
    .Q(\trgg.trigg_channel.mem.mem_regs[1][23] ));
 sg13g2_dfrbp_1 _1016_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net162),
    .D(\trgg.trigg_channel.mem.shift_gen[2].mem.if_will_be_data ),
    .Q_N(_0342_),
    .Q(\trgg.trigg_channel.mem.shift_gen[1].mem.is_in ));
 sg13g2_dfrbp_1 _1017_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net119),
    .D(_0072_),
    .Q_N(_0341_),
    .Q(\trgg.shft.word_to_tx[0] ));
 sg13g2_dfrbp_1 _1018_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net118),
    .D(net462),
    .Q_N(_0340_),
    .Q(\trgg.shft.word_to_tx[1] ));
 sg13g2_dfrbp_1 _1019_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net117),
    .D(net440),
    .Q_N(_0339_),
    .Q(\trgg.shft.word_to_tx[2] ));
 sg13g2_dfrbp_1 _1020_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net116),
    .D(net365),
    .Q_N(_0338_),
    .Q(\trgg.shft.word_to_tx[3] ));
 sg13g2_dfrbp_1 _1021_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net115),
    .D(_0076_),
    .Q_N(_0337_),
    .Q(\trgg.shft.word_to_tx[4] ));
 sg13g2_dfrbp_1 _1022_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net114),
    .D(net414),
    .Q_N(_0336_),
    .Q(\trgg.shft.word_to_tx[5] ));
 sg13g2_dfrbp_1 _1023_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net113),
    .D(net329),
    .Q_N(_0335_),
    .Q(\trgg.shft.word_to_tx[6] ));
 sg13g2_dfrbp_1 _1024_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net112),
    .D(net350),
    .Q_N(_0334_),
    .Q(\trgg.shft.word_to_tx[7] ));
 sg13g2_dfrbp_1 _1025_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net111),
    .D(net376),
    .Q_N(_0333_),
    .Q(\trgg.shft.word_to_tx[8] ));
 sg13g2_dfrbp_1 _1026_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net110),
    .D(net434),
    .Q_N(_0332_),
    .Q(\trgg.shft.word_to_tx[9] ));
 sg13g2_dfrbp_1 _1027_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net109),
    .D(net361),
    .Q_N(_0331_),
    .Q(\trgg.shft.word_to_tx[10] ));
 sg13g2_dfrbp_1 _1028_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net108),
    .D(net324),
    .Q_N(_0330_),
    .Q(\trgg.shft.word_to_tx[11] ));
 sg13g2_dfrbp_1 _1029_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net107),
    .D(net383),
    .Q_N(_0329_),
    .Q(\trgg.shft.word_to_tx[12] ));
 sg13g2_dfrbp_1 _1030_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net106),
    .D(net396),
    .Q_N(_0328_),
    .Q(\trgg.shft.word_to_tx[13] ));
 sg13g2_dfrbp_1 _1031_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net105),
    .D(net312),
    .Q_N(_0327_),
    .Q(\trgg.shft.word_to_tx[14] ));
 sg13g2_dfrbp_1 _1032_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net104),
    .D(net316),
    .Q_N(_0326_),
    .Q(\trgg.shft.word_to_tx[15] ));
 sg13g2_dfrbp_1 _1033_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net103),
    .D(_0088_),
    .Q_N(_0325_),
    .Q(\trgg.shft.word_to_tx[16] ));
 sg13g2_dfrbp_1 _1034_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net101),
    .D(_0089_),
    .Q_N(_0324_),
    .Q(\trgg.shft.word_to_tx[17] ));
 sg13g2_dfrbp_1 _1035_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net100),
    .D(net296),
    .Q_N(_0323_),
    .Q(\trgg.shft.word_to_tx[18] ));
 sg13g2_dfrbp_1 _1036_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net99),
    .D(net372),
    .Q_N(_0322_),
    .Q(\trgg.shft.word_to_tx[19] ));
 sg13g2_dfrbp_1 _1037_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net98),
    .D(net452),
    .Q_N(_0321_),
    .Q(\trgg.shft.word_to_tx[20] ));
 sg13g2_dfrbp_1 _1038_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net97),
    .D(net302),
    .Q_N(_0320_),
    .Q(\trgg.shft.word_to_tx[21] ));
 sg13g2_dfrbp_1 _1039_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net96),
    .D(_0094_),
    .Q_N(_0319_),
    .Q(\trgg.shft.word_to_tx[22] ));
 sg13g2_dfrbp_1 _1040_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net216),
    .D(net442),
    .Q_N(_0444_),
    .Q(\trgg.shft.word_to_tx[23] ));
 sg13g2_dfrbp_1 _1041_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net162),
    .D(\trgg.trigg_channel.mem.shift_gen[1].mem.if_will_be_data ),
    .Q_N(_0318_),
    .Q(\trgg.trigg_channel.mem.shift_gen[0].mem.is_in ));
 sg13g2_dfrbp_1 _1042_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net95),
    .D(_0096_),
    .Q_N(_0317_),
    .Q(\trgg.trigg_channel.ltch.latched_time[0] ));
 sg13g2_dfrbp_1 _1043_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net94),
    .D(net265),
    .Q_N(_0316_),
    .Q(\trgg.trigg_channel.ltch.latched_time[1] ));
 sg13g2_dfrbp_1 _1044_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net93),
    .D(_0098_),
    .Q_N(_0315_),
    .Q(\trgg.trigg_channel.ltch.latched_time[2] ));
 sg13g2_dfrbp_1 _1045_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net92),
    .D(_0099_),
    .Q_N(_0314_),
    .Q(\trgg.trigg_channel.ltch.latched_time[3] ));
 sg13g2_dfrbp_1 _1046_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net91),
    .D(net340),
    .Q_N(_0313_),
    .Q(\trgg.trigg_channel.ltch.latched_time[4] ));
 sg13g2_dfrbp_1 _1047_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net90),
    .D(net275),
    .Q_N(_0312_),
    .Q(\trgg.trigg_channel.ltch.latched_time[5] ));
 sg13g2_dfrbp_1 _1048_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net89),
    .D(net278),
    .Q_N(_0311_),
    .Q(\trgg.trigg_channel.ltch.latched_time[6] ));
 sg13g2_dfrbp_1 _1049_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net88),
    .D(net253),
    .Q_N(_0310_),
    .Q(\trgg.trigg_channel.ltch.latched_time[7] ));
 sg13g2_dfrbp_1 _1050_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net87),
    .D(_0104_),
    .Q_N(_0309_),
    .Q(\trgg.trigg_channel.ltch.latched_time[8] ));
 sg13g2_dfrbp_1 _1051_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net86),
    .D(_0105_),
    .Q_N(_0308_),
    .Q(\trgg.trigg_channel.ltch.latched_time[9] ));
 sg13g2_dfrbp_1 _1052_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net85),
    .D(_0106_),
    .Q_N(_0307_),
    .Q(\trgg.trigg_channel.ltch.latched_time[10] ));
 sg13g2_dfrbp_1 _1053_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net84),
    .D(_0107_),
    .Q_N(_0306_),
    .Q(\trgg.trigg_channel.ltch.latched_time[11] ));
 sg13g2_dfrbp_1 _1054_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net83),
    .D(net242),
    .Q_N(_0305_),
    .Q(\trgg.trigg_channel.ltch.latched_time[12] ));
 sg13g2_dfrbp_1 _1055_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net82),
    .D(_0109_),
    .Q_N(_0304_),
    .Q(\trgg.trigg_channel.ltch.latched_time[13] ));
 sg13g2_dfrbp_1 _1056_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net81),
    .D(net246),
    .Q_N(_0303_),
    .Q(\trgg.trigg_channel.ltch.latched_time[14] ));
 sg13g2_dfrbp_1 _1057_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net80),
    .D(net263),
    .Q_N(_0302_),
    .Q(\trgg.trigg_channel.ltch.latched_time[15] ));
 sg13g2_dfrbp_1 _1058_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net79),
    .D(net240),
    .Q_N(_0301_),
    .Q(\trgg.trigg_channel.ltch.latched_time[16] ));
 sg13g2_dfrbp_1 _1059_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net78),
    .D(net256),
    .Q_N(_0300_),
    .Q(\trgg.trigg_channel.ltch.latched_time[17] ));
 sg13g2_dfrbp_1 _1060_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net73),
    .D(_0114_),
    .Q_N(_0299_),
    .Q(\trgg.trigg_channel.ltch.latched_time[18] ));
 sg13g2_dfrbp_1 _1061_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net72),
    .D(net236),
    .Q_N(_0298_),
    .Q(\trgg.trigg_channel.ltch.latched_time[19] ));
 sg13g2_dfrbp_1 _1062_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net71),
    .D(net251),
    .Q_N(_0297_),
    .Q(\trgg.trigg_channel.ltch.latched_time[20] ));
 sg13g2_dfrbp_1 _1063_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net70),
    .D(net260),
    .Q_N(_0296_),
    .Q(\trgg.trigg_channel.ltch.latched_time[21] ));
 sg13g2_dfrbp_1 _1064_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net69),
    .D(_0118_),
    .Q_N(_0295_),
    .Q(\trgg.trigg_channel.ltch.latched_time[22] ));
 sg13g2_dfrbp_1 _1065_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net217),
    .D(_0119_),
    .Q_N(_0445_),
    .Q(\trgg.trigg_channel.ltch.latched_time[23] ));
 sg13g2_dfrbp_1 _1066_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net162),
    .D(net220),
    .Q_N(_0446_),
    .Q(DAT_RDY));
 sg13g2_dfrbp_1 _1067_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net162),
    .D(net218),
    .Q_N(_0293_),
    .Q(\trgg.cnt0.cnt[0] ));
 sg13g2_dfrbp_1 _1068_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net161),
    .D(_0011_),
    .Q_N(_0447_),
    .Q(\trgg.cnt0.cnt[1] ));
 sg13g2_dfrbp_1 _1069_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net161),
    .D(_0016_),
    .Q_N(_0448_),
    .Q(\trgg.cnt0.cnt[2] ));
 sg13g2_dfrbp_1 _1070_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net161),
    .D(_0017_),
    .Q_N(_0449_),
    .Q(\trgg.cnt0.cnt[3] ));
 sg13g2_dfrbp_1 _1071_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net160),
    .D(net448),
    .Q_N(_0450_),
    .Q(\trgg.cnt0.cnt[4] ));
 sg13g2_dfrbp_1 _1072_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net160),
    .D(_0019_),
    .Q_N(_0451_),
    .Q(\trgg.cnt0.cnt[5] ));
 sg13g2_dfrbp_1 _1073_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net160),
    .D(net318),
    .Q_N(_0452_),
    .Q(\trgg.cnt0.cnt[6] ));
 sg13g2_dfrbp_1 _1074_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net160),
    .D(net347),
    .Q_N(_0453_),
    .Q(\trgg.cnt0.cnt[7] ));
 sg13g2_dfrbp_1 _1075_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net159),
    .D(_0022_),
    .Q_N(_0454_),
    .Q(\trgg.cnt0.cnt[8] ));
 sg13g2_dfrbp_1 _1076_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net159),
    .D(_0023_),
    .Q_N(_0455_),
    .Q(\trgg.cnt0.cnt[9] ));
 sg13g2_dfrbp_1 _1077_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net159),
    .D(_0001_),
    .Q_N(_0456_),
    .Q(\trgg.cnt0.cnt[10] ));
 sg13g2_dfrbp_1 _1078_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net159),
    .D(_0002_),
    .Q_N(_0457_),
    .Q(\trgg.cnt0.cnt[11] ));
 sg13g2_dfrbp_1 _1079_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net159),
    .D(_0003_),
    .Q_N(_0458_),
    .Q(\trgg.cnt0.cnt[12] ));
 sg13g2_dfrbp_1 _1080_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net159),
    .D(_0004_),
    .Q_N(_0459_),
    .Q(\trgg.cnt0.cnt[13] ));
 sg13g2_dfrbp_1 _1081_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net159),
    .D(net410),
    .Q_N(_0460_),
    .Q(\trgg.cnt0.cnt[14] ));
 sg13g2_dfrbp_1 _1082_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net159),
    .D(net412),
    .Q_N(_0461_),
    .Q(\trgg.cnt0.cnt[15] ));
 sg13g2_dfrbp_1 _1083_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net160),
    .D(_0007_),
    .Q_N(_0462_),
    .Q(\trgg.cnt0.cnt[16] ));
 sg13g2_dfrbp_1 _1084_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net160),
    .D(net459),
    .Q_N(_0463_),
    .Q(\trgg.cnt0.cnt[17] ));
 sg13g2_dfrbp_1 _1085_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net160),
    .D(_0009_),
    .Q_N(_0464_),
    .Q(\trgg.cnt0.cnt[18] ));
 sg13g2_dfrbp_1 _1086_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net161),
    .D(net470),
    .Q_N(_0465_),
    .Q(\trgg.cnt0.cnt[19] ));
 sg13g2_dfrbp_1 _1087_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net161),
    .D(_0012_),
    .Q_N(_0466_),
    .Q(\trgg.cnt0.cnt[20] ));
 sg13g2_dfrbp_1 _1088_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net161),
    .D(net456),
    .Q_N(_0467_),
    .Q(\trgg.cnt0.cnt[21] ));
 sg13g2_dfrbp_1 _1089_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net161),
    .D(_0014_),
    .Q_N(_0468_),
    .Q(\trgg.cnt0.cnt[22] ));
 sg13g2_dfrbp_1 _1090_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net161),
    .D(net238),
    .Q_N(_0294_),
    .Q(\trgg.cnt0.cnt[23] ));
 sg13g2_tiehi _0955__28 (.L_HI(net28));
 sg13g2_tiehi _0954__29 (.L_HI(net29));
 sg13g2_tiehi _0953__30 (.L_HI(net30));
 sg13g2_tiehi _0952__31 (.L_HI(net31));
 sg13g2_tiehi _0951__32 (.L_HI(net32));
 sg13g2_tiehi _0950__33 (.L_HI(net33));
 sg13g2_tiehi _0949__34 (.L_HI(net34));
 sg13g2_tiehi _0948__35 (.L_HI(net35));
 sg13g2_tiehi _0947__36 (.L_HI(net36));
 sg13g2_tiehi _0946__37 (.L_HI(net37));
 sg13g2_tiehi _0945__38 (.L_HI(net38));
 sg13g2_tiehi _0944__39 (.L_HI(net39));
 sg13g2_tiehi _0943__40 (.L_HI(net40));
 sg13g2_tiehi _0942__41 (.L_HI(net41));
 sg13g2_tiehi _0941__42 (.L_HI(net42));
 sg13g2_tiehi _0940__43 (.L_HI(net43));
 sg13g2_tiehi _0939__44 (.L_HI(net44));
 sg13g2_tiehi _0938__45 (.L_HI(net45));
 sg13g2_tiehi _0937__46 (.L_HI(net46));
 sg13g2_tiehi _0936__47 (.L_HI(net47));
 sg13g2_tiehi _0935__48 (.L_HI(net48));
 sg13g2_tiehi _0934__49 (.L_HI(net49));
 sg13g2_tiehi _0933__50 (.L_HI(net50));
 sg13g2_tiehi _0932__51 (.L_HI(net51));
 sg13g2_tiehi _0931__52 (.L_HI(net52));
 sg13g2_tiehi _0930__53 (.L_HI(net53));
 sg13g2_tiehi _0929__54 (.L_HI(net54));
 sg13g2_tiehi _0928__55 (.L_HI(net55));
 sg13g2_tiehi _0927__56 (.L_HI(net56));
 sg13g2_tiehi _0926__57 (.L_HI(net57));
 sg13g2_tiehi _0925__58 (.L_HI(net58));
 sg13g2_tiehi _0924__59 (.L_HI(net59));
 sg13g2_tiehi _0923__60 (.L_HI(net60));
 sg13g2_tiehi _0922__61 (.L_HI(net61));
 sg13g2_tiehi _0921__62 (.L_HI(net62));
 sg13g2_tiehi _0920__63 (.L_HI(net63));
 sg13g2_tiehi _0919__64 (.L_HI(net64));
 sg13g2_tiehi _0918__65 (.L_HI(net65));
 sg13g2_tiehi _0917__66 (.L_HI(net66));
 sg13g2_tiehi _0916__67 (.L_HI(net67));
 sg13g2_tiehi _0915__68 (.L_HI(net68));
 sg13g2_tiehi _1064__69 (.L_HI(net69));
 sg13g2_tiehi _1063__70 (.L_HI(net70));
 sg13g2_tiehi _1062__71 (.L_HI(net71));
 sg13g2_tiehi _1061__72 (.L_HI(net72));
 sg13g2_tiehi _1060__73 (.L_HI(net73));
 sg13g2_tiehi _0914__74 (.L_HI(net74));
 sg13g2_tiehi _0961__75 (.L_HI(net75));
 sg13g2_tiehi _0962__76 (.L_HI(net76));
 sg13g2_tiehi _0963__77 (.L_HI(net77));
 sg13g2_tiehi _1059__78 (.L_HI(net78));
 sg13g2_tiehi _1058__79 (.L_HI(net79));
 sg13g2_tiehi _1057__80 (.L_HI(net80));
 sg13g2_tiehi _1056__81 (.L_HI(net81));
 sg13g2_tiehi _1055__82 (.L_HI(net82));
 sg13g2_tiehi _1054__83 (.L_HI(net83));
 sg13g2_tiehi _1053__84 (.L_HI(net84));
 sg13g2_tiehi _1052__85 (.L_HI(net85));
 sg13g2_tiehi _1051__86 (.L_HI(net86));
 sg13g2_tiehi _1050__87 (.L_HI(net87));
 sg13g2_tiehi _1049__88 (.L_HI(net88));
 sg13g2_tiehi _1048__89 (.L_HI(net89));
 sg13g2_tiehi _1047__90 (.L_HI(net90));
 sg13g2_tiehi _1046__91 (.L_HI(net91));
 sg13g2_tiehi _1045__92 (.L_HI(net92));
 sg13g2_tiehi _1044__93 (.L_HI(net93));
 sg13g2_tiehi _1043__94 (.L_HI(net94));
 sg13g2_tiehi _1042__95 (.L_HI(net95));
 sg13g2_tiehi _1039__96 (.L_HI(net96));
 sg13g2_tiehi _1038__97 (.L_HI(net97));
 sg13g2_tiehi _1037__98 (.L_HI(net98));
 sg13g2_tiehi _1036__99 (.L_HI(net99));
 sg13g2_tiehi _1035__100 (.L_HI(net100));
 sg13g2_tiehi _1034__101 (.L_HI(net101));
 sg13g2_tiehi _0964__102 (.L_HI(net102));
 sg13g2_tiehi _1033__103 (.L_HI(net103));
 sg13g2_tiehi _1032__104 (.L_HI(net104));
 sg13g2_tiehi _1031__105 (.L_HI(net105));
 sg13g2_tiehi _1030__106 (.L_HI(net106));
 sg13g2_tiehi _1029__107 (.L_HI(net107));
 sg13g2_tiehi _1028__108 (.L_HI(net108));
 sg13g2_tiehi _1027__109 (.L_HI(net109));
 sg13g2_tiehi _1026__110 (.L_HI(net110));
 sg13g2_tiehi _1025__111 (.L_HI(net111));
 sg13g2_tiehi _1024__112 (.L_HI(net112));
 sg13g2_tiehi _1023__113 (.L_HI(net113));
 sg13g2_tiehi _1022__114 (.L_HI(net114));
 sg13g2_tiehi _1021__115 (.L_HI(net115));
 sg13g2_tiehi _1020__116 (.L_HI(net116));
 sg13g2_tiehi _1019__117 (.L_HI(net117));
 sg13g2_tiehi _1018__118 (.L_HI(net118));
 sg13g2_tiehi _1017__119 (.L_HI(net119));
 sg13g2_tiehi _1014__120 (.L_HI(net120));
 sg13g2_tiehi _1013__121 (.L_HI(net163));
 sg13g2_tiehi _1012__122 (.L_HI(net164));
 sg13g2_tiehi _1011__123 (.L_HI(net165));
 sg13g2_tiehi _1010__124 (.L_HI(net166));
 sg13g2_tiehi _1009__125 (.L_HI(net167));
 sg13g2_tiehi _0990__126 (.L_HI(net168));
 sg13g2_tiehi _1008__127 (.L_HI(net169));
 sg13g2_tiehi _1007__128 (.L_HI(net170));
 sg13g2_tiehi _1006__129 (.L_HI(net171));
 sg13g2_tiehi _1005__130 (.L_HI(net172));
 sg13g2_tiehi _1004__131 (.L_HI(net173));
 sg13g2_tiehi _1003__132 (.L_HI(net174));
 sg13g2_tiehi _1002__133 (.L_HI(net175));
 sg13g2_tiehi _1001__134 (.L_HI(net176));
 sg13g2_tiehi _1000__135 (.L_HI(net177));
 sg13g2_tiehi _0999__136 (.L_HI(net178));
 sg13g2_tiehi _0998__137 (.L_HI(net179));
 sg13g2_tiehi _0997__138 (.L_HI(net180));
 sg13g2_tiehi _0996__139 (.L_HI(net181));
 sg13g2_tiehi _0995__140 (.L_HI(net182));
 sg13g2_tiehi _0994__141 (.L_HI(net183));
 sg13g2_tiehi _0993__142 (.L_HI(net184));
 sg13g2_tiehi _0992__143 (.L_HI(net185));
 sg13g2_tiehi _0989__144 (.L_HI(net186));
 sg13g2_tiehi _0988__145 (.L_HI(net187));
 sg13g2_tiehi _0987__146 (.L_HI(net188));
 sg13g2_tiehi _0986__147 (.L_HI(net189));
 sg13g2_tiehi _0985__148 (.L_HI(net190));
 sg13g2_tiehi _0984__149 (.L_HI(net191));
 sg13g2_tiehi _1015__150 (.L_HI(net192));
 sg13g2_tiehi _0983__151 (.L_HI(net193));
 sg13g2_tiehi _0982__152 (.L_HI(net194));
 sg13g2_tiehi _0981__153 (.L_HI(net195));
 sg13g2_tiehi _0980__154 (.L_HI(net196));
 sg13g2_tiehi _0979__155 (.L_HI(net197));
 sg13g2_tiehi _0978__156 (.L_HI(net198));
 sg13g2_tiehi _0977__157 (.L_HI(net199));
 sg13g2_tiehi _0976__158 (.L_HI(net200));
 sg13g2_tiehi _0975__159 (.L_HI(net201));
 sg13g2_tiehi _0974__160 (.L_HI(net202));
 sg13g2_tiehi _0973__161 (.L_HI(net203));
 sg13g2_tiehi _0972__162 (.L_HI(net204));
 sg13g2_tiehi _0971__163 (.L_HI(net205));
 sg13g2_tiehi _0970__164 (.L_HI(net206));
 sg13g2_tiehi _0969__165 (.L_HI(net207));
 sg13g2_tiehi _0968__166 (.L_HI(net208));
 sg13g2_tiehi _0967__167 (.L_HI(net209));
 sg13g2_tiehi _0966__168 (.L_HI(net210));
 sg13g2_tiehi _0965__169 (.L_HI(net211));
 sg13g2_tiehi _0960__170 (.L_HI(net212));
 sg13g2_tiehi _0959__171 (.L_HI(net213));
 sg13g2_tiehi _0958__172 (.L_HI(net214));
 sg13g2_tiehi _0957__173 (.L_HI(net215));
 sg13g2_tiehi _1040__174 (.L_HI(net216));
 sg13g2_tiehi _1065__175 (.L_HI(net217));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_tetrap_triggerer_6 (.L_LO(net6));
 sg13g2_tielo tt_um_tetrap_triggerer_7 (.L_LO(net7));
 sg13g2_tielo tt_um_tetrap_triggerer_8 (.L_LO(net8));
 sg13g2_tielo tt_um_tetrap_triggerer_9 (.L_LO(net9));
 sg13g2_tielo tt_um_tetrap_triggerer_10 (.L_LO(net10));
 sg13g2_tielo tt_um_tetrap_triggerer_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tetrap_triggerer_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tetrap_triggerer_13 (.L_LO(net13));
 sg13g2_tielo tt_um_tetrap_triggerer_14 (.L_LO(net14));
 sg13g2_tielo tt_um_tetrap_triggerer_15 (.L_LO(net15));
 sg13g2_tielo tt_um_tetrap_triggerer_16 (.L_LO(net16));
 sg13g2_tielo tt_um_tetrap_triggerer_17 (.L_LO(net17));
 sg13g2_tielo tt_um_tetrap_triggerer_18 (.L_LO(net18));
 sg13g2_tielo tt_um_tetrap_triggerer_19 (.L_LO(net19));
 sg13g2_tielo tt_um_tetrap_triggerer_20 (.L_LO(net20));
 sg13g2_tielo tt_um_tetrap_triggerer_21 (.L_LO(net21));
 sg13g2_tielo tt_um_tetrap_triggerer_22 (.L_LO(net22));
 sg13g2_tielo tt_um_tetrap_triggerer_23 (.L_LO(net23));
 sg13g2_tielo tt_um_tetrap_triggerer_24 (.L_LO(net24));
 sg13g2_tielo tt_um_tetrap_triggerer_25 (.L_LO(net25));
 sg13g2_tielo tt_um_tetrap_triggerer_26 (.L_LO(net26));
 sg13g2_tiehi _0956__27 (.L_HI(net27));
 sg13g2_buf_1 _1262_ (.A(DAT_OUT),
    .X(uo_out[0]));
 sg13g2_buf_1 _1263_ (.A(DAT_RDY),
    .X(uo_out[1]));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(net125));
 sg13g2_buf_2 fanout122 (.A(net125),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(net125));
 sg13g2_buf_2 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0287_),
    .X(net125));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(net130));
 sg13g2_buf_2 fanout127 (.A(net130),
    .X(net127));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(net130));
 sg13g2_buf_2 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0286_),
    .X(net130));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(net135));
 sg13g2_buf_2 fanout132 (.A(net135),
    .X(net132));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(net135));
 sg13g2_buf_2 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_0285_),
    .X(net135));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(net140));
 sg13g2_buf_2 fanout137 (.A(net140),
    .X(net137));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(net140));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_0283_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(net144),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_1 fanout144 (.A(_0215_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(net146),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(net148),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_1 fanout148 (.A(_0211_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_0201_),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(net151));
 sg13g2_buf_2 fanout151 (.A(net154),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net154),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net281),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_0179_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_0179_),
    .X(net157));
 sg13g2_buf_1 fanout158 (.A(_0179_),
    .X(net158));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(net160));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(net162));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(net162));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(net1));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_tielo tt_um_tetrap_triggerer_5 (.L_LO(net5));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0293_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0024_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold3 (.A(\trgg.trigg_channel.mem.shift_gen[0].mem.if_will_be_data ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold4 (.A(\trgg.trigg_channel.ltch.latched_time[8] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0152_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold6 (.A(\trgg.trigg_channel.ltch.latched_time[9] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0153_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold8 (.A(\trgg.cnt0.cnt[22] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold9 (.A(\trgg.trigg_channel.ltch.latched_time[13] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0157_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold11 (.A(\trgg.cnt0.cnt[13] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold12 (.A(\trgg.trigg_channel.ltch.latched_time[3] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0147_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold14 (.A(\trgg.trigg_channel.ltch.latched_time[11] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0155_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold16 (.A(\trgg.cnt0.cnt[8] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold17 (.A(\trgg.cnt0.cnt[3] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold18 (.A(\trgg.trigg_channel.ltch.latched_time[19] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0115_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold20 (.A(\trgg.cnt0.cnt[23] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0015_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold22 (.A(\trgg.trigg_channel.ltch.latched_time[16] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0112_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold24 (.A(\trgg.trigg_channel.ltch.latched_time[12] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0108_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold26 (.A(\trgg.trigg_channel.ltch.latched_time[10] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0154_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold28 (.A(\trgg.trigg_channel.ltch.latched_time[14] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0110_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold30 (.A(\trgg.trigg_channel.mem.mem_regs[3][16] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold31 (.A(\trgg.trigg_channel.ltch.latched_time[22] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0166_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold33 (.A(\trgg.trigg_channel.ltch.latched_time[20] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0116_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold35 (.A(\trgg.trigg_channel.ltch.latched_time[7] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0103_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold37 (.A(\trgg.trigg_channel.mem.mem_regs[3][12] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold38 (.A(\trgg.trigg_channel.ltch.latched_time[17] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0113_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold40 (.A(\trgg.cnt0.cnt[2] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0184_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold42 (.A(\trgg.trigg_channel.ltch.latched_time[21] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0117_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold44 (.A(\trgg.cnt0.cnt[9] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold45 (.A(\trgg.trigg_channel.ltch.latched_time[15] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0111_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold47 (.A(\trgg.trigg_channel.ltch.latched_time[1] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0097_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold49 (.A(\trgg.trigg_channel.ltch.latched_time[23] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold50 (.A(\trgg.trigg_channel.mem.mem_regs[3][20] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold51 (.A(\trgg.cnt0.cnt[10] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold52 (.A(\trgg.shft.word_to_tx[0] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0120_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold54 (.A(\trgg.trigg_channel.ltch.latched_time[18] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0162_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold56 (.A(\trgg.trigg_channel.mem.mem_regs[3][17] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold57 (.A(\trgg.trigg_channel.ltch.latched_time[5] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0101_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold59 (.A(\trgg.trigg_channel.mem.mem_regs[3][7] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold60 (.A(\trgg.trigg_channel.ltch.latched_time[6] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0102_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold62 (.A(\trgg.trigg_channel.ltch.latched_time[2] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold63 (.A(\trgg.trigg_channel.ltch.prev_trigger ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0284_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold65 (.A(\trgg.cnt0.cnt[11] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold66 (.A(\trgg.cnt0.cnt[18] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold67 (.A(\trgg.trigg_channel.mem.mem_regs[3][14] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold68 (.A(\trgg.trigg_channel.mem.mem_regs[3][23] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold69 (.A(\trgg.trigg_channel.mem.mem_regs[2][8] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0056_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold71 (.A(\trgg.trigg_channel.mem.mem_regs[2][9] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0057_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold73 (.A(\trgg.trigg_channel.mem.mem_regs[3][1] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold74 (.A(\trgg.trigg_channel.mem.mem_regs[2][20] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0068_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold76 (.A(\trgg.trigg_channel.mem.mem_regs[3][5] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold77 (.A(\trgg.trigg_channel.mem.mem_regs[2][7] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold78 (.A(\trgg.trigg_channel.mem.mem_regs[1][18] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0090_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold80 (.A(\trgg.trigg_channel.mem.mem_regs[3][6] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold81 (.A(\trgg.trigg_channel.mem.mem_regs[2][11] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0059_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold83 (.A(\trgg.trigg_channel.mem.mem_regs[3][2] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold84 (.A(\trgg.trigg_channel.mem.mem_regs[1][21] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0093_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold86 (.A(\trgg.trigg_channel.mem.mem_regs[3][18] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0042_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold88 (.A(\trgg.trigg_channel.mem.mem_regs[2][23] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0071_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold90 (.A(\trgg.trigg_channel.mem.mem_regs[2][1] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0049_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold92 (.A(\trgg.trigg_channel.mem.mem_regs[2][6] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0054_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold94 (.A(\trgg.trigg_channel.mem.mem_regs[1][14] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0086_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold96 (.A(\trgg.trigg_channel.mem.mem_regs[2][15] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0063_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold98 (.A(\trgg.trigg_channel.mem.mem_regs[1][15] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0087_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold100 (.A(\trgg.cnt0.cnt[6] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0020_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold102 (.A(\trgg.trigg_channel.ltch.latched_time[0] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0144_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold104 (.A(\trgg.trigg_channel.mem.mem_regs[2][5] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0053_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold106 (.A(\trgg.trigg_channel.mem.mem_regs[1][11] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0083_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold108 (.A(\trgg.trigg_channel.mem.mem_regs[3][19] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold109 (.A(\trgg.shft.word_to_tx[17] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0137_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold111 (.A(\trgg.trigg_channel.mem.mem_regs[1][6] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0078_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold113 (.A(\trgg.trigg_channel.mem.mem_regs[2][21] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold114 (.A(\trgg.trigg_channel.mem.mem_regs[2][22] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0070_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold116 (.A(\trgg.shft.word_to_tx[6] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0126_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold118 (.A(\trgg.trigg_channel.mem.mem_regs[2][17] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold119 (.A(\trgg.shft.word_to_tx[16] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0136_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold121 (.A(\trgg.cnt0.cnt[0] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold122 (.A(\trgg.trigg_channel.ltch.latched_time[4] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0100_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold124 (.A(\trgg.trigg_channel.mem.mem_regs[2][3] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0051_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold126 (.A(\trgg.trigg_channel.mem.mem_regs[2][16] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0064_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold128 (.A(\trgg.cnt0.cnt[7] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0191_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0021_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold131 (.A(\trgg.trigg_channel.mem.mem_regs[3][3] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold132 (.A(\trgg.trigg_channel.mem.mem_regs[1][7] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0079_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold134 (.A(\trgg.trigg_channel.mem.shift_gen[1].mem.is_in ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0180_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold136 (.A(\trgg.trigg_channel.mem.mem_regs[2][18] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold137 (.A(\trgg.trigg_channel.mem.mem_regs[3][4] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0028_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold139 (.A(\trgg.trigg_channel.mem.mem_regs[2][19] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0067_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold141 (.A(\trgg.trigg_channel.mem.mem_regs[3][15] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold142 (.A(\trgg.trigg_channel.mem.mem_regs[3][21] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold143 (.A(\trgg.trigg_channel.mem.mem_regs[1][10] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0082_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold145 (.A(\trgg.trigg_channel.mem.mem_regs[3][0] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0169_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold147 (.A(\trgg.trigg_channel.mem.mem_regs[1][3] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0075_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold149 (.A(\trgg.trigg_channel.is_mem_full ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold150 (.A(\trgg.trigg_channel.mem.mem_regs[2][14] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold151 (.A(\trgg.trigg_channel.mem.mem_regs[2][12] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0060_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold153 (.A(\trgg.trigg_channel.mem.shift_gen[0].mem.is_in ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold154 (.A(\trgg.trigg_channel.mem.mem_regs[1][19] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0091_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold156 (.A(\trgg.trigg_channel.mem.mem_regs[1][16] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold157 (.A(\trgg.trigg_channel.mem.mem_regs[1][17] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold158 (.A(\trgg.trigg_channel.mem.mem_regs[1][8] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0080_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold160 (.A(\trgg.trigg_channel.mem.mem_regs[2][10] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold161 (.A(\trgg.shft.tx_word[14] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0135_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold163 (.A(\trgg.trigg_channel.mem.mem_regs[1][4] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0052_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold165 (.A(\trgg.trigg_channel.mem.mem_regs[1][12] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0084_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold167 (.A(\trgg.shft.tx_word[13] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0134_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold169 (.A(\trgg.shft.tx_word[12] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0132_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold171 (.A(\trgg.shft.word_to_tx[8] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0128_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold173 (.A(\trgg.trigg_channel.mem.mem_regs[2][13] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0061_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold175 (.A(\trgg.trigg_channel.mem.mem_regs[3][22] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold176 (.A(\trgg.trigg_channel.mem.mem_regs[3][9] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold177 (.A(\trgg.trigg_channel.mem.mem_regs[3][13] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold178 (.A(\trgg.trigg_channel.mem.mem_regs[1][13] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0085_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold180 (.A(\trgg.trigg_channel.mem.mem_regs[3][8] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold181 (.A(\trgg.trigg_channel.is_timestamp_present ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold182 (.A(\trgg.shft.tx_word[4] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0125_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold184 (.A(\trgg.trigg_channel.mem.mem_regs[3][11] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold185 (.A(\trgg.trigg_channel.mem.mem_regs[2][2] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0050_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold187 (.A(\trgg.shft.word_to_tx[7] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0127_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold189 (.A(\trgg.shft.tx_word[0] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0121_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold191 (.A(\trgg.shft.word_to_tx[4] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold192 (.A(\trgg.cnt0.cnt[14] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0005_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold194 (.A(\trgg.cnt0.cnt[15] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0006_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold196 (.A(\trgg.trigg_channel.mem.mem_regs[1][5] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0077_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold198 (.A(\trgg.shft.word_to_tx[22] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0142_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold200 (.A(\trgg.shft.word_to_tx[13] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold201 (.A(\trgg.trigg_channel.mem.mem_regs[3][10] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold202 (.A(\trgg.shft.tx_word[2] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0123_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold204 (.A(\trgg.cnt0.cnt[20] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0206_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold206 (.A(\trgg.shft.tx_word[22] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0143_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold208 (.A(\trgg.shft.tx_word[19] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0140_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold210 (.A(\trgg.shft.word_to_tx[21] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0141_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold212 (.A(\trgg.shft.tx_word[18] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0139_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold214 (.A(\trgg.trigg_channel.mem.mem_regs[2][0] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0048_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold216 (.A(\trgg.trigg_channel.mem.mem_regs[1][9] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0081_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold218 (.A(\trgg.shft.word_to_tx[18] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0138_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold220 (.A(\trgg.cnt0.cnt[5] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold221 (.A(\trgg.cnt0.cnt[8] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold222 (.A(\trgg.shft.word_to_tx[2] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0074_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold224 (.A(\trgg.trigg_channel.mem.mem_regs[1][23] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0095_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold226 (.A(\trgg.shft.tx_word[1] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold227 (.A(\trgg.trigg_channel.mem.mem_regs[1][0] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold228 (.A(\trgg.shft.word_to_tx[10] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0130_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold230 (.A(\trgg.cnt0.cnt[4] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0018_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold232 (.A(\trgg.shft.word_to_tx[11] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0131_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold234 (.A(\trgg.shft.word_to_tx[20] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0092_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold236 (.A(\trgg.shft.tx_word[9] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0129_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold238 (.A(\trgg.cnt0.cnt[21] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0013_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold240 (.A(\trgg.cnt0.cnt[17] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0202_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0008_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold243 (.A(\trgg.cnt0.cnt[16] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold244 (.A(\trgg.trigg_channel.mem.mem_regs[1][1] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0073_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold246 (.A(\trgg.cnt0.cnt[1] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold247 (.A(\trgg.cnt0.cnt[12] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold248 (.A(\trgg.trigg_channel.mem.mem_regs[1][22] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold249 (.A(DAT_RDY),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold250 (.A(\trgg.shft.tx_word[3] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold251 (.A(\trgg.cnt0.cnt[4] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold252 (.A(\trgg.cnt0.cnt[19] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0010_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold254 (.A(\trgg.shft.prev_ena ),
    .X(net471));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_fill_2 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_272 ();
 sg13g2_decap_8 FILLER_3_279 ();
 sg13g2_decap_8 FILLER_3_286 ();
 sg13g2_decap_8 FILLER_3_293 ();
 sg13g2_decap_8 FILLER_3_300 ();
 sg13g2_decap_8 FILLER_3_307 ();
 sg13g2_decap_8 FILLER_3_314 ();
 sg13g2_decap_8 FILLER_3_321 ();
 sg13g2_decap_8 FILLER_3_328 ();
 sg13g2_decap_8 FILLER_3_335 ();
 sg13g2_decap_8 FILLER_3_342 ();
 sg13g2_decap_8 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_356 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_156 ();
 sg13g2_decap_4 FILLER_4_163 ();
 sg13g2_decap_8 FILLER_4_171 ();
 sg13g2_fill_1 FILLER_4_178 ();
 sg13g2_fill_1 FILLER_4_183 ();
 sg13g2_fill_2 FILLER_4_193 ();
 sg13g2_fill_1 FILLER_4_195 ();
 sg13g2_decap_8 FILLER_4_214 ();
 sg13g2_fill_2 FILLER_4_221 ();
 sg13g2_fill_1 FILLER_4_223 ();
 sg13g2_decap_4 FILLER_4_242 ();
 sg13g2_fill_2 FILLER_4_246 ();
 sg13g2_decap_4 FILLER_4_260 ();
 sg13g2_decap_4 FILLER_4_282 ();
 sg13g2_fill_2 FILLER_4_286 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_fill_2 FILLER_4_303 ();
 sg13g2_decap_4 FILLER_4_335 ();
 sg13g2_fill_1 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_2 FILLER_5_130 ();
 sg13g2_fill_2 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_152 ();
 sg13g2_fill_2 FILLER_5_183 ();
 sg13g2_fill_2 FILLER_5_221 ();
 sg13g2_fill_1 FILLER_5_223 ();
 sg13g2_fill_2 FILLER_5_260 ();
 sg13g2_fill_1 FILLER_5_262 ();
 sg13g2_fill_2 FILLER_5_299 ();
 sg13g2_fill_1 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_fill_2 FILLER_6_112 ();
 sg13g2_fill_1 FILLER_6_114 ();
 sg13g2_fill_2 FILLER_6_141 ();
 sg13g2_fill_2 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_185 ();
 sg13g2_fill_2 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_261 ();
 sg13g2_fill_1 FILLER_6_299 ();
 sg13g2_fill_2 FILLER_6_336 ();
 sg13g2_fill_1 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_157 ();
 sg13g2_fill_1 FILLER_7_184 ();
 sg13g2_fill_2 FILLER_7_260 ();
 sg13g2_fill_1 FILLER_7_262 ();
 sg13g2_fill_2 FILLER_7_299 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_4 FILLER_8_98 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_fill_2 FILLER_8_184 ();
 sg13g2_fill_1 FILLER_8_186 ();
 sg13g2_fill_2 FILLER_8_246 ();
 sg13g2_fill_2 FILLER_8_336 ();
 sg13g2_fill_2 FILLER_8_343 ();
 sg13g2_fill_1 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_4 FILLER_9_91 ();
 sg13g2_fill_1 FILLER_9_95 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_4 FILLER_10_105 ();
 sg13g2_fill_2 FILLER_10_109 ();
 sg13g2_fill_1 FILLER_10_148 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_fill_1 FILLER_10_174 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_1 FILLER_10_223 ();
 sg13g2_fill_2 FILLER_10_251 ();
 sg13g2_fill_1 FILLER_10_253 ();
 sg13g2_fill_1 FILLER_10_292 ();
 sg13g2_fill_2 FILLER_10_325 ();
 sg13g2_fill_2 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_fill_2 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_300 ();
 sg13g2_fill_2 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_4 FILLER_12_91 ();
 sg13g2_fill_2 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_260 ();
 sg13g2_fill_2 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_4 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_102 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_fill_2 FILLER_14_134 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_fill_2 FILLER_14_190 ();
 sg13g2_fill_2 FILLER_14_202 ();
 sg13g2_fill_1 FILLER_14_204 ();
 sg13g2_fill_2 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_226 ();
 sg13g2_decap_4 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_fill_2 FILLER_14_261 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_188 ();
 sg13g2_fill_1 FILLER_15_202 ();
 sg13g2_decap_8 FILLER_15_220 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_234 ();
 sg13g2_fill_2 FILLER_15_241 ();
 sg13g2_decap_4 FILLER_15_256 ();
 sg13g2_fill_2 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_277 ();
 sg13g2_fill_1 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_4 FILLER_16_77 ();
 sg13g2_fill_1 FILLER_16_81 ();
 sg13g2_fill_1 FILLER_16_176 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_86 ();
 sg13g2_decap_4 FILLER_17_255 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_fill_2 FILLER_17_297 ();
 sg13g2_fill_1 FILLER_17_299 ();
 sg13g2_fill_1 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_4 FILLER_18_84 ();
 sg13g2_fill_1 FILLER_18_164 ();
 sg13g2_fill_2 FILLER_18_174 ();
 sg13g2_fill_2 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_218 ();
 sg13g2_decap_4 FILLER_18_255 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_fill_1 FILLER_19_164 ();
 sg13g2_fill_2 FILLER_19_215 ();
 sg13g2_decap_4 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_235 ();
 sg13g2_fill_2 FILLER_19_249 ();
 sg13g2_fill_2 FILLER_19_269 ();
 sg13g2_decap_4 FILLER_19_311 ();
 sg13g2_fill_2 FILLER_19_350 ();
 sg13g2_fill_2 FILLER_19_357 ();
 sg13g2_fill_1 FILLER_19_359 ();
 sg13g2_fill_1 FILLER_19_398 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_4 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_113 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_209 ();
 sg13g2_fill_2 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_399 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_decap_4 FILLER_21_203 ();
 sg13g2_decap_4 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_4 FILLER_21_302 ();
 sg13g2_fill_2 FILLER_21_342 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_fill_1 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_96 ();
 sg13g2_fill_1 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_2 FILLER_23_128 ();
 sg13g2_fill_2 FILLER_23_178 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_272 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_fill_1 FILLER_23_400 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_95 ();
 sg13g2_fill_2 FILLER_24_216 ();
 sg13g2_fill_2 FILLER_24_254 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_decap_4 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_fill_2 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_165 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_2 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_310 ();
 sg13g2_fill_2 FILLER_25_348 ();
 sg13g2_fill_2 FILLER_25_369 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_1 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_fill_2 FILLER_27_353 ();
 sg13g2_fill_1 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_2 FILLER_28_350 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_4 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_fill_2 FILLER_29_350 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_168 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_138 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_155 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_100 ();
 sg13g2_fill_1 FILLER_32_157 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_fill_1 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_359 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_fill_1 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_167 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_277 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_fill_1 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_177 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_fill_2 FILLER_35_395 ();
 sg13g2_fill_1 FILLER_35_397 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_fill_2 FILLER_36_194 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_356 ();
 sg13g2_fill_1 FILLER_36_358 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_4 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_88 ();
 sg13g2_fill_1 FILLER_37_157 ();
 sg13g2_fill_1 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_392 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_fill_1 FILLER_38_261 ();
 sg13g2_fill_2 FILLER_38_346 ();
 sg13g2_fill_1 FILLER_38_348 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net5;
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
 assign uo_out[2] = net21;
 assign uo_out[3] = net22;
 assign uo_out[4] = net23;
 assign uo_out[5] = net24;
 assign uo_out[6] = net25;
 assign uo_out[7] = net26;
endmodule

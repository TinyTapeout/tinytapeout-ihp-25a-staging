module tt_um_rte_sine_synth (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire \delta[0] ;
 wire \delta[1] ;
 wire \delta[2] ;
 wire \delta[3] ;
 wire \event_count[0] ;
 wire \event_count[1] ;
 wire \event_count[2] ;
 wire \event_count[3] ;
 wire \event_count[4] ;
 wire \event_count[5] ;
 wire \event_count[6] ;
 wire \event_count[7] ;
 wire \event_count[8] ;
 wire \last_input[0] ;
 wire \last_input[1] ;
 wire \last_input[2] ;
 wire \last_input[3] ;
 wire \last_input[4] ;
 wire \last_input[5] ;
 wire \last_input[6] ;
 wire \last_input[7] ;
 wire \new_input[0] ;
 wire \new_input[1] ;
 wire \new_input[2] ;
 wire \new_input[3] ;
 wire \new_input[4] ;
 wire \new_input[5] ;
 wire \new_input[6] ;
 wire \new_input[7] ;
 wire \next_limit[0] ;
 wire \next_limit[1] ;
 wire \next_limit[2] ;
 wire \next_limit[3] ;
 wire \next_limit[4] ;
 wire \next_limit[5] ;
 wire \next_limit[6] ;
 wire \next_limit[7] ;
 wire \next_limit[8] ;
 wire \out_val[0] ;
 wire \out_val[1] ;
 wire \out_val[2] ;
 wire \out_val[3] ;
 wire \out_val[4] ;
 wire \out_val[5] ;
 wire \out_val[6] ;
 wire \out_val[7] ;
 wire \out_val[8] ;
 wire \out_val[9] ;
 wire \phase_check[0] ;
 wire \phase_check[1] ;
 wire \phase_check[2] ;
 wire \phase_check[3] ;
 wire \phase_check[4] ;
 wire \phase_check[5] ;
 wire \phase_count[0] ;
 wire \phase_count[1] ;
 wire \phase_count[2] ;
 wire \phase_count[3] ;
 wire \phase_count[4] ;
 wire \phase_count[5] ;
 wire \phase_limit[0] ;
 wire \phase_limit[1] ;
 wire \phase_limit[2] ;
 wire \phase_limit[3] ;
 wire \phase_limit[4] ;
 wire \phase_limit[5] ;
 wire \phase_limit[6] ;
 wire \phase_limit[7] ;
 wire \phase_limit[8] ;
 wire \pwm.count[0] ;
 wire \pwm.count[1] ;
 wire \pwm.count[2] ;
 wire \pwm.count[3] ;
 wire \pwm.count[4] ;
 wire \pwm.count[5] ;
 wire \pwm.count[6] ;
 wire \pwm.count[7] ;
 wire \pwm.count[8] ;
 wire \pwm.count[9] ;
 wire \pwm.pwm ;
 wire \qtr_count[0] ;
 wire \qtr_count[1] ;
 wire rst_n_i;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;

 sg13g2_inv_1 _405_ (.Y(_079_),
    .A(net132));
 sg13g2_inv_1 _406_ (.Y(_080_),
    .A(\pwm.count[0] ));
 sg13g2_inv_1 _407_ (.Y(_081_),
    .A(\pwm.count[7] ));
 sg13g2_inv_1 _408_ (.Y(_082_),
    .A(\pwm.count[6] ));
 sg13g2_inv_1 _409_ (.Y(_083_),
    .A(\pwm.count[8] ));
 sg13g2_inv_2 _410_ (.Y(_084_),
    .A(net170));
 sg13g2_inv_1 _411_ (.Y(_085_),
    .A(net168));
 sg13g2_inv_1 _412_ (.Y(_086_),
    .A(net126));
 sg13g2_inv_1 _413_ (.Y(_087_),
    .A(net120));
 sg13g2_inv_1 _414_ (.Y(_088_),
    .A(\out_val[8] ));
 sg13g2_inv_1 _415_ (.Y(_089_),
    .A(\out_val[7] ));
 sg13g2_inv_1 _416_ (.Y(_090_),
    .A(\out_val[4] ));
 sg13g2_inv_1 _417_ (.Y(_091_),
    .A(\out_val[3] ));
 sg13g2_inv_1 _418_ (.Y(_092_),
    .A(net160));
 sg13g2_inv_1 _419_ (.Y(_093_),
    .A(\delta[3] ));
 sg13g2_inv_1 _420_ (.Y(_094_),
    .A(net65));
 sg13g2_inv_1 _421_ (.Y(_095_),
    .A(net90));
 sg13g2_inv_1 _422_ (.Y(_096_),
    .A(net111));
 sg13g2_inv_1 _423_ (.Y(_097_),
    .A(net94));
 sg13g2_nor2_2 _424_ (.A(\event_count[1] ),
    .B(net97),
    .Y(_098_));
 sg13g2_or2_1 _425_ (.X(_099_),
    .B(net97),
    .A(\event_count[1] ));
 sg13g2_or3_1 _426_ (.A(\event_count[5] ),
    .B(\event_count[4] ),
    .C(\event_count[6] ),
    .X(_100_));
 sg13g2_nor3_1 _427_ (.A(\event_count[3] ),
    .B(\event_count[7] ),
    .C(_100_),
    .Y(_101_));
 sg13g2_nor4_2 _428_ (.A(net106),
    .B(net114),
    .C(net116),
    .Y(_102_),
    .D(_100_));
 sg13g2_nand2_1 _429_ (.Y(_103_),
    .A(_098_),
    .B(_102_));
 sg13g2_nand2_1 _430_ (.Y(_104_),
    .A(_009_),
    .B(net100));
 sg13g2_o21ai_1 _431_ (.B1(_104_),
    .Y(_105_),
    .A1(net132),
    .A2(_009_));
 sg13g2_nor2_1 _432_ (.A(_103_),
    .B(_105_),
    .Y(_106_));
 sg13g2_a21oi_1 _433_ (.A1(_079_),
    .A2(_103_),
    .Y(_008_),
    .B1(_106_));
 sg13g2_nand3_1 _434_ (.B(_098_),
    .C(_102_),
    .A(_009_),
    .Y(_107_));
 sg13g2_mux2_1 _435_ (.A0(\phase_limit[0] ),
    .A1(net45),
    .S(net72),
    .X(_000_));
 sg13g2_nand2_1 _436_ (.Y(_108_),
    .A(\event_count[1] ),
    .B(net97));
 sg13g2_nor2_1 _437_ (.A(net93),
    .B(_107_),
    .Y(_109_));
 sg13g2_a21oi_1 _438_ (.A1(_099_),
    .A2(net98),
    .Y(_001_),
    .B1(_109_));
 sg13g2_xnor2_1 _439_ (.Y(_110_),
    .A(net114),
    .B(_098_));
 sg13g2_nor2_1 _440_ (.A(net87),
    .B(net72),
    .Y(_111_));
 sg13g2_nor2_1 _441_ (.A(net115),
    .B(_111_),
    .Y(_002_));
 sg13g2_nor2_1 _442_ (.A(net104),
    .B(net72),
    .Y(_112_));
 sg13g2_or3_2 _443_ (.A(net106),
    .B(\event_count[2] ),
    .C(_099_),
    .X(_113_));
 sg13g2_o21ai_1 _444_ (.B1(net106),
    .Y(_114_),
    .A1(\event_count[2] ),
    .A2(_099_));
 sg13g2_a21oi_1 _445_ (.A1(_113_),
    .A2(net107),
    .Y(_003_),
    .B1(_112_));
 sg13g2_xnor2_1 _446_ (.Y(_115_),
    .A(net156),
    .B(_113_));
 sg13g2_o21ai_1 _447_ (.B1(_115_),
    .Y(_116_),
    .A1(net103),
    .A2(net72));
 sg13g2_inv_1 _448_ (.Y(_004_),
    .A(_116_));
 sg13g2_nor3_1 _449_ (.A(net143),
    .B(\event_count[4] ),
    .C(_113_),
    .Y(_117_));
 sg13g2_o21ai_1 _450_ (.B1(net143),
    .Y(_118_),
    .A1(\event_count[4] ),
    .A2(_113_));
 sg13g2_nand2b_1 _451_ (.Y(_119_),
    .B(net144),
    .A_N(_117_));
 sg13g2_o21ai_1 _452_ (.B1(net145),
    .Y(_120_),
    .A1(net113),
    .A2(net72));
 sg13g2_inv_1 _453_ (.Y(_005_),
    .A(_120_));
 sg13g2_xor2_1 _454_ (.B(_117_),
    .A(net137),
    .X(_121_));
 sg13g2_o21ai_1 _455_ (.B1(net138),
    .Y(_122_),
    .A1(net61),
    .A2(net72));
 sg13g2_inv_1 _456_ (.Y(_006_),
    .A(_122_));
 sg13g2_o21ai_1 _457_ (.B1(net116),
    .Y(_123_),
    .A1(_100_),
    .A2(_113_));
 sg13g2_nor2b_1 _458_ (.A(\phase_limit[7] ),
    .B_N(_009_),
    .Y(_124_));
 sg13g2_o21ai_1 _459_ (.B1(net117),
    .Y(_007_),
    .A1(_103_),
    .A2(_124_));
 sg13g2_nand3_1 _460_ (.B(net157),
    .C(net123),
    .A(net176),
    .Y(_125_));
 sg13g2_and4_1 _461_ (.A(\pwm.count[1] ),
    .B(\pwm.count[2] ),
    .C(\pwm.count[7] ),
    .D(\pwm.count[8] ),
    .X(_126_));
 sg13g2_nand4_1 _462_ (.B(\pwm.count[6] ),
    .C(\pwm.count[9] ),
    .A(_080_),
    .Y(_127_),
    .D(_126_));
 sg13g2_o21ai_1 _463_ (.B1(net81),
    .Y(_128_),
    .A1(_125_),
    .A2(_127_));
 sg13g2_inv_1 _464_ (.Y(_129_),
    .A(_128_));
 sg13g2_and2_1 _465_ (.A(net42),
    .B(_129_),
    .X(_022_));
 sg13g2_o21ai_1 _466_ (.B1(_129_),
    .Y(_130_),
    .A1(net146),
    .A2(\pwm.count[1] ));
 sg13g2_a21oi_1 _467_ (.A1(net146),
    .A2(\pwm.count[1] ),
    .Y(_023_),
    .B1(_130_));
 sg13g2_and3_2 _468_ (.X(_131_),
    .A(net146),
    .B(\pwm.count[1] ),
    .C(net134));
 sg13g2_a21oi_1 _469_ (.A1(\pwm.count[0] ),
    .A2(\pwm.count[1] ),
    .Y(_132_),
    .B1(net134));
 sg13g2_nor3_1 _470_ (.A(_128_),
    .B(_131_),
    .C(net135),
    .Y(_024_));
 sg13g2_o21ai_1 _471_ (.B1(_129_),
    .Y(_133_),
    .A1(net165),
    .A2(_131_));
 sg13g2_a21oi_1 _472_ (.A1(net165),
    .A2(_131_),
    .Y(_025_),
    .B1(_133_));
 sg13g2_and3_1 _473_ (.X(_134_),
    .A(\pwm.count[3] ),
    .B(net123),
    .C(_131_));
 sg13g2_a21oi_1 _474_ (.A1(\pwm.count[3] ),
    .A2(_131_),
    .Y(_135_),
    .B1(net123));
 sg13g2_nor3_1 _475_ (.A(_128_),
    .B(_134_),
    .C(net124),
    .Y(_026_));
 sg13g2_nor2_1 _476_ (.A(net157),
    .B(_134_),
    .Y(_136_));
 sg13g2_nor2b_1 _477_ (.A(_125_),
    .B_N(_131_),
    .Y(_137_));
 sg13g2_nor3_1 _478_ (.A(_128_),
    .B(net158),
    .C(_137_),
    .Y(_027_));
 sg13g2_nor2_1 _479_ (.A(net154),
    .B(_137_),
    .Y(_138_));
 sg13g2_and2_1 _480_ (.A(net154),
    .B(_137_),
    .X(_139_));
 sg13g2_nor3_1 _481_ (.A(_128_),
    .B(net155),
    .C(_139_),
    .Y(_028_));
 sg13g2_nor2_1 _482_ (.A(net164),
    .B(_139_),
    .Y(_140_));
 sg13g2_and2_1 _483_ (.A(net164),
    .B(_139_),
    .X(_141_));
 sg13g2_nor3_1 _484_ (.A(_128_),
    .B(_140_),
    .C(_141_),
    .Y(_029_));
 sg13g2_and2_1 _485_ (.A(net172),
    .B(_141_),
    .X(_142_));
 sg13g2_o21ai_1 _486_ (.B1(_129_),
    .Y(_143_),
    .A1(net172),
    .A2(_141_));
 sg13g2_nor2_1 _487_ (.A(_142_),
    .B(_143_),
    .Y(_030_));
 sg13g2_o21ai_1 _488_ (.B1(_129_),
    .Y(_144_),
    .A1(net130),
    .A2(_142_));
 sg13g2_a21oi_1 _489_ (.A1(net130),
    .A2(_142_),
    .Y(_031_),
    .B1(_144_));
 sg13g2_nand4_1 _490_ (.B(_079_),
    .C(_098_),
    .A(\event_count[2] ),
    .Y(_145_),
    .D(_101_));
 sg13g2_nand2_1 _491_ (.Y(_146_),
    .A(net141),
    .B(net71));
 sg13g2_xnor2_1 _492_ (.Y(_147_),
    .A(net120),
    .B(\qtr_count[0] ));
 sg13g2_o21ai_1 _493_ (.B1(_146_),
    .Y(_032_),
    .A1(net71),
    .A2(_147_));
 sg13g2_nand2_1 _494_ (.Y(_148_),
    .A(net128),
    .B(net71));
 sg13g2_xnor2_1 _495_ (.Y(_149_),
    .A(\phase_count[1] ),
    .B(\qtr_count[0] ));
 sg13g2_o21ai_1 _496_ (.B1(_148_),
    .Y(_033_),
    .A1(net70),
    .A2(_149_));
 sg13g2_nand2_1 _497_ (.Y(_150_),
    .A(net162),
    .B(net71));
 sg13g2_xnor2_1 _498_ (.Y(_151_),
    .A(\phase_count[2] ),
    .B(net79));
 sg13g2_o21ai_1 _499_ (.B1(_150_),
    .Y(_034_),
    .A1(net70),
    .A2(_151_));
 sg13g2_nand2_1 _500_ (.Y(_152_),
    .A(net150),
    .B(net70));
 sg13g2_xnor2_1 _501_ (.Y(_153_),
    .A(net126),
    .B(net79));
 sg13g2_o21ai_1 _502_ (.B1(_152_),
    .Y(_035_),
    .A1(net70),
    .A2(_153_));
 sg13g2_xor2_1 _503_ (.B(net79),
    .A(net152),
    .X(_154_));
 sg13g2_nor2_1 _504_ (.A(net70),
    .B(_154_),
    .Y(_155_));
 sg13g2_a21oi_1 _505_ (.A1(_085_),
    .A2(net70),
    .Y(_036_),
    .B1(_155_));
 sg13g2_xor2_1 _506_ (.B(net79),
    .A(net166),
    .X(_156_));
 sg13g2_nor2_1 _507_ (.A(net70),
    .B(_156_),
    .Y(_157_));
 sg13g2_a21oi_1 _508_ (.A1(_084_),
    .A2(net70),
    .Y(_037_),
    .B1(_157_));
 sg13g2_nor2_1 _509_ (.A(\event_count[0] ),
    .B(net132),
    .Y(_158_));
 sg13g2_nand3_1 _510_ (.B(_102_),
    .C(_158_),
    .A(\event_count[1] ),
    .Y(_159_));
 sg13g2_nand2_1 _511_ (.Y(_160_),
    .A(\out_val[0] ),
    .B(\delta[0] ));
 sg13g2_xor2_1 _512_ (.B(\delta[0] ),
    .A(\out_val[0] ),
    .X(_161_));
 sg13g2_nand2_1 _513_ (.Y(_162_),
    .A(net51),
    .B(net68));
 sg13g2_o21ai_1 _514_ (.B1(_162_),
    .Y(_038_),
    .A1(net68),
    .A2(_161_));
 sg13g2_xor2_1 _515_ (.B(\qtr_count[1] ),
    .A(net79),
    .X(_163_));
 sg13g2_xnor2_1 _516_ (.Y(_164_),
    .A(net79),
    .B(\qtr_count[1] ));
 sg13g2_or2_1 _517_ (.X(_165_),
    .B(\delta[0] ),
    .A(\delta[1] ));
 sg13g2_nand2_1 _518_ (.Y(_166_),
    .A(\delta[1] ),
    .B(\delta[0] ));
 sg13g2_nand2_1 _519_ (.Y(_167_),
    .A(_011_),
    .B(_164_));
 sg13g2_a21o_1 _520_ (.A2(_166_),
    .A1(_165_),
    .B1(_164_),
    .X(_168_));
 sg13g2_and3_1 _521_ (.X(_169_),
    .A(\out_val[1] ),
    .B(_167_),
    .C(_168_));
 sg13g2_nand3_1 _522_ (.B(_167_),
    .C(_168_),
    .A(\out_val[1] ),
    .Y(_170_));
 sg13g2_a21oi_1 _523_ (.A1(_167_),
    .A2(_168_),
    .Y(_171_),
    .B1(\out_val[1] ));
 sg13g2_nor2_1 _524_ (.A(_169_),
    .B(_171_),
    .Y(_172_));
 sg13g2_xnor2_1 _525_ (.Y(_173_),
    .A(_160_),
    .B(_172_));
 sg13g2_nor2_1 _526_ (.A(net68),
    .B(_173_),
    .Y(_174_));
 sg13g2_a21oi_1 _527_ (.A1(_092_),
    .A2(net68),
    .Y(_039_),
    .B1(_174_));
 sg13g2_o21ai_1 _528_ (.B1(_170_),
    .Y(_175_),
    .A1(_160_),
    .A2(_171_));
 sg13g2_a21o_1 _529_ (.A2(_165_),
    .A1(_163_),
    .B1(\delta[2] ),
    .X(_176_));
 sg13g2_nand3_1 _530_ (.B(_163_),
    .C(_165_),
    .A(\delta[2] ),
    .Y(_177_));
 sg13g2_and3_1 _531_ (.X(_178_),
    .A(\out_val[2] ),
    .B(_176_),
    .C(_177_));
 sg13g2_nand3_1 _532_ (.B(_176_),
    .C(_177_),
    .A(\out_val[2] ),
    .Y(_179_));
 sg13g2_a21oi_1 _533_ (.A1(_176_),
    .A2(_177_),
    .Y(_180_),
    .B1(\out_val[2] ));
 sg13g2_nor2_1 _534_ (.A(_178_),
    .B(_180_),
    .Y(_181_));
 sg13g2_xnor2_1 _535_ (.Y(_182_),
    .A(_175_),
    .B(_181_));
 sg13g2_nand2_1 _536_ (.Y(_183_),
    .A(net148),
    .B(_159_));
 sg13g2_o21ai_1 _537_ (.B1(_183_),
    .Y(_040_),
    .A1(_159_),
    .A2(_182_));
 sg13g2_nor3_1 _538_ (.A(\delta[1] ),
    .B(\delta[0] ),
    .C(\delta[2] ),
    .Y(_184_));
 sg13g2_o21ai_1 _539_ (.B1(_093_),
    .Y(_185_),
    .A1(_164_),
    .A2(_184_));
 sg13g2_nand3b_1 _540_ (.B(_163_),
    .C(\delta[3] ),
    .Y(_186_),
    .A_N(_184_));
 sg13g2_and3_1 _541_ (.X(_187_),
    .A(\out_val[3] ),
    .B(_185_),
    .C(_186_));
 sg13g2_nand3_1 _542_ (.B(_185_),
    .C(_186_),
    .A(\out_val[3] ),
    .Y(_188_));
 sg13g2_a21oi_1 _543_ (.A1(_185_),
    .A2(_186_),
    .Y(_189_),
    .B1(\out_val[3] ));
 sg13g2_nor2_1 _544_ (.A(_187_),
    .B(_189_),
    .Y(_190_));
 sg13g2_a21oi_1 _545_ (.A1(_175_),
    .A2(_181_),
    .Y(_191_),
    .B1(_178_));
 sg13g2_xor2_1 _546_ (.B(_191_),
    .A(_190_),
    .X(_192_));
 sg13g2_mux2_1 _547_ (.A0(_192_),
    .A1(net96),
    .S(_159_),
    .X(_041_));
 sg13g2_nor4_1 _548_ (.A(_178_),
    .B(_180_),
    .C(_187_),
    .D(_189_),
    .Y(_193_));
 sg13g2_a21oi_1 _549_ (.A1(_179_),
    .A2(_188_),
    .Y(_194_),
    .B1(_189_));
 sg13g2_a21oi_2 _550_ (.B1(_194_),
    .Y(_195_),
    .A2(_193_),
    .A1(_175_));
 sg13g2_a21oi_1 _551_ (.A1(_093_),
    .A2(_184_),
    .Y(_196_),
    .B1(_164_));
 sg13g2_xnor2_1 _552_ (.Y(_197_),
    .A(_090_),
    .B(net74));
 sg13g2_nor2b_1 _553_ (.A(_195_),
    .B_N(_197_),
    .Y(_198_));
 sg13g2_nand2_1 _554_ (.Y(_199_),
    .A(net55),
    .B(net69));
 sg13g2_xnor2_1 _555_ (.Y(_200_),
    .A(_195_),
    .B(_197_));
 sg13g2_o21ai_1 _556_ (.B1(_199_),
    .Y(_042_),
    .A1(net69),
    .A2(_200_));
 sg13g2_xor2_1 _557_ (.B(net74),
    .A(\out_val[5] ),
    .X(_201_));
 sg13g2_a21oi_1 _558_ (.A1(\out_val[4] ),
    .A2(net73),
    .Y(_202_),
    .B1(_198_));
 sg13g2_xor2_1 _559_ (.B(_202_),
    .A(_201_),
    .X(_203_));
 sg13g2_mux2_1 _560_ (.A0(_203_),
    .A1(net101),
    .S(net69),
    .X(_043_));
 sg13g2_nand2_1 _561_ (.Y(_204_),
    .A(net47),
    .B(net69));
 sg13g2_and2_1 _562_ (.A(\out_val[6] ),
    .B(net74),
    .X(_205_));
 sg13g2_xor2_1 _563_ (.B(net74),
    .A(\out_val[6] ),
    .X(_206_));
 sg13g2_o21ai_1 _564_ (.B1(net73),
    .Y(_207_),
    .A1(\out_val[5] ),
    .A2(\out_val[4] ));
 sg13g2_nand2_1 _565_ (.Y(_208_),
    .A(_197_),
    .B(_201_));
 sg13g2_o21ai_1 _566_ (.B1(_207_),
    .Y(_209_),
    .A1(_195_),
    .A2(_208_));
 sg13g2_xor2_1 _567_ (.B(_209_),
    .A(_206_),
    .X(_210_));
 sg13g2_o21ai_1 _568_ (.B1(_204_),
    .Y(_044_),
    .A1(net69),
    .A2(_210_));
 sg13g2_xnor2_1 _569_ (.Y(_211_),
    .A(_089_),
    .B(net73));
 sg13g2_a21oi_1 _570_ (.A1(_206_),
    .A2(_209_),
    .Y(_212_),
    .B1(_205_));
 sg13g2_xnor2_1 _571_ (.Y(_213_),
    .A(_211_),
    .B(_212_));
 sg13g2_nand2_1 _572_ (.Y(_214_),
    .A(net48),
    .B(net68));
 sg13g2_o21ai_1 _573_ (.B1(_214_),
    .Y(_045_),
    .A1(net69),
    .A2(_213_));
 sg13g2_nand2_1 _574_ (.Y(_215_),
    .A(net53),
    .B(net68));
 sg13g2_nand2b_1 _575_ (.Y(_216_),
    .B(_088_),
    .A_N(net73));
 sg13g2_and2_1 _576_ (.A(\out_val[8] ),
    .B(net73),
    .X(_217_));
 sg13g2_xnor2_1 _577_ (.Y(_218_),
    .A(\out_val[8] ),
    .B(net73));
 sg13g2_nand4_1 _578_ (.B(_201_),
    .C(_206_),
    .A(_197_),
    .Y(_219_),
    .D(_211_));
 sg13g2_o21ai_1 _579_ (.B1(net73),
    .Y(_220_),
    .A1(\out_val[7] ),
    .A2(\out_val[6] ));
 sg13g2_and2_1 _580_ (.A(_207_),
    .B(_220_),
    .X(_221_));
 sg13g2_o21ai_1 _581_ (.B1(_221_),
    .Y(_222_),
    .A1(_195_),
    .A2(_219_));
 sg13g2_xnor2_1 _582_ (.Y(_223_),
    .A(_218_),
    .B(_222_));
 sg13g2_o21ai_1 _583_ (.B1(_215_),
    .Y(_046_),
    .A1(net69),
    .A2(_223_));
 sg13g2_a21oi_1 _584_ (.A1(_216_),
    .A2(_222_),
    .Y(_224_),
    .B1(_217_));
 sg13g2_xnor2_1 _585_ (.Y(_225_),
    .A(net119),
    .B(net73));
 sg13g2_xnor2_1 _586_ (.Y(_226_),
    .A(_224_),
    .B(_225_));
 sg13g2_nand2_1 _587_ (.Y(_227_),
    .A(net119),
    .B(net68));
 sg13g2_o21ai_1 _588_ (.B1(_227_),
    .Y(_047_),
    .A1(net68),
    .A2(_226_));
 sg13g2_nand2b_1 _589_ (.Y(_228_),
    .B(net38),
    .A_N(\last_input[0] ));
 sg13g2_nand2b_1 _590_ (.Y(_229_),
    .B(net39),
    .A_N(\last_input[1] ));
 sg13g2_and2_2 _591_ (.A(_228_),
    .B(_229_),
    .X(_230_));
 sg13g2_inv_1 _592_ (.Y(_231_),
    .A(_230_));
 sg13g2_nor2b_1 _593_ (.A(\last_input[2] ),
    .B_N(\new_input[2] ),
    .Y(_232_));
 sg13g2_nand2b_2 _594_ (.Y(_233_),
    .B(net44),
    .A_N(\last_input[2] ));
 sg13g2_nand2b_2 _595_ (.Y(_234_),
    .B(net40),
    .A_N(\last_input[3] ));
 sg13g2_nand2_1 _596_ (.Y(_235_),
    .A(_233_),
    .B(_234_));
 sg13g2_o21ai_1 _597_ (.B1(net77),
    .Y(_236_),
    .A1(_231_),
    .A2(_235_));
 sg13g2_nor4_1 _598_ (.A(\new_input[4] ),
    .B(\new_input[5] ),
    .C(\new_input[6] ),
    .D(\new_input[7] ),
    .Y(_237_));
 sg13g2_nor4_1 _599_ (.A(\new_input[0] ),
    .B(\new_input[1] ),
    .C(\new_input[2] ),
    .D(\new_input[3] ),
    .Y(_238_));
 sg13g2_nor2b_1 _600_ (.A(\last_input[4] ),
    .B_N(\new_input[4] ),
    .Y(_239_));
 sg13g2_nand2b_1 _601_ (.Y(_240_),
    .B(net43),
    .A_N(\last_input[4] ));
 sg13g2_nand2b_1 _602_ (.Y(_241_),
    .B(\new_input[5] ),
    .A_N(\last_input[5] ));
 sg13g2_nand2b_1 _603_ (.Y(_242_),
    .B(\new_input[6] ),
    .A_N(\last_input[6] ));
 sg13g2_nand2_1 _604_ (.Y(_243_),
    .A(_241_),
    .B(_242_));
 sg13g2_nor2b_2 _605_ (.A(\last_input[7] ),
    .B_N(net37),
    .Y(_244_));
 sg13g2_nor3_1 _606_ (.A(_239_),
    .B(_243_),
    .C(_244_),
    .Y(_245_));
 sg13g2_nand4_1 _607_ (.B(_233_),
    .C(_234_),
    .A(_230_),
    .Y(_246_),
    .D(_245_));
 sg13g2_a21oi_1 _608_ (.A1(_237_),
    .A2(_238_),
    .Y(_247_),
    .B1(_246_));
 sg13g2_nor2b_2 _609_ (.A(_247_),
    .B_N(net76),
    .Y(_248_));
 sg13g2_inv_1 _610_ (.Y(_249_),
    .A(_248_));
 sg13g2_nand2_1 _611_ (.Y(_250_),
    .A(_240_),
    .B(_243_));
 sg13g2_o21ai_1 _612_ (.B1(_234_),
    .Y(_251_),
    .A1(_239_),
    .A2(_244_));
 sg13g2_nand2b_1 _613_ (.Y(_252_),
    .B(_250_),
    .A_N(_251_));
 sg13g2_o21ai_1 _614_ (.B1(_230_),
    .Y(_253_),
    .A1(_232_),
    .A2(_252_));
 sg13g2_mux2_1 _615_ (.A0(net88),
    .A1(_253_),
    .S(_248_),
    .X(_048_));
 sg13g2_nand2_1 _616_ (.Y(_254_),
    .A(net56),
    .B(_249_));
 sg13g2_nand4_1 _617_ (.B(_230_),
    .C(_233_),
    .A(net76),
    .Y(_255_),
    .D(_234_));
 sg13g2_o21ai_1 _618_ (.B1(_240_),
    .Y(_256_),
    .A1(_243_),
    .A2(_244_));
 sg13g2_o21ai_1 _619_ (.B1(_254_),
    .Y(_049_),
    .A1(_255_),
    .A2(_256_));
 sg13g2_o21ai_1 _620_ (.B1(_230_),
    .Y(_257_),
    .A1(_235_),
    .A2(_250_));
 sg13g2_mux2_1 _621_ (.A0(net62),
    .A1(_257_),
    .S(_248_),
    .X(_050_));
 sg13g2_nand2_1 _622_ (.Y(_258_),
    .A(_242_),
    .B(_244_));
 sg13g2_nand4_1 _623_ (.B(_240_),
    .C(_241_),
    .A(_234_),
    .Y(_259_),
    .D(_258_));
 sg13g2_nand2_1 _624_ (.Y(_260_),
    .A(_229_),
    .B(_233_));
 sg13g2_and2_1 _625_ (.A(_228_),
    .B(_248_),
    .X(_261_));
 sg13g2_o21ai_1 _626_ (.B1(_261_),
    .Y(_262_),
    .A1(_259_),
    .A2(_260_));
 sg13g2_o21ai_1 _627_ (.B1(_262_),
    .Y(_051_),
    .A1(_094_),
    .A2(_248_));
 sg13g2_nand2b_1 _628_ (.Y(_263_),
    .B(_259_),
    .A_N(_260_));
 sg13g2_a22oi_1 _629_ (.Y(_052_),
    .B1(_261_),
    .B2(_263_),
    .A2(_249_),
    .A1(_095_));
 sg13g2_nand2_1 _630_ (.Y(_264_),
    .A(_233_),
    .B(_252_));
 sg13g2_nand2_1 _631_ (.Y(_265_),
    .A(_229_),
    .B(_264_));
 sg13g2_a22oi_1 _632_ (.Y(_053_),
    .B1(_261_),
    .B2(_265_),
    .A2(_249_),
    .A1(_096_));
 sg13g2_nor2_1 _633_ (.A(_239_),
    .B(_243_),
    .Y(_266_));
 sg13g2_o21ai_1 _634_ (.B1(_230_),
    .Y(_267_),
    .A1(_235_),
    .A2(_266_));
 sg13g2_mux2_1 _635_ (.A0(net60),
    .A1(_267_),
    .S(_248_),
    .X(_054_));
 sg13g2_nand2_1 _636_ (.Y(_268_),
    .A(net58),
    .B(_249_));
 sg13g2_o21ai_1 _637_ (.B1(_268_),
    .Y(_055_),
    .A1(_245_),
    .A2(_255_));
 sg13g2_o21ai_1 _638_ (.B1(_236_),
    .Y(_056_),
    .A1(_097_),
    .A2(_248_));
 sg13g2_nor2_1 _639_ (.A(_087_),
    .B(net72),
    .Y(_269_));
 sg13g2_nand3_1 _640_ (.B(net136),
    .C(_269_),
    .A(net174),
    .Y(_270_));
 sg13g2_nor2_2 _641_ (.A(_086_),
    .B(_270_),
    .Y(_271_));
 sg13g2_nand3_1 _642_ (.B(net152),
    .C(_271_),
    .A(net166),
    .Y(_272_));
 sg13g2_and4_1 _643_ (.A(\phase_count[5] ),
    .B(\phase_count[4] ),
    .C(net79),
    .D(_271_),
    .X(_273_));
 sg13g2_xnor2_1 _644_ (.Y(_057_),
    .A(net79),
    .B(_272_));
 sg13g2_nand2_1 _645_ (.Y(_274_),
    .A(\qtr_count[1] ),
    .B(_273_));
 sg13g2_xor2_1 _646_ (.B(_273_),
    .A(net139),
    .X(_058_));
 sg13g2_xnor2_1 _647_ (.Y(_059_),
    .A(net120),
    .B(net72));
 sg13g2_xor2_1 _648_ (.B(_269_),
    .A(net136),
    .X(_060_));
 sg13g2_a21o_1 _649_ (.A2(_269_),
    .A1(net136),
    .B1(net174),
    .X(_275_));
 sg13g2_and2_1 _650_ (.A(_270_),
    .B(_275_),
    .X(_061_));
 sg13g2_xnor2_1 _651_ (.Y(_062_),
    .A(net126),
    .B(_270_));
 sg13g2_xor2_1 _652_ (.B(_271_),
    .A(net152),
    .X(_063_));
 sg13g2_a21o_1 _653_ (.A2(_271_),
    .A1(net152),
    .B1(net166),
    .X(_276_));
 sg13g2_and2_1 _654_ (.A(_272_),
    .B(_276_),
    .X(_064_));
 sg13g2_nand2b_1 _655_ (.Y(_277_),
    .B(net63),
    .A_N(net81));
 sg13g2_nand2b_1 _656_ (.Y(_278_),
    .B(\pwm.count[2] ),
    .A_N(\out_val[2] ));
 sg13g2_nand2b_1 _657_ (.Y(_279_),
    .B(\pwm.count[9] ),
    .A_N(\out_val[9] ));
 sg13g2_nand2b_1 _658_ (.Y(_280_),
    .B(\out_val[0] ),
    .A_N(\pwm.count[0] ));
 sg13g2_nor2b_1 _659_ (.A(\out_val[0] ),
    .B_N(\pwm.count[0] ),
    .Y(_281_));
 sg13g2_a221oi_1 _660_ (.B2(_280_),
    .C1(_281_),
    .B1(_279_),
    .A1(\pwm.count[1] ),
    .Y(_282_),
    .A2(_092_));
 sg13g2_nand2b_1 _661_ (.Y(_283_),
    .B(\out_val[2] ),
    .A_N(\pwm.count[2] ));
 sg13g2_o21ai_1 _662_ (.B1(_283_),
    .Y(_284_),
    .A1(\pwm.count[1] ),
    .A2(_092_));
 sg13g2_o21ai_1 _663_ (.B1(_278_),
    .Y(_285_),
    .A1(_282_),
    .A2(_284_));
 sg13g2_o21ai_1 _664_ (.B1(_285_),
    .Y(_286_),
    .A1(\pwm.count[3] ),
    .A2(_091_));
 sg13g2_a22oi_1 _665_ (.Y(_287_),
    .B1(_091_),
    .B2(\pwm.count[3] ),
    .A2(_090_),
    .A1(\pwm.count[4] ));
 sg13g2_nand2b_1 _666_ (.Y(_288_),
    .B(\out_val[5] ),
    .A_N(\pwm.count[5] ));
 sg13g2_o21ai_1 _667_ (.B1(_288_),
    .Y(_289_),
    .A1(\pwm.count[4] ),
    .A2(_090_));
 sg13g2_a21oi_1 _668_ (.A1(_286_),
    .A2(_287_),
    .Y(_290_),
    .B1(_289_));
 sg13g2_nand2b_1 _669_ (.Y(_291_),
    .B(\pwm.count[5] ),
    .A_N(\out_val[5] ));
 sg13g2_o21ai_1 _670_ (.B1(_291_),
    .Y(_292_),
    .A1(_082_),
    .A2(\out_val[6] ));
 sg13g2_a22oi_1 _671_ (.Y(_293_),
    .B1(\out_val[6] ),
    .B2(_082_),
    .A2(\out_val[7] ),
    .A1(_081_));
 sg13g2_o21ai_1 _672_ (.B1(_293_),
    .Y(_294_),
    .A1(_290_),
    .A2(_292_));
 sg13g2_a22oi_1 _673_ (.Y(_295_),
    .B1(_089_),
    .B2(\pwm.count[7] ),
    .A2(_088_),
    .A1(\pwm.count[8] ));
 sg13g2_nor2b_1 _674_ (.A(\pwm.count[9] ),
    .B_N(\out_val[9] ),
    .Y(_296_));
 sg13g2_a221oi_1 _675_ (.B2(_295_),
    .C1(_296_),
    .B1(_294_),
    .A1(_083_),
    .Y(_297_),
    .A2(\out_val[8] ));
 sg13g2_nand2_1 _676_ (.Y(_298_),
    .A(net81),
    .B(_279_));
 sg13g2_o21ai_1 _677_ (.B1(_277_),
    .Y(_065_),
    .A1(_297_),
    .A2(_298_));
 sg13g2_mux2_1 _678_ (.A0(net88),
    .A1(net92),
    .S(net67),
    .X(_066_));
 sg13g2_mux2_1 _679_ (.A0(net56),
    .A1(net93),
    .S(net67),
    .X(_067_));
 sg13g2_mux2_1 _680_ (.A0(net62),
    .A1(net87),
    .S(net67),
    .X(_068_));
 sg13g2_mux2_1 _681_ (.A0(net65),
    .A1(net104),
    .S(_274_),
    .X(_069_));
 sg13g2_mux2_1 _682_ (.A0(net90),
    .A1(net103),
    .S(net67),
    .X(_070_));
 sg13g2_mux2_1 _683_ (.A0(net111),
    .A1(net113),
    .S(net67),
    .X(_071_));
 sg13g2_mux2_1 _684_ (.A0(net60),
    .A1(net61),
    .S(net67),
    .X(_072_));
 sg13g2_mux2_1 _685_ (.A0(net58),
    .A1(net122),
    .S(net67),
    .X(_073_));
 sg13g2_mux2_1 _686_ (.A0(net94),
    .A1(net100),
    .S(net67),
    .X(_074_));
 sg13g2_nand2b_1 _687_ (.Y(_299_),
    .B(\phase_check[3] ),
    .A_N(\phase_check[2] ));
 sg13g2_nor2_1 _688_ (.A(\phase_check[0] ),
    .B(\phase_check[1] ),
    .Y(_300_));
 sg13g2_nand2_1 _689_ (.Y(_301_),
    .A(\phase_check[1] ),
    .B(\phase_check[3] ));
 sg13g2_a21oi_1 _690_ (.A1(\phase_check[0] ),
    .A2(_299_),
    .Y(_302_),
    .B1(_300_));
 sg13g2_nand3_1 _691_ (.B(\phase_check[2] ),
    .C(_300_),
    .A(\phase_check[3] ),
    .Y(_303_));
 sg13g2_a21oi_1 _692_ (.A1(_301_),
    .A2(_302_),
    .Y(_304_),
    .B1(_084_));
 sg13g2_nor3_1 _693_ (.A(\phase_check[0] ),
    .B(\phase_check[1] ),
    .C(\phase_check[3] ),
    .Y(_305_));
 sg13g2_or3_1 _694_ (.A(\phase_check[0] ),
    .B(\phase_check[2] ),
    .C(_301_),
    .X(_306_));
 sg13g2_a21oi_1 _695_ (.A1(\phase_check[2] ),
    .A2(_305_),
    .Y(_307_),
    .B1(\phase_check[5] ));
 sg13g2_a221oi_1 _696_ (.B2(_307_),
    .C1(_085_),
    .B1(_306_),
    .A1(_303_),
    .Y(_308_),
    .A2(_304_));
 sg13g2_nand4_1 _697_ (.B(\phase_check[2] ),
    .C(_084_),
    .A(\phase_check[3] ),
    .Y(_309_),
    .D(\phase_check[4] ));
 sg13g2_o21ai_1 _698_ (.B1(_309_),
    .Y(_310_),
    .A1(_084_),
    .A2(\phase_check[4] ));
 sg13g2_nand3_1 _699_ (.B(\phase_check[1] ),
    .C(_310_),
    .A(\phase_check[0] ),
    .Y(_311_));
 sg13g2_nor3_1 _700_ (.A(\phase_check[2] ),
    .B(\phase_check[5] ),
    .C(\phase_check[4] ),
    .Y(_312_));
 sg13g2_and2_1 _701_ (.A(_305_),
    .B(_312_),
    .X(_313_));
 sg13g2_nand3b_1 _702_ (.B(_085_),
    .C(_084_),
    .Y(_314_),
    .A_N(_303_));
 sg13g2_nand2_1 _703_ (.Y(_315_),
    .A(_311_),
    .B(_314_));
 sg13g2_nor3_1 _704_ (.A(_308_),
    .B(_313_),
    .C(_315_),
    .Y(_316_));
 sg13g2_nand4_1 _705_ (.B(\event_count[0] ),
    .C(_009_),
    .A(\event_count[1] ),
    .Y(_317_),
    .D(_102_));
 sg13g2_or2_2 _706_ (.X(_318_),
    .B(_317_),
    .A(_316_));
 sg13g2_a21oi_1 _707_ (.A1(net162),
    .A2(_314_),
    .Y(_319_),
    .B1(_313_));
 sg13g2_mux2_1 _708_ (.A0(_319_),
    .A1(net173),
    .S(_318_),
    .X(_075_));
 sg13g2_a21oi_1 _709_ (.A1(net150),
    .A2(_314_),
    .Y(_320_),
    .B1(_313_));
 sg13g2_mux2_1 _710_ (.A0(_320_),
    .A1(net159),
    .S(_318_),
    .X(_076_));
 sg13g2_a21oi_1 _711_ (.A1(\phase_check[5] ),
    .A2(_085_),
    .Y(_321_),
    .B1(_313_));
 sg13g2_mux2_1 _712_ (.A0(_321_),
    .A1(net109),
    .S(_318_),
    .X(_077_));
 sg13g2_nand2_1 _713_ (.Y(_322_),
    .A(net49),
    .B(_318_));
 sg13g2_o21ai_1 _714_ (.B1(_322_),
    .Y(_078_),
    .A1(_084_),
    .A2(_318_));
 sg13g2_dfrbp_1 _715_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net32),
    .D(_022_),
    .Q_N(_012_),
    .Q(\pwm.count[0] ));
 sg13g2_dfrbp_1 _716_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net29),
    .D(net147),
    .Q_N(_367_),
    .Q(\pwm.count[1] ));
 sg13g2_dfrbp_1 _717_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net28),
    .D(_024_),
    .Q_N(_366_),
    .Q(\pwm.count[2] ));
 sg13g2_dfrbp_1 _718_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net27),
    .D(_025_),
    .Q_N(_365_),
    .Q(\pwm.count[3] ));
 sg13g2_dfrbp_1 _719_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net26),
    .D(net125),
    .Q_N(_364_),
    .Q(\pwm.count[4] ));
 sg13g2_dfrbp_1 _720_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net25),
    .D(_027_),
    .Q_N(_363_),
    .Q(\pwm.count[5] ));
 sg13g2_dfrbp_1 _721_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net24),
    .D(_028_),
    .Q_N(_362_),
    .Q(\pwm.count[6] ));
 sg13g2_dfrbp_1 _722_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net23),
    .D(_029_),
    .Q_N(_361_),
    .Q(\pwm.count[7] ));
 sg13g2_dfrbp_1 _723_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net34),
    .D(_030_),
    .Q_N(_360_),
    .Q(\pwm.count[8] ));
 sg13g2_dfrbp_1 _724_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net33),
    .D(net131),
    .Q_N(_359_),
    .Q(\pwm.count[9] ));
 sg13g2_dfrbp_1 _725_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net86),
    .D(net142),
    .Q_N(_358_),
    .Q(\phase_check[0] ));
 sg13g2_dfrbp_1 _726_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net82),
    .D(net129),
    .Q_N(_357_),
    .Q(\phase_check[1] ));
 sg13g2_dfrbp_1 _727_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net82),
    .D(net163),
    .Q_N(_356_),
    .Q(\phase_check[2] ));
 sg13g2_dfrbp_1 _728_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net82),
    .D(net151),
    .Q_N(_355_),
    .Q(\phase_check[3] ));
 sg13g2_dfrbp_1 _729_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net80),
    .D(net169),
    .Q_N(_354_),
    .Q(\phase_check[4] ));
 sg13g2_dfrbp_1 _730_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net80),
    .D(net171),
    .Q_N(_353_),
    .Q(\phase_check[5] ));
 sg13g2_dfrbp_1 _731_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net80),
    .D(net52),
    .Q_N(\out_val[0] ),
    .Q(_013_));
 sg13g2_dfrbp_1 _732_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net80),
    .D(net161),
    .Q_N(_352_),
    .Q(\out_val[1] ));
 sg13g2_dfrbp_1 _733_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net82),
    .D(net149),
    .Q_N(_351_),
    .Q(\out_val[2] ));
 sg13g2_dfrbp_1 _734_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net81),
    .D(_041_),
    .Q_N(\out_val[3] ),
    .Q(_014_));
 sg13g2_dfrbp_1 _735_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net81),
    .D(_042_),
    .Q_N(\out_val[4] ),
    .Q(_015_));
 sg13g2_dfrbp_1 _736_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net82),
    .D(net102),
    .Q_N(\out_val[5] ),
    .Q(_016_));
 sg13g2_dfrbp_1 _737_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net82),
    .D(_044_),
    .Q_N(\out_val[6] ),
    .Q(_017_));
 sg13g2_dfrbp_1 _738_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net81),
    .D(_045_),
    .Q_N(\out_val[7] ),
    .Q(_018_));
 sg13g2_dfrbp_1 _739_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net81),
    .D(net54),
    .Q_N(\out_val[8] ),
    .Q(_019_));
 sg13g2_dfrbp_1 _740_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net81),
    .D(_047_),
    .Q_N(_368_),
    .Q(\out_val[9] ));
 sg13g2_dfrbp_1 _741_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net84),
    .D(net38),
    .Q_N(_369_),
    .Q(\last_input[0] ));
 sg13g2_dfrbp_1 _742_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net84),
    .D(net39),
    .Q_N(_370_),
    .Q(\last_input[1] ));
 sg13g2_dfrbp_1 _743_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net83),
    .D(net44),
    .Q_N(_371_),
    .Q(\last_input[2] ));
 sg13g2_dfrbp_1 _744_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net84),
    .D(net40),
    .Q_N(_372_),
    .Q(\last_input[3] ));
 sg13g2_dfrbp_1 _745_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net85),
    .D(net43),
    .Q_N(_373_),
    .Q(\last_input[4] ));
 sg13g2_dfrbp_1 _746_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net83),
    .D(net36),
    .Q_N(_374_),
    .Q(\last_input[5] ));
 sg13g2_dfrbp_1 _747_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net85),
    .D(net41),
    .Q_N(_375_),
    .Q(\last_input[6] ));
 sg13g2_dfrbp_1 _748_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net85),
    .D(net37),
    .Q_N(_376_),
    .Q(\last_input[7] ));
 sg13g2_dfrbp_1 _749_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net83),
    .D(net1),
    .Q_N(_377_),
    .Q(\new_input[0] ));
 sg13g2_dfrbp_1 _750_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net83),
    .D(net2),
    .Q_N(_378_),
    .Q(\new_input[1] ));
 sg13g2_dfrbp_1 _751_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net83),
    .D(net3),
    .Q_N(_379_),
    .Q(\new_input[2] ));
 sg13g2_dfrbp_1 _752_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net83),
    .D(net4),
    .Q_N(_380_),
    .Q(\new_input[3] ));
 sg13g2_dfrbp_1 _753_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net83),
    .D(net5),
    .Q_N(_381_),
    .Q(\new_input[4] ));
 sg13g2_dfrbp_1 _754_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net83),
    .D(net6),
    .Q_N(_382_),
    .Q(\new_input[5] ));
 sg13g2_dfrbp_1 _755_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net85),
    .D(net7),
    .Q_N(_383_),
    .Q(\new_input[6] ));
 sg13g2_dfrbp_1 _756_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net85),
    .D(net8),
    .Q_N(_384_),
    .Q(\new_input[7] ));
 sg13g2_dfrbp_1 _757_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net77),
    .D(net46),
    .Q_N(_010_),
    .Q(\event_count[0] ));
 sg13g2_dfrbp_1 _758_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net75),
    .D(net99),
    .Q_N(_385_),
    .Q(\event_count[1] ));
 sg13g2_dfrbp_1 _759_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net77),
    .D(_002_),
    .Q_N(_386_),
    .Q(\event_count[2] ));
 sg13g2_dfrbp_1 _760_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net75),
    .D(net108),
    .Q_N(_387_),
    .Q(\event_count[3] ));
 sg13g2_dfrbp_1 _761_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net75),
    .D(_004_),
    .Q_N(_388_),
    .Q(\event_count[4] ));
 sg13g2_dfrbp_1 _762_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net75),
    .D(_005_),
    .Q_N(_389_),
    .Q(\event_count[5] ));
 sg13g2_dfrbp_1 _763_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net75),
    .D(_006_),
    .Q_N(_390_),
    .Q(\event_count[6] ));
 sg13g2_dfrbp_1 _764_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net75),
    .D(net118),
    .Q_N(_391_),
    .Q(\event_count[7] ));
 sg13g2_dfrbp_1 _765_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net77),
    .D(net133),
    .Q_N(_009_),
    .Q(\event_count[8] ));
 sg13g2_dfrbp_1 _766_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net85),
    .D(net89),
    .Q_N(_350_),
    .Q(\next_limit[0] ));
 sg13g2_dfrbp_1 _767_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net86),
    .D(net57),
    .Q_N(_349_),
    .Q(\next_limit[1] ));
 sg13g2_dfrbp_1 _768_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net86),
    .D(_050_),
    .Q_N(_348_),
    .Q(\next_limit[2] ));
 sg13g2_dfrbp_1 _769_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net86),
    .D(net66),
    .Q_N(_347_),
    .Q(\next_limit[3] ));
 sg13g2_dfrbp_1 _770_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net84),
    .D(net91),
    .Q_N(_346_),
    .Q(\next_limit[4] ));
 sg13g2_dfrbp_1 _771_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net84),
    .D(net112),
    .Q_N(_345_),
    .Q(\next_limit[5] ));
 sg13g2_dfrbp_1 _772_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net86),
    .D(_054_),
    .Q_N(_344_),
    .Q(\next_limit[6] ));
 sg13g2_dfrbp_1 _773_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net84),
    .D(net59),
    .Q_N(_343_),
    .Q(\next_limit[7] ));
 sg13g2_dfrbp_1 _774_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net86),
    .D(net95),
    .Q_N(_342_),
    .Q(\next_limit[8] ));
 sg13g2_dfrbp_1 _775_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net78),
    .D(net167),
    .Q_N(_341_),
    .Q(\qtr_count[0] ));
 sg13g2_dfrbp_1 _776_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net78),
    .D(net140),
    .Q_N(_340_),
    .Q(\qtr_count[1] ));
 sg13g2_dfrbp_1 _777_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net78),
    .D(net121),
    .Q_N(_339_),
    .Q(\phase_count[0] ));
 sg13g2_dfrbp_1 _778_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net78),
    .D(_060_),
    .Q_N(_338_),
    .Q(\phase_count[1] ));
 sg13g2_dfrbp_1 _779_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net78),
    .D(_061_),
    .Q_N(_337_),
    .Q(\phase_count[2] ));
 sg13g2_dfrbp_1 _780_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net78),
    .D(net127),
    .Q_N(_336_),
    .Q(\phase_count[3] ));
 sg13g2_dfrbp_1 _781_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net78),
    .D(net153),
    .Q_N(_335_),
    .Q(\phase_count[4] ));
 sg13g2_dfrbp_1 _782_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net78),
    .D(_064_),
    .Q_N(_392_),
    .Q(\phase_count[5] ));
 sg13g2_dfrbp_1 _783_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net85),
    .D(net31),
    .Q_N(_334_),
    .Q(rst_n_i));
 sg13g2_dfrbp_1 _784_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net30),
    .D(net64),
    .Q_N(_333_),
    .Q(\pwm.pwm ));
 sg13g2_dfrbp_1 _785_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net77),
    .D(_066_),
    .Q_N(_332_),
    .Q(\phase_limit[0] ));
 sg13g2_dfrbp_1 _786_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net76),
    .D(_067_),
    .Q_N(_331_),
    .Q(\phase_limit[1] ));
 sg13g2_dfrbp_1 _787_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net77),
    .D(_068_),
    .Q_N(_330_),
    .Q(\phase_limit[2] ));
 sg13g2_dfrbp_1 _788_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net75),
    .D(net105),
    .Q_N(_329_),
    .Q(\phase_limit[3] ));
 sg13g2_dfrbp_1 _789_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net76),
    .D(_070_),
    .Q_N(_328_),
    .Q(\phase_limit[4] ));
 sg13g2_dfrbp_1 _790_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net76),
    .D(_071_),
    .Q_N(_327_),
    .Q(\phase_limit[5] ));
 sg13g2_dfrbp_1 _791_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net75),
    .D(_072_),
    .Q_N(_326_),
    .Q(\phase_limit[6] ));
 sg13g2_dfrbp_1 _792_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net77),
    .D(_073_),
    .Q_N(_325_),
    .Q(\phase_limit[7] ));
 sg13g2_dfrbp_1 _793_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net77),
    .D(_074_),
    .Q_N(_324_),
    .Q(\phase_limit[8] ));
 sg13g2_dfrbp_1 _794_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net80),
    .D(_075_),
    .Q_N(_323_),
    .Q(\delta[0] ));
 sg13g2_dfrbp_1 _795_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net80),
    .D(_076_),
    .Q_N(_011_),
    .Q(\delta[1] ));
 sg13g2_dfrbp_1 _796_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net80),
    .D(net110),
    .Q_N(\delta[2] ),
    .Q(_020_));
 sg13g2_dfrbp_1 _797_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net80),
    .D(net50),
    .Q_N(\delta[3] ),
    .Q(_021_));
 sg13g2_tiehi _721__24 (.L_HI(net24));
 sg13g2_tiehi _720__25 (.L_HI(net25));
 sg13g2_tiehi _719__26 (.L_HI(net26));
 sg13g2_tiehi _718__27 (.L_HI(net27));
 sg13g2_tiehi _717__28 (.L_HI(net28));
 sg13g2_tiehi _716__29 (.L_HI(net29));
 sg13g2_tiehi _784__30 (.L_HI(net30));
 sg13g2_tiehi _783__31 (.L_HI(net31));
 sg13g2_tiehi _715__32 (.L_HI(net32));
 sg13g2_tiehi _724__33 (.L_HI(net33));
 sg13g2_tiehi _723__34 (.L_HI(net34));
 sg13g2_tiehi tt_um_rte_sine_synth_35 (.L_HI(net35));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rte_sine_synth_10 (.L_LO(net10));
 sg13g2_tielo tt_um_rte_sine_synth_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rte_sine_synth_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rte_sine_synth_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rte_sine_synth_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rte_sine_synth_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rte_sine_synth_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rte_sine_synth_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rte_sine_synth_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rte_sine_synth_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rte_sine_synth_20 (.L_LO(net20));
 sg13g2_tielo tt_um_rte_sine_synth_21 (.L_LO(net21));
 sg13g2_tielo tt_um_rte_sine_synth_22 (.L_LO(net22));
 sg13g2_tiehi _722__23 (.L_HI(net23));
 sg13g2_buf_1 _825_ (.A(\pwm.pwm ),
    .X(uio_out[7]));
 sg13g2_buf_1 _826_ (.A(\out_val[2] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _827_ (.A(\out_val[3] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _828_ (.A(\out_val[4] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _829_ (.A(\out_val[5] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _830_ (.A(\out_val[6] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _831_ (.A(\out_val[7] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _832_ (.A(\out_val[8] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _833_ (.A(\out_val[9] ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(_274_));
 sg13g2_buf_2 fanout68 (.A(net69),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_159_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_145_),
    .X(net70));
 sg13g2_buf_1 fanout71 (.A(_145_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_107_));
 sg13g2_buf_2 fanout73 (.A(_196_),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(_196_),
    .X(net74));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(rst_n_i));
 sg13g2_buf_2 fanout76 (.A(net175),
    .X(net76));
 sg13g2_buf_4 fanout77 (.X(net77),
    .A(rst_n_i));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(rst_n_i));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(\qtr_count[0] ));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(net82));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(net82));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(rst_n));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(net84));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(net85));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(net86));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_rte_sine_synth_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\new_input[5] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold2 (.A(\new_input[7] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold3 (.A(\new_input[0] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold4 (.A(\new_input[1] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold5 (.A(\new_input[3] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold6 (.A(\new_input[6] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold7 (.A(_012_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold8 (.A(\new_input[4] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold9 (.A(\new_input[2] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold10 (.A(_010_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold11 (.A(_000_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold12 (.A(_017_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold13 (.A(_018_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold14 (.A(_021_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold15 (.A(_078_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold16 (.A(_013_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold17 (.A(_038_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold18 (.A(_019_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold19 (.A(_046_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold20 (.A(_015_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold21 (.A(\next_limit[1] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold22 (.A(_049_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold23 (.A(\next_limit[7] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold24 (.A(_055_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold25 (.A(\next_limit[6] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold26 (.A(\phase_limit[6] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold27 (.A(\next_limit[2] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold28 (.A(\pwm.pwm ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold29 (.A(_065_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold30 (.A(\next_limit[3] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold31 (.A(_051_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold32 (.A(\phase_limit[2] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold33 (.A(\next_limit[0] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold34 (.A(_048_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold35 (.A(\next_limit[4] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold36 (.A(_052_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold37 (.A(\phase_limit[0] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold38 (.A(\phase_limit[1] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold39 (.A(\next_limit[8] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold40 (.A(_056_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold41 (.A(_014_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold42 (.A(\event_count[0] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold43 (.A(_108_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold44 (.A(_001_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold45 (.A(\phase_limit[8] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold46 (.A(_016_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold47 (.A(_043_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold48 (.A(\phase_limit[4] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold49 (.A(\phase_limit[3] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold50 (.A(_069_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold51 (.A(\event_count[3] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold52 (.A(_114_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold53 (.A(_003_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold54 (.A(_020_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold55 (.A(_077_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold56 (.A(\next_limit[5] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold57 (.A(_053_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold58 (.A(\phase_limit[5] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold59 (.A(\event_count[2] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold60 (.A(_110_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold61 (.A(\event_count[7] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold62 (.A(_123_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold63 (.A(_007_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold64 (.A(\out_val[9] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold65 (.A(\phase_count[0] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold66 (.A(_059_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold67 (.A(\phase_limit[7] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold68 (.A(\pwm.count[4] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold69 (.A(_135_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold70 (.A(_026_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold71 (.A(\phase_count[3] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold72 (.A(_062_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold73 (.A(\phase_check[1] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold74 (.A(_033_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold75 (.A(\pwm.count[9] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold76 (.A(_031_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold77 (.A(\event_count[8] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold78 (.A(_008_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold79 (.A(\pwm.count[2] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold80 (.A(_132_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold81 (.A(\phase_count[1] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold82 (.A(\event_count[6] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold83 (.A(_121_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold84 (.A(\qtr_count[1] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold85 (.A(_058_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold86 (.A(\phase_check[0] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold87 (.A(_032_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold88 (.A(\event_count[5] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold89 (.A(_118_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold90 (.A(_119_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold91 (.A(\pwm.count[0] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold92 (.A(_023_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold93 (.A(\out_val[2] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold94 (.A(_040_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold95 (.A(\phase_check[3] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold96 (.A(_035_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold97 (.A(\phase_count[4] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold98 (.A(_063_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold99 (.A(\pwm.count[6] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold100 (.A(_138_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold101 (.A(\event_count[4] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold102 (.A(\pwm.count[5] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold103 (.A(_136_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold104 (.A(\delta[1] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold105 (.A(\out_val[1] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold106 (.A(_039_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold107 (.A(\phase_check[2] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold108 (.A(_034_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold109 (.A(\pwm.count[7] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold110 (.A(\pwm.count[3] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold111 (.A(\phase_count[5] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold112 (.A(_057_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold113 (.A(\phase_check[4] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold114 (.A(_036_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold115 (.A(\phase_check[5] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold116 (.A(_037_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold117 (.A(\pwm.count[8] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold118 (.A(\delta[0] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold119 (.A(\phase_count[2] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold120 (.A(rst_n_i),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold121 (.A(\pwm.count[3] ),
    .X(net176));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_205 ();
 sg13g2_fill_1 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_fill_1 FILLER_17_184 ();
 sg13g2_decap_4 FILLER_17_194 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_fill_2 FILLER_17_208 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_decap_4 FILLER_17_220 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_fill_2 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_decap_4 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_258 ();
 sg13g2_decap_4 FILLER_17_264 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_175 ();
 sg13g2_decap_4 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_decap_8 FILLER_18_316 ();
 sg13g2_decap_8 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_18_337 ();
 sg13g2_decap_8 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_decap_4 FILLER_19_249 ();
 sg13g2_fill_2 FILLER_19_253 ();
 sg13g2_decap_4 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_4 FILLER_20_168 ();
 sg13g2_decap_4 FILLER_20_207 ();
 sg13g2_fill_1 FILLER_20_211 ();
 sg13g2_fill_1 FILLER_20_220 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_fill_2 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_247 ();
 sg13g2_fill_2 FILLER_20_272 ();
 sg13g2_fill_2 FILLER_20_282 ();
 sg13g2_decap_8 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_decap_4 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_256 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_fill_1 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_fill_1 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_250 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_fill_1 FILLER_22_282 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_fill_1 FILLER_22_383 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_fill_1 FILLER_22_394 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_fill_2 FILLER_23_229 ();
 sg13g2_fill_1 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_304 ();
 sg13g2_fill_1 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_315 ();
 sg13g2_fill_1 FILLER_23_317 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_4 FILLER_24_133 ();
 sg13g2_fill_2 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_313 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_250 ();
 sg13g2_fill_2 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_180 ();
 sg13g2_decap_4 FILLER_26_208 ();
 sg13g2_fill_2 FILLER_26_212 ();
 sg13g2_decap_4 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_262 ();
 sg13g2_fill_2 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_118 ();
 sg13g2_decap_4 FILLER_27_125 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_decap_4 FILLER_27_215 ();
 sg13g2_fill_1 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_4 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_146 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_176 ();
 sg13g2_decap_4 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_282 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_123 ();
 sg13g2_fill_2 FILLER_29_127 ();
 sg13g2_decap_4 FILLER_29_147 ();
 sg13g2_fill_1 FILLER_29_151 ();
 sg13g2_decap_8 FILLER_29_166 ();
 sg13g2_fill_2 FILLER_29_173 ();
 sg13g2_fill_1 FILLER_29_183 ();
 sg13g2_decap_4 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_decap_4 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_90 ();
 sg13g2_fill_2 FILLER_30_130 ();
 sg13g2_fill_2 FILLER_30_136 ();
 sg13g2_decap_8 FILLER_30_142 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_decap_8 FILLER_30_216 ();
 sg13g2_fill_2 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_fill_2 FILLER_30_243 ();
 sg13g2_decap_8 FILLER_30_271 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_317 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_4 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_60 ();
 sg13g2_fill_2 FILLER_31_110 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_decap_4 FILLER_31_172 ();
 sg13g2_fill_2 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_197 ();
 sg13g2_decap_4 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_4 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_58 ();
 sg13g2_fill_2 FILLER_32_99 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_139 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_fill_2 FILLER_32_226 ();
 sg13g2_fill_1 FILLER_32_246 ();
 sg13g2_decap_8 FILLER_32_268 ();
 sg13g2_decap_4 FILLER_32_275 ();
 sg13g2_fill_2 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_357 ();
 sg13g2_fill_1 FILLER_32_376 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_decap_4 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_324 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_fill_1 FILLER_34_85 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_fill_2 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_fill_2 FILLER_34_152 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_fill_1 FILLER_34_177 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_2 FILLER_34_233 ();
 sg13g2_fill_1 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_262 ();
 sg13g2_fill_2 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_347 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_4 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_67 ();
 sg13g2_decap_4 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_282 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_106 ();
 sg13g2_fill_1 FILLER_36_110 ();
 sg13g2_fill_2 FILLER_36_146 ();
 sg13g2_fill_1 FILLER_36_148 ();
 sg13g2_fill_2 FILLER_36_162 ();
 sg13g2_fill_1 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_4 FILLER_36_232 ();
 sg13g2_fill_2 FILLER_36_236 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_4 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_143 ();
 sg13g2_fill_1 FILLER_37_153 ();
 sg13g2_decap_4 FILLER_37_232 ();
 sg13g2_fill_2 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_fill_2 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_163 ();
 sg13g2_fill_2 FILLER_38_173 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_318 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net35;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
endmodule

module tt_um_MichaelBell_hd_8b10b (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire clknet_0_clk;
 wire \i_decoder_a.count[0] ;
 wire \i_decoder_a.count[1] ;
 wire \i_decoder_a.count[2] ;
 wire \i_decoder_a.count[3] ;
 wire \i_decoder_a.data_out[0] ;
 wire \i_decoder_a.data_out[1] ;
 wire \i_decoder_a.data_out[2] ;
 wire \i_decoder_a.data_out[3] ;
 wire \i_decoder_a.data_out[4] ;
 wire \i_decoder_a.data_out[5] ;
 wire \i_decoder_a.data_out[6] ;
 wire \i_decoder_a.data_out[7] ;
 wire \i_decoder_a.i_raw_data.data_out[0] ;
 wire \i_decoder_a.i_raw_data.data_out[1] ;
 wire \i_decoder_a.i_raw_data.data_out[2] ;
 wire \i_decoder_a.i_raw_data.data_out[3] ;
 wire \i_decoder_a.i_raw_data.data_out[4] ;
 wire \i_decoder_a.i_raw_data.data_out[5] ;
 wire \i_decoder_a.i_raw_data.data_out[6] ;
 wire \i_decoder_a.i_raw_data.data_out[7] ;
 wire \i_decoder_a.i_raw_data.data_out[8] ;
 wire \i_decoder_a.i_raw_data.data_out[9] ;
 wire \i_decoder_a.updated ;
 wire \i_decoder_a.valid ;
 wire \i_decoder_b.count[0] ;
 wire \i_decoder_b.count[1] ;
 wire \i_decoder_b.count[2] ;
 wire \i_decoder_b.count[3] ;
 wire \i_decoder_b.data_out[0] ;
 wire \i_decoder_b.data_out[1] ;
 wire \i_decoder_b.data_out[2] ;
 wire \i_decoder_b.data_out[3] ;
 wire \i_decoder_b.data_out[4] ;
 wire \i_decoder_b.data_out[5] ;
 wire \i_decoder_b.data_out[6] ;
 wire \i_decoder_b.data_out[7] ;
 wire \i_decoder_b.i_raw_data.data_out[0] ;
 wire \i_decoder_b.i_raw_data.data_out[1] ;
 wire \i_decoder_b.i_raw_data.data_out[2] ;
 wire \i_decoder_b.i_raw_data.data_out[3] ;
 wire \i_decoder_b.i_raw_data.data_out[4] ;
 wire \i_decoder_b.i_raw_data.data_out[5] ;
 wire \i_decoder_b.i_raw_data.data_out[6] ;
 wire \i_decoder_b.i_raw_data.data_out[7] ;
 wire \i_decoder_b.i_raw_data.data_out[8] ;
 wire \i_decoder_b.i_raw_data.data_out[9] ;
 wire \i_decoder_b.updated ;
 wire \i_decoder_b.valid ;
 wire \result[0] ;
 wire \result[10] ;
 wire \result[11] ;
 wire \result[12] ;
 wire \result[13] ;
 wire \result[14] ;
 wire \result[15] ;
 wire \result[1] ;
 wire \result[2] ;
 wire \result[3] ;
 wire \result[4] ;
 wire \result[5] ;
 wire \result[6] ;
 wire \result[7] ;
 wire \result[8] ;
 wire \result[9] ;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;

 sg13g2_inv_1 _0905_ (.Y(_0056_),
    .A(net154));
 sg13g2_inv_1 _0906_ (.Y(_0057_),
    .A(net138));
 sg13g2_inv_1 _0907_ (.Y(_0058_),
    .A(\i_decoder_a.i_raw_data.data_out[5] ));
 sg13g2_inv_1 _0908_ (.Y(_0059_),
    .A(_0000_));
 sg13g2_inv_1 _0909_ (.Y(_0060_),
    .A(_0001_));
 sg13g2_inv_1 _0910_ (.Y(_0061_),
    .A(\i_decoder_a.i_raw_data.data_out[3] ));
 sg13g2_inv_1 _0911_ (.Y(_0062_),
    .A(\i_decoder_a.i_raw_data.data_out[0] ));
 sg13g2_inv_1 _0912_ (.Y(_0063_),
    .A(net267));
 sg13g2_inv_2 _0913_ (.Y(_0064_),
    .A(net116));
 sg13g2_inv_1 _0914_ (.Y(_0065_),
    .A(_0006_));
 sg13g2_inv_1 _0915_ (.Y(_0066_),
    .A(\i_decoder_b.i_raw_data.data_out[3] ));
 sg13g2_inv_1 _0916_ (.Y(_0067_),
    .A(\i_decoder_b.i_raw_data.data_out[0] ));
 sg13g2_inv_2 _0917_ (.Y(_0068_),
    .A(net124));
 sg13g2_inv_1 _0918_ (.Y(_0069_),
    .A(net262));
 sg13g2_inv_1 _0919_ (.Y(_0070_),
    .A(net252));
 sg13g2_inv_1 _0920_ (.Y(_0071_),
    .A(net239));
 sg13g2_inv_1 _0921_ (.Y(_0072_),
    .A(net229));
 sg13g2_inv_1 _0922_ (.Y(_0073_),
    .A(net224));
 sg13g2_inv_1 _0923_ (.Y(_0074_),
    .A(net216));
 sg13g2_nand2b_2 _0924_ (.Y(uio_oe[7]),
    .B(net265),
    .A_N(net8));
 sg13g2_nand2_1 _0925_ (.Y(_0075_),
    .A(net254),
    .B(net264));
 sg13g2_nor2_2 _0926_ (.A(net257),
    .B(net4),
    .Y(_0076_));
 sg13g2_nand2b_2 _0927_ (.Y(_0077_),
    .B(net266),
    .A_N(net4));
 sg13g2_a21oi_1 _0928_ (.A1(\result[0] ),
    .A2(net255),
    .Y(_0078_),
    .B1(_0077_));
 sg13g2_nor2_1 _0929_ (.A(net267),
    .B(net2),
    .Y(_0079_));
 sg13g2_or2_1 _0930_ (.X(_0080_),
    .B(net2),
    .A(net267));
 sg13g2_and2_2 _0931_ (.A(net266),
    .B(net4),
    .X(_0081_));
 sg13g2_a221oi_1 _0932_ (.B2(_0064_),
    .C1(_0079_),
    .B1(_0081_),
    .A1(_0075_),
    .Y(uo_out[0]),
    .A2(_0078_));
 sg13g2_a21oi_1 _0933_ (.A1(net263),
    .A2(_0070_),
    .Y(_0082_),
    .B1(_0077_));
 sg13g2_o21ai_1 _0934_ (.B1(_0082_),
    .Y(_0083_),
    .A1(\result[1] ),
    .A2(net263));
 sg13g2_nand2_1 _0935_ (.Y(_0084_),
    .A(\i_decoder_a.updated ),
    .B(_0081_));
 sg13g2_nand3_1 _0936_ (.B(_0083_),
    .C(_0084_),
    .A(_0080_),
    .Y(uo_out[1]));
 sg13g2_nand2_1 _0937_ (.Y(_0085_),
    .A(net264),
    .B(net251));
 sg13g2_a21oi_1 _0938_ (.A1(\result[2] ),
    .A2(net255),
    .Y(_0086_),
    .B1(_0077_));
 sg13g2_nor2_1 _0939_ (.A(net267),
    .B(net3),
    .Y(_0087_));
 sg13g2_a221oi_1 _0940_ (.B2(_0086_),
    .C1(_0087_),
    .B1(_0085_),
    .A1(_0068_),
    .Y(uo_out[2]),
    .A2(_0081_));
 sg13g2_nor2_1 _0941_ (.A(net255),
    .B(net249),
    .Y(_0088_));
 sg13g2_o21ai_1 _0942_ (.B1(_0076_),
    .Y(_0089_),
    .A1(\result[3] ),
    .A2(net263));
 sg13g2_a21oi_1 _0943_ (.A1(\i_decoder_b.updated ),
    .A2(_0081_),
    .Y(_0090_),
    .B1(_0087_));
 sg13g2_o21ai_1 _0944_ (.B1(_0090_),
    .Y(uo_out[3]),
    .A1(_0088_),
    .A2(_0089_));
 sg13g2_nand2_1 _0945_ (.Y(_0091_),
    .A(net257),
    .B(net4));
 sg13g2_nor2_1 _0946_ (.A(\result[4] ),
    .B(net263),
    .Y(_0092_));
 sg13g2_o21ai_1 _0947_ (.B1(_0076_),
    .Y(_0093_),
    .A1(_0069_),
    .A2(net247));
 sg13g2_o21ai_1 _0948_ (.B1(_0091_),
    .Y(uo_out[4]),
    .A1(_0092_),
    .A2(_0093_));
 sg13g2_and2_1 _0949_ (.A(net263),
    .B(net245),
    .X(_0094_));
 sg13g2_a21oi_1 _0950_ (.A1(\result[5] ),
    .A2(_0069_),
    .Y(_0095_),
    .B1(_0094_));
 sg13g2_a21oi_2 _0951_ (.B1(net4),
    .Y(uo_out[5]),
    .A2(_0095_),
    .A1(net266));
 sg13g2_nand2_1 _0952_ (.Y(_0096_),
    .A(net257),
    .B(net5));
 sg13g2_nor2_1 _0953_ (.A(\result[6] ),
    .B(net263),
    .Y(_0097_));
 sg13g2_o21ai_1 _0954_ (.B1(_0076_),
    .Y(_0098_),
    .A1(_0069_),
    .A2(net242));
 sg13g2_o21ai_1 _0955_ (.B1(_0096_),
    .Y(uo_out[6]),
    .A1(_0097_),
    .A2(_0098_));
 sg13g2_a21oi_1 _0956_ (.A1(net263),
    .A2(_0071_),
    .Y(_0099_),
    .B1(_0077_));
 sg13g2_o21ai_1 _0957_ (.B1(_0099_),
    .Y(_0100_),
    .A1(\result[7] ),
    .A2(net263));
 sg13g2_o21ai_1 _0958_ (.B1(_0100_),
    .Y(uo_out[7]),
    .A1(net266),
    .A2(net5));
 sg13g2_nand2_1 _0959_ (.Y(_0101_),
    .A(net257),
    .B(net6));
 sg13g2_nor2_1 _0960_ (.A(\result[8] ),
    .B(net262),
    .Y(_0102_));
 sg13g2_o21ai_1 _0961_ (.B1(_0076_),
    .Y(_0103_),
    .A1(net255),
    .A2(net234));
 sg13g2_o21ai_1 _0962_ (.B1(_0101_),
    .Y(uio_out[0]),
    .A1(_0102_),
    .A2(_0103_));
 sg13g2_a21oi_1 _0963_ (.A1(net262),
    .A2(_0072_),
    .Y(_0104_),
    .B1(_0077_));
 sg13g2_o21ai_1 _0964_ (.B1(_0104_),
    .Y(_0105_),
    .A1(\result[9] ),
    .A2(net262));
 sg13g2_o21ai_1 _0965_ (.B1(_0105_),
    .Y(uio_out[1]),
    .A1(net265),
    .A2(net6));
 sg13g2_nand2_1 _0966_ (.Y(_0106_),
    .A(net257),
    .B(net7));
 sg13g2_nor2_1 _0967_ (.A(\result[10] ),
    .B(net261),
    .Y(_0107_));
 sg13g2_o21ai_1 _0968_ (.B1(_0076_),
    .Y(_0108_),
    .A1(net255),
    .A2(\i_decoder_b.data_out[2] ));
 sg13g2_o21ai_1 _0969_ (.B1(_0106_),
    .Y(uio_out[2]),
    .A1(_0107_),
    .A2(_0108_));
 sg13g2_a21oi_1 _0970_ (.A1(net261),
    .A2(_0073_),
    .Y(_0109_),
    .B1(_0077_));
 sg13g2_o21ai_1 _0971_ (.B1(_0109_),
    .Y(_0110_),
    .A1(\result[11] ),
    .A2(net261));
 sg13g2_o21ai_1 _0972_ (.B1(_0110_),
    .Y(uio_out[3]),
    .A1(net265),
    .A2(net7));
 sg13g2_a21oi_1 _0973_ (.A1(\result[12] ),
    .A2(net265),
    .Y(_0111_),
    .B1(net261));
 sg13g2_nor3_1 _0974_ (.A(net256),
    .B(net255),
    .C(net222),
    .Y(_0112_));
 sg13g2_nor3_2 _0975_ (.A(_0081_),
    .B(_0111_),
    .C(_0112_),
    .Y(uio_out[4]));
 sg13g2_o21ai_1 _0976_ (.B1(net255),
    .Y(_0113_),
    .A1(\result[13] ),
    .A2(net256));
 sg13g2_nand3_1 _0977_ (.B(net261),
    .C(net219),
    .A(net265),
    .Y(_0114_));
 sg13g2_a21oi_1 _0978_ (.A1(_0113_),
    .A2(_0114_),
    .Y(uio_out[5]),
    .B1(_0081_));
 sg13g2_nand2_1 _0979_ (.Y(_0115_),
    .A(net258),
    .B(net8));
 sg13g2_nor2_1 _0980_ (.A(\result[14] ),
    .B(net261),
    .Y(_0116_));
 sg13g2_o21ai_1 _0981_ (.B1(_0076_),
    .Y(_0117_),
    .A1(net255),
    .A2(net218));
 sg13g2_o21ai_1 _0982_ (.B1(_0115_),
    .Y(uio_out[6]),
    .A1(_0116_),
    .A2(_0117_));
 sg13g2_a21oi_1 _0983_ (.A1(net261),
    .A2(_0074_),
    .Y(_0118_),
    .B1(_0077_));
 sg13g2_o21ai_1 _0984_ (.B1(_0118_),
    .Y(_0119_),
    .A1(\result[15] ),
    .A2(net261));
 sg13g2_o21ai_1 _0985_ (.B1(_0119_),
    .Y(uio_out[7]),
    .A1(net265),
    .A2(net8));
 sg13g2_nand2_2 _0986_ (.Y(_0120_),
    .A(\i_decoder_a.i_raw_data.data_out[8] ),
    .B(\i_decoder_a.i_raw_data.data_out[9] ));
 sg13g2_xnor2_1 _0987_ (.Y(_0121_),
    .A(\i_decoder_a.i_raw_data.data_out[8] ),
    .B(\i_decoder_a.i_raw_data.data_out[9] ));
 sg13g2_xor2_1 _0988_ (.B(_0121_),
    .A(\i_decoder_a.i_raw_data.data_out[4] ),
    .X(_0122_));
 sg13g2_nor2b_1 _0989_ (.A(_0122_),
    .B_N(\i_decoder_a.i_raw_data.data_out[6] ),
    .Y(_0123_));
 sg13g2_nor2b_1 _0990_ (.A(net236),
    .B_N(_0122_),
    .Y(_0124_));
 sg13g2_xnor2_1 _0991_ (.Y(_0125_),
    .A(net236),
    .B(_0122_));
 sg13g2_xor2_1 _0992_ (.B(_0125_),
    .A(\i_decoder_a.i_raw_data.data_out[7] ),
    .X(_0126_));
 sg13g2_nor2_1 _0993_ (.A(_0000_),
    .B(_0121_),
    .Y(_0127_));
 sg13g2_a21oi_1 _0994_ (.A1(\i_decoder_a.i_raw_data.data_out[4] ),
    .A2(net236),
    .Y(_0128_),
    .B1(_0120_));
 sg13g2_nor2_1 _0995_ (.A(_0127_),
    .B(_0128_),
    .Y(_0129_));
 sg13g2_or2_1 _0996_ (.X(_0130_),
    .B(_0128_),
    .A(_0127_));
 sg13g2_a21oi_1 _0997_ (.A1(_0120_),
    .A2(_0123_),
    .Y(_0131_),
    .B1(_0130_));
 sg13g2_nand3_1 _0998_ (.B(net236),
    .C(\i_decoder_a.i_raw_data.data_out[7] ),
    .A(\i_decoder_a.i_raw_data.data_out[4] ),
    .Y(_0132_));
 sg13g2_and4_2 _0999_ (.A(\i_decoder_a.i_raw_data.data_out[5] ),
    .B(_0126_),
    .C(_0131_),
    .D(_0132_),
    .X(_0133_));
 sg13g2_nor4_2 _1000_ (.A(_0001_),
    .B(_0123_),
    .C(_0124_),
    .Y(_0134_),
    .D(_0129_));
 sg13g2_a221oi_1 _1001_ (.B2(_0060_),
    .C1(_0130_),
    .B1(_0125_),
    .A1(_0120_),
    .Y(_0135_),
    .A2(_0123_));
 sg13g2_or3_1 _1002_ (.A(_0126_),
    .B(_0134_),
    .C(_0135_),
    .X(_0136_));
 sg13g2_nor4_2 _1003_ (.A(\i_decoder_a.i_raw_data.data_out[5] ),
    .B(_0126_),
    .C(_0134_),
    .Y(_0137_),
    .D(_0135_));
 sg13g2_nor2_2 _1004_ (.A(_0133_),
    .B(_0137_),
    .Y(_0138_));
 sg13g2_xor2_1 _1005_ (.B(_0138_),
    .A(\i_decoder_a.i_raw_data.data_out[8] ),
    .X(_0139_));
 sg13g2_o21ai_1 _1006_ (.B1(_0059_),
    .Y(_0140_),
    .A1(_0133_),
    .A2(_0137_));
 sg13g2_or3_1 _1007_ (.A(_0059_),
    .B(_0133_),
    .C(_0137_),
    .X(_0141_));
 sg13g2_and2_1 _1008_ (.A(_0140_),
    .B(_0141_),
    .X(_0142_));
 sg13g2_a21oi_2 _1009_ (.B1(_0133_),
    .Y(_0143_),
    .A2(_0136_),
    .A1(_0058_));
 sg13g2_nand3_1 _1010_ (.B(_0141_),
    .C(_0143_),
    .A(_0140_),
    .Y(_0144_));
 sg13g2_xor2_1 _1011_ (.B(_0138_),
    .A(net236),
    .X(_0145_));
 sg13g2_xnor2_1 _1012_ (.Y(_0146_),
    .A(net236),
    .B(_0138_));
 sg13g2_nand2_2 _1013_ (.Y(_0147_),
    .A(_0144_),
    .B(_0145_));
 sg13g2_a21o_1 _1014_ (.A2(_0141_),
    .A1(_0140_),
    .B1(_0143_),
    .X(_0148_));
 sg13g2_inv_1 _1015_ (.Y(_0149_),
    .A(_0148_));
 sg13g2_xnor2_1 _1016_ (.Y(_0150_),
    .A(_0060_),
    .B(_0138_));
 sg13g2_xnor2_1 _1017_ (.Y(_0151_),
    .A(_0001_),
    .B(_0138_));
 sg13g2_and2_1 _1018_ (.A(_0148_),
    .B(_0151_),
    .X(_0152_));
 sg13g2_mux2_1 _1019_ (.A0(_0144_),
    .A1(_0148_),
    .S(_0145_),
    .X(_0153_));
 sg13g2_a22oi_1 _1020_ (.Y(_0154_),
    .B1(_0153_),
    .B2(_0150_),
    .A2(_0152_),
    .A1(_0147_));
 sg13g2_nand2_1 _1021_ (.Y(_0155_),
    .A(_0142_),
    .B(net206));
 sg13g2_nand4_1 _1022_ (.B(_0143_),
    .C(_0146_),
    .A(_0142_),
    .Y(_0156_),
    .D(_0151_));
 sg13g2_nand2_1 _1023_ (.Y(_0157_),
    .A(_0139_),
    .B(_0156_));
 sg13g2_mux2_1 _1024_ (.A0(_0154_),
    .A1(_0156_),
    .S(net207),
    .X(_0158_));
 sg13g2_and3_1 _1025_ (.X(_0159_),
    .A(_0144_),
    .B(_0146_),
    .C(_0148_));
 sg13g2_nand2b_1 _1026_ (.Y(_0160_),
    .B(_0145_),
    .A_N(_0144_));
 sg13g2_nand2b_1 _1027_ (.Y(_0161_),
    .B(_0160_),
    .A_N(_0159_));
 sg13g2_and2_1 _1028_ (.A(net207),
    .B(_0150_),
    .X(_0162_));
 sg13g2_nand2_1 _1029_ (.Y(_0163_),
    .A(_0161_),
    .B(_0162_));
 sg13g2_xor2_1 _1030_ (.B(_0138_),
    .A(\i_decoder_a.i_raw_data.data_out[9] ),
    .X(_0164_));
 sg13g2_xnor2_1 _1031_ (.Y(_0165_),
    .A(\i_decoder_a.i_raw_data.data_out[9] ),
    .B(_0138_));
 sg13g2_a21oi_1 _1032_ (.A1(_0161_),
    .A2(_0162_),
    .Y(_0166_),
    .B1(_0165_));
 sg13g2_nor2_1 _1033_ (.A(\i_decoder_a.i_raw_data.data_out[3] ),
    .B(\i_decoder_a.i_raw_data.data_out[2] ),
    .Y(_0167_));
 sg13g2_nand2_1 _1034_ (.Y(_0168_),
    .A(\i_decoder_a.i_raw_data.data_out[3] ),
    .B(\i_decoder_a.i_raw_data.data_out[2] ));
 sg13g2_nand2_1 _1035_ (.Y(_0169_),
    .A(_0003_),
    .B(_0168_));
 sg13g2_a21oi_1 _1036_ (.A1(_0003_),
    .A2(_0168_),
    .Y(_0170_),
    .B1(_0167_));
 sg13g2_xnor2_1 _1037_ (.Y(_0171_),
    .A(\i_decoder_a.i_raw_data.data_out[3] ),
    .B(\i_decoder_a.i_raw_data.data_out[2] ));
 sg13g2_xnor2_1 _1038_ (.Y(_0172_),
    .A(\i_decoder_a.i_raw_data.data_out[0] ),
    .B(_0171_));
 sg13g2_nand2b_1 _1039_ (.Y(_0173_),
    .B(_0002_),
    .A_N(\i_decoder_a.i_raw_data.data_out[1] ));
 sg13g2_nand2_1 _1040_ (.Y(_0174_),
    .A(_0002_),
    .B(_0172_));
 sg13g2_or3_1 _1041_ (.A(\i_decoder_a.i_raw_data.data_out[1] ),
    .B(_0170_),
    .C(_0174_),
    .X(_0175_));
 sg13g2_mux2_1 _1042_ (.A0(_0002_),
    .A1(_0173_),
    .S(_0172_),
    .X(_0176_));
 sg13g2_nor2_2 _1043_ (.A(_0170_),
    .B(_0176_),
    .Y(_0177_));
 sg13g2_o21ai_1 _1044_ (.B1(_0175_),
    .Y(_0178_),
    .A1(_0002_),
    .A2(_0177_));
 sg13g2_xnor2_1 _1045_ (.Y(_0179_),
    .A(_0062_),
    .B(_0177_));
 sg13g2_nor2_1 _1046_ (.A(_0178_),
    .B(_0179_),
    .Y(_0180_));
 sg13g2_xnor2_1 _1047_ (.Y(_0181_),
    .A(\i_decoder_a.i_raw_data.data_out[3] ),
    .B(_0177_));
 sg13g2_xnor2_1 _1048_ (.Y(_0182_),
    .A(\i_decoder_a.i_raw_data.data_out[2] ),
    .B(_0177_));
 sg13g2_a21oi_1 _1049_ (.A1(_0002_),
    .A2(_0182_),
    .Y(_0183_),
    .B1(_0180_));
 sg13g2_nand2_1 _1050_ (.Y(_0184_),
    .A(_0181_),
    .B(_0183_));
 sg13g2_and2_1 _1051_ (.A(_0178_),
    .B(_0179_),
    .X(_0185_));
 sg13g2_mux2_1 _1052_ (.A0(_0185_),
    .A1(_0180_),
    .S(_0182_),
    .X(_0186_));
 sg13g2_o21ai_1 _1053_ (.B1(_0184_),
    .Y(_0187_),
    .A1(_0181_),
    .A2(_0186_));
 sg13g2_inv_1 _1054_ (.Y(_0188_),
    .A(_0187_));
 sg13g2_nand2b_1 _1055_ (.Y(_0189_),
    .B(net207),
    .A_N(_0154_));
 sg13g2_nor2_1 _1056_ (.A(_0139_),
    .B(_0150_),
    .Y(_0190_));
 sg13g2_nor2_1 _1057_ (.A(net207),
    .B(_0151_),
    .Y(_0191_));
 sg13g2_nand2b_2 _1058_ (.Y(_0192_),
    .B(_0150_),
    .A_N(net207));
 sg13g2_o21ai_1 _1059_ (.B1(_0165_),
    .Y(_0193_),
    .A1(_0147_),
    .A2(_0192_));
 sg13g2_a21oi_1 _1060_ (.A1(_0153_),
    .A2(_0190_),
    .Y(_0194_),
    .B1(_0193_));
 sg13g2_a221oi_1 _1061_ (.B2(_0194_),
    .C1(_0188_),
    .B1(_0189_),
    .A1(_0158_),
    .Y(_0195_),
    .A2(_0166_));
 sg13g2_inv_1 _1062_ (.Y(_0196_),
    .A(_0195_));
 sg13g2_nor4_1 _1063_ (.A(\i_decoder_a.i_raw_data.data_out[4] ),
    .B(net236),
    .C(\i_decoder_a.i_raw_data.data_out[7] ),
    .D(\i_decoder_a.i_raw_data.data_out[5] ),
    .Y(_0197_));
 sg13g2_nor3_1 _1064_ (.A(\i_decoder_a.i_raw_data.data_out[1] ),
    .B(_0062_),
    .C(_0120_),
    .Y(_0198_));
 sg13g2_nand4_1 _1065_ (.B(\i_decoder_a.i_raw_data.data_out[2] ),
    .C(_0197_),
    .A(_0061_),
    .Y(_0199_),
    .D(_0198_));
 sg13g2_nor4_1 _1066_ (.A(\i_decoder_a.i_raw_data.data_out[8] ),
    .B(\i_decoder_a.i_raw_data.data_out[9] ),
    .C(_0061_),
    .D(\i_decoder_a.i_raw_data.data_out[2] ),
    .Y(_0200_));
 sg13g2_nand4_1 _1067_ (.B(\i_decoder_a.i_raw_data.data_out[1] ),
    .C(_0062_),
    .A(\i_decoder_a.i_raw_data.data_out[5] ),
    .Y(_0201_),
    .D(_0200_));
 sg13g2_o21ai_1 _1068_ (.B1(_0199_),
    .Y(_0202_),
    .A1(_0132_),
    .A2(_0201_));
 sg13g2_nor2_1 _1069_ (.A(_0057_),
    .B(\i_decoder_a.count[2] ),
    .Y(_0203_));
 sg13g2_nor2b_1 _1070_ (.A(\i_decoder_a.count[1] ),
    .B_N(net131),
    .Y(_0204_));
 sg13g2_nand2_2 _1071_ (.Y(_0205_),
    .A(_0203_),
    .B(_0204_));
 sg13g2_nor3_1 _1072_ (.A(_0195_),
    .B(_0202_),
    .C(_0205_),
    .Y(_0206_));
 sg13g2_nor2_1 _1073_ (.A(_0064_),
    .B(_0206_),
    .Y(_0207_));
 sg13g2_nand3_1 _1074_ (.B(\i_decoder_a.count[1] ),
    .C(net131),
    .A(net144),
    .Y(_0208_));
 sg13g2_nor2_1 _1075_ (.A(_0057_),
    .B(net145),
    .Y(_0209_));
 sg13g2_a21oi_1 _1076_ (.A1(_0202_),
    .A2(_0209_),
    .Y(_0210_),
    .B1(_0207_));
 sg13g2_nor2_1 _1077_ (.A(net259),
    .B(_0210_),
    .Y(_0012_));
 sg13g2_or4_1 _1078_ (.A(net259),
    .B(_0064_),
    .C(_0196_),
    .D(_0205_),
    .X(_0211_));
 sg13g2_nand2_1 _1079_ (.Y(_0212_),
    .A(net101),
    .B(net204));
 sg13g2_nand2_1 _1080_ (.Y(_0213_),
    .A(_0156_),
    .B(_0164_));
 sg13g2_nor2b_1 _1081_ (.A(_0143_),
    .B_N(_0142_),
    .Y(_0214_));
 sg13g2_nand2_1 _1082_ (.Y(_0215_),
    .A(net206),
    .B(_0214_));
 sg13g2_nor2_1 _1083_ (.A(net207),
    .B(_0145_),
    .Y(_0216_));
 sg13g2_nor2_1 _1084_ (.A(_0192_),
    .B(_0215_),
    .Y(_0217_));
 sg13g2_xnor2_1 _1085_ (.Y(_0218_),
    .A(\i_decoder_a.i_raw_data.data_out[4] ),
    .B(_0138_));
 sg13g2_nand2b_1 _1086_ (.Y(_0219_),
    .B(net206),
    .A_N(_0218_));
 sg13g2_o21ai_1 _1087_ (.B1(_0219_),
    .Y(_0220_),
    .A1(net206),
    .A2(_0149_));
 sg13g2_nor2_1 _1088_ (.A(net206),
    .B(_0192_),
    .Y(_0221_));
 sg13g2_nor2_1 _1089_ (.A(_0151_),
    .B(_0218_),
    .Y(_0222_));
 sg13g2_nor3_1 _1090_ (.A(net206),
    .B(_0192_),
    .C(_0218_),
    .Y(_0223_));
 sg13g2_o21ai_1 _1091_ (.B1(_0219_),
    .Y(_0224_),
    .A1(_0147_),
    .A2(_0149_));
 sg13g2_and2_1 _1092_ (.A(net207),
    .B(_0151_),
    .X(_0225_));
 sg13g2_inv_1 _1093_ (.Y(_0226_),
    .A(_0225_));
 sg13g2_nand2_1 _1094_ (.Y(_0227_),
    .A(_0161_),
    .B(_0225_));
 sg13g2_a21oi_1 _1095_ (.A1(_0162_),
    .A2(_0220_),
    .Y(_0228_),
    .B1(_0164_));
 sg13g2_a21oi_1 _1096_ (.A1(_0190_),
    .A2(_0224_),
    .Y(_0229_),
    .B1(_0223_));
 sg13g2_nand3_1 _1097_ (.B(_0228_),
    .C(_0229_),
    .A(_0227_),
    .Y(_0230_));
 sg13g2_o21ai_1 _1098_ (.B1(_0230_),
    .Y(_0231_),
    .A1(_0213_),
    .A2(_0217_));
 sg13g2_o21ai_1 _1099_ (.B1(_0212_),
    .Y(_0013_),
    .A1(net204),
    .A2(_0231_));
 sg13g2_a21oi_1 _1100_ (.A1(_0191_),
    .A2(_0224_),
    .Y(_0232_),
    .B1(_0213_));
 sg13g2_nand3_1 _1101_ (.B(_0152_),
    .C(_0157_),
    .A(_0147_),
    .Y(_0233_));
 sg13g2_o21ai_1 _1102_ (.B1(_0162_),
    .Y(_0234_),
    .A1(_0145_),
    .A2(_0214_));
 sg13g2_inv_1 _1103_ (.Y(_0235_),
    .A(_0234_));
 sg13g2_a21oi_1 _1104_ (.A1(_0147_),
    .A2(_0235_),
    .Y(_0236_),
    .B1(_0164_));
 sg13g2_a221oi_1 _1105_ (.B2(_0229_),
    .C1(net203),
    .B1(_0236_),
    .A1(_0232_),
    .Y(_0237_),
    .A2(_0233_));
 sg13g2_a21o_1 _1106_ (.A2(net203),
    .A1(net252),
    .B1(_0237_),
    .X(_0014_));
 sg13g2_nor3_1 _1107_ (.A(net207),
    .B(_0150_),
    .C(_0215_),
    .Y(_0238_));
 sg13g2_nor2_1 _1108_ (.A(_0223_),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_a221oi_1 _1109_ (.B2(_0228_),
    .C1(net203),
    .B1(_0239_),
    .A1(_0163_),
    .Y(_0240_),
    .A2(_0232_));
 sg13g2_a21o_1 _1110_ (.A2(net203),
    .A1(net250),
    .B1(_0240_),
    .X(_0015_));
 sg13g2_nand2_1 _1111_ (.Y(_0241_),
    .A(_0160_),
    .B(_0219_));
 sg13g2_nand3_1 _1112_ (.B(_0226_),
    .C(_0241_),
    .A(_0192_),
    .Y(_0242_));
 sg13g2_a221oi_1 _1113_ (.B2(_0159_),
    .C1(_0164_),
    .B1(_0225_),
    .A1(_0214_),
    .Y(_0243_),
    .A2(_0221_));
 sg13g2_o21ai_1 _1114_ (.B1(_0216_),
    .Y(_0244_),
    .A1(_0152_),
    .A2(_0222_));
 sg13g2_a21oi_1 _1115_ (.A1(_0159_),
    .A2(_0162_),
    .Y(_0245_),
    .B1(_0165_));
 sg13g2_a221oi_1 _1116_ (.B2(_0245_),
    .C1(net203),
    .B1(_0244_),
    .A1(_0242_),
    .Y(_0246_),
    .A2(_0243_));
 sg13g2_a21o_1 _1117_ (.A2(net203),
    .A1(net248),
    .B1(_0246_),
    .X(_0016_));
 sg13g2_o21ai_1 _1118_ (.B1(_0165_),
    .Y(_0247_),
    .A1(_0142_),
    .A2(net206));
 sg13g2_nand2_1 _1119_ (.Y(_0248_),
    .A(_0225_),
    .B(_0247_));
 sg13g2_nor4_1 _1120_ (.A(_0142_),
    .B(net206),
    .C(_0165_),
    .D(_0191_),
    .Y(_0249_));
 sg13g2_or2_1 _1121_ (.X(_0250_),
    .B(_0247_),
    .A(_0192_));
 sg13g2_nand4_1 _1122_ (.B(_0155_),
    .C(_0248_),
    .A(_0143_),
    .Y(_0251_),
    .D(_0250_));
 sg13g2_nor3_1 _1123_ (.A(net203),
    .B(_0249_),
    .C(_0251_),
    .Y(_0252_));
 sg13g2_a21o_1 _1124_ (.A2(net203),
    .A1(net246),
    .B1(_0252_),
    .X(_0017_));
 sg13g2_xnor2_1 _1125_ (.Y(_0253_),
    .A(\i_decoder_a.i_raw_data.data_out[1] ),
    .B(\i_decoder_a.i_raw_data.data_out[0] ));
 sg13g2_nor2_1 _1126_ (.A(_0181_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_nor2b_1 _1127_ (.A(_0176_),
    .B_N(_0167_),
    .Y(_0255_));
 sg13g2_o21ai_1 _1128_ (.B1(_0169_),
    .Y(_0256_),
    .A1(_0003_),
    .A2(_0255_));
 sg13g2_a22oi_1 _1129_ (.Y(_0257_),
    .B1(_0254_),
    .B2(_0182_),
    .A2(_0185_),
    .A1(_0181_));
 sg13g2_nand2_1 _1130_ (.Y(_0258_),
    .A(_0256_),
    .B(_0257_));
 sg13g2_mux2_1 _1131_ (.A0(_0258_),
    .A1(net245),
    .S(net204),
    .X(_0018_));
 sg13g2_nand2_1 _1132_ (.Y(_0259_),
    .A(_0184_),
    .B(_0256_));
 sg13g2_mux2_1 _1133_ (.A0(_0259_),
    .A1(net242),
    .S(net204),
    .X(_0019_));
 sg13g2_a21oi_1 _1134_ (.A1(_0178_),
    .A2(_0181_),
    .Y(_0260_),
    .B1(_0254_));
 sg13g2_nor2_1 _1135_ (.A(_0182_),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_nor4_1 _1136_ (.A(_0061_),
    .B(\i_decoder_a.i_raw_data.data_out[2] ),
    .C(net80),
    .D(net152),
    .Y(_0262_));
 sg13g2_nor3_1 _1137_ (.A(net204),
    .B(_0261_),
    .C(_0262_),
    .Y(_0263_));
 sg13g2_a21oi_1 _1138_ (.A1(_0071_),
    .A2(net204),
    .Y(_0020_),
    .B1(_0263_));
 sg13g2_nand2_1 _1139_ (.Y(_0264_),
    .A(net99),
    .B(_0205_));
 sg13g2_a22oi_1 _1140_ (.Y(_0265_),
    .B1(_0207_),
    .B2(_0264_),
    .A2(_0064_),
    .A1(\i_decoder_a.count[0] ));
 sg13g2_nand3b_1 _1141_ (.B(_0209_),
    .C(_0064_),
    .Y(_0266_),
    .A_N(_0202_));
 sg13g2_and2_1 _1142_ (.A(net267),
    .B(_0266_),
    .X(_0267_));
 sg13g2_nand2b_1 _1143_ (.Y(_0021_),
    .B(_0267_),
    .A_N(net100));
 sg13g2_nor2b_1 _1144_ (.A(net131),
    .B_N(\i_decoder_a.count[1] ),
    .Y(_0268_));
 sg13g2_nand2_1 _1145_ (.Y(_0269_),
    .A(net116),
    .B(_0203_));
 sg13g2_a21oi_1 _1146_ (.A1(_0204_),
    .A2(_0269_),
    .Y(_0270_),
    .B1(net132));
 sg13g2_a21oi_1 _1147_ (.A1(_0266_),
    .A2(net133),
    .Y(_0022_),
    .B1(net259));
 sg13g2_nand2_1 _1148_ (.Y(_0271_),
    .A(net116),
    .B(_0206_));
 sg13g2_a21o_1 _1149_ (.A2(\i_decoder_a.count[0] ),
    .A1(\i_decoder_a.count[1] ),
    .B1(\i_decoder_a.count[2] ),
    .X(_0272_));
 sg13g2_nand2_1 _1150_ (.Y(_0273_),
    .A(_0208_),
    .B(_0272_));
 sg13g2_nand3_1 _1151_ (.B(_0271_),
    .C(_0273_),
    .A(_0267_),
    .Y(_0023_));
 sg13g2_xnor2_1 _1152_ (.Y(_0274_),
    .A(net138),
    .B(_0208_));
 sg13g2_a22oi_1 _1153_ (.Y(_0275_),
    .B1(_0205_),
    .B2(net139),
    .A2(_0203_),
    .A1(_0064_));
 sg13g2_a21oi_1 _1154_ (.A1(_0266_),
    .A2(net140),
    .Y(_0024_),
    .B1(net259));
 sg13g2_nor4_1 _1155_ (.A(net259),
    .B(net75),
    .C(_0196_),
    .D(_0205_),
    .Y(_0025_));
 sg13g2_nand2_2 _1156_ (.Y(_0276_),
    .A(\i_decoder_b.i_raw_data.data_out[8] ),
    .B(\i_decoder_b.i_raw_data.data_out[9] ));
 sg13g2_xnor2_1 _1157_ (.Y(_0277_),
    .A(\i_decoder_b.i_raw_data.data_out[8] ),
    .B(\i_decoder_b.i_raw_data.data_out[9] ));
 sg13g2_xor2_1 _1158_ (.B(_0277_),
    .A(\i_decoder_b.i_raw_data.data_out[4] ),
    .X(_0278_));
 sg13g2_nor2b_1 _1159_ (.A(_0278_),
    .B_N(\i_decoder_b.i_raw_data.data_out[6] ),
    .Y(_0279_));
 sg13g2_xnor2_1 _1160_ (.Y(_0280_),
    .A(\i_decoder_b.i_raw_data.data_out[6] ),
    .B(_0278_));
 sg13g2_xor2_1 _1161_ (.B(_0280_),
    .A(\i_decoder_b.i_raw_data.data_out[7] ),
    .X(_0281_));
 sg13g2_nand2_1 _1162_ (.Y(_0282_),
    .A(\i_decoder_b.i_raw_data.data_out[5] ),
    .B(_0281_));
 sg13g2_and4_1 _1163_ (.A(\i_decoder_b.i_raw_data.data_out[4] ),
    .B(\i_decoder_b.i_raw_data.data_out[6] ),
    .C(\i_decoder_b.i_raw_data.data_out[7] ),
    .D(\i_decoder_b.i_raw_data.data_out[5] ),
    .X(_0283_));
 sg13g2_a21o_1 _1164_ (.A2(\i_decoder_b.i_raw_data.data_out[6] ),
    .A1(\i_decoder_b.i_raw_data.data_out[4] ),
    .B1(_0276_),
    .X(_0284_));
 sg13g2_o21ai_1 _1165_ (.B1(_0284_),
    .Y(_0285_),
    .A1(_0005_),
    .A2(_0277_));
 sg13g2_a21o_1 _1166_ (.A2(_0279_),
    .A1(_0276_),
    .B1(_0285_),
    .X(_0286_));
 sg13g2_and2_1 _1167_ (.A(_0065_),
    .B(_0280_),
    .X(_0287_));
 sg13g2_a21o_1 _1168_ (.A2(_0281_),
    .A1(\i_decoder_b.i_raw_data.data_out[5] ),
    .B1(_0287_),
    .X(_0288_));
 sg13g2_or3_1 _1169_ (.A(_0282_),
    .B(_0283_),
    .C(_0286_),
    .X(_0289_));
 sg13g2_a221oi_1 _1170_ (.B2(_0065_),
    .C1(_0285_),
    .B1(_0280_),
    .A1(_0276_),
    .Y(_0290_),
    .A2(_0279_));
 sg13g2_or3_1 _1171_ (.A(\i_decoder_b.i_raw_data.data_out[5] ),
    .B(_0281_),
    .C(_0290_),
    .X(_0291_));
 sg13g2_a221oi_1 _1172_ (.B2(_0282_),
    .C1(_0283_),
    .B1(_0291_),
    .A1(_0286_),
    .Y(_0292_),
    .A2(_0288_));
 sg13g2_xnor2_1 _1173_ (.Y(_0293_),
    .A(\i_decoder_b.i_raw_data.data_out[8] ),
    .B(_0292_));
 sg13g2_xor2_1 _1174_ (.B(net208),
    .A(_0005_),
    .X(_0294_));
 sg13g2_o21ai_1 _1175_ (.B1(_0289_),
    .Y(_0295_),
    .A1(\i_decoder_b.i_raw_data.data_out[5] ),
    .A2(net208));
 sg13g2_nor2_1 _1176_ (.A(_0294_),
    .B(_0295_),
    .Y(_0296_));
 sg13g2_xnor2_1 _1177_ (.Y(_0297_),
    .A(\i_decoder_b.i_raw_data.data_out[6] ),
    .B(net208));
 sg13g2_xor2_1 _1178_ (.B(net208),
    .A(\i_decoder_b.i_raw_data.data_out[6] ),
    .X(_0298_));
 sg13g2_xnor2_1 _1179_ (.Y(_0299_),
    .A(_0065_),
    .B(net208));
 sg13g2_xnor2_1 _1180_ (.Y(_0300_),
    .A(_0006_),
    .B(net208));
 sg13g2_nor2_1 _1181_ (.A(_0294_),
    .B(net205),
    .Y(_0301_));
 sg13g2_nor4_2 _1182_ (.A(_0294_),
    .B(_0295_),
    .C(_0297_),
    .Y(_0302_),
    .D(_0300_));
 sg13g2_nand2b_1 _1183_ (.Y(_0303_),
    .B(_0293_),
    .A_N(_0302_));
 sg13g2_o21ai_1 _1184_ (.B1(net205),
    .Y(_0304_),
    .A1(_0294_),
    .A2(_0295_));
 sg13g2_and2_2 _1185_ (.A(_0294_),
    .B(_0295_),
    .X(_0305_));
 sg13g2_nor2_1 _1186_ (.A(_0300_),
    .B(_0305_),
    .Y(_0306_));
 sg13g2_nand3b_1 _1187_ (.B(_0299_),
    .C(_0304_),
    .Y(_0307_),
    .A_N(_0305_));
 sg13g2_o21ai_1 _1188_ (.B1(_0298_),
    .Y(_0308_),
    .A1(_0294_),
    .A2(_0295_));
 sg13g2_mux2_1 _1189_ (.A0(_0296_),
    .A1(_0305_),
    .S(net205),
    .X(_0309_));
 sg13g2_o21ai_1 _1190_ (.B1(_0308_),
    .Y(_0310_),
    .A1(_0298_),
    .A2(_0305_));
 sg13g2_o21ai_1 _1191_ (.B1(_0307_),
    .Y(_0311_),
    .A1(_0299_),
    .A2(_0309_));
 sg13g2_o21ai_1 _1192_ (.B1(_0303_),
    .Y(_0312_),
    .A1(_0293_),
    .A2(_0311_));
 sg13g2_xor2_1 _1193_ (.B(net208),
    .A(\i_decoder_b.i_raw_data.data_out[9] ),
    .X(_0313_));
 sg13g2_and2_2 _1194_ (.A(_0293_),
    .B(_0300_),
    .X(_0314_));
 sg13g2_nand2_1 _1195_ (.Y(_0315_),
    .A(_0296_),
    .B(net205));
 sg13g2_nor2_1 _1196_ (.A(_0305_),
    .B(_0308_),
    .Y(_0316_));
 sg13g2_o21ai_1 _1197_ (.B1(_0315_),
    .Y(_0317_),
    .A1(_0305_),
    .A2(_0308_));
 sg13g2_nand2_1 _1198_ (.Y(_0318_),
    .A(_0314_),
    .B(_0317_));
 sg13g2_a21oi_1 _1199_ (.A1(_0314_),
    .A2(_0317_),
    .Y(_0319_),
    .B1(_0313_));
 sg13g2_nor2_2 _1200_ (.A(_0293_),
    .B(_0300_),
    .Y(_0320_));
 sg13g2_nor2_2 _1201_ (.A(_0293_),
    .B(_0299_),
    .Y(_0321_));
 sg13g2_nand2b_1 _1202_ (.Y(_0322_),
    .B(_0321_),
    .A_N(_0304_));
 sg13g2_nand2_1 _1203_ (.Y(_0323_),
    .A(_0313_),
    .B(_0322_));
 sg13g2_a221oi_1 _1204_ (.B2(_0310_),
    .C1(_0323_),
    .B1(_0320_),
    .A1(_0293_),
    .Y(_0324_),
    .A2(_0311_));
 sg13g2_nor2_1 _1205_ (.A(\i_decoder_b.i_raw_data.data_out[3] ),
    .B(\i_decoder_b.i_raw_data.data_out[2] ),
    .Y(_0325_));
 sg13g2_nand2_1 _1206_ (.Y(_0326_),
    .A(\i_decoder_b.i_raw_data.data_out[3] ),
    .B(\i_decoder_b.i_raw_data.data_out[2] ));
 sg13g2_nand2_1 _1207_ (.Y(_0327_),
    .A(_0008_),
    .B(_0326_));
 sg13g2_a21oi_1 _1208_ (.A1(_0008_),
    .A2(_0326_),
    .Y(_0328_),
    .B1(_0325_));
 sg13g2_xnor2_1 _1209_ (.Y(_0329_),
    .A(\i_decoder_b.i_raw_data.data_out[3] ),
    .B(\i_decoder_b.i_raw_data.data_out[2] ));
 sg13g2_xnor2_1 _1210_ (.Y(_0330_),
    .A(\i_decoder_b.i_raw_data.data_out[0] ),
    .B(_0329_));
 sg13g2_nor2b_1 _1211_ (.A(\i_decoder_b.i_raw_data.data_out[1] ),
    .B_N(_0007_),
    .Y(_0331_));
 sg13g2_nor2_1 _1212_ (.A(_0007_),
    .B(_0330_),
    .Y(_0332_));
 sg13g2_a21oi_1 _1213_ (.A1(_0330_),
    .A2(_0331_),
    .Y(_0333_),
    .B1(_0332_));
 sg13g2_nor2_2 _1214_ (.A(_0328_),
    .B(_0333_),
    .Y(_0334_));
 sg13g2_xnor2_1 _1215_ (.Y(_0335_),
    .A(\i_decoder_b.i_raw_data.data_out[2] ),
    .B(_0334_));
 sg13g2_nand2_1 _1216_ (.Y(_0336_),
    .A(_0007_),
    .B(_0335_));
 sg13g2_nand3b_1 _1217_ (.B(_0330_),
    .C(_0331_),
    .Y(_0337_),
    .A_N(_0328_));
 sg13g2_o21ai_1 _1218_ (.B1(_0337_),
    .Y(_0338_),
    .A1(_0007_),
    .A2(_0334_));
 sg13g2_xnor2_1 _1219_ (.Y(_0339_),
    .A(_0067_),
    .B(_0334_));
 sg13g2_or2_1 _1220_ (.X(_0340_),
    .B(_0339_),
    .A(_0338_));
 sg13g2_xnor2_1 _1221_ (.Y(_0341_),
    .A(\i_decoder_b.i_raw_data.data_out[3] ),
    .B(_0334_));
 sg13g2_nand3_1 _1222_ (.B(_0340_),
    .C(_0341_),
    .A(_0336_),
    .Y(_0342_));
 sg13g2_nor2b_1 _1223_ (.A(_0341_),
    .B_N(_0335_),
    .Y(_0343_));
 sg13g2_nand2_1 _1224_ (.Y(_0344_),
    .A(_0338_),
    .B(_0339_));
 sg13g2_nor2_1 _1225_ (.A(_0335_),
    .B(_0341_),
    .Y(_0345_));
 sg13g2_a22oi_1 _1226_ (.Y(_0346_),
    .B1(_0344_),
    .B2(_0345_),
    .A2(_0343_),
    .A1(_0340_));
 sg13g2_a221oi_1 _1227_ (.B2(_0346_),
    .C1(_0324_),
    .B1(_0342_),
    .A1(_0312_),
    .Y(_0347_),
    .A2(_0319_));
 sg13g2_inv_1 _1228_ (.Y(_0348_),
    .A(_0347_));
 sg13g2_nor4_1 _1229_ (.A(\i_decoder_b.i_raw_data.data_out[4] ),
    .B(\i_decoder_b.i_raw_data.data_out[6] ),
    .C(\i_decoder_b.i_raw_data.data_out[7] ),
    .D(\i_decoder_b.i_raw_data.data_out[5] ),
    .Y(_0349_));
 sg13g2_nor2_1 _1230_ (.A(\i_decoder_b.i_raw_data.data_out[1] ),
    .B(_0067_),
    .Y(_0350_));
 sg13g2_nand4_1 _1231_ (.B(\i_decoder_b.i_raw_data.data_out[2] ),
    .C(_0349_),
    .A(_0066_),
    .Y(_0351_),
    .D(_0350_));
 sg13g2_nor4_1 _1232_ (.A(\i_decoder_b.i_raw_data.data_out[8] ),
    .B(\i_decoder_b.i_raw_data.data_out[9] ),
    .C(_0066_),
    .D(\i_decoder_b.i_raw_data.data_out[2] ),
    .Y(_0352_));
 sg13g2_nand4_1 _1233_ (.B(_0067_),
    .C(_0283_),
    .A(\i_decoder_b.i_raw_data.data_out[1] ),
    .Y(_0353_),
    .D(_0352_));
 sg13g2_o21ai_1 _1234_ (.B1(_0353_),
    .Y(_0354_),
    .A1(_0276_),
    .A2(_0351_));
 sg13g2_nor2b_1 _1235_ (.A(\i_decoder_b.count[1] ),
    .B_N(net125),
    .Y(_0355_));
 sg13g2_nor2_2 _1236_ (.A(_0056_),
    .B(net149),
    .Y(_0356_));
 sg13g2_nand2_2 _1237_ (.Y(_0357_),
    .A(_0355_),
    .B(_0356_));
 sg13g2_or2_1 _1238_ (.X(_0358_),
    .B(_0357_),
    .A(_0354_));
 sg13g2_o21ai_1 _1239_ (.B1(net124),
    .Y(_0359_),
    .A1(_0347_),
    .A2(_0358_));
 sg13g2_nand3_1 _1240_ (.B(\i_decoder_b.count[1] ),
    .C(net125),
    .A(net149),
    .Y(_0360_));
 sg13g2_or2_1 _1241_ (.X(_0361_),
    .B(_0360_),
    .A(_0056_));
 sg13g2_nand2b_1 _1242_ (.Y(_0362_),
    .B(_0354_),
    .A_N(_0361_));
 sg13g2_a21oi_1 _1243_ (.A1(_0359_),
    .A2(_0362_),
    .Y(_0026_),
    .B1(net259));
 sg13g2_nor4_2 _1244_ (.A(net259),
    .B(_0068_),
    .C(_0348_),
    .Y(_0363_),
    .D(_0357_));
 sg13g2_nor2b_1 _1245_ (.A(_0294_),
    .B_N(_0295_),
    .Y(_0364_));
 sg13g2_and2_1 _1246_ (.A(_0298_),
    .B(_0364_),
    .X(_0365_));
 sg13g2_nand2_1 _1247_ (.Y(_0366_),
    .A(_0321_),
    .B(_0365_));
 sg13g2_nor2_1 _1248_ (.A(_0302_),
    .B(_0313_),
    .Y(_0367_));
 sg13g2_xnor2_1 _1249_ (.Y(_0368_),
    .A(\i_decoder_b.i_raw_data.data_out[4] ),
    .B(net208));
 sg13g2_nand2_1 _1250_ (.Y(_0369_),
    .A(_0298_),
    .B(_0368_));
 sg13g2_o21ai_1 _1251_ (.B1(_0369_),
    .Y(_0370_),
    .A1(_0298_),
    .A2(_0305_));
 sg13g2_nand3_1 _1252_ (.B(_0321_),
    .C(_0368_),
    .A(net205),
    .Y(_0371_));
 sg13g2_nand2_1 _1253_ (.Y(_0372_),
    .A(_0313_),
    .B(_0371_));
 sg13g2_a21oi_1 _1254_ (.A1(_0314_),
    .A2(_0370_),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_o21ai_1 _1255_ (.B1(_0369_),
    .Y(_0374_),
    .A1(_0304_),
    .A2(_0305_));
 sg13g2_and2_1 _1256_ (.A(_0293_),
    .B(_0299_),
    .X(_0375_));
 sg13g2_a22oi_1 _1257_ (.Y(_0376_),
    .B1(_0375_),
    .B2(_0317_),
    .A2(_0374_),
    .A1(_0320_));
 sg13g2_a22oi_1 _1258_ (.Y(_0377_),
    .B1(_0373_),
    .B2(_0376_),
    .A2(_0367_),
    .A1(_0366_));
 sg13g2_mux2_1 _1259_ (.A0(net234),
    .A1(_0377_),
    .S(_0363_),
    .X(_0027_));
 sg13g2_nand2_1 _1260_ (.Y(_0378_),
    .A(_0321_),
    .B(_0374_));
 sg13g2_and2_1 _1261_ (.A(_0367_),
    .B(_0378_),
    .X(_0379_));
 sg13g2_nand2b_1 _1262_ (.Y(_0380_),
    .B(_0303_),
    .A_N(_0307_));
 sg13g2_a21o_1 _1263_ (.A2(net205),
    .A1(_0296_),
    .B1(_0365_),
    .X(_0381_));
 sg13g2_a221oi_1 _1264_ (.B2(_0314_),
    .C1(_0372_),
    .B1(_0381_),
    .A1(_0320_),
    .Y(_0382_),
    .A2(_0374_));
 sg13g2_a21oi_1 _1265_ (.A1(_0379_),
    .A2(_0380_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_mux2_1 _1266_ (.A0(net230),
    .A1(_0383_),
    .S(_0363_),
    .X(_0028_));
 sg13g2_nand2_1 _1267_ (.Y(_0384_),
    .A(_0320_),
    .B(_0365_));
 sg13g2_a22oi_1 _1268_ (.Y(_0385_),
    .B1(_0384_),
    .B2(_0373_),
    .A2(_0379_),
    .A1(_0318_));
 sg13g2_mux2_1 _1269_ (.A0(net226),
    .A1(_0385_),
    .S(_0363_),
    .X(_0029_));
 sg13g2_a21oi_1 _1270_ (.A1(_0300_),
    .A2(_0368_),
    .Y(_0386_),
    .B1(_0306_));
 sg13g2_or3_1 _1271_ (.A(_0293_),
    .B(_0297_),
    .C(_0386_),
    .X(_0387_));
 sg13g2_a21oi_1 _1272_ (.A1(_0314_),
    .A2(_0316_),
    .Y(_0388_),
    .B1(_0313_));
 sg13g2_nand3_1 _1273_ (.B(_0321_),
    .C(_0364_),
    .A(net205),
    .Y(_0389_));
 sg13g2_nand2_1 _1274_ (.Y(_0390_),
    .A(_0313_),
    .B(_0389_));
 sg13g2_nand2_1 _1275_ (.Y(_0391_),
    .A(_0315_),
    .B(_0369_));
 sg13g2_o21ai_1 _1276_ (.B1(_0391_),
    .Y(_0392_),
    .A1(_0314_),
    .A2(_0320_));
 sg13g2_a21oi_1 _1277_ (.A1(_0316_),
    .A2(_0375_),
    .Y(_0393_),
    .B1(_0390_));
 sg13g2_a22oi_1 _1278_ (.Y(_0394_),
    .B1(_0392_),
    .B2(_0393_),
    .A2(_0388_),
    .A1(_0387_));
 sg13g2_mux2_1 _1279_ (.A0(net225),
    .A1(_0394_),
    .S(_0363_),
    .X(_0030_));
 sg13g2_nand2_1 _1280_ (.Y(_0395_),
    .A(_0294_),
    .B(net205));
 sg13g2_nand2_1 _1281_ (.Y(_0396_),
    .A(_0313_),
    .B(_0395_));
 sg13g2_nor3_1 _1282_ (.A(_0313_),
    .B(_0321_),
    .C(_0395_),
    .Y(_0397_));
 sg13g2_mux2_1 _1283_ (.A0(_0321_),
    .A1(_0375_),
    .S(_0396_),
    .X(_0398_));
 sg13g2_nor4_1 _1284_ (.A(_0295_),
    .B(_0301_),
    .C(_0397_),
    .D(_0398_),
    .Y(_0399_));
 sg13g2_mux2_1 _1285_ (.A0(net222),
    .A1(_0399_),
    .S(_0363_),
    .X(_0031_));
 sg13g2_xor2_1 _1286_ (.B(\i_decoder_b.i_raw_data.data_out[0] ),
    .A(\i_decoder_b.i_raw_data.data_out[1] ),
    .X(_0400_));
 sg13g2_nor2b_1 _1287_ (.A(_0333_),
    .B_N(_0325_),
    .Y(_0401_));
 sg13g2_o21ai_1 _1288_ (.B1(_0327_),
    .Y(_0402_),
    .A1(_0008_),
    .A2(_0401_));
 sg13g2_nand3_1 _1289_ (.B(_0339_),
    .C(_0341_),
    .A(_0338_),
    .Y(_0403_));
 sg13g2_nand2_1 _1290_ (.Y(_0404_),
    .A(_0402_),
    .B(_0403_));
 sg13g2_a21o_1 _1291_ (.A2(_0400_),
    .A1(_0343_),
    .B1(_0404_),
    .X(_0405_));
 sg13g2_mux2_1 _1292_ (.A0(net220),
    .A1(_0405_),
    .S(_0363_),
    .X(_0032_));
 sg13g2_nand2_1 _1293_ (.Y(_0406_),
    .A(_0342_),
    .B(_0402_));
 sg13g2_mux2_1 _1294_ (.A0(net97),
    .A1(_0406_),
    .S(_0363_),
    .X(_0033_));
 sg13g2_o21ai_1 _1295_ (.B1(_0335_),
    .Y(_0407_),
    .A1(_0339_),
    .A2(_0341_));
 sg13g2_nand2_1 _1296_ (.Y(_0408_),
    .A(_0338_),
    .B(_0407_));
 sg13g2_nand2_1 _1297_ (.Y(_0409_),
    .A(_0345_),
    .B(_0400_));
 sg13g2_o21ai_1 _1298_ (.B1(_0409_),
    .Y(_0410_),
    .A1(_0345_),
    .A2(_0408_));
 sg13g2_mux2_1 _1299_ (.A0(net216),
    .A1(_0410_),
    .S(_0363_),
    .X(_0034_));
 sg13g2_a21oi_1 _1300_ (.A1(net93),
    .A2(_0357_),
    .Y(_0411_),
    .B1(_0359_));
 sg13g2_nor2b_1 _1301_ (.A(\i_decoder_b.valid ),
    .B_N(\i_decoder_b.count[0] ),
    .Y(_0412_));
 sg13g2_or3_1 _1302_ (.A(net124),
    .B(_0354_),
    .C(_0361_),
    .X(_0413_));
 sg13g2_and2_1 _1303_ (.A(net267),
    .B(_0413_),
    .X(_0414_));
 sg13g2_o21ai_1 _1304_ (.B1(_0414_),
    .Y(_0035_),
    .A1(net94),
    .A2(_0412_));
 sg13g2_nor2b_1 _1305_ (.A(net125),
    .B_N(\i_decoder_b.count[1] ),
    .Y(_0415_));
 sg13g2_nand2_1 _1306_ (.Y(_0416_),
    .A(net124),
    .B(_0356_));
 sg13g2_a21oi_1 _1307_ (.A1(_0355_),
    .A2(_0416_),
    .Y(_0417_),
    .B1(net126));
 sg13g2_a21oi_1 _1308_ (.A1(_0413_),
    .A2(net127),
    .Y(_0036_),
    .B1(net259));
 sg13g2_nor3_1 _1309_ (.A(_0068_),
    .B(_0347_),
    .C(_0358_),
    .Y(_0418_));
 sg13g2_a21o_1 _1310_ (.A2(net125),
    .A1(\i_decoder_b.count[1] ),
    .B1(net149),
    .X(_0419_));
 sg13g2_nand2b_1 _1311_ (.Y(_0420_),
    .B(_0414_),
    .A_N(_0418_));
 sg13g2_a21o_1 _1312_ (.A2(net150),
    .A1(_0360_),
    .B1(_0420_),
    .X(_0037_));
 sg13g2_a22oi_1 _1313_ (.Y(_0421_),
    .B1(_0360_),
    .B2(_0056_),
    .A2(_0356_),
    .A1(_0355_));
 sg13g2_a22oi_1 _1314_ (.Y(_0422_),
    .B1(_0361_),
    .B2(net155),
    .A2(_0356_),
    .A1(_0068_));
 sg13g2_a21oi_1 _1315_ (.A1(_0413_),
    .A2(_0422_),
    .Y(_0038_),
    .B1(net260));
 sg13g2_nand3_1 _1316_ (.B(net6),
    .C(\i_decoder_b.updated ),
    .A(\i_decoder_a.updated ),
    .Y(_0423_));
 sg13g2_nor2b_1 _1317_ (.A(net5),
    .B_N(_0423_),
    .Y(_0424_));
 sg13g2_nand2b_1 _1318_ (.Y(_0425_),
    .B(_0423_),
    .A_N(net5));
 sg13g2_nor2_1 _1319_ (.A(net7),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_nor3_1 _1320_ (.A(net123),
    .B(net7),
    .C(net213),
    .Y(_0427_));
 sg13g2_o21ai_1 _1321_ (.B1(net1),
    .Y(_0428_),
    .A1(net234),
    .A2(_0424_));
 sg13g2_nor2_1 _1322_ (.A(net254),
    .B(net212),
    .Y(_0429_));
 sg13g2_nor3_1 _1323_ (.A(_0427_),
    .B(_0428_),
    .C(_0429_),
    .Y(_0039_));
 sg13g2_and2_1 _1324_ (.A(net7),
    .B(_0424_),
    .X(_0430_));
 sg13g2_and4_1 _1325_ (.A(net254),
    .B(net252),
    .C(net234),
    .D(net230),
    .X(_0431_));
 sg13g2_a22oi_1 _1326_ (.Y(_0432_),
    .B1(net229),
    .B2(net254),
    .A2(net234),
    .A1(net252));
 sg13g2_o21ai_1 _1327_ (.B1(net213),
    .Y(_0433_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_nand2b_1 _1328_ (.Y(_0434_),
    .B(net212),
    .A_N(net122));
 sg13g2_nand3_1 _1329_ (.B(_0433_),
    .C(_0434_),
    .A(net266),
    .Y(_0435_));
 sg13g2_a21oi_1 _1330_ (.A1(_0070_),
    .A2(net210),
    .Y(_0040_),
    .B1(_0435_));
 sg13g2_nand2_1 _1331_ (.Y(_0436_),
    .A(\i_decoder_a.data_out[0] ),
    .B(net226));
 sg13g2_and4_1 _1332_ (.A(net252),
    .B(net250),
    .C(net233),
    .D(net230),
    .X(_0437_));
 sg13g2_a22oi_1 _1333_ (.Y(_0438_),
    .B1(net230),
    .B2(net253),
    .A2(net233),
    .A1(net250));
 sg13g2_nor3_1 _1334_ (.A(_0436_),
    .B(_0437_),
    .C(_0438_),
    .Y(_0439_));
 sg13g2_o21ai_1 _1335_ (.B1(_0436_),
    .Y(_0440_),
    .A1(_0437_),
    .A2(_0438_));
 sg13g2_nor2b_1 _1336_ (.A(_0439_),
    .B_N(_0440_),
    .Y(_0441_));
 sg13g2_nand2_1 _1337_ (.Y(_0442_),
    .A(_0431_),
    .B(_0441_));
 sg13g2_o21ai_1 _1338_ (.B1(net213),
    .Y(_0443_),
    .A1(_0431_),
    .A2(_0441_));
 sg13g2_nand2b_1 _1339_ (.Y(_0444_),
    .B(_0442_),
    .A_N(_0443_));
 sg13g2_a22oi_1 _1340_ (.Y(_0445_),
    .B1(net210),
    .B2(net250),
    .A2(net212),
    .A1(net115));
 sg13g2_a21oi_1 _1341_ (.A1(_0444_),
    .A2(_0445_),
    .Y(_0041_),
    .B1(net258));
 sg13g2_nand2_2 _1342_ (.Y(_0446_),
    .A(\i_decoder_a.data_out[0] ),
    .B(net225));
 sg13g2_or2_1 _1343_ (.X(_0447_),
    .B(_0439_),
    .A(_0437_));
 sg13g2_nand2_1 _1344_ (.Y(_0448_),
    .A(net252),
    .B(\i_decoder_b.data_out[2] ));
 sg13g2_and4_1 _1345_ (.A(net250),
    .B(net248),
    .C(net233),
    .D(net229),
    .X(_0449_));
 sg13g2_nand4_1 _1346_ (.B(net248),
    .C(net233),
    .A(net250),
    .Y(_0450_),
    .D(net229));
 sg13g2_a22oi_1 _1347_ (.Y(_0451_),
    .B1(net229),
    .B2(net250),
    .A2(net233),
    .A1(net248));
 sg13g2_nor3_1 _1348_ (.A(_0448_),
    .B(_0449_),
    .C(_0451_),
    .Y(_0452_));
 sg13g2_o21ai_1 _1349_ (.B1(_0448_),
    .Y(_0453_),
    .A1(_0449_),
    .A2(_0451_));
 sg13g2_nor2b_1 _1350_ (.A(_0452_),
    .B_N(_0453_),
    .Y(_0454_));
 sg13g2_nand2_1 _1351_ (.Y(_0455_),
    .A(_0447_),
    .B(_0454_));
 sg13g2_xnor2_1 _1352_ (.Y(_0456_),
    .A(_0447_),
    .B(_0454_));
 sg13g2_xnor2_1 _1353_ (.Y(_0457_),
    .A(_0446_),
    .B(_0456_));
 sg13g2_or2_1 _1354_ (.X(_0458_),
    .B(_0457_),
    .A(_0442_));
 sg13g2_a21oi_1 _1355_ (.A1(_0442_),
    .A2(_0457_),
    .Y(_0459_),
    .B1(net214));
 sg13g2_nand2_1 _1356_ (.Y(_0460_),
    .A(_0458_),
    .B(_0459_));
 sg13g2_a22oi_1 _1357_ (.Y(_0461_),
    .B1(net210),
    .B2(net249),
    .A2(net212),
    .A1(net108));
 sg13g2_a21oi_1 _1358_ (.A1(_0460_),
    .A2(net109),
    .Y(_0042_),
    .B1(net258));
 sg13g2_nand2_2 _1359_ (.Y(_0462_),
    .A(net252),
    .B(net222));
 sg13g2_nor2_1 _1360_ (.A(_0446_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_or2_1 _1361_ (.X(_0464_),
    .B(_0462_),
    .A(_0446_));
 sg13g2_a22oi_1 _1362_ (.Y(_0465_),
    .B1(net222),
    .B2(net254),
    .A2(net225),
    .A1(net252));
 sg13g2_or2_1 _1363_ (.X(_0466_),
    .B(_0465_),
    .A(_0463_));
 sg13g2_o21ai_1 _1364_ (.B1(_0450_),
    .Y(_0467_),
    .A1(_0448_),
    .A2(_0451_));
 sg13g2_nand2_1 _1365_ (.Y(_0468_),
    .A(net250),
    .B(\i_decoder_b.data_out[2] ));
 sg13g2_and4_1 _1366_ (.A(net248),
    .B(net246),
    .C(net233),
    .D(net229),
    .X(_0469_));
 sg13g2_nand4_1 _1367_ (.B(net246),
    .C(net233),
    .A(net248),
    .Y(_0470_),
    .D(net229));
 sg13g2_a22oi_1 _1368_ (.Y(_0471_),
    .B1(net229),
    .B2(net248),
    .A2(net233),
    .A1(net246));
 sg13g2_or3_1 _1369_ (.A(_0468_),
    .B(_0469_),
    .C(_0471_),
    .X(_0472_));
 sg13g2_o21ai_1 _1370_ (.B1(_0468_),
    .Y(_0473_),
    .A1(_0469_),
    .A2(_0471_));
 sg13g2_nand3_1 _1371_ (.B(_0472_),
    .C(_0473_),
    .A(_0467_),
    .Y(_0474_));
 sg13g2_a21oi_1 _1372_ (.A1(_0472_),
    .A2(_0473_),
    .Y(_0475_),
    .B1(_0467_));
 sg13g2_a21o_1 _1373_ (.A2(_0473_),
    .A1(_0472_),
    .B1(_0467_),
    .X(_0476_));
 sg13g2_nand2_1 _1374_ (.Y(_0477_),
    .A(_0474_),
    .B(_0476_));
 sg13g2_xnor2_1 _1375_ (.Y(_0478_),
    .A(_0466_),
    .B(_0477_));
 sg13g2_o21ai_1 _1376_ (.B1(_0455_),
    .Y(_0479_),
    .A1(_0446_),
    .A2(_0456_));
 sg13g2_nand2b_1 _1377_ (.Y(_0480_),
    .B(_0479_),
    .A_N(_0478_));
 sg13g2_xor2_1 _1378_ (.B(_0479_),
    .A(_0478_),
    .X(_0481_));
 sg13g2_and2_1 _1379_ (.A(_0458_),
    .B(_0481_),
    .X(_0482_));
 sg13g2_nor2_1 _1380_ (.A(_0458_),
    .B(_0481_),
    .Y(_0483_));
 sg13g2_or3_1 _1381_ (.A(net214),
    .B(_0482_),
    .C(_0483_),
    .X(_0484_));
 sg13g2_a22oi_1 _1382_ (.Y(_0485_),
    .B1(net210),
    .B2(net246),
    .A2(net212),
    .A1(net114));
 sg13g2_a21oi_1 _1383_ (.A1(_0484_),
    .A2(_0485_),
    .Y(_0043_),
    .B1(net257));
 sg13g2_o21ai_1 _1384_ (.B1(_0474_),
    .Y(_0486_),
    .A1(_0466_),
    .A2(_0475_));
 sg13g2_nand2_1 _1385_ (.Y(_0487_),
    .A(net254),
    .B(net220));
 sg13g2_nand2_1 _1386_ (.Y(_0488_),
    .A(net251),
    .B(net222));
 sg13g2_nand2_1 _1387_ (.Y(_0489_),
    .A(net251),
    .B(net224));
 sg13g2_xor2_1 _1388_ (.B(_0489_),
    .A(_0462_),
    .X(_0490_));
 sg13g2_nand2b_1 _1389_ (.Y(_0491_),
    .B(_0490_),
    .A_N(_0487_));
 sg13g2_xor2_1 _1390_ (.B(_0490_),
    .A(_0487_),
    .X(_0492_));
 sg13g2_o21ai_1 _1391_ (.B1(_0470_),
    .Y(_0493_),
    .A1(_0468_),
    .A2(_0471_));
 sg13g2_nand2_1 _1392_ (.Y(_0494_),
    .A(net248),
    .B(net226));
 sg13g2_and4_1 _1393_ (.A(net246),
    .B(net245),
    .C(net235),
    .D(net228),
    .X(_0495_));
 sg13g2_nand4_1 _1394_ (.B(net244),
    .C(net232),
    .A(net246),
    .Y(_0496_),
    .D(net228));
 sg13g2_a22oi_1 _1395_ (.Y(_0497_),
    .B1(net228),
    .B2(net246),
    .A2(net232),
    .A1(net245));
 sg13g2_or3_1 _1396_ (.A(_0494_),
    .B(_0495_),
    .C(_0497_),
    .X(_0498_));
 sg13g2_o21ai_1 _1397_ (.B1(_0494_),
    .Y(_0499_),
    .A1(_0495_),
    .A2(_0497_));
 sg13g2_and3_1 _1398_ (.X(_0500_),
    .A(_0493_),
    .B(_0498_),
    .C(_0499_));
 sg13g2_nand3_1 _1399_ (.B(_0498_),
    .C(_0499_),
    .A(_0493_),
    .Y(_0501_));
 sg13g2_a21oi_1 _1400_ (.A1(_0498_),
    .A2(_0499_),
    .Y(_0502_),
    .B1(_0493_));
 sg13g2_or3_1 _1401_ (.A(_0492_),
    .B(_0500_),
    .C(_0502_),
    .X(_0503_));
 sg13g2_o21ai_1 _1402_ (.B1(_0492_),
    .Y(_0504_),
    .A1(_0500_),
    .A2(_0502_));
 sg13g2_nand3_1 _1403_ (.B(_0503_),
    .C(_0504_),
    .A(_0486_),
    .Y(_0505_));
 sg13g2_a21oi_1 _1404_ (.A1(_0503_),
    .A2(_0504_),
    .Y(_0506_),
    .B1(_0486_));
 sg13g2_a21o_1 _1405_ (.A2(_0504_),
    .A1(_0503_),
    .B1(_0486_),
    .X(_0507_));
 sg13g2_and3_1 _1406_ (.X(_0508_),
    .A(_0463_),
    .B(_0505_),
    .C(_0507_));
 sg13g2_a21oi_1 _1407_ (.A1(_0505_),
    .A2(_0507_),
    .Y(_0509_),
    .B1(_0463_));
 sg13g2_nor3_1 _1408_ (.A(_0480_),
    .B(_0508_),
    .C(_0509_),
    .Y(_0510_));
 sg13g2_or3_1 _1409_ (.A(_0480_),
    .B(_0508_),
    .C(_0509_),
    .X(_0511_));
 sg13g2_o21ai_1 _1410_ (.B1(_0480_),
    .Y(_0512_),
    .A1(_0508_),
    .A2(_0509_));
 sg13g2_nand3_1 _1411_ (.B(_0511_),
    .C(_0512_),
    .A(_0483_),
    .Y(_0513_));
 sg13g2_a21o_1 _1412_ (.A2(_0512_),
    .A1(_0511_),
    .B1(_0483_),
    .X(_0514_));
 sg13g2_nand3_1 _1413_ (.B(_0513_),
    .C(_0514_),
    .A(net213),
    .Y(_0515_));
 sg13g2_a22oi_1 _1414_ (.Y(_0516_),
    .B1(net210),
    .B2(net245),
    .A2(net212),
    .A1(net102));
 sg13g2_a21oi_1 _1415_ (.A1(_0515_),
    .A2(net103),
    .Y(_0044_),
    .B1(net257));
 sg13g2_o21ai_1 _1416_ (.B1(_0505_),
    .Y(_0517_),
    .A1(_0464_),
    .A2(_0506_));
 sg13g2_o21ai_1 _1417_ (.B1(_0491_),
    .Y(_0518_),
    .A1(_0462_),
    .A2(_0489_));
 sg13g2_nand2_1 _1418_ (.Y(_0519_),
    .A(net254),
    .B(net218));
 sg13g2_nor2b_1 _1419_ (.A(_0519_),
    .B_N(_0518_),
    .Y(_0520_));
 sg13g2_xor2_1 _1420_ (.B(_0519_),
    .A(_0518_),
    .X(_0521_));
 sg13g2_o21ai_1 _1421_ (.B1(_0501_),
    .Y(_0522_),
    .A1(_0492_),
    .A2(_0502_));
 sg13g2_nand2_1 _1422_ (.Y(_0523_),
    .A(net253),
    .B(net220));
 sg13g2_nand2_1 _1423_ (.Y(_0524_),
    .A(net249),
    .B(net222));
 sg13g2_nand2_1 _1424_ (.Y(_0525_),
    .A(net249),
    .B(net223));
 sg13g2_or2_1 _1425_ (.X(_0526_),
    .B(_0524_),
    .A(_0489_));
 sg13g2_xnor2_1 _1426_ (.Y(_0527_),
    .A(_0488_),
    .B(_0525_));
 sg13g2_xnor2_1 _1427_ (.Y(_0528_),
    .A(_0523_),
    .B(_0527_));
 sg13g2_o21ai_1 _1428_ (.B1(_0496_),
    .Y(_0529_),
    .A1(_0494_),
    .A2(_0497_));
 sg13g2_nand2_1 _1429_ (.Y(_0530_),
    .A(net247),
    .B(net226));
 sg13g2_and4_1 _1430_ (.A(net243),
    .B(net241),
    .C(net232),
    .D(net228),
    .X(_0531_));
 sg13g2_nand4_1 _1431_ (.B(net241),
    .C(net232),
    .A(net243),
    .Y(_0532_),
    .D(net227));
 sg13g2_a22oi_1 _1432_ (.Y(_0533_),
    .B1(net227),
    .B2(net243),
    .A2(net232),
    .A1(net241));
 sg13g2_or3_1 _1433_ (.A(_0530_),
    .B(_0531_),
    .C(_0533_),
    .X(_0534_));
 sg13g2_o21ai_1 _1434_ (.B1(_0530_),
    .Y(_0535_),
    .A1(_0531_),
    .A2(_0533_));
 sg13g2_and3_1 _1435_ (.X(_0536_),
    .A(_0529_),
    .B(_0534_),
    .C(_0535_));
 sg13g2_nand3_1 _1436_ (.B(_0534_),
    .C(_0535_),
    .A(_0529_),
    .Y(_0537_));
 sg13g2_a21oi_1 _1437_ (.A1(_0534_),
    .A2(_0535_),
    .Y(_0538_),
    .B1(_0529_));
 sg13g2_or3_1 _1438_ (.A(_0528_),
    .B(_0536_),
    .C(_0538_),
    .X(_0539_));
 sg13g2_o21ai_1 _1439_ (.B1(_0528_),
    .Y(_0540_),
    .A1(_0536_),
    .A2(_0538_));
 sg13g2_and3_1 _1440_ (.X(_0541_),
    .A(_0522_),
    .B(_0539_),
    .C(_0540_));
 sg13g2_nand3_1 _1441_ (.B(_0539_),
    .C(_0540_),
    .A(_0522_),
    .Y(_0542_));
 sg13g2_a21oi_1 _1442_ (.A1(_0539_),
    .A2(_0540_),
    .Y(_0543_),
    .B1(_0522_));
 sg13g2_or3_1 _1443_ (.A(_0521_),
    .B(_0541_),
    .C(_0543_),
    .X(_0544_));
 sg13g2_o21ai_1 _1444_ (.B1(_0521_),
    .Y(_0545_),
    .A1(_0541_),
    .A2(_0543_));
 sg13g2_a21o_1 _1445_ (.A2(_0545_),
    .A1(_0544_),
    .B1(_0517_),
    .X(_0546_));
 sg13g2_and3_1 _1446_ (.X(_0547_),
    .A(_0517_),
    .B(_0544_),
    .C(_0545_));
 sg13g2_nand3_1 _1447_ (.B(_0544_),
    .C(_0545_),
    .A(_0517_),
    .Y(_0548_));
 sg13g2_nand3_1 _1448_ (.B(_0546_),
    .C(_0548_),
    .A(_0510_),
    .Y(_0549_));
 sg13g2_a21oi_1 _1449_ (.A1(_0546_),
    .A2(_0548_),
    .Y(_0550_),
    .B1(_0510_));
 sg13g2_a21o_1 _1450_ (.A2(_0548_),
    .A1(_0546_),
    .B1(_0510_),
    .X(_0551_));
 sg13g2_nand2_1 _1451_ (.Y(_0552_),
    .A(_0549_),
    .B(_0551_));
 sg13g2_a21oi_1 _1452_ (.A1(_0513_),
    .A2(_0552_),
    .Y(_0553_),
    .B1(net214));
 sg13g2_o21ai_1 _1453_ (.B1(_0553_),
    .Y(_0554_),
    .A1(_0513_),
    .A2(_0552_));
 sg13g2_a22oi_1 _1454_ (.Y(_0555_),
    .B1(net210),
    .B2(net242),
    .A2(net212),
    .A1(net120));
 sg13g2_a21oi_1 _1455_ (.A1(_0554_),
    .A2(net121),
    .Y(_0045_),
    .B1(net257));
 sg13g2_o21ai_1 _1456_ (.B1(_0542_),
    .Y(_0556_),
    .A1(_0521_),
    .A2(_0543_));
 sg13g2_nand2_1 _1457_ (.Y(_0557_),
    .A(net254),
    .B(net216));
 sg13g2_o21ai_1 _1458_ (.B1(_0526_),
    .Y(_0558_),
    .A1(_0523_),
    .A2(_0527_));
 sg13g2_nand2_1 _1459_ (.Y(_0559_),
    .A(net253),
    .B(net218));
 sg13g2_nand2b_1 _1460_ (.Y(_0560_),
    .B(_0558_),
    .A_N(_0559_));
 sg13g2_xnor2_1 _1461_ (.Y(_0561_),
    .A(_0558_),
    .B(_0559_));
 sg13g2_nand2b_1 _1462_ (.Y(_0562_),
    .B(_0561_),
    .A_N(_0557_));
 sg13g2_xor2_1 _1463_ (.B(_0561_),
    .A(_0557_),
    .X(_0563_));
 sg13g2_o21ai_1 _1464_ (.B1(_0537_),
    .Y(_0564_),
    .A1(_0528_),
    .A2(_0538_));
 sg13g2_nand2_1 _1465_ (.Y(_0565_),
    .A(net251),
    .B(net219));
 sg13g2_nand2_1 _1466_ (.Y(_0566_),
    .A(net247),
    .B(net221));
 sg13g2_nand2_1 _1467_ (.Y(_0567_),
    .A(net247),
    .B(net224));
 sg13g2_or2_1 _1468_ (.X(_0568_),
    .B(_0566_),
    .A(_0525_));
 sg13g2_xnor2_1 _1469_ (.Y(_0569_),
    .A(_0524_),
    .B(_0567_));
 sg13g2_xnor2_1 _1470_ (.Y(_0570_),
    .A(_0565_),
    .B(_0569_));
 sg13g2_o21ai_1 _1471_ (.B1(_0532_),
    .Y(_0571_),
    .A1(_0530_),
    .A2(_0533_));
 sg13g2_nand2_1 _1472_ (.Y(_0572_),
    .A(net243),
    .B(net226));
 sg13g2_nand2_1 _1473_ (.Y(_0573_),
    .A(net237),
    .B(net227));
 sg13g2_and4_1 _1474_ (.A(net240),
    .B(net237),
    .C(net232),
    .D(net227),
    .X(_0574_));
 sg13g2_nand4_1 _1475_ (.B(net237),
    .C(net232),
    .A(net240),
    .Y(_0575_),
    .D(net227));
 sg13g2_a22oi_1 _1476_ (.Y(_0576_),
    .B1(net227),
    .B2(net240),
    .A2(net232),
    .A1(net237));
 sg13g2_or3_1 _1477_ (.A(_0572_),
    .B(_0574_),
    .C(_0576_),
    .X(_0577_));
 sg13g2_o21ai_1 _1478_ (.B1(_0572_),
    .Y(_0578_),
    .A1(_0574_),
    .A2(_0576_));
 sg13g2_and3_1 _1479_ (.X(_0579_),
    .A(_0571_),
    .B(_0577_),
    .C(_0578_));
 sg13g2_nand3_1 _1480_ (.B(_0577_),
    .C(_0578_),
    .A(_0571_),
    .Y(_0580_));
 sg13g2_a21oi_1 _1481_ (.A1(_0577_),
    .A2(_0578_),
    .Y(_0581_),
    .B1(_0571_));
 sg13g2_or3_1 _1482_ (.A(_0570_),
    .B(_0579_),
    .C(_0581_),
    .X(_0582_));
 sg13g2_o21ai_1 _1483_ (.B1(_0570_),
    .Y(_0583_),
    .A1(_0579_),
    .A2(_0581_));
 sg13g2_and3_1 _1484_ (.X(_0584_),
    .A(_0564_),
    .B(_0582_),
    .C(_0583_));
 sg13g2_nand3_1 _1485_ (.B(_0582_),
    .C(_0583_),
    .A(_0564_),
    .Y(_0585_));
 sg13g2_a21oi_1 _1486_ (.A1(_0582_),
    .A2(_0583_),
    .Y(_0586_),
    .B1(_0564_));
 sg13g2_or3_1 _1487_ (.A(_0563_),
    .B(_0584_),
    .C(_0586_),
    .X(_0587_));
 sg13g2_o21ai_1 _1488_ (.B1(_0563_),
    .Y(_0588_),
    .A1(_0584_),
    .A2(_0586_));
 sg13g2_and3_1 _1489_ (.X(_0589_),
    .A(_0556_),
    .B(_0587_),
    .C(_0588_));
 sg13g2_nand3_1 _1490_ (.B(_0587_),
    .C(_0588_),
    .A(_0556_),
    .Y(_0590_));
 sg13g2_a21o_1 _1491_ (.A2(_0588_),
    .A1(_0587_),
    .B1(_0556_),
    .X(_0591_));
 sg13g2_nand3_1 _1492_ (.B(_0590_),
    .C(_0591_),
    .A(_0520_),
    .Y(_0592_));
 sg13g2_a21o_1 _1493_ (.A2(_0591_),
    .A1(_0590_),
    .B1(_0520_),
    .X(_0593_));
 sg13g2_and3_1 _1494_ (.X(_0594_),
    .A(_0547_),
    .B(_0592_),
    .C(_0593_));
 sg13g2_nand3_1 _1495_ (.B(_0592_),
    .C(_0593_),
    .A(_0547_),
    .Y(_0595_));
 sg13g2_a21o_1 _1496_ (.A2(_0593_),
    .A1(_0592_),
    .B1(_0547_),
    .X(_0596_));
 sg13g2_o21ai_1 _1497_ (.B1(_0549_),
    .Y(_0597_),
    .A1(_0513_),
    .A2(_0550_));
 sg13g2_a21oi_1 _1498_ (.A1(_0595_),
    .A2(_0596_),
    .Y(_0598_),
    .B1(_0597_));
 sg13g2_nand3_1 _1499_ (.B(_0596_),
    .C(_0597_),
    .A(_0595_),
    .Y(_0599_));
 sg13g2_nand2_1 _1500_ (.Y(_0600_),
    .A(net213),
    .B(_0599_));
 sg13g2_a22oi_1 _1501_ (.Y(_0601_),
    .B1(net210),
    .B2(net239),
    .A2(net212),
    .A1(net128));
 sg13g2_o21ai_1 _1502_ (.B1(net129),
    .Y(_0602_),
    .A1(_0598_),
    .A2(_0600_));
 sg13g2_and2_1 _1503_ (.A(net265),
    .B(_0602_),
    .X(_0046_));
 sg13g2_a21oi_1 _1504_ (.A1(_0520_),
    .A2(_0591_),
    .Y(_0603_),
    .B1(_0589_));
 sg13g2_nand2_1 _1505_ (.Y(_0604_),
    .A(_0560_),
    .B(_0562_));
 sg13g2_o21ai_1 _1506_ (.B1(_0585_),
    .Y(_0605_),
    .A1(_0563_),
    .A2(_0586_));
 sg13g2_nand2_1 _1507_ (.Y(_0606_),
    .A(net253),
    .B(net215));
 sg13g2_o21ai_1 _1508_ (.B1(_0568_),
    .Y(_0607_),
    .A1(_0565_),
    .A2(_0569_));
 sg13g2_nand2_1 _1509_ (.Y(_0608_),
    .A(net251),
    .B(net217));
 sg13g2_nand2b_1 _1510_ (.Y(_0609_),
    .B(_0607_),
    .A_N(_0608_));
 sg13g2_xnor2_1 _1511_ (.Y(_0610_),
    .A(_0607_),
    .B(_0608_));
 sg13g2_nand2b_1 _1512_ (.Y(_0611_),
    .B(_0610_),
    .A_N(_0606_));
 sg13g2_xor2_1 _1513_ (.B(_0610_),
    .A(_0606_),
    .X(_0612_));
 sg13g2_o21ai_1 _1514_ (.B1(_0580_),
    .Y(_0613_),
    .A1(_0570_),
    .A2(_0581_));
 sg13g2_nand2_1 _1515_ (.Y(_0614_),
    .A(net249),
    .B(net219));
 sg13g2_nand2_1 _1516_ (.Y(_0615_),
    .A(net243),
    .B(net223));
 sg13g2_or2_1 _1517_ (.X(_0616_),
    .B(_0615_),
    .A(_0566_));
 sg13g2_xnor2_1 _1518_ (.Y(_0617_),
    .A(_0566_),
    .B(_0615_));
 sg13g2_xnor2_1 _1519_ (.Y(_0618_),
    .A(_0614_),
    .B(_0617_));
 sg13g2_o21ai_1 _1520_ (.B1(_0575_),
    .Y(_0619_),
    .A1(_0572_),
    .A2(_0576_));
 sg13g2_nand2_1 _1521_ (.Y(_0620_),
    .A(net240),
    .B(net226));
 sg13g2_nand2_1 _1522_ (.Y(_0621_),
    .A(net237),
    .B(net226));
 sg13g2_or2_1 _1523_ (.X(_0622_),
    .B(_0620_),
    .A(_0573_));
 sg13g2_xor2_1 _1524_ (.B(_0620_),
    .A(_0573_),
    .X(_0623_));
 sg13g2_nand2_1 _1525_ (.Y(_0624_),
    .A(_0619_),
    .B(_0623_));
 sg13g2_xnor2_1 _1526_ (.Y(_0625_),
    .A(_0619_),
    .B(_0623_));
 sg13g2_xnor2_1 _1527_ (.Y(_0626_),
    .A(_0618_),
    .B(_0625_));
 sg13g2_nand2b_1 _1528_ (.Y(_0627_),
    .B(_0613_),
    .A_N(_0626_));
 sg13g2_xor2_1 _1529_ (.B(_0626_),
    .A(_0613_),
    .X(_0628_));
 sg13g2_xnor2_1 _1530_ (.Y(_0629_),
    .A(_0612_),
    .B(_0628_));
 sg13g2_nor2b_1 _1531_ (.A(_0629_),
    .B_N(_0605_),
    .Y(_0630_));
 sg13g2_xnor2_1 _1532_ (.Y(_0631_),
    .A(_0605_),
    .B(_0629_));
 sg13g2_xnor2_1 _1533_ (.Y(_0632_),
    .A(_0604_),
    .B(_0631_));
 sg13g2_nor2_1 _1534_ (.A(_0603_),
    .B(_0632_),
    .Y(_0633_));
 sg13g2_xnor2_1 _1535_ (.Y(_0634_),
    .A(_0603_),
    .B(_0632_));
 sg13g2_a21oi_2 _1536_ (.B1(_0594_),
    .Y(_0635_),
    .A2(_0597_),
    .A1(_0596_));
 sg13g2_and2_1 _1537_ (.A(_0634_),
    .B(_0635_),
    .X(_0636_));
 sg13g2_nor2_1 _1538_ (.A(_0634_),
    .B(_0635_),
    .Y(_0637_));
 sg13g2_or3_1 _1539_ (.A(net214),
    .B(_0636_),
    .C(_0637_),
    .X(_0638_));
 sg13g2_a22oi_1 _1540_ (.Y(_0639_),
    .B1(net209),
    .B2(net235),
    .A2(net211),
    .A1(net106));
 sg13g2_a21oi_1 _1541_ (.A1(_0638_),
    .A2(net107),
    .Y(_0047_),
    .B1(net258));
 sg13g2_nor2_1 _1542_ (.A(_0633_),
    .B(_0637_),
    .Y(_0640_));
 sg13g2_a21oi_2 _1543_ (.B1(_0630_),
    .Y(_0641_),
    .A2(_0631_),
    .A1(_0604_));
 sg13g2_nand2_1 _1544_ (.Y(_0642_),
    .A(_0609_),
    .B(_0611_));
 sg13g2_o21ai_1 _1545_ (.B1(_0627_),
    .Y(_0643_),
    .A1(_0612_),
    .A2(_0628_));
 sg13g2_nand2_1 _1546_ (.Y(_0644_),
    .A(net251),
    .B(net215));
 sg13g2_o21ai_1 _1547_ (.B1(_0616_),
    .Y(_0645_),
    .A1(_0614_),
    .A2(_0617_));
 sg13g2_nand2_1 _1548_ (.Y(_0646_),
    .A(net249),
    .B(net217));
 sg13g2_nand2b_1 _1549_ (.Y(_0647_),
    .B(_0645_),
    .A_N(_0646_));
 sg13g2_xnor2_1 _1550_ (.Y(_0648_),
    .A(_0645_),
    .B(_0646_));
 sg13g2_nand2b_1 _1551_ (.Y(_0649_),
    .B(_0648_),
    .A_N(_0644_));
 sg13g2_xnor2_1 _1552_ (.Y(_0650_),
    .A(_0644_),
    .B(_0648_));
 sg13g2_o21ai_1 _1553_ (.B1(_0624_),
    .Y(_0651_),
    .A1(_0618_),
    .A2(_0625_));
 sg13g2_a21oi_1 _1554_ (.A1(net240),
    .A2(net227),
    .Y(_0652_),
    .B1(_0621_));
 sg13g2_nand2_1 _1555_ (.Y(_0653_),
    .A(net247),
    .B(net219));
 sg13g2_nand2_1 _1556_ (.Y(_0654_),
    .A(net241),
    .B(net221));
 sg13g2_and4_1 _1557_ (.A(net243),
    .B(net240),
    .C(net223),
    .D(net221),
    .X(_0655_));
 sg13g2_nand4_1 _1558_ (.B(net240),
    .C(net223),
    .A(net243),
    .Y(_0656_),
    .D(net221));
 sg13g2_a22oi_1 _1559_ (.Y(_0657_),
    .B1(net221),
    .B2(net243),
    .A2(net223),
    .A1(net240));
 sg13g2_or3_1 _1560_ (.A(_0653_),
    .B(_0655_),
    .C(_0657_),
    .X(_0658_));
 sg13g2_o21ai_1 _1561_ (.B1(_0653_),
    .Y(_0659_),
    .A1(_0655_),
    .A2(_0657_));
 sg13g2_nand3_1 _1562_ (.B(_0658_),
    .C(_0659_),
    .A(_0652_),
    .Y(_0660_));
 sg13g2_a21o_1 _1563_ (.A2(_0659_),
    .A1(_0658_),
    .B1(_0652_),
    .X(_0661_));
 sg13g2_nand2_1 _1564_ (.Y(_0662_),
    .A(_0660_),
    .B(_0661_));
 sg13g2_nor2b_1 _1565_ (.A(_0662_),
    .B_N(_0651_),
    .Y(_0663_));
 sg13g2_xnor2_1 _1566_ (.Y(_0664_),
    .A(_0651_),
    .B(_0662_));
 sg13g2_xnor2_1 _1567_ (.Y(_0665_),
    .A(_0650_),
    .B(_0664_));
 sg13g2_nor2b_1 _1568_ (.A(_0665_),
    .B_N(_0643_),
    .Y(_0666_));
 sg13g2_xnor2_1 _1569_ (.Y(_0667_),
    .A(_0643_),
    .B(_0665_));
 sg13g2_xnor2_1 _1570_ (.Y(_0668_),
    .A(_0642_),
    .B(_0667_));
 sg13g2_nor2_1 _1571_ (.A(_0641_),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_xnor2_1 _1572_ (.Y(_0670_),
    .A(_0641_),
    .B(_0668_));
 sg13g2_a21oi_1 _1573_ (.A1(_0640_),
    .A2(_0670_),
    .Y(_0671_),
    .B1(net214));
 sg13g2_o21ai_1 _1574_ (.B1(_0671_),
    .Y(_0672_),
    .A1(_0640_),
    .A2(_0670_));
 sg13g2_a22oi_1 _1575_ (.Y(_0673_),
    .B1(net209),
    .B2(net227),
    .A2(net211),
    .A1(net110));
 sg13g2_a21oi_1 _1576_ (.A1(_0672_),
    .A2(_0673_),
    .Y(_0048_),
    .B1(net256));
 sg13g2_a21oi_1 _1577_ (.A1(_0642_),
    .A2(_0667_),
    .Y(_0674_),
    .B1(_0666_));
 sg13g2_nand2_1 _1578_ (.Y(_0675_),
    .A(_0647_),
    .B(_0649_));
 sg13g2_a21oi_1 _1579_ (.A1(_0650_),
    .A2(_0664_),
    .Y(_0676_),
    .B1(_0663_));
 sg13g2_nand2_1 _1580_ (.Y(_0677_),
    .A(net249),
    .B(net215));
 sg13g2_o21ai_1 _1581_ (.B1(_0656_),
    .Y(_0678_),
    .A1(_0653_),
    .A2(_0657_));
 sg13g2_nand2_1 _1582_ (.Y(_0679_),
    .A(net247),
    .B(net217));
 sg13g2_nand2b_1 _1583_ (.Y(_0680_),
    .B(_0678_),
    .A_N(_0679_));
 sg13g2_xnor2_1 _1584_ (.Y(_0681_),
    .A(_0678_),
    .B(_0679_));
 sg13g2_nand2b_1 _1585_ (.Y(_0682_),
    .B(_0681_),
    .A_N(_0677_));
 sg13g2_xnor2_1 _1586_ (.Y(_0683_),
    .A(_0677_),
    .B(_0681_));
 sg13g2_nand2_1 _1587_ (.Y(_0684_),
    .A(net244),
    .B(net219));
 sg13g2_nand2_1 _1588_ (.Y(_0685_),
    .A(net238),
    .B(net223));
 sg13g2_nand4_1 _1589_ (.B(net238),
    .C(net223),
    .A(net241),
    .Y(_0686_),
    .D(net221));
 sg13g2_a22oi_1 _1590_ (.Y(_0687_),
    .B1(net221),
    .B2(net241),
    .A2(net223),
    .A1(net238));
 sg13g2_xnor2_1 _1591_ (.Y(_0688_),
    .A(_0654_),
    .B(_0685_));
 sg13g2_xnor2_1 _1592_ (.Y(_0689_),
    .A(_0684_),
    .B(_0688_));
 sg13g2_a21oi_1 _1593_ (.A1(_0622_),
    .A2(_0660_),
    .Y(_0690_),
    .B1(_0689_));
 sg13g2_nand3_1 _1594_ (.B(_0660_),
    .C(_0689_),
    .A(_0622_),
    .Y(_0691_));
 sg13g2_nand2b_1 _1595_ (.Y(_0692_),
    .B(_0691_),
    .A_N(_0690_));
 sg13g2_xor2_1 _1596_ (.B(_0692_),
    .A(_0683_),
    .X(_0693_));
 sg13g2_nor2_1 _1597_ (.A(_0676_),
    .B(_0693_),
    .Y(_0694_));
 sg13g2_xor2_1 _1598_ (.B(_0693_),
    .A(_0676_),
    .X(_0695_));
 sg13g2_xnor2_1 _1599_ (.Y(_0696_),
    .A(_0675_),
    .B(_0695_));
 sg13g2_nand2_1 _1600_ (.Y(_0697_),
    .A(_0674_),
    .B(_0696_));
 sg13g2_or2_1 _1601_ (.X(_0698_),
    .B(_0696_),
    .A(_0674_));
 sg13g2_and2_1 _1602_ (.A(_0697_),
    .B(_0698_),
    .X(_0699_));
 sg13g2_or2_1 _1603_ (.X(_0700_),
    .B(_0670_),
    .A(_0634_));
 sg13g2_nor2_1 _1604_ (.A(_0635_),
    .B(_0700_),
    .Y(_0701_));
 sg13g2_a221oi_1 _1605_ (.B2(_0668_),
    .C1(_0632_),
    .B1(_0641_),
    .A1(_0590_),
    .Y(_0702_),
    .A2(_0592_));
 sg13g2_or2_1 _1606_ (.X(_0703_),
    .B(_0702_),
    .A(_0669_));
 sg13g2_o21ai_1 _1607_ (.B1(_0699_),
    .Y(_0704_),
    .A1(_0701_),
    .A2(_0703_));
 sg13g2_nor3_1 _1608_ (.A(_0699_),
    .B(_0701_),
    .C(_0703_),
    .Y(_0705_));
 sg13g2_nor2_1 _1609_ (.A(net214),
    .B(_0705_),
    .Y(_0706_));
 sg13g2_nand2_1 _1610_ (.Y(_0707_),
    .A(_0704_),
    .B(_0706_));
 sg13g2_a22oi_1 _1611_ (.Y(_0708_),
    .B1(net209),
    .B2(net226),
    .A2(net211),
    .A1(net113));
 sg13g2_a21oi_1 _1612_ (.A1(_0707_),
    .A2(_0708_),
    .Y(_0049_),
    .B1(net256));
 sg13g2_a21oi_1 _1613_ (.A1(_0675_),
    .A2(_0695_),
    .Y(_0709_),
    .B1(_0694_));
 sg13g2_nand2_1 _1614_ (.Y(_0710_),
    .A(_0680_),
    .B(_0682_));
 sg13g2_nand2_1 _1615_ (.Y(_0711_),
    .A(net237),
    .B(net219));
 sg13g2_nor2_1 _1616_ (.A(_0654_),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_a22oi_1 _1617_ (.Y(_0713_),
    .B1(net219),
    .B2(net242),
    .A2(net221),
    .A1(net237));
 sg13g2_nor2_1 _1618_ (.A(_0712_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_nand2_1 _1619_ (.Y(_0715_),
    .A(net247),
    .B(net215));
 sg13g2_o21ai_1 _1620_ (.B1(_0686_),
    .Y(_0716_),
    .A1(_0684_),
    .A2(_0687_));
 sg13g2_nand2_1 _1621_ (.Y(_0717_),
    .A(net244),
    .B(net217));
 sg13g2_nand2b_1 _1622_ (.Y(_0718_),
    .B(_0716_),
    .A_N(_0717_));
 sg13g2_xnor2_1 _1623_ (.Y(_0719_),
    .A(_0716_),
    .B(_0717_));
 sg13g2_nand2b_1 _1624_ (.Y(_0720_),
    .B(_0719_),
    .A_N(_0715_));
 sg13g2_xnor2_1 _1625_ (.Y(_0721_),
    .A(_0715_),
    .B(_0719_));
 sg13g2_nand2_1 _1626_ (.Y(_0722_),
    .A(_0714_),
    .B(_0721_));
 sg13g2_xnor2_1 _1627_ (.Y(_0723_),
    .A(_0714_),
    .B(_0721_));
 sg13g2_a21oi_1 _1628_ (.A1(_0683_),
    .A2(_0691_),
    .Y(_0724_),
    .B1(_0690_));
 sg13g2_nor2_1 _1629_ (.A(_0723_),
    .B(_0724_),
    .Y(_0725_));
 sg13g2_xnor2_1 _1630_ (.Y(_0726_),
    .A(_0723_),
    .B(_0724_));
 sg13g2_nand2b_1 _1631_ (.Y(_0727_),
    .B(_0710_),
    .A_N(_0726_));
 sg13g2_nand2b_1 _1632_ (.Y(_0728_),
    .B(_0726_),
    .A_N(_0710_));
 sg13g2_nand2_1 _1633_ (.Y(_0729_),
    .A(_0727_),
    .B(_0728_));
 sg13g2_a221oi_1 _1634_ (.B2(_0728_),
    .C1(_0694_),
    .B1(_0727_),
    .A1(_0675_),
    .Y(_0730_),
    .A2(_0695_));
 sg13g2_nor2_1 _1635_ (.A(_0709_),
    .B(_0729_),
    .Y(_0731_));
 sg13g2_or2_1 _1636_ (.X(_0732_),
    .B(_0731_),
    .A(_0730_));
 sg13g2_nand3_1 _1637_ (.B(_0704_),
    .C(_0732_),
    .A(_0698_),
    .Y(_0733_));
 sg13g2_a21o_1 _1638_ (.A2(_0704_),
    .A1(_0698_),
    .B1(_0732_),
    .X(_0734_));
 sg13g2_nand3_1 _1639_ (.B(_0733_),
    .C(_0734_),
    .A(net213),
    .Y(_0735_));
 sg13g2_a22oi_1 _1640_ (.Y(_0736_),
    .B1(net209),
    .B2(net224),
    .A2(net211),
    .A1(net111));
 sg13g2_a21oi_1 _1641_ (.A1(_0735_),
    .A2(_0736_),
    .Y(_0050_),
    .B1(net256));
 sg13g2_nor2b_1 _1642_ (.A(_0725_),
    .B_N(_0727_),
    .Y(_0737_));
 sg13g2_nand2_1 _1643_ (.Y(_0738_),
    .A(net242),
    .B(net218));
 sg13g2_mux2_1 _1644_ (.A0(_0738_),
    .A1(net217),
    .S(_0712_),
    .X(_0739_));
 sg13g2_nand2_1 _1645_ (.Y(_0740_),
    .A(net244),
    .B(net215));
 sg13g2_nor2_1 _1646_ (.A(_0739_),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_xor2_1 _1647_ (.B(_0740_),
    .A(_0739_),
    .X(_0742_));
 sg13g2_nand2b_1 _1648_ (.Y(_0743_),
    .B(_0742_),
    .A_N(_0711_));
 sg13g2_xnor2_1 _1649_ (.Y(_0744_),
    .A(_0711_),
    .B(_0742_));
 sg13g2_nand2b_1 _1650_ (.Y(_0745_),
    .B(_0744_),
    .A_N(_0722_));
 sg13g2_xnor2_1 _1651_ (.Y(_0746_),
    .A(_0722_),
    .B(_0744_));
 sg13g2_nand2_1 _1652_ (.Y(_0747_),
    .A(_0718_),
    .B(_0720_));
 sg13g2_nand2_1 _1653_ (.Y(_0748_),
    .A(_0746_),
    .B(_0747_));
 sg13g2_xor2_1 _1654_ (.B(_0747_),
    .A(_0746_),
    .X(_0749_));
 sg13g2_nor2b_1 _1655_ (.A(_0737_),
    .B_N(_0749_),
    .Y(_0750_));
 sg13g2_xnor2_1 _1656_ (.Y(_0751_),
    .A(_0737_),
    .B(_0749_));
 sg13g2_nor3_1 _1657_ (.A(_0674_),
    .B(_0696_),
    .C(_0730_),
    .Y(_0752_));
 sg13g2_nor4_1 _1658_ (.A(_0669_),
    .B(_0702_),
    .C(_0731_),
    .D(_0752_),
    .Y(_0753_));
 sg13g2_o21ai_1 _1659_ (.B1(_0753_),
    .Y(_0754_),
    .A1(_0635_),
    .A2(_0700_));
 sg13g2_nor2_1 _1660_ (.A(_0697_),
    .B(_0731_),
    .Y(_0755_));
 sg13g2_nor2_1 _1661_ (.A(_0730_),
    .B(_0755_),
    .Y(_0756_));
 sg13g2_a21oi_1 _1662_ (.A1(_0754_),
    .A2(_0756_),
    .Y(_0757_),
    .B1(_0751_));
 sg13g2_and3_1 _1663_ (.X(_0758_),
    .A(_0751_),
    .B(_0754_),
    .C(_0756_));
 sg13g2_nor3_1 _1664_ (.A(net214),
    .B(_0757_),
    .C(_0758_),
    .Y(_0759_));
 sg13g2_a22oi_1 _1665_ (.Y(_0760_),
    .B1(net209),
    .B2(net222),
    .A2(net211),
    .A1(net137));
 sg13g2_nand2b_1 _1666_ (.Y(_0761_),
    .B(_0760_),
    .A_N(_0759_));
 sg13g2_and2_1 _1667_ (.A(net265),
    .B(_0761_),
    .X(_0051_));
 sg13g2_a21oi_1 _1668_ (.A1(net217),
    .A2(_0712_),
    .Y(_0762_),
    .B1(_0741_));
 sg13g2_a22oi_1 _1669_ (.Y(_0763_),
    .B1(net215),
    .B2(net242),
    .A2(net217),
    .A1(net237));
 sg13g2_nand4_1 _1670_ (.B(net238),
    .C(net217),
    .A(net241),
    .Y(_0764_),
    .D(net215));
 sg13g2_nor2b_1 _1671_ (.A(_0763_),
    .B_N(_0764_),
    .Y(_0765_));
 sg13g2_nand2b_1 _1672_ (.Y(_0766_),
    .B(_0765_),
    .A_N(_0743_));
 sg13g2_xor2_1 _1673_ (.B(_0765_),
    .A(_0743_),
    .X(_0767_));
 sg13g2_xnor2_1 _1674_ (.Y(_0768_),
    .A(_0762_),
    .B(_0767_));
 sg13g2_a21oi_1 _1675_ (.A1(_0745_),
    .A2(_0748_),
    .Y(_0769_),
    .B1(_0768_));
 sg13g2_nand3_1 _1676_ (.B(_0748_),
    .C(_0768_),
    .A(_0745_),
    .Y(_0770_));
 sg13g2_nor2b_1 _1677_ (.A(_0769_),
    .B_N(_0770_),
    .Y(_0771_));
 sg13g2_or3_1 _1678_ (.A(_0750_),
    .B(_0758_),
    .C(_0771_),
    .X(_0772_));
 sg13g2_o21ai_1 _1679_ (.B1(_0771_),
    .Y(_0773_),
    .A1(_0750_),
    .A2(_0758_));
 sg13g2_nand3_1 _1680_ (.B(_0772_),
    .C(_0773_),
    .A(net213),
    .Y(_0774_));
 sg13g2_a22oi_1 _1681_ (.Y(_0775_),
    .B1(net209),
    .B2(net219),
    .A2(net211),
    .A1(net105));
 sg13g2_a21oi_1 _1682_ (.A1(_0774_),
    .A2(_0775_),
    .Y(_0052_),
    .B1(net256));
 sg13g2_nand3_1 _1683_ (.B(net215),
    .C(_0738_),
    .A(net238),
    .Y(_0776_));
 sg13g2_o21ai_1 _1684_ (.B1(_0766_),
    .Y(_0777_),
    .A1(_0762_),
    .A2(_0767_));
 sg13g2_nand2b_1 _1685_ (.Y(_0778_),
    .B(_0777_),
    .A_N(_0776_));
 sg13g2_xor2_1 _1686_ (.B(_0777_),
    .A(_0776_),
    .X(_0779_));
 sg13g2_nand4_1 _1687_ (.B(_0754_),
    .C(_0756_),
    .A(_0751_),
    .Y(_0780_),
    .D(_0771_));
 sg13g2_a21oi_1 _1688_ (.A1(_0750_),
    .A2(_0770_),
    .Y(_0781_),
    .B1(_0769_));
 sg13g2_a21oi_1 _1689_ (.A1(_0780_),
    .A2(_0781_),
    .Y(_0782_),
    .B1(_0779_));
 sg13g2_and3_1 _1690_ (.X(_0783_),
    .A(_0779_),
    .B(_0780_),
    .C(_0781_));
 sg13g2_or3_1 _1691_ (.A(net214),
    .B(_0782_),
    .C(_0783_),
    .X(_0784_));
 sg13g2_a22oi_1 _1692_ (.Y(_0785_),
    .B1(net209),
    .B2(net218),
    .A2(net211),
    .A1(net104));
 sg13g2_a21oi_1 _1693_ (.A1(_0784_),
    .A2(_0785_),
    .Y(_0053_),
    .B1(net256));
 sg13g2_nand2_1 _1694_ (.Y(_0786_),
    .A(_0764_),
    .B(_0778_));
 sg13g2_o21ai_1 _1695_ (.B1(net213),
    .Y(_0787_),
    .A1(_0782_),
    .A2(_0786_));
 sg13g2_a22oi_1 _1696_ (.Y(_0788_),
    .B1(net209),
    .B2(net216),
    .A2(net211),
    .A1(net118));
 sg13g2_a21oi_1 _1697_ (.A1(_0787_),
    .A2(net119),
    .Y(_0054_),
    .B1(net256));
 sg13g2_nor4_1 _1698_ (.A(net260),
    .B(net73),
    .C(_0348_),
    .D(_0357_),
    .Y(_0055_));
 sg13g2_dfrbp_1 _1699_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net22),
    .D(_0012_),
    .Q_N(_0004_),
    .Q(\i_decoder_a.valid ));
 sg13g2_dfrbp_1 _1700_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net60),
    .D(_0013_),
    .Q_N(_0828_),
    .Q(\i_decoder_a.data_out[0] ));
 sg13g2_dfrbp_1 _1701_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net59),
    .D(_0014_),
    .Q_N(_0827_),
    .Q(\i_decoder_a.data_out[1] ));
 sg13g2_dfrbp_1 _1702_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net58),
    .D(_0015_),
    .Q_N(_0826_),
    .Q(\i_decoder_a.data_out[2] ));
 sg13g2_dfrbp_1 _1703_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net57),
    .D(_0016_),
    .Q_N(_0825_),
    .Q(\i_decoder_a.data_out[3] ));
 sg13g2_dfrbp_1 _1704_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net56),
    .D(_0017_),
    .Q_N(_0824_),
    .Q(\i_decoder_a.data_out[4] ));
 sg13g2_dfrbp_1 _1705_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net45),
    .D(net148),
    .Q_N(_0823_),
    .Q(\i_decoder_a.data_out[5] ));
 sg13g2_dfrbp_1 _1706_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net44),
    .D(net143),
    .Q_N(_0822_),
    .Q(\i_decoder_a.data_out[6] ));
 sg13g2_dfrbp_1 _1707_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net43),
    .D(net153),
    .Q_N(_0821_),
    .Q(\i_decoder_a.data_out[7] ));
 sg13g2_dfrbp_1 _1708_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net42),
    .D(_0021_),
    .Q_N(_0010_),
    .Q(\i_decoder_a.count[0] ));
 sg13g2_dfrbp_1 _1709_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net40),
    .D(net134),
    .Q_N(_0820_),
    .Q(\i_decoder_a.count[1] ));
 sg13g2_dfrbp_1 _1710_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net38),
    .D(net117),
    .Q_N(_0819_),
    .Q(\i_decoder_a.count[2] ));
 sg13g2_dfrbp_1 _1711_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net23),
    .D(net141),
    .Q_N(_0829_),
    .Q(\i_decoder_a.count[3] ));
 sg13g2_dfrbp_1 _1712_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net24),
    .D(net2),
    .Q_N(_0003_),
    .Q(\i_decoder_a.i_raw_data.data_out[0] ));
 sg13g2_dfrbp_1 _1713_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net25),
    .D(net80),
    .Q_N(_0002_),
    .Q(\i_decoder_a.i_raw_data.data_out[1] ));
 sg13g2_dfrbp_1 _1714_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net26),
    .D(net83),
    .Q_N(_0830_),
    .Q(\i_decoder_a.i_raw_data.data_out[2] ));
 sg13g2_dfrbp_1 _1715_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net27),
    .D(net92),
    .Q_N(_0831_),
    .Q(\i_decoder_a.i_raw_data.data_out[3] ));
 sg13g2_dfrbp_1 _1716_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net28),
    .D(net87),
    .Q_N(_0000_),
    .Q(\i_decoder_a.i_raw_data.data_out[4] ));
 sg13g2_dfrbp_1 _1717_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net29),
    .D(net85),
    .Q_N(_0832_),
    .Q(\i_decoder_a.i_raw_data.data_out[5] ));
 sg13g2_dfrbp_1 _1718_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net30),
    .D(net84),
    .Q_N(_0833_),
    .Q(\i_decoder_a.i_raw_data.data_out[6] ));
 sg13g2_dfrbp_1 _1719_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net31),
    .D(net236),
    .Q_N(_0001_),
    .Q(\i_decoder_a.i_raw_data.data_out[7] ));
 sg13g2_dfrbp_1 _1720_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net46),
    .D(net78),
    .Q_N(_0834_),
    .Q(\i_decoder_a.i_raw_data.data_out[8] ));
 sg13g2_dfrbp_1 _1721_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net36),
    .D(net86),
    .Q_N(_0818_),
    .Q(\i_decoder_a.i_raw_data.data_out[9] ));
 sg13g2_dfrbp_1 _1722_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net34),
    .D(net76),
    .Q_N(_0817_),
    .Q(\i_decoder_a.updated ));
 sg13g2_dfrbp_1 _1723_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net33),
    .D(_0026_),
    .Q_N(_0009_),
    .Q(\i_decoder_b.valid ));
 sg13g2_dfrbp_1 _1724_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net32),
    .D(_0027_),
    .Q_N(_0816_),
    .Q(\i_decoder_b.data_out[0] ));
 sg13g2_dfrbp_1 _1725_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net21),
    .D(_0028_),
    .Q_N(_0815_),
    .Q(\i_decoder_b.data_out[1] ));
 sg13g2_dfrbp_1 _1726_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net20),
    .D(_0029_),
    .Q_N(_0814_),
    .Q(\i_decoder_b.data_out[2] ));
 sg13g2_dfrbp_1 _1727_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net19),
    .D(_0030_),
    .Q_N(_0813_),
    .Q(\i_decoder_b.data_out[3] ));
 sg13g2_dfrbp_1 _1728_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net18),
    .D(_0031_),
    .Q_N(_0812_),
    .Q(\i_decoder_b.data_out[4] ));
 sg13g2_dfrbp_1 _1729_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net17),
    .D(_0032_),
    .Q_N(_0811_),
    .Q(\i_decoder_b.data_out[5] ));
 sg13g2_dfrbp_1 _1730_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net16),
    .D(net98),
    .Q_N(_0810_),
    .Q(\i_decoder_b.data_out[6] ));
 sg13g2_dfrbp_1 _1731_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net15),
    .D(_0034_),
    .Q_N(_0809_),
    .Q(\i_decoder_b.data_out[7] ));
 sg13g2_dfrbp_1 _1732_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net14),
    .D(net95),
    .Q_N(_0011_),
    .Q(\i_decoder_b.count[0] ));
 sg13g2_dfrbp_1 _1733_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net12),
    .D(_0036_),
    .Q_N(_0808_),
    .Q(\i_decoder_b.count[1] ));
 sg13g2_dfrbp_1 _1734_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net10),
    .D(net151),
    .Q_N(_0807_),
    .Q(\i_decoder_b.count[2] ));
 sg13g2_dfrbp_1 _1735_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net47),
    .D(_0038_),
    .Q_N(_0835_),
    .Q(\i_decoder_b.count[3] ));
 sg13g2_dfrbp_1 _1736_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net48),
    .D(net3),
    .Q_N(_0008_),
    .Q(\i_decoder_b.i_raw_data.data_out[0] ));
 sg13g2_dfrbp_1 _1737_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net49),
    .D(net81),
    .Q_N(_0007_),
    .Q(\i_decoder_b.i_raw_data.data_out[1] ));
 sg13g2_dfrbp_1 _1738_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net50),
    .D(net79),
    .Q_N(_0836_),
    .Q(\i_decoder_b.i_raw_data.data_out[2] ));
 sg13g2_dfrbp_1 _1739_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net51),
    .D(net91),
    .Q_N(_0837_),
    .Q(\i_decoder_b.i_raw_data.data_out[3] ));
 sg13g2_dfrbp_1 _1740_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net52),
    .D(net90),
    .Q_N(_0005_),
    .Q(\i_decoder_b.i_raw_data.data_out[4] ));
 sg13g2_dfrbp_1 _1741_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net53),
    .D(net89),
    .Q_N(_0838_),
    .Q(\i_decoder_b.i_raw_data.data_out[5] ));
 sg13g2_dfrbp_1 _1742_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net54),
    .D(net82),
    .Q_N(_0839_),
    .Q(\i_decoder_b.i_raw_data.data_out[6] ));
 sg13g2_dfrbp_1 _1743_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net55),
    .D(net96),
    .Q_N(_0006_),
    .Q(\i_decoder_b.i_raw_data.data_out[7] ));
 sg13g2_dfrbp_1 _1744_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net67),
    .D(net77),
    .Q_N(_0840_),
    .Q(\i_decoder_b.i_raw_data.data_out[8] ));
 sg13g2_dfrbp_1 _1745_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net72),
    .D(net88),
    .Q_N(_0806_),
    .Q(\i_decoder_b.i_raw_data.data_out[9] ));
 sg13g2_dfrbp_1 _1746_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net70),
    .D(_0039_),
    .Q_N(_0805_),
    .Q(\result[0] ));
 sg13g2_dfrbp_1 _1747_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net68),
    .D(_0040_),
    .Q_N(_0804_),
    .Q(\result[1] ));
 sg13g2_dfrbp_1 _1748_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net66),
    .D(_0041_),
    .Q_N(_0803_),
    .Q(\result[2] ));
 sg13g2_dfrbp_1 _1749_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net64),
    .D(_0042_),
    .Q_N(_0802_),
    .Q(\result[3] ));
 sg13g2_dfrbp_1 _1750_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net62),
    .D(_0043_),
    .Q_N(_0801_),
    .Q(\result[4] ));
 sg13g2_dfrbp_1 _1751_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net41),
    .D(_0044_),
    .Q_N(_0800_),
    .Q(\result[5] ));
 sg13g2_dfrbp_1 _1752_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net37),
    .D(_0045_),
    .Q_N(_0799_),
    .Q(\result[6] ));
 sg13g2_dfrbp_1 _1753_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net13),
    .D(_0046_),
    .Q_N(_0798_),
    .Q(\result[7] ));
 sg13g2_dfrbp_1 _1754_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net9),
    .D(_0047_),
    .Q_N(_0797_),
    .Q(\result[8] ));
 sg13g2_dfrbp_1 _1755_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net69),
    .D(_0048_),
    .Q_N(_0796_),
    .Q(\result[9] ));
 sg13g2_dfrbp_1 _1756_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net65),
    .D(_0049_),
    .Q_N(_0795_),
    .Q(\result[10] ));
 sg13g2_dfrbp_1 _1757_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net61),
    .D(_0050_),
    .Q_N(_0794_),
    .Q(\result[11] ));
 sg13g2_dfrbp_1 _1758_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net35),
    .D(_0051_),
    .Q_N(_0793_),
    .Q(\result[12] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net71),
    .D(_0052_),
    .Q_N(_0792_),
    .Q(\result[13] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net63),
    .D(_0053_),
    .Q_N(_0791_),
    .Q(\result[14] ));
 sg13g2_dfrbp_1 _1761_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net11),
    .D(_0054_),
    .Q_N(_0790_),
    .Q(\result[15] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net39),
    .D(net74),
    .Q_N(_0789_),
    .Q(\i_decoder_b.updated ));
 sg13g2_tiehi _1734__10 (.L_HI(net10));
 sg13g2_tiehi _1761__11 (.L_HI(net11));
 sg13g2_tiehi _1733__12 (.L_HI(net12));
 sg13g2_tiehi _1753__13 (.L_HI(net13));
 sg13g2_tiehi _1732__14 (.L_HI(net14));
 sg13g2_tiehi _1731__15 (.L_HI(net15));
 sg13g2_tiehi _1730__16 (.L_HI(net16));
 sg13g2_tiehi _1729__17 (.L_HI(net17));
 sg13g2_tiehi _1728__18 (.L_HI(net18));
 sg13g2_tiehi _1727__19 (.L_HI(net19));
 sg13g2_tiehi _1726__20 (.L_HI(net20));
 sg13g2_tiehi _1725__21 (.L_HI(net21));
 sg13g2_tiehi _1699__22 (.L_HI(net22));
 sg13g2_tiehi _1711__23 (.L_HI(net23));
 sg13g2_tiehi _1712__24 (.L_HI(net24));
 sg13g2_tiehi _1713__25 (.L_HI(net25));
 sg13g2_tiehi _1714__26 (.L_HI(net26));
 sg13g2_tiehi _1715__27 (.L_HI(net27));
 sg13g2_tiehi _1716__28 (.L_HI(net28));
 sg13g2_tiehi _1717__29 (.L_HI(net29));
 sg13g2_tiehi _1718__30 (.L_HI(net30));
 sg13g2_tiehi _1719__31 (.L_HI(net31));
 sg13g2_tiehi _1724__32 (.L_HI(net32));
 sg13g2_tiehi _1723__33 (.L_HI(net33));
 sg13g2_tiehi _1722__34 (.L_HI(net34));
 sg13g2_tiehi _1758__35 (.L_HI(net35));
 sg13g2_tiehi _1721__36 (.L_HI(net36));
 sg13g2_tiehi _1752__37 (.L_HI(net37));
 sg13g2_tiehi _1710__38 (.L_HI(net38));
 sg13g2_tiehi _1762__39 (.L_HI(net39));
 sg13g2_tiehi _1709__40 (.L_HI(net40));
 sg13g2_tiehi _1751__41 (.L_HI(net41));
 sg13g2_tiehi _1708__42 (.L_HI(net42));
 sg13g2_tiehi _1707__43 (.L_HI(net43));
 sg13g2_tiehi _1706__44 (.L_HI(net44));
 sg13g2_tiehi _1705__45 (.L_HI(net45));
 sg13g2_tiehi _1720__46 (.L_HI(net46));
 sg13g2_tiehi _1735__47 (.L_HI(net47));
 sg13g2_tiehi _1736__48 (.L_HI(net48));
 sg13g2_tiehi _1737__49 (.L_HI(net49));
 sg13g2_tiehi _1738__50 (.L_HI(net50));
 sg13g2_tiehi _1739__51 (.L_HI(net51));
 sg13g2_tiehi _1740__52 (.L_HI(net52));
 sg13g2_tiehi _1741__53 (.L_HI(net53));
 sg13g2_tiehi _1742__54 (.L_HI(net54));
 sg13g2_tiehi _1743__55 (.L_HI(net55));
 sg13g2_tiehi _1704__56 (.L_HI(net56));
 sg13g2_tiehi _1703__57 (.L_HI(net57));
 sg13g2_tiehi _1702__58 (.L_HI(net58));
 sg13g2_tiehi _1701__59 (.L_HI(net59));
 sg13g2_tiehi _1700__60 (.L_HI(net60));
 sg13g2_tiehi _1757__61 (.L_HI(net61));
 sg13g2_tiehi _1750__62 (.L_HI(net62));
 sg13g2_tiehi _1760__63 (.L_HI(net63));
 sg13g2_tiehi _1749__64 (.L_HI(net64));
 sg13g2_tiehi _1756__65 (.L_HI(net65));
 sg13g2_tiehi _1748__66 (.L_HI(net66));
 sg13g2_tiehi _1744__67 (.L_HI(net67));
 sg13g2_tiehi _1747__68 (.L_HI(net68));
 sg13g2_tiehi _1755__69 (.L_HI(net69));
 sg13g2_tiehi _1746__70 (.L_HI(net70));
 sg13g2_tiehi _1759__71 (.L_HI(net71));
 sg13g2_tiehi _1745__72 (.L_HI(net72));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _1827_ (.A(uio_oe[7]),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1828_ (.A(uio_oe[7]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1829_ (.A(uio_oe[7]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1830_ (.A(uio_oe[7]),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1831_ (.A(uio_oe[7]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1832_ (.A(uio_oe[7]),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1833_ (.A(uio_oe[7]),
    .X(uio_oe[6]));
 sg13g2_buf_2 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_0211_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_0297_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_0146_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_0139_),
    .X(net207));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(_0292_));
 sg13g2_buf_2 fanout209 (.A(_0430_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_0430_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_0426_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_0426_),
    .X(net212));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(_0425_));
 sg13g2_buf_2 fanout214 (.A(_0424_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(net216),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(net146),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(net218),
    .X(net217));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(net97));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(net220));
 sg13g2_buf_2 fanout220 (.A(net135),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(net222),
    .X(net221));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(net136));
 sg13g2_buf_2 fanout223 (.A(net225),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(net225),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(net130),
    .X(net225));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(net156));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(net231));
 sg13g2_buf_1 fanout228 (.A(net231),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(net231),
    .X(net229));
 sg13g2_buf_1 fanout230 (.A(net231),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(\i_decoder_b.data_out[1] ),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(net235),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(net234),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(net235),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(\i_decoder_b.data_out[0] ),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net112),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(net239),
    .X(net237));
 sg13g2_buf_1 fanout238 (.A(net239),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(\i_decoder_a.data_out[7] ),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(net242));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(net142));
 sg13g2_buf_2 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(net245),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(net147),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(net247),
    .X(net246));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(\i_decoder_a.data_out[4] ));
 sg13g2_buf_2 fanout248 (.A(net249),
    .X(net248));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(\i_decoder_a.data_out[3] ));
 sg13g2_buf_2 fanout250 (.A(net251),
    .X(net250));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(\i_decoder_a.data_out[2] ));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(\i_decoder_a.data_out[1] ),
    .X(net253));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(net101));
 sg13g2_buf_2 fanout255 (.A(_0069_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(net258),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(net258),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net260),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(net260),
    .X(net259));
 sg13g2_buf_1 fanout260 (.A(_0063_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(net264),
    .X(net261));
 sg13g2_buf_1 fanout262 (.A(net264),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(net264),
    .X(net263));
 sg13g2_buf_1 fanout264 (.A(ui_in[6]),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(net267),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(net267),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(net1),
    .X(net267));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tiehi _1754__9 (.L_HI(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0009_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0055_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0004_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0025_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i_decoder_b.i_raw_data.data_out[7] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_decoder_a.i_raw_data.data_out[7] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_decoder_b.i_raw_data.data_out[1] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_decoder_a.i_raw_data.data_out[0] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_decoder_b.i_raw_data.data_out[0] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_decoder_b.i_raw_data.data_out[5] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_decoder_a.i_raw_data.data_out[1] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_decoder_a.i_raw_data.data_out[5] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_decoder_a.i_raw_data.data_out[4] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_decoder_a.i_raw_data.data_out[8] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_decoder_a.i_raw_data.data_out[3] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_decoder_b.i_raw_data.data_out[8] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_decoder_b.i_raw_data.data_out[4] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_decoder_b.i_raw_data.data_out[3] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_decoder_b.i_raw_data.data_out[2] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_decoder_a.i_raw_data.data_out[2] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0011_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0411_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0035_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_decoder_b.i_raw_data.data_out[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_decoder_b.data_out[6] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0033_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0010_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0265_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i_decoder_a.data_out[0] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold30 (.A(\result[5] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0516_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold32 (.A(\result[14] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold33 (.A(\result[13] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold34 (.A(\result[8] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0639_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold36 (.A(\result[3] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0461_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold38 (.A(\result[9] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold39 (.A(\result[11] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_decoder_a.i_raw_data.data_out[6] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold41 (.A(\result[10] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold42 (.A(\result[4] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold43 (.A(\result[2] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_decoder_a.valid ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0023_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold46 (.A(\result[15] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0788_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold48 (.A(\result[6] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0555_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold50 (.A(\result[1] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold51 (.A(\result[0] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_decoder_b.valid ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_decoder_b.count[0] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0415_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0417_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold56 (.A(\result[7] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0601_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_decoder_b.data_out[3] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_decoder_a.count[0] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0268_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0270_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0022_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_decoder_b.data_out[5] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold64 (.A(\i_decoder_b.data_out[4] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold65 (.A(\result[12] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_decoder_a.count[3] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0274_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0275_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0024_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_decoder_a.data_out[6] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0019_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_decoder_a.count[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0208_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_decoder_b.data_out[7] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_decoder_a.data_out[5] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0018_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold77 (.A(\i_decoder_b.count[2] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0419_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0037_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0002_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0020_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_decoder_b.count[3] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0421_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_decoder_b.data_out[2] ),
    .X(net156));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_174 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_196 ();
 sg13g2_fill_1 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_215 ();
 sg13g2_decap_8 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_233 ();
 sg13g2_decap_8 FILLER_9_240 ();
 sg13g2_decap_8 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_decap_8 FILLER_9_268 ();
 sg13g2_decap_8 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_310 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_fill_1 FILLER_10_147 ();
 sg13g2_fill_1 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_decap_8 FILLER_10_253 ();
 sg13g2_decap_8 FILLER_10_260 ();
 sg13g2_decap_8 FILLER_10_267 ();
 sg13g2_decap_8 FILLER_10_274 ();
 sg13g2_decap_8 FILLER_10_281 ();
 sg13g2_decap_8 FILLER_10_288 ();
 sg13g2_decap_8 FILLER_10_295 ();
 sg13g2_decap_8 FILLER_10_302 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_10_337 ();
 sg13g2_decap_8 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_4 FILLER_11_133 ();
 sg13g2_decap_4 FILLER_11_163 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_fill_1 FILLER_11_194 ();
 sg13g2_fill_2 FILLER_11_203 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_4 FILLER_11_266 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_283 ();
 sg13g2_decap_8 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_fill_2 FILLER_12_140 ();
 sg13g2_fill_2 FILLER_12_161 ();
 sg13g2_fill_1 FILLER_12_163 ();
 sg13g2_fill_2 FILLER_12_172 ();
 sg13g2_fill_1 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_201 ();
 sg13g2_fill_1 FILLER_12_229 ();
 sg13g2_fill_1 FILLER_12_236 ();
 sg13g2_fill_2 FILLER_12_243 ();
 sg13g2_fill_2 FILLER_12_258 ();
 sg13g2_fill_1 FILLER_12_260 ();
 sg13g2_decap_4 FILLER_12_287 ();
 sg13g2_fill_2 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_157 ();
 sg13g2_fill_2 FILLER_13_164 ();
 sg13g2_fill_1 FILLER_13_166 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_fill_1 FILLER_13_186 ();
 sg13g2_fill_1 FILLER_13_210 ();
 sg13g2_decap_4 FILLER_13_223 ();
 sg13g2_fill_2 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_4 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_137 ();
 sg13g2_decap_4 FILLER_14_151 ();
 sg13g2_fill_1 FILLER_14_155 ();
 sg13g2_fill_2 FILLER_14_164 ();
 sg13g2_decap_4 FILLER_14_174 ();
 sg13g2_fill_2 FILLER_14_178 ();
 sg13g2_decap_4 FILLER_14_204 ();
 sg13g2_fill_2 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_fill_2 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_253 ();
 sg13g2_fill_2 FILLER_14_267 ();
 sg13g2_fill_1 FILLER_14_269 ();
 sg13g2_fill_2 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_4 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_2 FILLER_15_167 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_187 ();
 sg13g2_fill_2 FILLER_15_199 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_234 ();
 sg13g2_fill_1 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_4 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_150 ();
 sg13g2_fill_1 FILLER_16_152 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_172 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_178 ();
 sg13g2_decap_4 FILLER_16_185 ();
 sg13g2_fill_2 FILLER_16_189 ();
 sg13g2_decap_4 FILLER_16_201 ();
 sg13g2_fill_1 FILLER_16_205 ();
 sg13g2_decap_4 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_fill_2 FILLER_16_273 ();
 sg13g2_fill_1 FILLER_16_275 ();
 sg13g2_decap_4 FILLER_16_289 ();
 sg13g2_fill_2 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_4 FILLER_16_374 ();
 sg13g2_fill_1 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_2 FILLER_17_150 ();
 sg13g2_fill_1 FILLER_17_152 ();
 sg13g2_fill_2 FILLER_17_183 ();
 sg13g2_fill_1 FILLER_17_185 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_decap_4 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_201 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_decap_4 FILLER_17_219 ();
 sg13g2_fill_2 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_fill_1 FILLER_17_235 ();
 sg13g2_fill_1 FILLER_17_241 ();
 sg13g2_decap_4 FILLER_17_246 ();
 sg13g2_fill_1 FILLER_17_256 ();
 sg13g2_fill_2 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_fill_2 FILLER_17_335 ();
 sg13g2_decap_4 FILLER_17_341 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_4 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_170 ();
 sg13g2_decap_8 FILLER_18_229 ();
 sg13g2_fill_2 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_4 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_274 ();
 sg13g2_fill_2 FILLER_18_285 ();
 sg13g2_decap_4 FILLER_18_322 ();
 sg13g2_decap_4 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_fill_1 FILLER_18_361 ();
 sg13g2_fill_2 FILLER_18_380 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_127 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_fill_2 FILLER_19_141 ();
 sg13g2_decap_4 FILLER_19_148 ();
 sg13g2_decap_4 FILLER_19_170 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_4 FILLER_19_196 ();
 sg13g2_fill_2 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_215 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_fill_1 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_decap_4 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_320 ();
 sg13g2_fill_2 FILLER_19_338 ();
 sg13g2_decap_4 FILLER_19_359 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_4 FILLER_20_146 ();
 sg13g2_decap_4 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_206 ();
 sg13g2_fill_1 FILLER_20_261 ();
 sg13g2_fill_2 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_fill_1 FILLER_20_287 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_330 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_360 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_78 ();
 sg13g2_fill_1 FILLER_21_83 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_decap_8 FILLER_21_96 ();
 sg13g2_decap_8 FILLER_21_103 ();
 sg13g2_decap_8 FILLER_21_110 ();
 sg13g2_decap_4 FILLER_21_117 ();
 sg13g2_fill_2 FILLER_21_121 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_decap_8 FILLER_21_141 ();
 sg13g2_fill_2 FILLER_21_148 ();
 sg13g2_decap_4 FILLER_21_155 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_fill_2 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_207 ();
 sg13g2_fill_2 FILLER_21_214 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_4 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_297 ();
 sg13g2_decap_8 FILLER_21_303 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_349 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_375 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_50 ();
 sg13g2_decap_4 FILLER_22_57 ();
 sg13g2_fill_1 FILLER_22_61 ();
 sg13g2_fill_2 FILLER_22_90 ();
 sg13g2_fill_1 FILLER_22_92 ();
 sg13g2_decap_8 FILLER_22_110 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_2 FILLER_22_146 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_4 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_4 FILLER_22_236 ();
 sg13g2_decap_8 FILLER_22_250 ();
 sg13g2_decap_8 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_269 ();
 sg13g2_decap_4 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_287 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_fill_2 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_24 ();
 sg13g2_fill_2 FILLER_23_31 ();
 sg13g2_fill_1 FILLER_23_33 ();
 sg13g2_fill_2 FILLER_23_60 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_8 FILLER_23_81 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_decap_4 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_4 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_132 ();
 sg13g2_decap_8 FILLER_23_138 ();
 sg13g2_decap_8 FILLER_23_145 ();
 sg13g2_fill_1 FILLER_23_152 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_fill_2 FILLER_23_164 ();
 sg13g2_fill_1 FILLER_23_166 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_decap_8 FILLER_23_186 ();
 sg13g2_fill_2 FILLER_23_193 ();
 sg13g2_fill_1 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_306 ();
 sg13g2_decap_4 FILLER_23_338 ();
 sg13g2_fill_1 FILLER_23_342 ();
 sg13g2_fill_2 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_fill_2 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_decap_4 FILLER_24_22 ();
 sg13g2_fill_1 FILLER_24_26 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_47 ();
 sg13g2_fill_2 FILLER_24_54 ();
 sg13g2_fill_2 FILLER_24_85 ();
 sg13g2_fill_2 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_136 ();
 sg13g2_decap_4 FILLER_24_164 ();
 sg13g2_fill_1 FILLER_24_168 ();
 sg13g2_decap_4 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_222 ();
 sg13g2_decap_4 FILLER_24_227 ();
 sg13g2_fill_2 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_316 ();
 sg13g2_fill_2 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_2 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_17 ();
 sg13g2_fill_1 FILLER_25_19 ();
 sg13g2_fill_2 FILLER_25_45 ();
 sg13g2_fill_1 FILLER_25_47 ();
 sg13g2_decap_4 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_64 ();
 sg13g2_fill_2 FILLER_25_71 ();
 sg13g2_fill_2 FILLER_25_116 ();
 sg13g2_fill_1 FILLER_25_118 ();
 sg13g2_fill_2 FILLER_25_127 ();
 sg13g2_decap_8 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_decap_8 FILLER_25_156 ();
 sg13g2_decap_4 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_193 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_fill_2 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_236 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_fill_1 FILLER_25_324 ();
 sg13g2_decap_4 FILLER_25_330 ();
 sg13g2_fill_1 FILLER_25_334 ();
 sg13g2_fill_1 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_23 ();
 sg13g2_fill_2 FILLER_26_30 ();
 sg13g2_fill_1 FILLER_26_66 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_102 ();
 sg13g2_decap_4 FILLER_26_120 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_fill_2 FILLER_26_158 ();
 sg13g2_decap_4 FILLER_26_173 ();
 sg13g2_fill_2 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_192 ();
 sg13g2_decap_4 FILLER_26_199 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_decap_4 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_fill_2 FILLER_26_334 ();
 sg13g2_fill_1 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_369 ();
 sg13g2_fill_1 FILLER_26_378 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_26 ();
 sg13g2_decap_8 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_46 ();
 sg13g2_fill_1 FILLER_27_53 ();
 sg13g2_decap_8 FILLER_27_59 ();
 sg13g2_decap_8 FILLER_27_66 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_decap_8 FILLER_27_88 ();
 sg13g2_fill_2 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_118 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_decap_4 FILLER_27_169 ();
 sg13g2_decap_8 FILLER_27_197 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_decap_4 FILLER_27_256 ();
 sg13g2_decap_4 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_272 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_25 ();
 sg13g2_fill_2 FILLER_28_32 ();
 sg13g2_fill_1 FILLER_28_34 ();
 sg13g2_decap_8 FILLER_28_48 ();
 sg13g2_fill_2 FILLER_28_55 ();
 sg13g2_fill_1 FILLER_28_57 ();
 sg13g2_decap_4 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_71 ();
 sg13g2_decap_4 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_fill_2 FILLER_28_130 ();
 sg13g2_fill_2 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_4 FILLER_28_154 ();
 sg13g2_fill_2 FILLER_28_183 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_decap_8 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_198 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_decap_4 FILLER_28_240 ();
 sg13g2_fill_2 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_301 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_fill_2 FILLER_28_348 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_395 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_18 ();
 sg13g2_decap_8 FILLER_29_30 ();
 sg13g2_decap_4 FILLER_29_37 ();
 sg13g2_fill_1 FILLER_29_54 ();
 sg13g2_fill_2 FILLER_29_79 ();
 sg13g2_decap_8 FILLER_29_90 ();
 sg13g2_decap_4 FILLER_29_97 ();
 sg13g2_decap_4 FILLER_29_125 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_2 FILLER_29_386 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_48 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_2 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_decap_8 FILLER_30_67 ();
 sg13g2_decap_4 FILLER_30_95 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_decap_4 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_153 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_decap_4 FILLER_30_239 ();
 sg13g2_fill_1 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_1 FILLER_30_309 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_23 ();
 sg13g2_fill_1 FILLER_31_30 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_fill_2 FILLER_31_79 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_151 ();
 sg13g2_fill_2 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_247 ();
 sg13g2_decap_4 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_2 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_389 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_32 ();
 sg13g2_fill_2 FILLER_32_38 ();
 sg13g2_fill_1 FILLER_32_40 ();
 sg13g2_decap_8 FILLER_32_46 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_fill_1 FILLER_32_70 ();
 sg13g2_decap_4 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_decap_8 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_127 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_135 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_209 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_decap_8 FILLER_32_241 ();
 sg13g2_decap_4 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_fill_1 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_317 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_11 ();
 sg13g2_fill_2 FILLER_33_26 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_41 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_decap_4 FILLER_33_64 ();
 sg13g2_decap_4 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_fill_2 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_decap_4 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_279 ();
 sg13g2_fill_2 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_388 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_decap_8 FILLER_34_57 ();
 sg13g2_fill_2 FILLER_34_64 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_decap_8 FILLER_34_72 ();
 sg13g2_fill_2 FILLER_34_79 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_fill_2 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_139 ();
 sg13g2_fill_2 FILLER_34_152 ();
 sg13g2_fill_1 FILLER_34_168 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_decap_4 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_11 ();
 sg13g2_decap_8 FILLER_35_26 ();
 sg13g2_fill_2 FILLER_35_33 ();
 sg13g2_fill_1 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_44 ();
 sg13g2_decap_8 FILLER_35_51 ();
 sg13g2_decap_4 FILLER_35_79 ();
 sg13g2_fill_1 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_110 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_fill_1 FILLER_35_158 ();
 sg13g2_fill_2 FILLER_35_189 ();
 sg13g2_fill_1 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_219 ();
 sg13g2_decap_8 FILLER_35_229 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_290 ();
 sg13g2_fill_1 FILLER_35_308 ();
 sg13g2_fill_2 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_fill_1 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_4 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_25 ();
 sg13g2_fill_2 FILLER_36_43 ();
 sg13g2_fill_1 FILLER_36_45 ();
 sg13g2_decap_4 FILLER_36_59 ();
 sg13g2_decap_4 FILLER_36_83 ();
 sg13g2_fill_2 FILLER_36_87 ();
 sg13g2_fill_1 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_fill_2 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_decap_4 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_45 ();
 sg13g2_decap_8 FILLER_37_52 ();
 sg13g2_decap_8 FILLER_37_59 ();
 sg13g2_decap_8 FILLER_37_71 ();
 sg13g2_decap_8 FILLER_37_78 ();
 sg13g2_fill_1 FILLER_37_85 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_4 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_197 ();
 sg13g2_fill_2 FILLER_37_204 ();
 sg13g2_fill_1 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_fill_2 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_4 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_fill_2 FILLER_38_134 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_1 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_329 ();
 sg13g2_fill_1 FILLER_38_393 ();
 sg13g2_fill_1 FILLER_38_408 ();
endmodule

module tt_um_schoeberl_wildcat (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \ChiselTop._cntReg_T_1[0] ;
 wire \ChiselTop.cntReg[0] ;
 wire \ChiselTop.cntReg[10] ;
 wire \ChiselTop.cntReg[11] ;
 wire \ChiselTop.cntReg[12] ;
 wire \ChiselTop.cntReg[13] ;
 wire \ChiselTop.cntReg[14] ;
 wire \ChiselTop.cntReg[15] ;
 wire \ChiselTop.cntReg[16] ;
 wire \ChiselTop.cntReg[17] ;
 wire \ChiselTop.cntReg[18] ;
 wire \ChiselTop.cntReg[19] ;
 wire \ChiselTop.cntReg[1] ;
 wire \ChiselTop.cntReg[20] ;
 wire \ChiselTop.cntReg[21] ;
 wire \ChiselTop.cntReg[22] ;
 wire \ChiselTop.cntReg[23] ;
 wire \ChiselTop.cntReg[24] ;
 wire \ChiselTop.cntReg[25] ;
 wire \ChiselTop.cntReg[26] ;
 wire \ChiselTop.cntReg[27] ;
 wire \ChiselTop.cntReg[28] ;
 wire \ChiselTop.cntReg[29] ;
 wire \ChiselTop.cntReg[2] ;
 wire \ChiselTop.cntReg[30] ;
 wire \ChiselTop.cntReg[31] ;
 wire \ChiselTop.cntReg[3] ;
 wire \ChiselTop.cntReg[4] ;
 wire \ChiselTop.cntReg[5] ;
 wire \ChiselTop.cntReg[6] ;
 wire \ChiselTop.cntReg[7] ;
 wire \ChiselTop.cntReg[8] ;
 wire \ChiselTop.cntReg[9] ;
 wire \ChiselTop.dec.counter[0] ;
 wire \ChiselTop.dec.counter[1] ;
 wire \ChiselTop.dec.counter[2] ;
 wire \ChiselTop.dec.counter[3] ;
 wire \ChiselTop.led ;
 wire \ChiselTop.ledReg ;
 wire \ChiselTop.wild.cpu._GEN_176[10] ;
 wire \ChiselTop.wild.cpu._GEN_176[1] ;
 wire \ChiselTop.wild.cpu._GEN_176[20] ;
 wire \ChiselTop.wild.cpu._GEN_176[2] ;
 wire \ChiselTop.wild.cpu._GEN_176[5] ;
 wire \ChiselTop.wild.cpu._GEN_176[6] ;
 wire \ChiselTop.wild.cpu._T_12 ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[0] ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[1] ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[2] ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[3] ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[4] ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_1[0] ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[13] ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[15] ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[16] ;
 wire \ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[17] ;
 wire \ChiselTop.wild.cpu._pcNext_T_1[0] ;
 wire \ChiselTop.wild.cpu._pcNext_T_1[1] ;
 wire \ChiselTop.wild.cpu._wbData_T_1[0] ;
 wire \ChiselTop.wild.cpu._wbData_T_1[1] ;
 wire \ChiselTop.wild.cpu.decExReg_csrVal[0] ;
 wire \ChiselTop.wild.cpu.decExReg_csrVal[1] ;
 wire \ChiselTop.wild.cpu.decExReg_csrVal[2] ;
 wire \ChiselTop.wild.cpu.decExReg_csrVal[3] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_aluOp[0] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_aluOp[1] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_aluOp[2] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[0] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[10] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[11] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[12] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[13] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[14] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[15] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[16] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[17] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[1] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[20] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[21] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[22] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[25] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[26] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[28] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[2] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[31] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[3] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[4] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[5] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_imm[6] ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_isAuiPc ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_isBranch ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_isCssrw ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_isImm ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_isLoad ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_isLui ;
 wire \ChiselTop.wild.cpu.decExReg_decOut_rfWrite ;
 wire \ChiselTop.wild.cpu.decExReg_func3[0] ;
 wire \ChiselTop.wild.cpu.decExReg_func3[1] ;
 wire \ChiselTop.wild.cpu.decExReg_memLow[0] ;
 wire \ChiselTop.wild.cpu.decExReg_memLow[1] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[10] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[11] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[12] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[13] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[14] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[15] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[16] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[17] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[18] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[19] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[20] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[21] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[22] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[23] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[24] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[25] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[26] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[27] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[28] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[29] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[2] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[30] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[31] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[3] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[4] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[5] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[6] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[7] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[8] ;
 wire \ChiselTop.wild.cpu.decExReg_pc[9] ;
 wire \ChiselTop.wild.cpu.decExReg_rd[0] ;
 wire \ChiselTop.wild.cpu.decExReg_rd[1] ;
 wire \ChiselTop.wild.cpu.decExReg_rd[2] ;
 wire \ChiselTop.wild.cpu.decExReg_rd[3] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[0] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[10] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[11] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[12] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[13] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[14] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[15] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[16] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[17] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[18] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[19] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[1] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[20] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[21] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[22] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[23] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[24] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[25] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[26] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[27] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[28] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[29] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[2] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[30] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[31] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[3] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[4] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[5] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[6] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[7] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[8] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1Val[9] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1[0] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1[1] ;
 wire \ChiselTop.wild.cpu.decExReg_rs1[2] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[0] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[10] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[11] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[12] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[13] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[14] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[15] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[16] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[17] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[18] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[19] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[1] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[20] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[21] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[22] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[23] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[24] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[25] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[26] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[27] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[28] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[29] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[2] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[30] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[31] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[3] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[4] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[5] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[6] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[7] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[8] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2Val[9] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2[0] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2[1] ;
 wire \ChiselTop.wild.cpu.decExReg_rs2[2] ;
 wire \ChiselTop.wild.cpu.decExReg_valid ;
 wire \ChiselTop.wild.cpu.decEx_memLow[0] ;
 wire \ChiselTop.wild.cpu.decEx_memLow[1] ;
 wire \ChiselTop.wild.cpu.decOut_opcode[2] ;
 wire \ChiselTop.wild.cpu.decOut_opcode[4] ;
 wire \ChiselTop.wild.cpu.decOut_opcode[5] ;
 wire \ChiselTop.wild.cpu.exFwdReg_valid ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[0] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[10] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[11] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[12] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[13] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[14] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[15] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[16] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[17] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[18] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[19] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[1] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[20] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[21] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[22] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[23] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[24] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[25] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[26] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[27] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[28] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[29] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[2] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[30] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[31] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[3] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[4] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[5] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[6] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[7] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[8] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbData[9] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbDest[0] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbDest[1] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbDest[2] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbDest[3] ;
 wire \ChiselTop.wild.cpu.exFwdReg_wbDest[4] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[16] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[17] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[18] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[19] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[28] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[29] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[2] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[30] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[31] ;
 wire \ChiselTop.wild.cpu.io_dmem_rdAddress[3] ;
 wire \ChiselTop.wild.cpu.io_imem_data[13] ;
 wire \ChiselTop.wild.cpu.io_imem_data[15] ;
 wire \ChiselTop.wild.cpu.io_imem_data[16] ;
 wire \ChiselTop.wild.cpu.io_imem_data[20] ;
 wire \ChiselTop.wild.cpu.io_imem_data[21] ;
 wire \ChiselTop.wild.cpu.io_imem_data[22] ;
 wire \ChiselTop.wild.cpu.pcRegReg[0] ;
 wire \ChiselTop.wild.cpu.pcRegReg[10] ;
 wire \ChiselTop.wild.cpu.pcRegReg[11] ;
 wire \ChiselTop.wild.cpu.pcRegReg[12] ;
 wire \ChiselTop.wild.cpu.pcRegReg[13] ;
 wire \ChiselTop.wild.cpu.pcRegReg[14] ;
 wire \ChiselTop.wild.cpu.pcRegReg[15] ;
 wire \ChiselTop.wild.cpu.pcRegReg[16] ;
 wire \ChiselTop.wild.cpu.pcRegReg[17] ;
 wire \ChiselTop.wild.cpu.pcRegReg[18] ;
 wire \ChiselTop.wild.cpu.pcRegReg[19] ;
 wire \ChiselTop.wild.cpu.pcRegReg[1] ;
 wire \ChiselTop.wild.cpu.pcRegReg[20] ;
 wire \ChiselTop.wild.cpu.pcRegReg[21] ;
 wire \ChiselTop.wild.cpu.pcRegReg[22] ;
 wire \ChiselTop.wild.cpu.pcRegReg[23] ;
 wire \ChiselTop.wild.cpu.pcRegReg[24] ;
 wire \ChiselTop.wild.cpu.pcRegReg[25] ;
 wire \ChiselTop.wild.cpu.pcRegReg[26] ;
 wire \ChiselTop.wild.cpu.pcRegReg[27] ;
 wire \ChiselTop.wild.cpu.pcRegReg[28] ;
 wire \ChiselTop.wild.cpu.pcRegReg[29] ;
 wire \ChiselTop.wild.cpu.pcRegReg[2] ;
 wire \ChiselTop.wild.cpu.pcRegReg[30] ;
 wire \ChiselTop.wild.cpu.pcRegReg[31] ;
 wire \ChiselTop.wild.cpu.pcRegReg[3] ;
 wire \ChiselTop.wild.cpu.pcRegReg[4] ;
 wire \ChiselTop.wild.cpu.pcRegReg[5] ;
 wire \ChiselTop.wild.cpu.pcRegReg[6] ;
 wire \ChiselTop.wild.cpu.pcRegReg[7] ;
 wire \ChiselTop.wild.cpu.pcRegReg[8] ;
 wire \ChiselTop.wild.cpu.pcRegReg[9] ;
 wire \ChiselTop.wild.cpu.pcReg[10] ;
 wire \ChiselTop.wild.cpu.pcReg[11] ;
 wire \ChiselTop.wild.cpu.pcReg[12] ;
 wire \ChiselTop.wild.cpu.pcReg[13] ;
 wire \ChiselTop.wild.cpu.pcReg[14] ;
 wire \ChiselTop.wild.cpu.pcReg[15] ;
 wire \ChiselTop.wild.cpu.pcReg[16] ;
 wire \ChiselTop.wild.cpu.pcReg[17] ;
 wire \ChiselTop.wild.cpu.pcReg[18] ;
 wire \ChiselTop.wild.cpu.pcReg[19] ;
 wire \ChiselTop.wild.cpu.pcReg[20] ;
 wire \ChiselTop.wild.cpu.pcReg[21] ;
 wire \ChiselTop.wild.cpu.pcReg[22] ;
 wire \ChiselTop.wild.cpu.pcReg[23] ;
 wire \ChiselTop.wild.cpu.pcReg[24] ;
 wire \ChiselTop.wild.cpu.pcReg[25] ;
 wire \ChiselTop.wild.cpu.pcReg[26] ;
 wire \ChiselTop.wild.cpu.pcReg[27] ;
 wire \ChiselTop.wild.cpu.pcReg[28] ;
 wire \ChiselTop.wild.cpu.pcReg[29] ;
 wire \ChiselTop.wild.cpu.pcReg[2] ;
 wire \ChiselTop.wild.cpu.pcReg[30] ;
 wire \ChiselTop.wild.cpu.pcReg[31] ;
 wire \ChiselTop.wild.cpu.pcReg[3] ;
 wire \ChiselTop.wild.cpu.pcReg[4] ;
 wire \ChiselTop.wild.cpu.pcReg[5] ;
 wire \ChiselTop.wild.cpu.pcReg[6] ;
 wire \ChiselTop.wild.cpu.pcReg[7] ;
 wire \ChiselTop.wild.cpu.pcReg[8] ;
 wire \ChiselTop.wild.cpu.pcReg[9] ;
 wire \ChiselTop.wild.cpu.regs[0][0] ;
 wire \ChiselTop.wild.cpu.regs[0][10] ;
 wire \ChiselTop.wild.cpu.regs[0][11] ;
 wire \ChiselTop.wild.cpu.regs[0][12] ;
 wire \ChiselTop.wild.cpu.regs[0][13] ;
 wire \ChiselTop.wild.cpu.regs[0][14] ;
 wire \ChiselTop.wild.cpu.regs[0][15] ;
 wire \ChiselTop.wild.cpu.regs[0][16] ;
 wire \ChiselTop.wild.cpu.regs[0][17] ;
 wire \ChiselTop.wild.cpu.regs[0][18] ;
 wire \ChiselTop.wild.cpu.regs[0][19] ;
 wire \ChiselTop.wild.cpu.regs[0][1] ;
 wire \ChiselTop.wild.cpu.regs[0][20] ;
 wire \ChiselTop.wild.cpu.regs[0][21] ;
 wire \ChiselTop.wild.cpu.regs[0][22] ;
 wire \ChiselTop.wild.cpu.regs[0][23] ;
 wire \ChiselTop.wild.cpu.regs[0][24] ;
 wire \ChiselTop.wild.cpu.regs[0][25] ;
 wire \ChiselTop.wild.cpu.regs[0][26] ;
 wire \ChiselTop.wild.cpu.regs[0][27] ;
 wire \ChiselTop.wild.cpu.regs[0][28] ;
 wire \ChiselTop.wild.cpu.regs[0][29] ;
 wire \ChiselTop.wild.cpu.regs[0][2] ;
 wire \ChiselTop.wild.cpu.regs[0][30] ;
 wire \ChiselTop.wild.cpu.regs[0][31] ;
 wire \ChiselTop.wild.cpu.regs[0][3] ;
 wire \ChiselTop.wild.cpu.regs[0][4] ;
 wire \ChiselTop.wild.cpu.regs[0][5] ;
 wire \ChiselTop.wild.cpu.regs[0][6] ;
 wire \ChiselTop.wild.cpu.regs[0][7] ;
 wire \ChiselTop.wild.cpu.regs[0][8] ;
 wire \ChiselTop.wild.cpu.regs[0][9] ;
 wire \ChiselTop.wild.cpu.regs[1][0] ;
 wire \ChiselTop.wild.cpu.regs[1][10] ;
 wire \ChiselTop.wild.cpu.regs[1][11] ;
 wire \ChiselTop.wild.cpu.regs[1][12] ;
 wire \ChiselTop.wild.cpu.regs[1][13] ;
 wire \ChiselTop.wild.cpu.regs[1][14] ;
 wire \ChiselTop.wild.cpu.regs[1][15] ;
 wire \ChiselTop.wild.cpu.regs[1][16] ;
 wire \ChiselTop.wild.cpu.regs[1][17] ;
 wire \ChiselTop.wild.cpu.regs[1][18] ;
 wire \ChiselTop.wild.cpu.regs[1][19] ;
 wire \ChiselTop.wild.cpu.regs[1][1] ;
 wire \ChiselTop.wild.cpu.regs[1][20] ;
 wire \ChiselTop.wild.cpu.regs[1][21] ;
 wire \ChiselTop.wild.cpu.regs[1][22] ;
 wire \ChiselTop.wild.cpu.regs[1][23] ;
 wire \ChiselTop.wild.cpu.regs[1][24] ;
 wire \ChiselTop.wild.cpu.regs[1][25] ;
 wire \ChiselTop.wild.cpu.regs[1][26] ;
 wire \ChiselTop.wild.cpu.regs[1][27] ;
 wire \ChiselTop.wild.cpu.regs[1][28] ;
 wire \ChiselTop.wild.cpu.regs[1][29] ;
 wire \ChiselTop.wild.cpu.regs[1][2] ;
 wire \ChiselTop.wild.cpu.regs[1][30] ;
 wire \ChiselTop.wild.cpu.regs[1][31] ;
 wire \ChiselTop.wild.cpu.regs[1][3] ;
 wire \ChiselTop.wild.cpu.regs[1][4] ;
 wire \ChiselTop.wild.cpu.regs[1][5] ;
 wire \ChiselTop.wild.cpu.regs[1][6] ;
 wire \ChiselTop.wild.cpu.regs[1][7] ;
 wire \ChiselTop.wild.cpu.regs[1][8] ;
 wire \ChiselTop.wild.cpu.regs[1][9] ;
 wire \ChiselTop.wild.cpu.regs[28][0] ;
 wire \ChiselTop.wild.cpu.regs[28][10] ;
 wire \ChiselTop.wild.cpu.regs[28][11] ;
 wire \ChiselTop.wild.cpu.regs[28][12] ;
 wire \ChiselTop.wild.cpu.regs[28][13] ;
 wire \ChiselTop.wild.cpu.regs[28][14] ;
 wire \ChiselTop.wild.cpu.regs[28][15] ;
 wire \ChiselTop.wild.cpu.regs[28][16] ;
 wire \ChiselTop.wild.cpu.regs[28][17] ;
 wire \ChiselTop.wild.cpu.regs[28][18] ;
 wire \ChiselTop.wild.cpu.regs[28][19] ;
 wire \ChiselTop.wild.cpu.regs[28][1] ;
 wire \ChiselTop.wild.cpu.regs[28][20] ;
 wire \ChiselTop.wild.cpu.regs[28][21] ;
 wire \ChiselTop.wild.cpu.regs[28][22] ;
 wire \ChiselTop.wild.cpu.regs[28][23] ;
 wire \ChiselTop.wild.cpu.regs[28][24] ;
 wire \ChiselTop.wild.cpu.regs[28][25] ;
 wire \ChiselTop.wild.cpu.regs[28][26] ;
 wire \ChiselTop.wild.cpu.regs[28][27] ;
 wire \ChiselTop.wild.cpu.regs[28][28] ;
 wire \ChiselTop.wild.cpu.regs[28][29] ;
 wire \ChiselTop.wild.cpu.regs[28][2] ;
 wire \ChiselTop.wild.cpu.regs[28][30] ;
 wire \ChiselTop.wild.cpu.regs[28][31] ;
 wire \ChiselTop.wild.cpu.regs[28][3] ;
 wire \ChiselTop.wild.cpu.regs[28][4] ;
 wire \ChiselTop.wild.cpu.regs[28][5] ;
 wire \ChiselTop.wild.cpu.regs[28][6] ;
 wire \ChiselTop.wild.cpu.regs[28][7] ;
 wire \ChiselTop.wild.cpu.regs[28][8] ;
 wire \ChiselTop.wild.cpu.regs[28][9] ;
 wire \ChiselTop.wild.cpu.regs[29][0] ;
 wire \ChiselTop.wild.cpu.regs[29][10] ;
 wire \ChiselTop.wild.cpu.regs[29][11] ;
 wire \ChiselTop.wild.cpu.regs[29][12] ;
 wire \ChiselTop.wild.cpu.regs[29][13] ;
 wire \ChiselTop.wild.cpu.regs[29][14] ;
 wire \ChiselTop.wild.cpu.regs[29][15] ;
 wire \ChiselTop.wild.cpu.regs[29][16] ;
 wire \ChiselTop.wild.cpu.regs[29][17] ;
 wire \ChiselTop.wild.cpu.regs[29][18] ;
 wire \ChiselTop.wild.cpu.regs[29][19] ;
 wire \ChiselTop.wild.cpu.regs[29][1] ;
 wire \ChiselTop.wild.cpu.regs[29][20] ;
 wire \ChiselTop.wild.cpu.regs[29][21] ;
 wire \ChiselTop.wild.cpu.regs[29][22] ;
 wire \ChiselTop.wild.cpu.regs[29][23] ;
 wire \ChiselTop.wild.cpu.regs[29][24] ;
 wire \ChiselTop.wild.cpu.regs[29][25] ;
 wire \ChiselTop.wild.cpu.regs[29][26] ;
 wire \ChiselTop.wild.cpu.regs[29][27] ;
 wire \ChiselTop.wild.cpu.regs[29][28] ;
 wire \ChiselTop.wild.cpu.regs[29][29] ;
 wire \ChiselTop.wild.cpu.regs[29][2] ;
 wire \ChiselTop.wild.cpu.regs[29][30] ;
 wire \ChiselTop.wild.cpu.regs[29][31] ;
 wire \ChiselTop.wild.cpu.regs[29][3] ;
 wire \ChiselTop.wild.cpu.regs[29][4] ;
 wire \ChiselTop.wild.cpu.regs[29][5] ;
 wire \ChiselTop.wild.cpu.regs[29][6] ;
 wire \ChiselTop.wild.cpu.regs[29][7] ;
 wire \ChiselTop.wild.cpu.regs[29][8] ;
 wire \ChiselTop.wild.cpu.regs[29][9] ;
 wire \ChiselTop.wild.cpu.regs[2][0] ;
 wire \ChiselTop.wild.cpu.regs[2][10] ;
 wire \ChiselTop.wild.cpu.regs[2][11] ;
 wire \ChiselTop.wild.cpu.regs[2][12] ;
 wire \ChiselTop.wild.cpu.regs[2][13] ;
 wire \ChiselTop.wild.cpu.regs[2][14] ;
 wire \ChiselTop.wild.cpu.regs[2][15] ;
 wire \ChiselTop.wild.cpu.regs[2][16] ;
 wire \ChiselTop.wild.cpu.regs[2][17] ;
 wire \ChiselTop.wild.cpu.regs[2][18] ;
 wire \ChiselTop.wild.cpu.regs[2][19] ;
 wire \ChiselTop.wild.cpu.regs[2][1] ;
 wire \ChiselTop.wild.cpu.regs[2][20] ;
 wire \ChiselTop.wild.cpu.regs[2][21] ;
 wire \ChiselTop.wild.cpu.regs[2][22] ;
 wire \ChiselTop.wild.cpu.regs[2][23] ;
 wire \ChiselTop.wild.cpu.regs[2][24] ;
 wire \ChiselTop.wild.cpu.regs[2][25] ;
 wire \ChiselTop.wild.cpu.regs[2][26] ;
 wire \ChiselTop.wild.cpu.regs[2][27] ;
 wire \ChiselTop.wild.cpu.regs[2][28] ;
 wire \ChiselTop.wild.cpu.regs[2][29] ;
 wire \ChiselTop.wild.cpu.regs[2][2] ;
 wire \ChiselTop.wild.cpu.regs[2][30] ;
 wire \ChiselTop.wild.cpu.regs[2][31] ;
 wire \ChiselTop.wild.cpu.regs[2][3] ;
 wire \ChiselTop.wild.cpu.regs[2][4] ;
 wire \ChiselTop.wild.cpu.regs[2][5] ;
 wire \ChiselTop.wild.cpu.regs[2][6] ;
 wire \ChiselTop.wild.cpu.regs[2][7] ;
 wire \ChiselTop.wild.cpu.regs[2][8] ;
 wire \ChiselTop.wild.cpu.regs[2][9] ;
 wire \ChiselTop.wild.cpu.regs[30][0] ;
 wire \ChiselTop.wild.cpu.regs[30][10] ;
 wire \ChiselTop.wild.cpu.regs[30][11] ;
 wire \ChiselTop.wild.cpu.regs[30][12] ;
 wire \ChiselTop.wild.cpu.regs[30][13] ;
 wire \ChiselTop.wild.cpu.regs[30][14] ;
 wire \ChiselTop.wild.cpu.regs[30][15] ;
 wire \ChiselTop.wild.cpu.regs[30][16] ;
 wire \ChiselTop.wild.cpu.regs[30][17] ;
 wire \ChiselTop.wild.cpu.regs[30][18] ;
 wire \ChiselTop.wild.cpu.regs[30][19] ;
 wire \ChiselTop.wild.cpu.regs[30][1] ;
 wire \ChiselTop.wild.cpu.regs[30][20] ;
 wire \ChiselTop.wild.cpu.regs[30][21] ;
 wire \ChiselTop.wild.cpu.regs[30][22] ;
 wire \ChiselTop.wild.cpu.regs[30][23] ;
 wire \ChiselTop.wild.cpu.regs[30][24] ;
 wire \ChiselTop.wild.cpu.regs[30][25] ;
 wire \ChiselTop.wild.cpu.regs[30][26] ;
 wire \ChiselTop.wild.cpu.regs[30][27] ;
 wire \ChiselTop.wild.cpu.regs[30][28] ;
 wire \ChiselTop.wild.cpu.regs[30][29] ;
 wire \ChiselTop.wild.cpu.regs[30][2] ;
 wire \ChiselTop.wild.cpu.regs[30][30] ;
 wire \ChiselTop.wild.cpu.regs[30][31] ;
 wire \ChiselTop.wild.cpu.regs[30][3] ;
 wire \ChiselTop.wild.cpu.regs[30][4] ;
 wire \ChiselTop.wild.cpu.regs[30][5] ;
 wire \ChiselTop.wild.cpu.regs[30][6] ;
 wire \ChiselTop.wild.cpu.regs[30][7] ;
 wire \ChiselTop.wild.cpu.regs[30][8] ;
 wire \ChiselTop.wild.cpu.regs[30][9] ;
 wire \ChiselTop.wild.cpu.regs[31][0] ;
 wire \ChiselTop.wild.cpu.regs[31][10] ;
 wire \ChiselTop.wild.cpu.regs[31][11] ;
 wire \ChiselTop.wild.cpu.regs[31][12] ;
 wire \ChiselTop.wild.cpu.regs[31][13] ;
 wire \ChiselTop.wild.cpu.regs[31][14] ;
 wire \ChiselTop.wild.cpu.regs[31][15] ;
 wire \ChiselTop.wild.cpu.regs[31][16] ;
 wire \ChiselTop.wild.cpu.regs[31][17] ;
 wire \ChiselTop.wild.cpu.regs[31][18] ;
 wire \ChiselTop.wild.cpu.regs[31][19] ;
 wire \ChiselTop.wild.cpu.regs[31][1] ;
 wire \ChiselTop.wild.cpu.regs[31][20] ;
 wire \ChiselTop.wild.cpu.regs[31][21] ;
 wire \ChiselTop.wild.cpu.regs[31][22] ;
 wire \ChiselTop.wild.cpu.regs[31][23] ;
 wire \ChiselTop.wild.cpu.regs[31][24] ;
 wire \ChiselTop.wild.cpu.regs[31][25] ;
 wire \ChiselTop.wild.cpu.regs[31][26] ;
 wire \ChiselTop.wild.cpu.regs[31][27] ;
 wire \ChiselTop.wild.cpu.regs[31][28] ;
 wire \ChiselTop.wild.cpu.regs[31][29] ;
 wire \ChiselTop.wild.cpu.regs[31][2] ;
 wire \ChiselTop.wild.cpu.regs[31][30] ;
 wire \ChiselTop.wild.cpu.regs[31][31] ;
 wire \ChiselTop.wild.cpu.regs[31][3] ;
 wire \ChiselTop.wild.cpu.regs[31][4] ;
 wire \ChiselTop.wild.cpu.regs[31][5] ;
 wire \ChiselTop.wild.cpu.regs[31][6] ;
 wire \ChiselTop.wild.cpu.regs[31][7] ;
 wire \ChiselTop.wild.cpu.regs[31][8] ;
 wire \ChiselTop.wild.cpu.regs[31][9] ;
 wire \ChiselTop.wild.cpu.regs[3][0] ;
 wire \ChiselTop.wild.cpu.regs[3][10] ;
 wire \ChiselTop.wild.cpu.regs[3][11] ;
 wire \ChiselTop.wild.cpu.regs[3][12] ;
 wire \ChiselTop.wild.cpu.regs[3][13] ;
 wire \ChiselTop.wild.cpu.regs[3][14] ;
 wire \ChiselTop.wild.cpu.regs[3][15] ;
 wire \ChiselTop.wild.cpu.regs[3][16] ;
 wire \ChiselTop.wild.cpu.regs[3][17] ;
 wire \ChiselTop.wild.cpu.regs[3][18] ;
 wire \ChiselTop.wild.cpu.regs[3][19] ;
 wire \ChiselTop.wild.cpu.regs[3][1] ;
 wire \ChiselTop.wild.cpu.regs[3][20] ;
 wire \ChiselTop.wild.cpu.regs[3][21] ;
 wire \ChiselTop.wild.cpu.regs[3][22] ;
 wire \ChiselTop.wild.cpu.regs[3][23] ;
 wire \ChiselTop.wild.cpu.regs[3][24] ;
 wire \ChiselTop.wild.cpu.regs[3][25] ;
 wire \ChiselTop.wild.cpu.regs[3][26] ;
 wire \ChiselTop.wild.cpu.regs[3][27] ;
 wire \ChiselTop.wild.cpu.regs[3][28] ;
 wire \ChiselTop.wild.cpu.regs[3][29] ;
 wire \ChiselTop.wild.cpu.regs[3][2] ;
 wire \ChiselTop.wild.cpu.regs[3][30] ;
 wire \ChiselTop.wild.cpu.regs[3][31] ;
 wire \ChiselTop.wild.cpu.regs[3][3] ;
 wire \ChiselTop.wild.cpu.regs[3][4] ;
 wire \ChiselTop.wild.cpu.regs[3][5] ;
 wire \ChiselTop.wild.cpu.regs[3][6] ;
 wire \ChiselTop.wild.cpu.regs[3][7] ;
 wire \ChiselTop.wild.cpu.regs[3][8] ;
 wire \ChiselTop.wild.cpu.regs[3][9] ;
 wire \ChiselTop.wild.cpu.regs[4][0] ;
 wire \ChiselTop.wild.cpu.regs[4][10] ;
 wire \ChiselTop.wild.cpu.regs[4][11] ;
 wire \ChiselTop.wild.cpu.regs[4][12] ;
 wire \ChiselTop.wild.cpu.regs[4][13] ;
 wire \ChiselTop.wild.cpu.regs[4][14] ;
 wire \ChiselTop.wild.cpu.regs[4][15] ;
 wire \ChiselTop.wild.cpu.regs[4][16] ;
 wire \ChiselTop.wild.cpu.regs[4][17] ;
 wire \ChiselTop.wild.cpu.regs[4][18] ;
 wire \ChiselTop.wild.cpu.regs[4][19] ;
 wire \ChiselTop.wild.cpu.regs[4][1] ;
 wire \ChiselTop.wild.cpu.regs[4][20] ;
 wire \ChiselTop.wild.cpu.regs[4][21] ;
 wire \ChiselTop.wild.cpu.regs[4][22] ;
 wire \ChiselTop.wild.cpu.regs[4][23] ;
 wire \ChiselTop.wild.cpu.regs[4][24] ;
 wire \ChiselTop.wild.cpu.regs[4][25] ;
 wire \ChiselTop.wild.cpu.regs[4][26] ;
 wire \ChiselTop.wild.cpu.regs[4][27] ;
 wire \ChiselTop.wild.cpu.regs[4][28] ;
 wire \ChiselTop.wild.cpu.regs[4][29] ;
 wire \ChiselTop.wild.cpu.regs[4][2] ;
 wire \ChiselTop.wild.cpu.regs[4][30] ;
 wire \ChiselTop.wild.cpu.regs[4][31] ;
 wire \ChiselTop.wild.cpu.regs[4][3] ;
 wire \ChiselTop.wild.cpu.regs[4][4] ;
 wire \ChiselTop.wild.cpu.regs[4][5] ;
 wire \ChiselTop.wild.cpu.regs[4][6] ;
 wire \ChiselTop.wild.cpu.regs[4][7] ;
 wire \ChiselTop.wild.cpu.regs[4][8] ;
 wire \ChiselTop.wild.cpu.regs[4][9] ;
 wire \ChiselTop.wild.cpu.regs[5][0] ;
 wire \ChiselTop.wild.cpu.regs[5][10] ;
 wire \ChiselTop.wild.cpu.regs[5][11] ;
 wire \ChiselTop.wild.cpu.regs[5][12] ;
 wire \ChiselTop.wild.cpu.regs[5][13] ;
 wire \ChiselTop.wild.cpu.regs[5][14] ;
 wire \ChiselTop.wild.cpu.regs[5][15] ;
 wire \ChiselTop.wild.cpu.regs[5][16] ;
 wire \ChiselTop.wild.cpu.regs[5][17] ;
 wire \ChiselTop.wild.cpu.regs[5][18] ;
 wire \ChiselTop.wild.cpu.regs[5][19] ;
 wire \ChiselTop.wild.cpu.regs[5][1] ;
 wire \ChiselTop.wild.cpu.regs[5][20] ;
 wire \ChiselTop.wild.cpu.regs[5][21] ;
 wire \ChiselTop.wild.cpu.regs[5][22] ;
 wire \ChiselTop.wild.cpu.regs[5][23] ;
 wire \ChiselTop.wild.cpu.regs[5][24] ;
 wire \ChiselTop.wild.cpu.regs[5][25] ;
 wire \ChiselTop.wild.cpu.regs[5][26] ;
 wire \ChiselTop.wild.cpu.regs[5][27] ;
 wire \ChiselTop.wild.cpu.regs[5][28] ;
 wire \ChiselTop.wild.cpu.regs[5][29] ;
 wire \ChiselTop.wild.cpu.regs[5][2] ;
 wire \ChiselTop.wild.cpu.regs[5][30] ;
 wire \ChiselTop.wild.cpu.regs[5][31] ;
 wire \ChiselTop.wild.cpu.regs[5][3] ;
 wire \ChiselTop.wild.cpu.regs[5][4] ;
 wire \ChiselTop.wild.cpu.regs[5][5] ;
 wire \ChiselTop.wild.cpu.regs[5][6] ;
 wire \ChiselTop.wild.cpu.regs[5][7] ;
 wire \ChiselTop.wild.cpu.regs[5][8] ;
 wire \ChiselTop.wild.cpu.regs[5][9] ;
 wire \ChiselTop.wild.cpu.regs[6][0] ;
 wire \ChiselTop.wild.cpu.regs[6][10] ;
 wire \ChiselTop.wild.cpu.regs[6][11] ;
 wire \ChiselTop.wild.cpu.regs[6][12] ;
 wire \ChiselTop.wild.cpu.regs[6][13] ;
 wire \ChiselTop.wild.cpu.regs[6][14] ;
 wire \ChiselTop.wild.cpu.regs[6][15] ;
 wire \ChiselTop.wild.cpu.regs[6][16] ;
 wire \ChiselTop.wild.cpu.regs[6][17] ;
 wire \ChiselTop.wild.cpu.regs[6][18] ;
 wire \ChiselTop.wild.cpu.regs[6][19] ;
 wire \ChiselTop.wild.cpu.regs[6][1] ;
 wire \ChiselTop.wild.cpu.regs[6][20] ;
 wire \ChiselTop.wild.cpu.regs[6][21] ;
 wire \ChiselTop.wild.cpu.regs[6][22] ;
 wire \ChiselTop.wild.cpu.regs[6][23] ;
 wire \ChiselTop.wild.cpu.regs[6][24] ;
 wire \ChiselTop.wild.cpu.regs[6][25] ;
 wire \ChiselTop.wild.cpu.regs[6][26] ;
 wire \ChiselTop.wild.cpu.regs[6][27] ;
 wire \ChiselTop.wild.cpu.regs[6][28] ;
 wire \ChiselTop.wild.cpu.regs[6][29] ;
 wire \ChiselTop.wild.cpu.regs[6][2] ;
 wire \ChiselTop.wild.cpu.regs[6][30] ;
 wire \ChiselTop.wild.cpu.regs[6][31] ;
 wire \ChiselTop.wild.cpu.regs[6][3] ;
 wire \ChiselTop.wild.cpu.regs[6][4] ;
 wire \ChiselTop.wild.cpu.regs[6][5] ;
 wire \ChiselTop.wild.cpu.regs[6][6] ;
 wire \ChiselTop.wild.cpu.regs[6][7] ;
 wire \ChiselTop.wild.cpu.regs[6][8] ;
 wire \ChiselTop.wild.cpu.regs[6][9] ;
 wire \ChiselTop.wild.cpu.regs[7][0] ;
 wire \ChiselTop.wild.cpu.regs[7][10] ;
 wire \ChiselTop.wild.cpu.regs[7][11] ;
 wire \ChiselTop.wild.cpu.regs[7][12] ;
 wire \ChiselTop.wild.cpu.regs[7][13] ;
 wire \ChiselTop.wild.cpu.regs[7][14] ;
 wire \ChiselTop.wild.cpu.regs[7][15] ;
 wire \ChiselTop.wild.cpu.regs[7][16] ;
 wire \ChiselTop.wild.cpu.regs[7][17] ;
 wire \ChiselTop.wild.cpu.regs[7][18] ;
 wire \ChiselTop.wild.cpu.regs[7][19] ;
 wire \ChiselTop.wild.cpu.regs[7][1] ;
 wire \ChiselTop.wild.cpu.regs[7][20] ;
 wire \ChiselTop.wild.cpu.regs[7][21] ;
 wire \ChiselTop.wild.cpu.regs[7][22] ;
 wire \ChiselTop.wild.cpu.regs[7][23] ;
 wire \ChiselTop.wild.cpu.regs[7][24] ;
 wire \ChiselTop.wild.cpu.regs[7][25] ;
 wire \ChiselTop.wild.cpu.regs[7][26] ;
 wire \ChiselTop.wild.cpu.regs[7][27] ;
 wire \ChiselTop.wild.cpu.regs[7][28] ;
 wire \ChiselTop.wild.cpu.regs[7][29] ;
 wire \ChiselTop.wild.cpu.regs[7][2] ;
 wire \ChiselTop.wild.cpu.regs[7][30] ;
 wire \ChiselTop.wild.cpu.regs[7][31] ;
 wire \ChiselTop.wild.cpu.regs[7][3] ;
 wire \ChiselTop.wild.cpu.regs[7][4] ;
 wire \ChiselTop.wild.cpu.regs[7][5] ;
 wire \ChiselTop.wild.cpu.regs[7][6] ;
 wire \ChiselTop.wild.cpu.regs[7][7] ;
 wire \ChiselTop.wild.cpu.regs[7][8] ;
 wire \ChiselTop.wild.cpu.regs[7][9] ;
 wire \ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[0] ;
 wire \ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[1] ;
 wire \ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[2] ;
 wire \ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[0] ;
 wire \ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[1] ;
 wire \ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[2] ;
 wire \ChiselTop.wild.dmem.MEM[0][0] ;
 wire \ChiselTop.wild.dmem.MEM[0][1] ;
 wire \ChiselTop.wild.dmem.MEM[0][2] ;
 wire \ChiselTop.wild.dmem.MEM[0][3] ;
 wire \ChiselTop.wild.dmem.MEM[0][4] ;
 wire \ChiselTop.wild.dmem.MEM[0][5] ;
 wire \ChiselTop.wild.dmem.MEM[0][6] ;
 wire \ChiselTop.wild.dmem.MEM[0][7] ;
 wire \ChiselTop.wild.dmem.MEM_1[0][0] ;
 wire \ChiselTop.wild.dmem.MEM_1[0][1] ;
 wire \ChiselTop.wild.dmem.MEM_1[0][2] ;
 wire \ChiselTop.wild.dmem.MEM_1[0][3] ;
 wire \ChiselTop.wild.dmem.MEM_1[0][4] ;
 wire \ChiselTop.wild.dmem.MEM_1[0][5] ;
 wire \ChiselTop.wild.dmem.MEM_1[0][6] ;
 wire \ChiselTop.wild.dmem.MEM_1[0][7] ;
 wire \ChiselTop.wild.dmem.MEM_2[0][0] ;
 wire \ChiselTop.wild.dmem.MEM_2[0][1] ;
 wire \ChiselTop.wild.dmem.MEM_2[0][2] ;
 wire \ChiselTop.wild.dmem.MEM_2[0][3] ;
 wire \ChiselTop.wild.dmem.MEM_2[0][4] ;
 wire \ChiselTop.wild.dmem.MEM_2[0][5] ;
 wire \ChiselTop.wild.dmem.MEM_2[0][6] ;
 wire \ChiselTop.wild.dmem.MEM_2[0][7] ;
 wire \ChiselTop.wild.dmem.MEM_3[0][0] ;
 wire \ChiselTop.wild.dmem.MEM_3[0][1] ;
 wire \ChiselTop.wild.dmem.MEM_3[0][2] ;
 wire \ChiselTop.wild.dmem.MEM_3[0][3] ;
 wire \ChiselTop.wild.dmem.MEM_3[0][4] ;
 wire \ChiselTop.wild.dmem.MEM_3[0][5] ;
 wire \ChiselTop.wild.dmem.MEM_3[0][6] ;
 wire \ChiselTop.wild.dmem.MEM_3[0][7] ;
 wire \ChiselTop.wild.ledReg[0] ;
 wire \ChiselTop.wild.ledReg[1] ;
 wire \ChiselTop.wild.ledReg[2] ;
 wire \ChiselTop.wild.ledReg[3] ;
 wire \ChiselTop.wild.memAddressReg[0] ;
 wire \ChiselTop.wild.memAddressReg[16] ;
 wire \ChiselTop.wild.memAddressReg[17] ;
 wire \ChiselTop.wild.memAddressReg[18] ;
 wire \ChiselTop.wild.memAddressReg[19] ;
 wire \ChiselTop.wild.memAddressReg[1] ;
 wire \ChiselTop.wild.memAddressReg[28] ;
 wire \ChiselTop.wild.memAddressReg[29] ;
 wire \ChiselTop.wild.memAddressReg[2] ;
 wire \ChiselTop.wild.memAddressReg[30] ;
 wire \ChiselTop.wild.memAddressReg[31] ;
 wire \ChiselTop.wild.memAddressReg[3] ;
 wire \ChiselTop.wild.rx._shiftReg_T_1[0] ;
 wire \ChiselTop.wild.rx._shiftReg_T_1[1] ;
 wire \ChiselTop.wild.rx._shiftReg_T_1[2] ;
 wire \ChiselTop.wild.rx._shiftReg_T_1[3] ;
 wire \ChiselTop.wild.rx._shiftReg_T_1[4] ;
 wire \ChiselTop.wild.rx._shiftReg_T_1[5] ;
 wire \ChiselTop.wild.rx._shiftReg_T_1[6] ;
 wire \ChiselTop.wild.rx._shiftReg_T_1[7] ;
 wire \ChiselTop.wild.rx.bitsReg[0] ;
 wire \ChiselTop.wild.rx.bitsReg[1] ;
 wire \ChiselTop.wild.rx.bitsReg[2] ;
 wire \ChiselTop.wild.rx.bitsReg[3] ;
 wire \ChiselTop.wild.rx.cntReg[0] ;
 wire \ChiselTop.wild.rx.cntReg[10] ;
 wire \ChiselTop.wild.rx.cntReg[11] ;
 wire \ChiselTop.wild.rx.cntReg[12] ;
 wire \ChiselTop.wild.rx.cntReg[13] ;
 wire \ChiselTop.wild.rx.cntReg[14] ;
 wire \ChiselTop.wild.rx.cntReg[15] ;
 wire \ChiselTop.wild.rx.cntReg[16] ;
 wire \ChiselTop.wild.rx.cntReg[17] ;
 wire \ChiselTop.wild.rx.cntReg[18] ;
 wire \ChiselTop.wild.rx.cntReg[19] ;
 wire \ChiselTop.wild.rx.cntReg[1] ;
 wire \ChiselTop.wild.rx.cntReg[2] ;
 wire \ChiselTop.wild.rx.cntReg[3] ;
 wire \ChiselTop.wild.rx.cntReg[4] ;
 wire \ChiselTop.wild.rx.cntReg[5] ;
 wire \ChiselTop.wild.rx.cntReg[6] ;
 wire \ChiselTop.wild.rx.cntReg[7] ;
 wire \ChiselTop.wild.rx.cntReg[8] ;
 wire \ChiselTop.wild.rx.cntReg[9] ;
 wire \ChiselTop.wild.rx.falling_REG ;
 wire \ChiselTop.wild.rx.io_channel_bits[0] ;
 wire \ChiselTop.wild.rx.io_channel_valid ;
 wire \ChiselTop.wild.rx.rxReg_REG ;
 wire \ChiselTop.wild.tx.buf_.io_in_ready ;
 wire \ChiselTop.wild.tx.buf_.io_out_valid ;
 wire \ChiselTop.wild.tx.tx.bitsReg[0] ;
 wire \ChiselTop.wild.tx.tx.bitsReg[1] ;
 wire \ChiselTop.wild.tx.tx.bitsReg[2] ;
 wire \ChiselTop.wild.tx.tx.bitsReg[3] ;
 wire \ChiselTop.wild.tx.tx.cntReg[0] ;
 wire \ChiselTop.wild.tx.tx.cntReg[10] ;
 wire \ChiselTop.wild.tx.tx.cntReg[11] ;
 wire \ChiselTop.wild.tx.tx.cntReg[12] ;
 wire \ChiselTop.wild.tx.tx.cntReg[13] ;
 wire \ChiselTop.wild.tx.tx.cntReg[14] ;
 wire \ChiselTop.wild.tx.tx.cntReg[15] ;
 wire \ChiselTop.wild.tx.tx.cntReg[16] ;
 wire \ChiselTop.wild.tx.tx.cntReg[17] ;
 wire \ChiselTop.wild.tx.tx.cntReg[18] ;
 wire \ChiselTop.wild.tx.tx.cntReg[19] ;
 wire \ChiselTop.wild.tx.tx.cntReg[1] ;
 wire \ChiselTop.wild.tx.tx.cntReg[2] ;
 wire \ChiselTop.wild.tx.tx.cntReg[3] ;
 wire \ChiselTop.wild.tx.tx.cntReg[4] ;
 wire \ChiselTop.wild.tx.tx.cntReg[5] ;
 wire \ChiselTop.wild.tx.tx.cntReg[6] ;
 wire \ChiselTop.wild.tx.tx.cntReg[7] ;
 wire \ChiselTop.wild.tx.tx.cntReg[8] ;
 wire \ChiselTop.wild.tx.tx.cntReg[9] ;
 wire \ChiselTop.wild.uartStatusReg[0] ;
 wire \ChiselTop.wild.uartStatusReg[1] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire clknet_leaf_0_clk;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;

 sg13g2_inv_1 _06133_ (.Y(_00893_),
    .A(net861));
 sg13g2_inv_1 _06134_ (.Y(_00894_),
    .A(net1220));
 sg13g2_inv_1 _06135_ (.Y(_00895_),
    .A(net1185));
 sg13g2_inv_1 _06136_ (.Y(_00896_),
    .A(net1387));
 sg13g2_inv_1 _06137_ (.Y(_00897_),
    .A(net1413));
 sg13g2_inv_1 _06138_ (.Y(_00898_),
    .A(net1383));
 sg13g2_inv_1 _06139_ (.Y(_00899_),
    .A(net1276));
 sg13g2_inv_1 _06140_ (.Y(_00900_),
    .A(net1279));
 sg13g2_inv_1 _06141_ (.Y(_00901_),
    .A(net1064));
 sg13g2_inv_1 _06142_ (.Y(_00902_),
    .A(\ChiselTop.wild.rx.bitsReg[0] ));
 sg13g2_inv_1 _06143_ (.Y(_00903_),
    .A(net827));
 sg13g2_inv_1 _06144_ (.Y(_00904_),
    .A(net831));
 sg13g2_inv_1 _06145_ (.Y(_00905_),
    .A(net830));
 sg13g2_inv_1 _06146_ (.Y(_00906_),
    .A(net834));
 sg13g2_inv_1 _06147_ (.Y(_00907_),
    .A(net2619));
 sg13g2_inv_1 _06148_ (.Y(_00908_),
    .A(net2643));
 sg13g2_inv_1 _06149_ (.Y(_00909_),
    .A(_00010_));
 sg13g2_inv_1 _06150_ (.Y(_00910_),
    .A(_00014_));
 sg13g2_inv_1 _06151_ (.Y(_00911_),
    .A(_00023_));
 sg13g2_inv_1 _06152_ (.Y(_00912_),
    .A(_00036_));
 sg13g2_inv_1 _06153_ (.Y(_00913_),
    .A(_00040_));
 sg13g2_inv_1 _06154_ (.Y(_00914_),
    .A(_00043_));
 sg13g2_inv_2 _06155_ (.Y(_00915_),
    .A(_00053_));
 sg13g2_inv_1 _06156_ (.Y(_00916_),
    .A(_00068_));
 sg13g2_inv_1 _06157_ (.Y(_00917_),
    .A(_00070_));
 sg13g2_inv_1 _06158_ (.Y(_00918_),
    .A(_00084_));
 sg13g2_inv_1 _06159_ (.Y(_00919_),
    .A(_00086_));
 sg13g2_inv_2 _06160_ (.Y(_00920_),
    .A(_00088_));
 sg13g2_inv_1 _06161_ (.Y(_00921_),
    .A(\ChiselTop.wild.cpu.decExReg_rs1Val[30] ));
 sg13g2_inv_1 _06162_ (.Y(_00922_),
    .A(\ChiselTop.wild.cpu.decExReg_rs1Val[31] ));
 sg13g2_inv_1 _06163_ (.Y(_00923_),
    .A(net2639));
 sg13g2_inv_1 _06164_ (.Y(_00924_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[10] ));
 sg13g2_inv_2 _06165_ (.Y(_00925_),
    .A(net2630));
 sg13g2_inv_1 _06166_ (.Y(_00926_),
    .A(\ChiselTop.wild.memAddressReg[2] ));
 sg13g2_inv_1 _06167_ (.Y(_00927_),
    .A(\ChiselTop.wild.cpu.decOut_opcode[5] ));
 sg13g2_inv_1 _06168_ (.Y(_00928_),
    .A(net2550));
 sg13g2_inv_2 _06169_ (.Y(_00929_),
    .A(net1521));
 sg13g2_inv_1 _06170_ (.Y(_00930_),
    .A(_00114_));
 sg13g2_inv_1 _06171_ (.Y(_00931_),
    .A(net1458));
 sg13g2_inv_1 _06172_ (.Y(_00932_),
    .A(net1337));
 sg13g2_inv_1 _06173_ (.Y(_00933_),
    .A(net1325));
 sg13g2_inv_1 _06174_ (.Y(_00934_),
    .A(_00126_));
 sg13g2_inv_1 _06175_ (.Y(_00935_),
    .A(_00132_));
 sg13g2_inv_1 _06176_ (.Y(_00936_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[17] ));
 sg13g2_inv_1 _06177_ (.Y(_00937_),
    .A(_00133_));
 sg13g2_inv_1 _06178_ (.Y(_00938_),
    .A(net1353));
 sg13g2_inv_1 _06179_ (.Y(_00939_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[20] ));
 sg13g2_inv_1 _06180_ (.Y(_00940_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[17] ));
 sg13g2_inv_1 _06181_ (.Y(_00941_),
    .A(net1478));
 sg13g2_inv_1 _06182_ (.Y(_00942_),
    .A(net1533));
 sg13g2_inv_1 _06183_ (.Y(_00943_),
    .A(net2743));
 sg13g2_inv_1 _06184_ (.Y(_00944_),
    .A(net930));
 sg13g2_inv_1 _06185_ (.Y(_00945_),
    .A(\ChiselTop.cntReg[11] ));
 sg13g2_inv_1 _06186_ (.Y(_00946_),
    .A(\ChiselTop.cntReg[15] ));
 sg13g2_inv_1 _06187_ (.Y(_00947_),
    .A(\ChiselTop.cntReg[18] ));
 sg13g2_inv_1 _06188_ (.Y(_00948_),
    .A(\ChiselTop.cntReg[24] ));
 sg13g2_inv_1 _06189_ (.Y(_00949_),
    .A(\ChiselTop.dec.counter[0] ));
 sg13g2_inv_1 _06190_ (.Y(_00950_),
    .A(\ChiselTop.dec.counter[3] ));
 sg13g2_inv_1 _06191_ (.Y(_00951_),
    .A(\ChiselTop.dec.counter[2] ));
 sg13g2_inv_1 _06192_ (.Y(_00952_),
    .A(net832));
 sg13g2_inv_1 _06193_ (.Y(_00953_),
    .A(net844));
 sg13g2_inv_1 _06194_ (.Y(_00954_),
    .A(net852));
 sg13g2_inv_1 _06195_ (.Y(_00955_),
    .A(net835));
 sg13g2_inv_1 _06196_ (.Y(_00956_),
    .A(net828));
 sg13g2_inv_1 _06197_ (.Y(_00957_),
    .A(net869));
 sg13g2_inv_1 _06198_ (.Y(_00958_),
    .A(net939));
 sg13g2_inv_1 _06199_ (.Y(_00959_),
    .A(net853));
 sg13g2_nand2_1 _06200_ (.Y(_00960_),
    .A(\ChiselTop.wild.cpu.decOut_opcode[4] ),
    .B(\ChiselTop.wild.cpu.decOut_opcode[2] ));
 sg13g2_nor2_2 _06201_ (.A(net2550),
    .B(_00960_),
    .Y(_00961_));
 sg13g2_nand2b_1 _06202_ (.Y(_00962_),
    .B(net2528),
    .A_N(_00960_));
 sg13g2_nor2_2 _06203_ (.A(_00110_),
    .B(_00961_),
    .Y(_00963_));
 sg13g2_nand2b_2 _06204_ (.Y(_00964_),
    .B(net2522),
    .A_N(_00110_));
 sg13g2_o21ai_1 _06205_ (.B1(_00964_),
    .Y(_00965_),
    .A1(_00111_),
    .A2(net2522));
 sg13g2_nor2_1 _06206_ (.A(\ChiselTop.wild.cpu.decExReg_rd[1] ),
    .B(\ChiselTop.wild.cpu.decExReg_rd[0] ),
    .Y(_00966_));
 sg13g2_nor2_2 _06207_ (.A(\ChiselTop.wild.cpu.decExReg_rd[3] ),
    .B(net2612),
    .Y(_00967_));
 sg13g2_nor3_1 _06208_ (.A(\ChiselTop.wild.cpu.decExReg_rd[2] ),
    .B(\ChiselTop.wild.cpu.decExReg_rd[3] ),
    .C(net2612),
    .Y(_00968_));
 sg13g2_nand2_1 _06209_ (.Y(_00969_),
    .A(_00966_),
    .B(_00968_));
 sg13g2_nand3_1 _06210_ (.B(net1488),
    .C(_00969_),
    .A(net1519),
    .Y(_00970_));
 sg13g2_xnor2_1 _06211_ (.Y(_00971_),
    .A(net2649),
    .B(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[15] ));
 sg13g2_xor2_1 _06212_ (.B(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[17] ),
    .A(\ChiselTop.wild.cpu.decExReg_rd[2] ),
    .X(_00972_));
 sg13g2_xnor2_1 _06213_ (.Y(_00973_),
    .A(net2648),
    .B(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[16] ));
 sg13g2_nand3_1 _06214_ (.B(_00971_),
    .C(_00973_),
    .A(_00967_),
    .Y(_00974_));
 sg13g2_nor3_2 _06215_ (.A(_00970_),
    .B(_00972_),
    .C(_00974_),
    .Y(_00975_));
 sg13g2_inv_2 _06216_ (.Y(_00976_),
    .A(net2441));
 sg13g2_nand3_1 _06217_ (.B(\ChiselTop.wild.cpu.decExReg_pc[3] ),
    .C(\ChiselTop.wild.cpu.decExReg_pc[2] ),
    .A(\ChiselTop.wild.cpu.decExReg_pc[4] ),
    .Y(_00977_));
 sg13g2_nand4_1 _06218_ (.B(\ChiselTop.wild.cpu.decExReg_pc[4] ),
    .C(\ChiselTop.wild.cpu.decExReg_pc[3] ),
    .A(\ChiselTop.wild.cpu.decExReg_pc[5] ),
    .Y(_00978_),
    .D(\ChiselTop.wild.cpu.decExReg_pc[2] ));
 sg13g2_nand2_1 _06219_ (.Y(_00979_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[7] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[6] ));
 sg13g2_nor2_1 _06220_ (.A(_00978_),
    .B(_00979_),
    .Y(_00980_));
 sg13g2_nand3_1 _06221_ (.B(\ChiselTop.wild.cpu.decExReg_pc[8] ),
    .C(_00980_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[9] ),
    .Y(_00981_));
 sg13g2_nor2_1 _06222_ (.A(_00924_),
    .B(_00981_),
    .Y(_00982_));
 sg13g2_and2_1 _06223_ (.A(\ChiselTop.wild.cpu.decExReg_pc[11] ),
    .B(_00982_),
    .X(_00983_));
 sg13g2_and2_1 _06224_ (.A(\ChiselTop.wild.cpu.decExReg_pc[12] ),
    .B(_00983_),
    .X(_00984_));
 sg13g2_and3_2 _06225_ (.X(_00985_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[14] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[13] ),
    .C(_00984_));
 sg13g2_nand3_1 _06226_ (.B(\ChiselTop.wild.cpu.decExReg_pc[15] ),
    .C(_00985_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[16] ),
    .Y(_00986_));
 sg13g2_a21oi_1 _06227_ (.A1(\ChiselTop.wild.cpu.decExReg_pc[15] ),
    .A2(_00985_),
    .Y(_00987_),
    .B1(\ChiselTop.wild.cpu.decExReg_pc[16] ));
 sg13g2_nor2_2 _06228_ (.A(\ChiselTop.wild.cpu.exFwdReg_wbDest[3] ),
    .B(\ChiselTop.wild.cpu.exFwdReg_wbDest[4] ),
    .Y(_00988_));
 sg13g2_and2_2 _06229_ (.A(\ChiselTop.wild.cpu.exFwdReg_valid ),
    .B(_00988_),
    .X(_00989_));
 sg13g2_nand2_2 _06230_ (.Y(_00990_),
    .A(\ChiselTop.wild.cpu.exFwdReg_valid ),
    .B(_00988_));
 sg13g2_xnor2_1 _06231_ (.Y(_00991_),
    .A(\ChiselTop.wild.cpu.exFwdReg_wbDest[1] ),
    .B(\ChiselTop.wild.cpu.decExReg_rs1[1] ));
 sg13g2_xnor2_1 _06232_ (.Y(_00992_),
    .A(\ChiselTop.wild.cpu.exFwdReg_wbDest[0] ),
    .B(\ChiselTop.wild.cpu.decExReg_rs1[0] ));
 sg13g2_xnor2_1 _06233_ (.Y(_00993_),
    .A(\ChiselTop.wild.cpu.exFwdReg_wbDest[2] ),
    .B(\ChiselTop.wild.cpu.decExReg_rs1[2] ));
 sg13g2_and3_2 _06234_ (.X(_00994_),
    .A(_00991_),
    .B(_00992_),
    .C(_00993_));
 sg13g2_nand3_1 _06235_ (.B(_00992_),
    .C(_00993_),
    .A(_00991_),
    .Y(_00995_));
 sg13g2_nor2_1 _06236_ (.A(_00990_),
    .B(_00995_),
    .Y(_00996_));
 sg13g2_a21oi_2 _06237_ (.B1(_00919_),
    .Y(_00997_),
    .A2(net2518),
    .A1(net2520));
 sg13g2_a21oi_2 _06238_ (.B1(_00997_),
    .Y(_00998_),
    .A2(net2456),
    .A1(_00085_));
 sg13g2_a21o_2 _06239_ (.A2(net2456),
    .A1(_00085_),
    .B1(_00997_),
    .X(_00999_));
 sg13g2_nand4_1 _06240_ (.B(\ChiselTop.wild.cpu.exFwdReg_wbDest[2] ),
    .C(\ChiselTop.wild.cpu.exFwdReg_wbDest[3] ),
    .A(\ChiselTop.wild.cpu.decExReg_rs2[2] ),
    .Y(_01000_),
    .D(\ChiselTop.wild.cpu.exFwdReg_wbDest[4] ));
 sg13g2_or4_1 _06241_ (.A(\ChiselTop.wild.cpu.decExReg_rs2[2] ),
    .B(\ChiselTop.wild.cpu.exFwdReg_wbDest[2] ),
    .C(\ChiselTop.wild.cpu.exFwdReg_wbDest[3] ),
    .D(\ChiselTop.wild.cpu.exFwdReg_wbDest[4] ),
    .X(_01001_));
 sg13g2_nand2b_1 _06242_ (.Y(_01002_),
    .B(\ChiselTop.wild.cpu.decExReg_rs2[0] ),
    .A_N(\ChiselTop.wild.cpu.exFwdReg_wbDest[0] ));
 sg13g2_nand2b_1 _06243_ (.Y(_01003_),
    .B(\ChiselTop.wild.cpu.exFwdReg_wbDest[0] ),
    .A_N(\ChiselTop.wild.cpu.decExReg_rs2[0] ));
 sg13g2_and3_1 _06244_ (.X(_01004_),
    .A(\ChiselTop.wild.cpu.exFwdReg_valid ),
    .B(_01002_),
    .C(_01003_));
 sg13g2_nand3_1 _06245_ (.B(_01002_),
    .C(_01003_),
    .A(\ChiselTop.wild.cpu.exFwdReg_valid ),
    .Y(_01005_));
 sg13g2_xor2_1 _06246_ (.B(\ChiselTop.wild.cpu.exFwdReg_wbDest[1] ),
    .A(\ChiselTop.wild.cpu.decExReg_rs2[1] ),
    .X(_01006_));
 sg13g2_a21oi_1 _06247_ (.A1(_01000_),
    .A2(_01001_),
    .Y(_01007_),
    .B1(_01006_));
 sg13g2_a21o_2 _06248_ (.A2(_01001_),
    .A1(_01000_),
    .B1(_01006_),
    .X(_01008_));
 sg13g2_nand2_1 _06249_ (.Y(_01009_),
    .A(net2514),
    .B(net2509));
 sg13g2_a21oi_2 _06250_ (.B1(_00100_),
    .Y(_01010_),
    .A2(net2512),
    .A1(net2517));
 sg13g2_nor3_1 _06251_ (.A(_00085_),
    .B(net2513),
    .C(net2508),
    .Y(_01011_));
 sg13g2_nor2_1 _06252_ (.A(_01010_),
    .B(_01011_),
    .Y(_01012_));
 sg13g2_xnor2_1 _06253_ (.Y(_01013_),
    .A(_00999_),
    .B(_01012_));
 sg13g2_mux2_1 _06254_ (.A0(_00074_),
    .A1(_00073_),
    .S(net2452),
    .X(_01014_));
 sg13g2_inv_2 _06255_ (.Y(_01015_),
    .A(_01014_));
 sg13g2_and3_1 _06256_ (.X(_01016_),
    .A(_00073_),
    .B(net2514),
    .C(net2509));
 sg13g2_a21oi_2 _06257_ (.B1(_01016_),
    .Y(_01017_),
    .A2(net2449),
    .A1(_00106_));
 sg13g2_a21oi_1 _06258_ (.A1(net2515),
    .A2(net2510),
    .Y(_01018_),
    .B1(_00038_));
 sg13g2_nor3_1 _06259_ (.A(_00039_),
    .B(net2513),
    .C(net2508),
    .Y(_01019_));
 sg13g2_nor2_1 _06260_ (.A(_01018_),
    .B(_01019_),
    .Y(_01020_));
 sg13g2_a21oi_2 _06261_ (.B1(_00913_),
    .Y(_01021_),
    .A2(net2519),
    .A1(net2521));
 sg13g2_a21oi_2 _06262_ (.B1(_01021_),
    .Y(_01022_),
    .A2(net2455),
    .A1(_00039_));
 sg13g2_a21o_2 _06263_ (.A2(net2455),
    .A1(_00039_),
    .B1(_01021_),
    .X(_01023_));
 sg13g2_mux2_2 _06264_ (.A0(_00057_),
    .A1(_00056_),
    .S(net2454),
    .X(_01024_));
 sg13g2_inv_2 _06265_ (.Y(_01025_),
    .A(_01024_));
 sg13g2_mux2_2 _06266_ (.A0(_00056_),
    .A1(_00055_),
    .S(net2450),
    .X(_01026_));
 sg13g2_mux2_2 _06267_ (.A0(_00047_),
    .A1(_00046_),
    .S(net2454),
    .X(_01027_));
 sg13g2_inv_1 _06268_ (.Y(_01028_),
    .A(net2435));
 sg13g2_nand3_1 _06269_ (.B(net2515),
    .C(net2510),
    .A(_00046_),
    .Y(_01029_));
 sg13g2_o21ai_1 _06270_ (.B1(_00045_),
    .Y(_01030_),
    .A1(net2513),
    .A2(net2508));
 sg13g2_nand2_1 _06271_ (.Y(_01031_),
    .A(_01029_),
    .B(_01030_));
 sg13g2_a21o_1 _06272_ (.A2(net2509),
    .A1(net2514),
    .B1(_00041_),
    .X(_01032_));
 sg13g2_nand3b_1 _06273_ (.B(net2514),
    .C(net2509),
    .Y(_01033_),
    .A_N(_00042_));
 sg13g2_nand2_1 _06274_ (.Y(_01034_),
    .A(_01032_),
    .B(_01033_));
 sg13g2_a21oi_1 _06275_ (.A1(net2521),
    .A2(net2519),
    .Y(_01035_),
    .B1(_00914_));
 sg13g2_a21oi_2 _06276_ (.B1(_01035_),
    .Y(_01036_),
    .A2(net2453),
    .A1(_00042_));
 sg13g2_a21o_2 _06277_ (.A2(net2453),
    .A1(_00042_),
    .B1(_01035_),
    .X(_01037_));
 sg13g2_a21o_1 _06278_ (.A2(net2511),
    .A1(net2516),
    .B1(_00028_),
    .X(_01038_));
 sg13g2_nand3b_1 _06279_ (.B(net2516),
    .C(net2511),
    .Y(_01039_),
    .A_N(_00029_));
 sg13g2_nand2_2 _06280_ (.Y(_01040_),
    .A(_01038_),
    .B(_01039_));
 sg13g2_nand3_1 _06281_ (.B(net2520),
    .C(net2518),
    .A(_00029_),
    .Y(_01041_));
 sg13g2_o21ai_1 _06282_ (.B1(_00030_),
    .Y(_01042_),
    .A1(_00990_),
    .A2(_00995_));
 sg13g2_nand2_1 _06283_ (.Y(_01043_),
    .A(_01041_),
    .B(_01042_));
 sg13g2_nand4_1 _06284_ (.B(_01039_),
    .C(_01041_),
    .A(_01038_),
    .Y(_01044_),
    .D(_01042_));
 sg13g2_nand3_1 _06285_ (.B(net2520),
    .C(net2518),
    .A(_00017_),
    .Y(_01045_));
 sg13g2_o21ai_1 _06286_ (.B1(_00018_),
    .Y(_01046_),
    .A1(_00990_),
    .A2(_00995_));
 sg13g2_nand2_2 _06287_ (.Y(_01047_),
    .A(_01045_),
    .B(_01046_));
 sg13g2_inv_2 _06288_ (.Y(_01048_),
    .A(_01047_));
 sg13g2_a21o_1 _06289_ (.A2(net2511),
    .A1(net2516),
    .B1(_00016_),
    .X(_01049_));
 sg13g2_nand3b_1 _06290_ (.B(net2516),
    .C(net2511),
    .Y(_01050_),
    .A_N(_00017_));
 sg13g2_nand2_2 _06291_ (.Y(_01051_),
    .A(_01049_),
    .B(_01050_));
 sg13g2_nand4_1 _06292_ (.B(_01046_),
    .C(_01049_),
    .A(_01045_),
    .Y(_01052_),
    .D(_01050_));
 sg13g2_a21oi_2 _06293_ (.B1(_00922_),
    .Y(_01053_),
    .A2(net2518),
    .A1(net2520));
 sg13g2_a21oi_2 _06294_ (.B1(_01053_),
    .Y(_01054_),
    .A2(net2457),
    .A1(\ChiselTop.wild.cpu.exFwdReg_wbData[31] ));
 sg13g2_a21o_1 _06295_ (.A2(net2456),
    .A1(\ChiselTop.wild.cpu.exFwdReg_wbData[31] ),
    .B1(_01053_),
    .X(_01055_));
 sg13g2_mux2_2 _06296_ (.A0(_00094_),
    .A1(_00093_),
    .S(net2451),
    .X(_01056_));
 sg13g2_a21oi_1 _06297_ (.A1(net2521),
    .A2(net2519),
    .Y(_01057_),
    .B1(_00916_));
 sg13g2_a21oi_2 _06298_ (.B1(_01057_),
    .Y(_01058_),
    .A2(net2454),
    .A1(_00067_));
 sg13g2_a21o_1 _06299_ (.A2(net2454),
    .A1(_00067_),
    .B1(_01057_),
    .X(_01059_));
 sg13g2_mux2_1 _06300_ (.A0(_00067_),
    .A1(_00109_),
    .S(net2451),
    .X(_01060_));
 sg13g2_nand3_1 _06301_ (.B(net2520),
    .C(net2518),
    .A(_00081_),
    .Y(_01061_));
 sg13g2_o21ai_1 _06302_ (.B1(_00082_),
    .Y(_01062_),
    .A1(_00990_),
    .A2(_00995_));
 sg13g2_and2_1 _06303_ (.A(_01061_),
    .B(_01062_),
    .X(_01063_));
 sg13g2_nand2_2 _06304_ (.Y(_01064_),
    .A(_01061_),
    .B(_01062_));
 sg13g2_and3_1 _06305_ (.X(_01065_),
    .A(_00081_),
    .B(net2516),
    .C(net2511));
 sg13g2_a21oi_2 _06306_ (.B1(_01065_),
    .Y(_01066_),
    .A2(net2450),
    .A1(_00102_));
 sg13g2_a21o_1 _06307_ (.A2(net2450),
    .A1(_00102_),
    .B1(_01065_),
    .X(_01067_));
 sg13g2_mux2_1 _06308_ (.A0(_00022_),
    .A1(_00021_),
    .S(net2452),
    .X(_01068_));
 sg13g2_and3_1 _06309_ (.X(_01069_),
    .A(_00021_),
    .B(net2514),
    .C(net2509));
 sg13g2_a21oi_2 _06310_ (.B1(_01069_),
    .Y(_01070_),
    .A2(net2449),
    .A1(_00020_));
 sg13g2_mux2_2 _06311_ (.A0(_00061_),
    .A1(_00060_),
    .S(net2454),
    .X(_01071_));
 sg13g2_nand3_1 _06312_ (.B(net2515),
    .C(net2510),
    .A(_00060_),
    .Y(_01072_));
 sg13g2_o21ai_1 _06313_ (.B1(_00059_),
    .Y(_01073_),
    .A1(net2513),
    .A2(net2508));
 sg13g2_nand2_1 _06314_ (.Y(_01074_),
    .A(_01072_),
    .B(_01073_));
 sg13g2_nand2b_1 _06315_ (.Y(_01075_),
    .B(net2427),
    .A_N(_01074_));
 sg13g2_nand3_1 _06316_ (.B(net2520),
    .C(net2518),
    .A(_00048_),
    .Y(_01076_));
 sg13g2_o21ai_1 _06317_ (.B1(_00049_),
    .Y(_01077_),
    .A1(_00990_),
    .A2(_00995_));
 sg13g2_nand2_2 _06318_ (.Y(_01078_),
    .A(_01076_),
    .B(_01077_));
 sg13g2_nand3_1 _06319_ (.B(net2516),
    .C(net2511),
    .A(\ChiselTop.wild.cpu.exFwdReg_wbData[4] ),
    .Y(_01079_));
 sg13g2_o21ai_1 _06320_ (.B1(\ChiselTop.wild.cpu.decExReg_rs2Val[4] ),
    .Y(_01080_),
    .A1(_01005_),
    .A2(_01008_));
 sg13g2_nand2_1 _06321_ (.Y(_01081_),
    .A(_01079_),
    .B(_01080_));
 sg13g2_mux2_2 _06322_ (.A0(_00072_),
    .A1(_00071_),
    .S(net2457),
    .X(_01082_));
 sg13g2_mux2_2 _06323_ (.A0(_00071_),
    .A1(_00107_),
    .S(net2450),
    .X(_01083_));
 sg13g2_xnor2_1 _06324_ (.Y(_01084_),
    .A(_01082_),
    .B(_01083_));
 sg13g2_mux2_1 _06325_ (.A0(_00080_),
    .A1(_00079_),
    .S(net2452),
    .X(_01085_));
 sg13g2_and3_1 _06326_ (.X(_01086_),
    .A(_00079_),
    .B(net2514),
    .C(net2509));
 sg13g2_a21oi_2 _06327_ (.B1(_01086_),
    .Y(_01087_),
    .A2(net2449),
    .A1(_00103_));
 sg13g2_mux2_1 _06328_ (.A0(_00006_),
    .A1(_00005_),
    .S(net2457),
    .X(_01088_));
 sg13g2_mux2_1 _06329_ (.A0(\ChiselTop.wild.cpu.exFwdReg_wbData[16] ),
    .A1(\ChiselTop.wild.cpu.decExReg_rs2Val[16] ),
    .S(net2451),
    .X(_01089_));
 sg13g2_xnor2_1 _06330_ (.Y(_01090_),
    .A(net2423),
    .B(_01089_));
 sg13g2_nor2b_1 _06331_ (.A(net2452),
    .B_N(_00026_),
    .Y(_01091_));
 sg13g2_a21oi_2 _06332_ (.B1(_01091_),
    .Y(_01092_),
    .A2(net2453),
    .A1(_00025_));
 sg13g2_mux2_2 _06333_ (.A0(_00026_),
    .A1(_00025_),
    .S(net2452),
    .X(_01093_));
 sg13g2_mux2_2 _06334_ (.A0(_00025_),
    .A1(_00024_),
    .S(net2449),
    .X(_01094_));
 sg13g2_xnor2_1 _06335_ (.Y(_01095_),
    .A(_01093_),
    .B(_01094_));
 sg13g2_mux2_2 _06336_ (.A0(_00065_),
    .A1(_00064_),
    .S(net2454),
    .X(_01096_));
 sg13g2_nand3_1 _06337_ (.B(net2515),
    .C(net2510),
    .A(_00064_),
    .Y(_01097_));
 sg13g2_o21ai_1 _06338_ (.B1(_00063_),
    .Y(_01098_),
    .A1(net2513),
    .A2(net2508));
 sg13g2_nand2_1 _06339_ (.Y(_01099_),
    .A(_01097_),
    .B(_01098_));
 sg13g2_nand2b_1 _06340_ (.Y(_01100_),
    .B(_01099_),
    .A_N(_01096_));
 sg13g2_mux2_2 _06341_ (.A0(_00013_),
    .A1(_00012_),
    .S(net2450),
    .X(_01101_));
 sg13g2_a21oi_1 _06342_ (.A1(net2521),
    .A2(net2519),
    .Y(_01102_),
    .B1(_00910_));
 sg13g2_a21oi_2 _06343_ (.B1(_01102_),
    .Y(_01103_),
    .A2(net2455),
    .A1(_00013_));
 sg13g2_a21o_2 _06344_ (.A2(net2455),
    .A1(_00013_),
    .B1(_01102_),
    .X(_01104_));
 sg13g2_mux2_2 _06345_ (.A0(_00078_),
    .A1(_00077_),
    .S(net2453),
    .X(_01105_));
 sg13g2_mux2_2 _06346_ (.A0(_00077_),
    .A1(_00104_),
    .S(net2449),
    .X(_01106_));
 sg13g2_mux2_2 _06347_ (.A0(_00032_),
    .A1(_00031_),
    .S(net2449),
    .X(_01107_));
 sg13g2_mux2_2 _06348_ (.A0(_00033_),
    .A1(_00032_),
    .S(net2452),
    .X(_01108_));
 sg13g2_inv_1 _06349_ (.Y(_01109_),
    .A(net2420));
 sg13g2_xnor2_1 _06350_ (.Y(_01110_),
    .A(_01107_),
    .B(net2420));
 sg13g2_a21oi_2 _06351_ (.B1(_00918_),
    .Y(_01111_),
    .A2(net2519),
    .A1(net2521));
 sg13g2_a21oi_2 _06352_ (.B1(_01111_),
    .Y(_01112_),
    .A2(net2456),
    .A1(_00083_));
 sg13g2_a21o_2 _06353_ (.A2(net2454),
    .A1(_00083_),
    .B1(_01111_),
    .X(_01113_));
 sg13g2_a21oi_2 _06354_ (.B1(_00101_),
    .Y(_01114_),
    .A2(net2510),
    .A1(net2515));
 sg13g2_nor3_2 _06355_ (.A(_00083_),
    .B(net2513),
    .C(net2508),
    .Y(_01115_));
 sg13g2_or2_1 _06356_ (.X(_01116_),
    .B(_01115_),
    .A(_01114_));
 sg13g2_nor2_1 _06357_ (.A(_01114_),
    .B(_01115_),
    .Y(_01117_));
 sg13g2_a21oi_2 _06358_ (.B1(_00915_),
    .Y(_01118_),
    .A2(net2519),
    .A1(net2521));
 sg13g2_a21oi_2 _06359_ (.B1(_01118_),
    .Y(_01119_),
    .A2(net2455),
    .A1(_00052_));
 sg13g2_a21o_2 _06360_ (.A2(net2454),
    .A1(_00052_),
    .B1(_01118_),
    .X(_01120_));
 sg13g2_a21oi_2 _06361_ (.B1(_00051_),
    .Y(_01121_),
    .A2(net2509),
    .A1(net2515));
 sg13g2_nor3_1 _06362_ (.A(_00052_),
    .B(net2513),
    .C(net2508),
    .Y(_01122_));
 sg13g2_nor2_1 _06363_ (.A(_01121_),
    .B(_01122_),
    .Y(_01123_));
 sg13g2_xnor2_1 _06364_ (.Y(_01124_),
    .A(_01120_),
    .B(_01123_));
 sg13g2_mux2_2 _06365_ (.A0(_00090_),
    .A1(_00089_),
    .S(net2452),
    .X(_01125_));
 sg13g2_inv_2 _06366_ (.Y(_01126_),
    .A(_01125_));
 sg13g2_mux2_2 _06367_ (.A0(_00089_),
    .A1(_00098_),
    .S(net2449),
    .X(_01127_));
 sg13g2_xnor2_1 _06368_ (.Y(_01128_),
    .A(net2419),
    .B(_01127_));
 sg13g2_a21oi_2 _06369_ (.B1(_00909_),
    .Y(_01129_),
    .A2(_00994_),
    .A1(_00989_));
 sg13g2_a21oi_2 _06370_ (.B1(_01129_),
    .Y(_01130_),
    .A2(net2456),
    .A1(_00009_));
 sg13g2_a21o_2 _06371_ (.A2(net2456),
    .A1(_00009_),
    .B1(_01129_),
    .X(_01131_));
 sg13g2_mux2_2 _06372_ (.A0(_00009_),
    .A1(_00008_),
    .S(net2451),
    .X(_01132_));
 sg13g2_nor2_1 _06373_ (.A(_01130_),
    .B(_01132_),
    .Y(_01133_));
 sg13g2_mux2_1 _06374_ (.A0(_00076_),
    .A1(_00075_),
    .S(net2452),
    .X(_01134_));
 sg13g2_and3_1 _06375_ (.X(_01135_),
    .A(_00075_),
    .B(net2514),
    .C(net2509));
 sg13g2_a21oi_2 _06376_ (.B1(_01135_),
    .Y(_01136_),
    .A2(net2449),
    .A1(_00105_));
 sg13g2_nor2_1 _06377_ (.A(net2429),
    .B(_01070_),
    .Y(_01137_));
 sg13g2_nor2_1 _06378_ (.A(net2437),
    .B(_01017_),
    .Y(_01138_));
 sg13g2_a21oi_2 _06379_ (.B1(_00920_),
    .Y(_01139_),
    .A2(_00994_),
    .A1(_00989_));
 sg13g2_a21oi_2 _06380_ (.B1(_01139_),
    .Y(_01140_),
    .A2(net2456),
    .A1(_00087_));
 sg13g2_a21o_2 _06381_ (.A2(net2456),
    .A1(_00087_),
    .B1(_01139_),
    .X(_01141_));
 sg13g2_a21oi_2 _06382_ (.B1(_00099_),
    .Y(_01142_),
    .A2(net2511),
    .A1(net2516));
 sg13g2_nor3_2 _06383_ (.A(_00087_),
    .B(_01005_),
    .C(_01008_),
    .Y(_01143_));
 sg13g2_nor2_2 _06384_ (.A(_01142_),
    .B(_01143_),
    .Y(_01144_));
 sg13g2_nand2_1 _06385_ (.Y(_01145_),
    .A(_01140_),
    .B(_01144_));
 sg13g2_and2_1 _06386_ (.A(_01047_),
    .B(_01051_),
    .X(_01146_));
 sg13g2_nor2_1 _06387_ (.A(net2417),
    .B(_01136_),
    .Y(_01147_));
 sg13g2_nor2b_1 _06388_ (.A(net2427),
    .B_N(_01074_),
    .Y(_01148_));
 sg13g2_nor2_1 _06389_ (.A(_01101_),
    .B(_01103_),
    .Y(_01149_));
 sg13g2_nand3_1 _06390_ (.B(net2520),
    .C(net2518),
    .A(_00091_),
    .Y(_01150_));
 sg13g2_o21ai_1 _06391_ (.B1(_00092_),
    .Y(_01151_),
    .A1(_00990_),
    .A2(_00995_));
 sg13g2_nand2_1 _06392_ (.Y(_01152_),
    .A(_01150_),
    .B(_01151_));
 sg13g2_inv_2 _06393_ (.Y(_01153_),
    .A(_01152_));
 sg13g2_a21o_1 _06394_ (.A2(net2511),
    .A1(net2516),
    .B1(_00097_),
    .X(_01154_));
 sg13g2_nand3b_1 _06395_ (.B(net2517),
    .C(net2512),
    .Y(_01155_),
    .A_N(_00091_));
 sg13g2_nand2_2 _06396_ (.Y(_01156_),
    .A(_01154_),
    .B(_01155_));
 sg13g2_nand4_1 _06397_ (.B(_01151_),
    .C(_01154_),
    .A(_01150_),
    .Y(_01157_),
    .D(_01155_));
 sg13g2_a21oi_1 _06398_ (.A1(net2521),
    .A2(net2519),
    .Y(_01158_),
    .B1(_00917_));
 sg13g2_a21oi_2 _06399_ (.B1(_01158_),
    .Y(_01159_),
    .A2(net2458),
    .A1(_00069_));
 sg13g2_a21o_1 _06400_ (.A2(net2453),
    .A1(_00069_),
    .B1(_01158_),
    .X(_01160_));
 sg13g2_a21oi_1 _06401_ (.A1(net2514),
    .A2(net2510),
    .Y(_01161_),
    .B1(_00108_));
 sg13g2_nor3_2 _06402_ (.A(_00069_),
    .B(net2513),
    .C(net2508),
    .Y(_01162_));
 sg13g2_or2_1 _06403_ (.X(_01163_),
    .B(_01162_),
    .A(_01161_));
 sg13g2_nor2_1 _06404_ (.A(net2415),
    .B(_01163_),
    .Y(_01164_));
 sg13g2_nand2b_1 _06405_ (.Y(_01165_),
    .B(_01096_),
    .A_N(_01099_));
 sg13g2_a21oi_1 _06406_ (.A1(net2520),
    .A2(net2518),
    .Y(_01166_),
    .B1(_00921_));
 sg13g2_a21oi_2 _06407_ (.B1(_01166_),
    .Y(_01167_),
    .A2(net2457),
    .A1(\ChiselTop.wild.cpu.exFwdReg_wbData[30] ));
 sg13g2_mux2_2 _06408_ (.A0(_00096_),
    .A1(_00095_),
    .S(net2450),
    .X(_01168_));
 sg13g2_mux2_2 _06409_ (.A0(_00035_),
    .A1(_00034_),
    .S(net2450),
    .X(_01169_));
 sg13g2_a21oi_1 _06410_ (.A1(net2521),
    .A2(net2519),
    .Y(_01170_),
    .B1(_00912_));
 sg13g2_a21oi_2 _06411_ (.B1(_01170_),
    .Y(_01171_),
    .A2(net2453),
    .A1(_00035_));
 sg13g2_a21o_2 _06412_ (.A2(net2453),
    .A1(_00035_),
    .B1(_01170_),
    .X(_01172_));
 sg13g2_nor2_1 _06413_ (.A(_01169_),
    .B(_01171_),
    .Y(_01173_));
 sg13g2_nand4_1 _06414_ (.B(_01077_),
    .C(_01079_),
    .A(_01076_),
    .Y(_01174_),
    .D(_01080_));
 sg13g2_nor2_1 _06415_ (.A(\ChiselTop.wild.cpu.decExReg_func3[0] ),
    .B(net2611),
    .Y(_01175_));
 sg13g2_or2_2 _06416_ (.X(_01176_),
    .B(net2611),
    .A(\ChiselTop.wild.cpu.decExReg_func3[0] ));
 sg13g2_nor2b_2 _06417_ (.A(net2611),
    .B_N(net2612),
    .Y(_01177_));
 sg13g2_nand2b_2 _06418_ (.Y(_01178_),
    .B(net2612),
    .A_N(net2611));
 sg13g2_o21ai_1 _06419_ (.B1(_01145_),
    .Y(_01179_),
    .A1(_01058_),
    .A2(_01060_));
 sg13g2_or4_1 _06420_ (.A(_01137_),
    .B(_01146_),
    .C(_01147_),
    .D(_01164_),
    .X(_01180_));
 sg13g2_xnor2_1 _06421_ (.Y(_01181_),
    .A(_01034_),
    .B(_01036_));
 sg13g2_xnor2_1 _06422_ (.Y(_01182_),
    .A(_01024_),
    .B(_01026_));
 sg13g2_nand4_1 _06423_ (.B(_01110_),
    .C(_01181_),
    .A(_01084_),
    .Y(_01183_),
    .D(_01182_));
 sg13g2_nor4_1 _06424_ (.A(_01090_),
    .B(_01179_),
    .C(_01180_),
    .D(_01183_),
    .Y(_01184_));
 sg13g2_a21oi_1 _06425_ (.A1(_01040_),
    .A2(net2434),
    .Y(_01185_),
    .B1(_01149_));
 sg13g2_nor4_1 _06426_ (.A(_01133_),
    .B(_01138_),
    .C(_01148_),
    .D(_01173_),
    .Y(_01186_));
 sg13g2_and3_1 _06427_ (.X(_01187_),
    .A(_01124_),
    .B(_01185_),
    .C(_01186_));
 sg13g2_o21ai_1 _06428_ (.B1(_01165_),
    .Y(_01188_),
    .A1(net2432),
    .A2(_01056_));
 sg13g2_xor2_1 _06429_ (.B(_01031_),
    .A(net2435),
    .X(_01189_));
 sg13g2_o21ai_1 _06430_ (.B1(_01100_),
    .Y(_01190_),
    .A1(net2425),
    .A2(_01087_));
 sg13g2_nand4_1 _06431_ (.B(_01052_),
    .C(_01157_),
    .A(_01044_),
    .Y(_01191_),
    .D(_01174_));
 sg13g2_a22oi_1 _06432_ (.Y(_01192_),
    .B1(net2424),
    .B2(_01087_),
    .A2(_01081_),
    .A1(_01078_));
 sg13g2_xnor2_1 _06433_ (.Y(_01193_),
    .A(_01167_),
    .B(_01168_));
 sg13g2_nand3b_1 _06434_ (.B(_01192_),
    .C(_01193_),
    .Y(_01194_),
    .A_N(_01191_));
 sg13g2_xnor2_1 _06435_ (.Y(_01195_),
    .A(_01105_),
    .B(_01106_));
 sg13g2_xnor2_1 _06436_ (.Y(_01196_),
    .A(_01020_),
    .B(net2436));
 sg13g2_a22oi_1 _06437_ (.Y(_01197_),
    .B1(_01160_),
    .B2(_01163_),
    .A2(_01056_),
    .A1(net2432));
 sg13g2_a22oi_1 _06438_ (.Y(_01198_),
    .B1(_01130_),
    .B2(_01132_),
    .A2(_01067_),
    .A1(_01063_));
 sg13g2_nand4_1 _06439_ (.B(_01095_),
    .C(_01197_),
    .A(_01013_),
    .Y(_01199_),
    .D(_01198_));
 sg13g2_a22oi_1 _06440_ (.Y(_01200_),
    .B1(_01064_),
    .B2(_01066_),
    .A2(_01017_),
    .A1(net2437));
 sg13g2_a22oi_1 _06441_ (.Y(_01201_),
    .B1(_01112_),
    .B2(_01117_),
    .A2(_01070_),
    .A1(net2429));
 sg13g2_a22oi_1 _06442_ (.Y(_01202_),
    .B1(_01169_),
    .B2(_01171_),
    .A2(_01156_),
    .A1(net2416));
 sg13g2_o21ai_1 _06443_ (.B1(_01075_),
    .Y(_01203_),
    .A1(_01140_),
    .A2(_01144_));
 sg13g2_nor4_1 _06444_ (.A(_01188_),
    .B(_01189_),
    .C(_01190_),
    .D(_01203_),
    .Y(_01204_));
 sg13g2_a22oi_1 _06445_ (.Y(_01205_),
    .B1(_01113_),
    .B2(_01116_),
    .A2(_01103_),
    .A1(_01101_));
 sg13g2_nand4_1 _06446_ (.B(_01200_),
    .C(_01202_),
    .A(_01128_),
    .Y(_01206_),
    .D(_01205_));
 sg13g2_a22oi_1 _06447_ (.Y(_01207_),
    .B1(net2417),
    .B2(_01136_),
    .A2(_01060_),
    .A1(_01058_));
 sg13g2_nand4_1 _06448_ (.B(_01196_),
    .C(_01201_),
    .A(_01195_),
    .Y(_01208_),
    .D(_01207_));
 sg13g2_nor4_1 _06449_ (.A(_01194_),
    .B(_01199_),
    .C(_01206_),
    .D(_01208_),
    .Y(_01209_));
 sg13g2_nand4_1 _06450_ (.B(_01187_),
    .C(_01204_),
    .A(_01184_),
    .Y(_01210_),
    .D(_01209_));
 sg13g2_and2_1 _06451_ (.A(_01178_),
    .B(_01210_),
    .X(_01211_));
 sg13g2_o21ai_1 _06452_ (.B1(\ChiselTop.wild.cpu.decExReg_decOut_isBranch ),
    .Y(_01212_),
    .A1(net2526),
    .A2(_01210_));
 sg13g2_o21ai_1 _06453_ (.B1(_00002_),
    .Y(_01213_),
    .A1(_01211_),
    .A2(_01212_));
 sg13g2_nand2_1 _06454_ (.Y(_01214_),
    .A(\ChiselTop.wild.cpu.decExReg_valid ),
    .B(_01213_));
 sg13g2_and2_1 _06455_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_isLoad ),
    .B(net2192),
    .X(_01215_));
 sg13g2_nor3_1 _06456_ (.A(\ChiselTop.wild.memAddressReg[1] ),
    .B(\ChiselTop.wild.memAddressReg[0] ),
    .C(\ChiselTop.wild.memAddressReg[3] ),
    .Y(_01216_));
 sg13g2_nor4_1 _06457_ (.A(\ChiselTop.wild.memAddressReg[17] ),
    .B(\ChiselTop.wild.memAddressReg[16] ),
    .C(\ChiselTop.wild.memAddressReg[19] ),
    .D(\ChiselTop.wild.memAddressReg[18] ),
    .Y(_01217_));
 sg13g2_and4_1 _06458_ (.A(\ChiselTop.wild.memAddressReg[28] ),
    .B(\ChiselTop.wild.memAddressReg[29] ),
    .C(\ChiselTop.wild.memAddressReg[30] ),
    .D(\ChiselTop.wild.memAddressReg[31] ),
    .X(_01218_));
 sg13g2_nand3_1 _06459_ (.B(_01217_),
    .C(_01218_),
    .A(_01216_),
    .Y(_01219_));
 sg13g2_nand2_1 _06460_ (.Y(_01220_),
    .A(\ChiselTop.wild.dmem.MEM_2[0][0] ),
    .B(net2500));
 sg13g2_nor2_1 _06461_ (.A(net2611),
    .B(net2621),
    .Y(_01221_));
 sg13g2_or2_1 _06462_ (.X(_01222_),
    .B(\ChiselTop.wild.cpu.decExReg_memLow[0] ),
    .A(\ChiselTop.wild.cpu.decExReg_func3[1] ));
 sg13g2_nor2_1 _06463_ (.A(net2525),
    .B(_01221_),
    .Y(_01223_));
 sg13g2_nand2_2 _06464_ (.Y(_01224_),
    .A(_01176_),
    .B(_01222_));
 sg13g2_nor2_2 _06465_ (.A(net2621),
    .B(\ChiselTop.wild.cpu.decExReg_memLow[1] ),
    .Y(_01225_));
 sg13g2_nor2_1 _06466_ (.A(_00926_),
    .B(net2506),
    .Y(_01226_));
 sg13g2_a22oi_1 _06467_ (.Y(_01227_),
    .B1(net2448),
    .B2(\ChiselTop.wild.rx._shiftReg_T_1[6] ),
    .A2(net2506),
    .A1(\ChiselTop.wild.dmem.MEM[0][7] ));
 sg13g2_nand2_1 _06468_ (.Y(_01228_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][7] ),
    .B(net2502));
 sg13g2_nor2b_2 _06469_ (.A(\ChiselTop.wild.cpu.decExReg_memLow[1] ),
    .B_N(net2621),
    .Y(_01229_));
 sg13g2_nand2_2 _06470_ (.Y(_01230_),
    .A(\ChiselTop.wild.dmem.MEM_3[0][7] ),
    .B(net2505));
 sg13g2_and2_1 _06471_ (.A(net2621),
    .B(\ChiselTop.wild.cpu.decExReg_memLow[1] ),
    .X(_01231_));
 sg13g2_nand2_1 _06472_ (.Y(_01232_),
    .A(net2621),
    .B(\ChiselTop.wild.cpu.decExReg_memLow[1] ));
 sg13g2_nor2b_2 _06473_ (.A(net2621),
    .B_N(\ChiselTop.wild.cpu.decExReg_memLow[1] ),
    .Y(_01233_));
 sg13g2_nand2b_2 _06474_ (.Y(_01234_),
    .B(\ChiselTop.wild.cpu.decExReg_memLow[1] ),
    .A_N(net2621));
 sg13g2_a21oi_1 _06475_ (.A1(\ChiselTop.wild.dmem.MEM_2[0][7] ),
    .A2(net2501),
    .Y(_01235_),
    .B1(_01234_));
 sg13g2_a21o_1 _06476_ (.A2(_01231_),
    .A1(_01230_),
    .B1(_01235_),
    .X(_01236_));
 sg13g2_a221oi_1 _06477_ (.B2(_01229_),
    .C1(_01236_),
    .B1(_01228_),
    .A1(_01225_),
    .Y(_01237_),
    .A2(_01227_));
 sg13g2_and2_1 _06478_ (.A(net2525),
    .B(_01237_),
    .X(_01238_));
 sg13g2_nand2_1 _06479_ (.Y(_01239_),
    .A(net2525),
    .B(_01237_));
 sg13g2_a22oi_1 _06480_ (.Y(_01240_),
    .B1(_01230_),
    .B2(_01233_),
    .A2(_01228_),
    .A1(_01225_));
 sg13g2_nor2_1 _06481_ (.A(net2621),
    .B(_01178_),
    .Y(_01241_));
 sg13g2_a21oi_2 _06482_ (.B1(_01238_),
    .Y(_01242_),
    .A2(_01241_),
    .A1(_01240_));
 sg13g2_o21ai_1 _06483_ (.B1(_01242_),
    .Y(_01243_),
    .A1(_01220_),
    .A2(_01224_));
 sg13g2_mux2_2 _06484_ (.A0(\ChiselTop.wild.cpu.decExReg_decOut_imm[16] ),
    .A1(_01089_),
    .S(net2533),
    .X(_01244_));
 sg13g2_nor2_1 _06485_ (.A(net2423),
    .B(_01244_),
    .Y(_01245_));
 sg13g2_xor2_1 _06486_ (.B(_01244_),
    .A(net2423),
    .X(_01246_));
 sg13g2_xnor2_1 _06487_ (.Y(_01247_),
    .A(net2422),
    .B(_01244_));
 sg13g2_nand2_1 _06488_ (.Y(_01248_),
    .A(net2645),
    .B(_00015_));
 sg13g2_o21ai_1 _06489_ (.B1(_01248_),
    .Y(_01249_),
    .A1(net2646),
    .A2(_01051_));
 sg13g2_nor2_1 _06490_ (.A(_01048_),
    .B(_01249_),
    .Y(_01250_));
 sg13g2_nand2_1 _06491_ (.Y(_01251_),
    .A(_01048_),
    .B(_01249_));
 sg13g2_xnor2_1 _06492_ (.Y(_01252_),
    .A(_01048_),
    .B(_01249_));
 sg13g2_and2_2 _06493_ (.A(net2641),
    .B(_00011_),
    .X(_01253_));
 sg13g2_a21o_2 _06494_ (.A2(_01101_),
    .A1(net2532),
    .B1(_01253_),
    .X(_01254_));
 sg13g2_and2_1 _06495_ (.A(_01103_),
    .B(_01254_),
    .X(_01255_));
 sg13g2_nor2_1 _06496_ (.A(_01103_),
    .B(_01254_),
    .Y(_01256_));
 sg13g2_xnor2_1 _06497_ (.Y(_01257_),
    .A(_01104_),
    .B(_01254_));
 sg13g2_mux2_2 _06498_ (.A0(_00007_),
    .A1(_01132_),
    .S(net2535),
    .X(_01258_));
 sg13g2_inv_1 _06499_ (.Y(_01259_),
    .A(_01258_));
 sg13g2_nor2_1 _06500_ (.A(_01130_),
    .B(_01258_),
    .Y(_01260_));
 sg13g2_nand2_1 _06501_ (.Y(_01261_),
    .A(_01130_),
    .B(_01258_));
 sg13g2_xnor2_1 _06502_ (.Y(_01262_),
    .A(_01131_),
    .B(_01258_));
 sg13g2_nand2b_2 _06503_ (.Y(_01263_),
    .B(_01261_),
    .A_N(_01260_));
 sg13g2_nor2_1 _06504_ (.A(_01257_),
    .B(_01262_),
    .Y(_01264_));
 sg13g2_nor2_1 _06505_ (.A(_01104_),
    .B(_01254_),
    .Y(_01265_));
 sg13g2_nand2b_1 _06506_ (.Y(_01266_),
    .B(_01048_),
    .A_N(_01249_));
 sg13g2_nand2_1 _06507_ (.Y(_01267_),
    .A(net2646),
    .B(_00019_));
 sg13g2_o21ai_1 _06508_ (.B1(_01267_),
    .Y(_01268_),
    .A1(net2645),
    .A2(_01070_));
 sg13g2_nand2b_1 _06509_ (.Y(_01269_),
    .B(_01268_),
    .A_N(net2428));
 sg13g2_nor2b_1 _06510_ (.A(_01268_),
    .B_N(net2428),
    .Y(_01270_));
 sg13g2_xnor2_1 _06511_ (.Y(_01271_),
    .A(net2428),
    .B(_01268_));
 sg13g2_xor2_1 _06512_ (.B(_01268_),
    .A(net2428),
    .X(_01272_));
 sg13g2_mux2_1 _06513_ (.A0(_00023_),
    .A1(_01094_),
    .S(net2534),
    .X(_01273_));
 sg13g2_nor2_1 _06514_ (.A(_01093_),
    .B(_01273_),
    .Y(_01274_));
 sg13g2_and2_1 _06515_ (.A(_01092_),
    .B(_01273_),
    .X(_01275_));
 sg13g2_or2_1 _06516_ (.X(_01276_),
    .B(_01273_),
    .A(_01092_));
 sg13g2_xnor2_1 _06517_ (.Y(_01277_),
    .A(_01092_),
    .B(_01273_));
 sg13g2_and2_1 _06518_ (.A(net2645),
    .B(_00027_),
    .X(_01278_));
 sg13g2_nand2_1 _06519_ (.Y(_01279_),
    .A(net2646),
    .B(_00027_));
 sg13g2_o21ai_1 _06520_ (.B1(_01279_),
    .Y(_01280_),
    .A1(net2645),
    .A2(_01040_));
 sg13g2_nor2_1 _06521_ (.A(net2434),
    .B(_01280_),
    .Y(_01281_));
 sg13g2_a21oi_2 _06522_ (.B1(_01274_),
    .Y(_01282_),
    .A2(_01281_),
    .A1(net2321));
 sg13g2_nand2b_1 _06523_ (.Y(_01283_),
    .B(_01280_),
    .A_N(net2433));
 sg13g2_nand2b_1 _06524_ (.Y(_01284_),
    .B(net2433),
    .A_N(_01280_));
 sg13g2_xnor2_1 _06525_ (.Y(_01285_),
    .A(net2433),
    .B(_01280_));
 sg13g2_xor2_1 _06526_ (.B(_01280_),
    .A(net2433),
    .X(_01286_));
 sg13g2_nand2_1 _06527_ (.Y(_01287_),
    .A(net2321),
    .B(_01286_));
 sg13g2_a21oi_2 _06528_ (.B1(_01278_),
    .Y(_01288_),
    .A2(_01107_),
    .A1(net2534));
 sg13g2_nor2_2 _06529_ (.A(net2420),
    .B(_01288_),
    .Y(_01289_));
 sg13g2_nand2_1 _06530_ (.Y(_01290_),
    .A(net2420),
    .B(_01288_));
 sg13g2_nor2b_2 _06531_ (.A(_01289_),
    .B_N(_01290_),
    .Y(_01291_));
 sg13g2_a21o_1 _06532_ (.A2(_01169_),
    .A1(net2534),
    .B1(_01278_),
    .X(_01292_));
 sg13g2_and2_1 _06533_ (.A(_01171_),
    .B(_01292_),
    .X(_01293_));
 sg13g2_nand2b_1 _06534_ (.Y(_01294_),
    .B(_01172_),
    .A_N(_01292_));
 sg13g2_xnor2_1 _06535_ (.Y(_01295_),
    .A(_01172_),
    .B(_01292_));
 sg13g2_nand2b_1 _06536_ (.Y(_01296_),
    .B(_01294_),
    .A_N(_01293_));
 sg13g2_nand2_2 _06537_ (.Y(_01297_),
    .A(net2645),
    .B(_00037_));
 sg13g2_or3_2 _06538_ (.A(net2641),
    .B(_01018_),
    .C(_01019_),
    .X(_01298_));
 sg13g2_and3_1 _06539_ (.X(_01299_),
    .A(_01022_),
    .B(_01297_),
    .C(_01298_));
 sg13g2_and3_1 _06540_ (.X(_01300_),
    .A(net2436),
    .B(_01297_),
    .C(_01298_));
 sg13g2_a21oi_1 _06541_ (.A1(_01297_),
    .A2(_01298_),
    .Y(_01301_),
    .B1(net2436));
 sg13g2_nor2_2 _06542_ (.A(_01300_),
    .B(_01301_),
    .Y(_01302_));
 sg13g2_nand3_1 _06543_ (.B(_01032_),
    .C(_01033_),
    .A(net2532),
    .Y(_01303_));
 sg13g2_nand3_1 _06544_ (.B(_01297_),
    .C(_01303_),
    .A(_01036_),
    .Y(_01304_));
 sg13g2_and3_1 _06545_ (.X(_01305_),
    .A(_01037_),
    .B(_01297_),
    .C(_01303_));
 sg13g2_a21oi_1 _06546_ (.A1(_01297_),
    .A2(_01303_),
    .Y(_01306_),
    .B1(_01037_));
 sg13g2_or2_2 _06547_ (.X(_01307_),
    .B(_01306_),
    .A(_01305_));
 sg13g2_and3_2 _06548_ (.X(_01308_),
    .A(net2533),
    .B(_01029_),
    .C(_01030_));
 sg13g2_nor2_1 _06549_ (.A(net2534),
    .B(_00044_),
    .Y(_01309_));
 sg13g2_nor2_1 _06550_ (.A(_01308_),
    .B(_01309_),
    .Y(_01310_));
 sg13g2_nor2_1 _06551_ (.A(net2435),
    .B(_01310_),
    .Y(_01311_));
 sg13g2_nor3_1 _06552_ (.A(net2435),
    .B(_01308_),
    .C(_01309_),
    .Y(_01312_));
 sg13g2_nand2_1 _06553_ (.Y(_01313_),
    .A(_01028_),
    .B(_01310_));
 sg13g2_nor2_1 _06554_ (.A(_01028_),
    .B(_01310_),
    .Y(_01314_));
 sg13g2_o21ai_1 _06555_ (.B1(net2435),
    .Y(_01315_),
    .A1(_01308_),
    .A2(_01309_));
 sg13g2_nor2b_2 _06556_ (.A(_01312_),
    .B_N(_01315_),
    .Y(_01316_));
 sg13g2_nand3_1 _06557_ (.B(_01079_),
    .C(_01080_),
    .A(net2533),
    .Y(_01317_));
 sg13g2_nand2b_1 _06558_ (.Y(_01318_),
    .B(net2645),
    .A_N(\ChiselTop.wild.cpu.decExReg_decOut_imm[4] ));
 sg13g2_and2_2 _06559_ (.A(_01317_),
    .B(_01318_),
    .X(_01319_));
 sg13g2_nand2_1 _06560_ (.Y(_01320_),
    .A(_01317_),
    .B(_01318_));
 sg13g2_nand2b_1 _06561_ (.Y(_01321_),
    .B(_01319_),
    .A_N(_01078_));
 sg13g2_nand3_1 _06562_ (.B(_01317_),
    .C(_01318_),
    .A(_01078_),
    .Y(_01322_));
 sg13g2_nand2b_1 _06563_ (.Y(_01323_),
    .B(net2401),
    .A_N(_01078_));
 sg13g2_xnor2_1 _06564_ (.Y(_01324_),
    .A(_01078_),
    .B(net2401));
 sg13g2_inv_1 _06565_ (.Y(_01325_),
    .A(_01324_));
 sg13g2_and2_2 _06566_ (.A(net2644),
    .B(_00050_),
    .X(_01326_));
 sg13g2_nor3_2 _06567_ (.A(net2641),
    .B(_01121_),
    .C(_01122_),
    .Y(_01327_));
 sg13g2_or2_1 _06568_ (.X(_01328_),
    .B(_01327_),
    .A(_01326_));
 sg13g2_nor2_1 _06569_ (.A(_01326_),
    .B(_01327_),
    .Y(_01329_));
 sg13g2_nand2_1 _06570_ (.Y(_01330_),
    .A(_01119_),
    .B(net2395));
 sg13g2_nor3_1 _06571_ (.A(_01119_),
    .B(_01326_),
    .C(_01327_),
    .Y(_01331_));
 sg13g2_xnor2_1 _06572_ (.Y(_01332_),
    .A(_01120_),
    .B(net2394));
 sg13g2_nand2b_1 _06573_ (.Y(_01333_),
    .B(net2641),
    .A_N(_00054_));
 sg13g2_mux2_1 _06574_ (.A0(_00054_),
    .A1(_01026_),
    .S(net2532),
    .X(_01334_));
 sg13g2_o21ai_1 _06575_ (.B1(_01333_),
    .Y(_01335_),
    .A1(net2641),
    .A2(_01026_));
 sg13g2_nand2_1 _06576_ (.Y(_01336_),
    .A(_01025_),
    .B(net2363));
 sg13g2_nor2_1 _06577_ (.A(_01024_),
    .B(net2363),
    .Y(_01337_));
 sg13g2_xnor2_1 _06578_ (.Y(_01338_),
    .A(_01024_),
    .B(net2372));
 sg13g2_xnor2_1 _06579_ (.Y(_01339_),
    .A(_01025_),
    .B(net2372));
 sg13g2_and3_1 _06580_ (.X(_01340_),
    .A(net2532),
    .B(_01072_),
    .C(_01073_));
 sg13g2_nand3_1 _06581_ (.B(_01072_),
    .C(_01073_),
    .A(net2532),
    .Y(_01341_));
 sg13g2_nor2_1 _06582_ (.A(net2534),
    .B(_00058_),
    .Y(_01342_));
 sg13g2_nand2b_1 _06583_ (.Y(_01343_),
    .B(net2645),
    .A_N(_00058_));
 sg13g2_nand2_1 _06584_ (.Y(_01344_),
    .A(_01341_),
    .B(_01343_));
 sg13g2_nor2_1 _06585_ (.A(_01340_),
    .B(_01342_),
    .Y(_01345_));
 sg13g2_nor2_1 _06586_ (.A(_01071_),
    .B(net2348),
    .Y(_01346_));
 sg13g2_nor3_1 _06587_ (.A(net2427),
    .B(_01340_),
    .C(_01342_),
    .Y(_01347_));
 sg13g2_nand3b_1 _06588_ (.B(_01341_),
    .C(_01343_),
    .Y(_01348_),
    .A_N(net2427));
 sg13g2_o21ai_1 _06589_ (.B1(net2427),
    .Y(_01349_),
    .A1(_01340_),
    .A2(_01342_));
 sg13g2_and2_2 _06590_ (.A(_01348_),
    .B(_01349_),
    .X(_01350_));
 sg13g2_and3_2 _06591_ (.X(_01351_),
    .A(net2532),
    .B(_01097_),
    .C(_01098_));
 sg13g2_nand3_1 _06592_ (.B(_01097_),
    .C(_01098_),
    .A(net2532),
    .Y(_01352_));
 sg13g2_nor2_2 _06593_ (.A(net2534),
    .B(_00062_),
    .Y(_01353_));
 sg13g2_nand2b_1 _06594_ (.Y(_01354_),
    .B(net2645),
    .A_N(_00062_));
 sg13g2_nor2_1 _06595_ (.A(_01351_),
    .B(_01353_),
    .Y(_01355_));
 sg13g2_nor2_1 _06596_ (.A(_01096_),
    .B(net2337),
    .Y(_01356_));
 sg13g2_a221oi_1 _06597_ (.B2(_01354_),
    .C1(_01096_),
    .B1(_01352_),
    .A1(_01348_),
    .Y(_01357_),
    .A2(_01349_));
 sg13g2_nor2_1 _06598_ (.A(_01346_),
    .B(_01357_),
    .Y(_01358_));
 sg13g2_o21ai_1 _06599_ (.B1(_01339_),
    .Y(_01359_),
    .A1(_01346_),
    .A2(_01357_));
 sg13g2_nand2_1 _06600_ (.Y(_01360_),
    .A(_01336_),
    .B(_01359_));
 sg13g2_a21oi_1 _06601_ (.A1(_01336_),
    .A2(_01359_),
    .Y(_01361_),
    .B1(_01332_));
 sg13g2_nor2_1 _06602_ (.A(_01120_),
    .B(net2394),
    .Y(_01362_));
 sg13g2_o21ai_1 _06603_ (.B1(_01325_),
    .Y(_01363_),
    .A1(_01361_),
    .A2(_01362_));
 sg13g2_a21oi_1 _06604_ (.A1(_01321_),
    .A2(_01363_),
    .Y(_01364_),
    .B1(_01316_));
 sg13g2_o21ai_1 _06605_ (.B1(_01307_),
    .Y(_01365_),
    .A1(_01311_),
    .A2(_01364_));
 sg13g2_a21oi_2 _06606_ (.B1(_01302_),
    .Y(_01366_),
    .A2(_01365_),
    .A1(_01304_));
 sg13g2_o21ai_1 _06607_ (.B1(_01296_),
    .Y(_01367_),
    .A1(_01299_),
    .A2(_01366_));
 sg13g2_nor2_1 _06608_ (.A(_01291_),
    .B(_01295_),
    .Y(_01368_));
 sg13g2_o21ai_1 _06609_ (.B1(_01368_),
    .Y(_01369_),
    .A1(_01299_),
    .A2(_01366_));
 sg13g2_or2_1 _06610_ (.X(_01370_),
    .B(_01292_),
    .A(_01172_));
 sg13g2_nor2_1 _06611_ (.A(_01291_),
    .B(_01370_),
    .Y(_01371_));
 sg13g2_a21oi_1 _06612_ (.A1(_01109_),
    .A2(_01288_),
    .Y(_01372_),
    .B1(_01371_));
 sg13g2_and2_1 _06613_ (.A(_01282_),
    .B(_01372_),
    .X(_01373_));
 sg13g2_a22oi_1 _06614_ (.Y(_01374_),
    .B1(_01369_),
    .B2(_01373_),
    .A2(_01287_),
    .A1(_01282_));
 sg13g2_a221oi_1 _06615_ (.B2(_01373_),
    .C1(_01271_),
    .B1(_01369_),
    .A1(_01282_),
    .Y(_01375_),
    .A2(_01287_));
 sg13g2_nor2_1 _06616_ (.A(net2429),
    .B(_01268_),
    .Y(_01376_));
 sg13g2_nand3_1 _06617_ (.B(_01264_),
    .C(_01272_),
    .A(_01252_),
    .Y(_01377_));
 sg13g2_a221oi_1 _06618_ (.B2(_01373_),
    .C1(_01377_),
    .B1(_01369_),
    .A1(_01282_),
    .Y(_01378_),
    .A2(_01287_));
 sg13g2_nand2_1 _06619_ (.Y(_01379_),
    .A(_01252_),
    .B(_01376_));
 sg13g2_a21oi_1 _06620_ (.A1(_01266_),
    .A2(_01379_),
    .Y(_01380_),
    .B1(_01257_));
 sg13g2_o21ai_1 _06621_ (.B1(_01263_),
    .Y(_01381_),
    .A1(_01265_),
    .A2(_01380_));
 sg13g2_o21ai_1 _06622_ (.B1(_01381_),
    .Y(_01382_),
    .A1(_01131_),
    .A2(_01258_));
 sg13g2_nor3_1 _06623_ (.A(_01247_),
    .B(_01378_),
    .C(_01382_),
    .Y(_01383_));
 sg13g2_o21ai_1 _06624_ (.B1(_01247_),
    .Y(_01384_),
    .A1(_01378_),
    .A2(_01382_));
 sg13g2_nor2b_2 _06625_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[1] ),
    .B_N(_00066_),
    .Y(_01385_));
 sg13g2_nand2b_2 _06626_ (.Y(_01386_),
    .B(_00066_),
    .A_N(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[1] ));
 sg13g2_nor2_1 _06627_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[0] ),
    .B(_01386_),
    .Y(_01387_));
 sg13g2_nand2b_1 _06628_ (.Y(_01388_),
    .B(_01385_),
    .A_N(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[0] ));
 sg13g2_nor2_1 _06629_ (.A(_01383_),
    .B(net2496),
    .Y(_01389_));
 sg13g2_nor2_1 _06630_ (.A(net2321),
    .B(_01286_),
    .Y(_01390_));
 sg13g2_nand2b_1 _06631_ (.Y(_01391_),
    .B(_01285_),
    .A_N(net2321));
 sg13g2_nor4_1 _06632_ (.A(_01300_),
    .B(_01301_),
    .C(_01305_),
    .D(_01306_),
    .Y(_01392_));
 sg13g2_nand3_1 _06633_ (.B(_01324_),
    .C(_01392_),
    .A(_01316_),
    .Y(_01393_));
 sg13g2_o21ai_1 _06634_ (.B1(_01096_),
    .Y(_01394_),
    .A1(_01351_),
    .A2(_01353_));
 sg13g2_nor3_2 _06635_ (.A(_01096_),
    .B(_01351_),
    .C(_01353_),
    .Y(_01395_));
 sg13g2_xnor2_1 _06636_ (.Y(_01396_),
    .A(_01096_),
    .B(net2339));
 sg13g2_and4_1 _06637_ (.A(_01332_),
    .B(_01338_),
    .C(_01350_),
    .D(_01396_),
    .X(_01397_));
 sg13g2_nand4_1 _06638_ (.B(_01338_),
    .C(_01350_),
    .A(_01332_),
    .Y(_01398_),
    .D(_01396_));
 sg13g2_nor2_1 _06639_ (.A(_01393_),
    .B(_01398_),
    .Y(_01399_));
 sg13g2_nand2b_1 _06640_ (.Y(_01400_),
    .B(_01397_),
    .A_N(_01393_));
 sg13g2_a221oi_1 _06641_ (.B2(_01395_),
    .C1(_01347_),
    .B1(_01349_),
    .A1(_01025_),
    .Y(_01401_),
    .A2(net2372));
 sg13g2_a21o_1 _06642_ (.A2(net2363),
    .A1(_01024_),
    .B1(_01331_),
    .X(_01402_));
 sg13g2_o21ai_1 _06643_ (.B1(_01330_),
    .Y(_01403_),
    .A1(_01401_),
    .A2(_01402_));
 sg13g2_a21oi_1 _06644_ (.A1(_01315_),
    .A2(_01322_),
    .Y(_01404_),
    .B1(_01312_));
 sg13g2_a221oi_1 _06645_ (.B2(_01404_),
    .C1(_01300_),
    .B1(_01392_),
    .A1(_01302_),
    .Y(_01405_),
    .A2(_01305_));
 sg13g2_o21ai_1 _06646_ (.B1(_01405_),
    .Y(_01406_),
    .A1(_01393_),
    .A2(_01403_));
 sg13g2_a21oi_1 _06647_ (.A1(_01400_),
    .A2(_01406_),
    .Y(_01407_),
    .B1(_01296_));
 sg13g2_or2_1 _06648_ (.X(_01408_),
    .B(_01407_),
    .A(_01293_));
 sg13g2_nand3b_1 _06649_ (.B(_01290_),
    .C(_01295_),
    .Y(_01409_),
    .A_N(_01289_));
 sg13g2_a21oi_1 _06650_ (.A1(_01400_),
    .A2(_01406_),
    .Y(_01410_),
    .B1(_01409_));
 sg13g2_a21o_1 _06651_ (.A2(_01293_),
    .A1(_01290_),
    .B1(_01289_),
    .X(_01411_));
 sg13g2_nor2_1 _06652_ (.A(_01410_),
    .B(_01411_),
    .Y(_01412_));
 sg13g2_o21ai_1 _06653_ (.B1(_01390_),
    .Y(_01413_),
    .A1(_01410_),
    .A2(_01411_));
 sg13g2_nand2b_1 _06654_ (.Y(_01414_),
    .B(_01283_),
    .A_N(_01275_));
 sg13g2_nand2_1 _06655_ (.Y(_01415_),
    .A(_01276_),
    .B(_01414_));
 sg13g2_nand2_1 _06656_ (.Y(_01416_),
    .A(_01413_),
    .B(_01415_));
 sg13g2_a21o_1 _06657_ (.A2(_01415_),
    .A1(_01413_),
    .B1(_01272_),
    .X(_01417_));
 sg13g2_and2_1 _06658_ (.A(_01269_),
    .B(_01417_),
    .X(_01418_));
 sg13g2_nand3_1 _06659_ (.B(_01269_),
    .C(_01417_),
    .A(_01251_),
    .Y(_01419_));
 sg13g2_nor2b_1 _06660_ (.A(_01250_),
    .B_N(_01419_),
    .Y(_01420_));
 sg13g2_nand3b_1 _06661_ (.B(_01257_),
    .C(_01419_),
    .Y(_01421_),
    .A_N(_01250_));
 sg13g2_nor2b_1 _06662_ (.A(_01255_),
    .B_N(_01421_),
    .Y(_01422_));
 sg13g2_nor2b_1 _06663_ (.A(_01255_),
    .B_N(_01261_),
    .Y(_01423_));
 sg13g2_a21oi_1 _06664_ (.A1(_01421_),
    .A2(_01423_),
    .Y(_01424_),
    .B1(_01260_));
 sg13g2_and2_1 _06665_ (.A(net2640),
    .B(_01385_),
    .X(_01425_));
 sg13g2_nand2_1 _06666_ (.Y(_01426_),
    .A(net2640),
    .B(_01385_));
 sg13g2_a221oi_1 _06667_ (.B2(_01423_),
    .C1(_01247_),
    .B1(_01421_),
    .A1(_01131_),
    .Y(_01427_),
    .A2(_01259_));
 sg13g2_nor2_1 _06668_ (.A(_01426_),
    .B(_01427_),
    .Y(_01428_));
 sg13g2_o21ai_1 _06669_ (.B1(_01428_),
    .Y(_01429_),
    .A1(_01246_),
    .A2(_01424_));
 sg13g2_mux4_1 _06670_ (.S0(net2342),
    .A0(_01141_),
    .A1(_01113_),
    .A2(_00999_),
    .A3(_01064_),
    .S1(net2329),
    .X(_01430_));
 sg13g2_nand2_1 _06671_ (.Y(_01431_),
    .A(net2370),
    .B(_01430_));
 sg13g2_nand2_1 _06672_ (.Y(_01432_),
    .A(net2419),
    .B(net2337));
 sg13g2_o21ai_1 _06673_ (.B1(_01432_),
    .Y(_01433_),
    .A1(_01153_),
    .A2(net2339));
 sg13g2_o21ai_1 _06674_ (.B1(_01054_),
    .Y(_01434_),
    .A1(_01351_),
    .A2(_01353_));
 sg13g2_nand3_1 _06675_ (.B(_01352_),
    .C(_01354_),
    .A(net2414),
    .Y(_01435_));
 sg13g2_nand3_1 _06676_ (.B(_01434_),
    .C(_01435_),
    .A(net2353),
    .Y(_01436_));
 sg13g2_o21ai_1 _06677_ (.B1(_01436_),
    .Y(_01437_),
    .A1(net2353),
    .A2(_01433_));
 sg13g2_o21ai_1 _06678_ (.B1(_01431_),
    .Y(_01438_),
    .A1(net2370),
    .A2(_01437_));
 sg13g2_nand2_1 _06679_ (.Y(_01439_),
    .A(_01160_),
    .B(net2337));
 sg13g2_mux4_1 _06680_ (.S0(net2350),
    .A0(net2430),
    .A1(net2426),
    .A2(net2422),
    .A3(net2415),
    .S1(net2332),
    .X(_01440_));
 sg13g2_nor2b_1 _06681_ (.A(net2336),
    .B_N(net2425),
    .Y(_01441_));
 sg13g2_mux4_1 _06682_ (.S0(net2328),
    .A0(net2424),
    .A1(net2421),
    .A2(net2417),
    .A3(net2437),
    .S1(net2342),
    .X(_01442_));
 sg13g2_mux2_1 _06683_ (.A0(_01440_),
    .A1(_01442_),
    .S(net2359),
    .X(_01443_));
 sg13g2_mux2_1 _06684_ (.A0(_01438_),
    .A1(_01443_),
    .S(net2392),
    .X(_01444_));
 sg13g2_nor2b_2 _06685_ (.A(net2640),
    .B_N(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[1] ),
    .Y(_01445_));
 sg13g2_and2_1 _06686_ (.A(_00066_),
    .B(_01445_),
    .X(_01446_));
 sg13g2_nand2_1 _06687_ (.Y(_01447_),
    .A(_00066_),
    .B(_01445_));
 sg13g2_nand2_1 _06688_ (.Y(_01448_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[1] ),
    .B(net2640));
 sg13g2_nor2_2 _06689_ (.A(_00066_),
    .B(_01448_),
    .Y(_01449_));
 sg13g2_or2_2 _06690_ (.X(_01450_),
    .B(_01448_),
    .A(_00066_));
 sg13g2_nand2_1 _06691_ (.Y(_01451_),
    .A(net2431),
    .B(_01449_));
 sg13g2_nand2_2 _06692_ (.Y(_01452_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[2] ),
    .B(_01445_));
 sg13g2_a22oi_1 _06693_ (.Y(_01453_),
    .B1(_01449_),
    .B2(net2400),
    .A2(_01445_),
    .A1(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[2] ));
 sg13g2_o21ai_1 _06694_ (.B1(_01452_),
    .Y(_01454_),
    .A1(net2403),
    .A2(_01450_));
 sg13g2_a21oi_1 _06695_ (.A1(_01451_),
    .A2(net2319),
    .Y(_01455_),
    .B1(net2484));
 sg13g2_nor2_1 _06696_ (.A(net2398),
    .B(_01452_),
    .Y(_01456_));
 sg13g2_or2_2 _06697_ (.X(_01457_),
    .B(_01452_),
    .A(net2398));
 sg13g2_a21oi_1 _06698_ (.A1(net2398),
    .A2(_01444_),
    .Y(_01458_),
    .B1(_01456_));
 sg13g2_nand2_1 _06699_ (.Y(_01459_),
    .A(_01455_),
    .B(_01458_));
 sg13g2_nor2_1 _06700_ (.A(net2427),
    .B(net2339),
    .Y(_01460_));
 sg13g2_a21oi_1 _06701_ (.A1(_01025_),
    .A2(net2339),
    .Y(_01461_),
    .B1(_01460_));
 sg13g2_nand2_1 _06702_ (.Y(_01462_),
    .A(_01078_),
    .B(net2340));
 sg13g2_o21ai_1 _06703_ (.B1(_01462_),
    .Y(_01463_),
    .A1(_01119_),
    .A2(net2340));
 sg13g2_mux2_1 _06704_ (.A0(_01461_),
    .A1(_01463_),
    .S(net2348),
    .X(_01464_));
 sg13g2_o21ai_1 _06705_ (.B1(_01027_),
    .Y(_01465_),
    .A1(_01351_),
    .A2(_01353_));
 sg13g2_nand2_1 _06706_ (.Y(_01466_),
    .A(_01037_),
    .B(net2340));
 sg13g2_o21ai_1 _06707_ (.B1(net2436),
    .Y(_01467_),
    .A1(_01351_),
    .A2(_01353_));
 sg13g2_mux4_1 _06708_ (.S0(net2355),
    .A0(_01022_),
    .A1(_01028_),
    .A2(_01171_),
    .A3(_01036_),
    .S1(net2340),
    .X(_01468_));
 sg13g2_nand2_1 _06709_ (.Y(_01469_),
    .A(net2373),
    .B(_01468_));
 sg13g2_o21ai_1 _06710_ (.B1(_01469_),
    .Y(_01470_),
    .A1(net2373),
    .A2(_01464_));
 sg13g2_nor2_1 _06711_ (.A(_01048_),
    .B(net2340),
    .Y(_01471_));
 sg13g2_a221oi_1 _06712_ (.B2(_01104_),
    .C1(_01471_),
    .B1(net2339),
    .A1(_01341_),
    .Y(_01472_),
    .A2(_01343_));
 sg13g2_nor2_1 _06713_ (.A(_01130_),
    .B(net2340),
    .Y(_01473_));
 sg13g2_a21oi_1 _06714_ (.A1(net2422),
    .A2(net2339),
    .Y(_01474_),
    .B1(_01473_));
 sg13g2_a21oi_1 _06715_ (.A1(net2348),
    .A2(_01474_),
    .Y(_01475_),
    .B1(_01472_));
 sg13g2_mux4_1 _06716_ (.S0(net2349),
    .A0(_01108_),
    .A1(_01093_),
    .A2(net2433),
    .A3(net2428),
    .S1(net2338),
    .X(_01476_));
 sg13g2_mux2_1 _06717_ (.A0(_01475_),
    .A1(_01476_),
    .S(net2363),
    .X(_01477_));
 sg13g2_nor2_1 _06718_ (.A(net2403),
    .B(net2483),
    .Y(_01478_));
 sg13g2_nand2_1 _06719_ (.Y(_01479_),
    .A(net2400),
    .B(net2486));
 sg13g2_a21oi_1 _06720_ (.A1(net2394),
    .A2(_01477_),
    .Y(_01480_),
    .B1(net2315));
 sg13g2_o21ai_1 _06721_ (.B1(_01480_),
    .Y(_01481_),
    .A1(net2396),
    .A2(_01470_));
 sg13g2_nand2_1 _06722_ (.Y(_01482_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[2] ),
    .B(net2640));
 sg13g2_nor2_2 _06723_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[1] ),
    .B(_01482_),
    .Y(_01483_));
 sg13g2_or2_1 _06724_ (.X(_01484_),
    .B(_01482_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[1] ));
 sg13g2_nor2_2 _06725_ (.A(net2400),
    .B(net2482),
    .Y(_01485_));
 sg13g2_nand2_2 _06726_ (.Y(_01486_),
    .A(net2403),
    .B(net2484));
 sg13g2_nand2_1 _06727_ (.Y(_01487_),
    .A(net2349),
    .B(_01395_));
 sg13g2_nand3_1 _06728_ (.B(net2348),
    .C(_01395_),
    .A(net2373),
    .Y(_01488_));
 sg13g2_nor2_1 _06729_ (.A(net2382),
    .B(_01488_),
    .Y(_01489_));
 sg13g2_a21oi_1 _06730_ (.A1(net2313),
    .A2(_01489_),
    .Y(_01490_),
    .B1(net2476));
 sg13g2_nand3_1 _06731_ (.B(_01481_),
    .C(_01490_),
    .A(_01459_),
    .Y(_01491_));
 sg13g2_a21oi_1 _06732_ (.A1(_01246_),
    .A2(net2479),
    .Y(_01492_),
    .B1(net2494));
 sg13g2_a221oi_1 _06733_ (.B2(_01492_),
    .C1(net2634),
    .B1(_01491_),
    .A1(_01384_),
    .Y(_01493_),
    .A2(_01389_));
 sg13g2_a22oi_1 _06734_ (.Y(_01494_),
    .B1(_01429_),
    .B2(_01493_),
    .A2(net2633),
    .A1(net1494));
 sg13g2_xnor2_1 _06735_ (.Y(_01495_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[16] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[16] ));
 sg13g2_nor2_1 _06736_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[15] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[15] ),
    .Y(_01496_));
 sg13g2_and2_1 _06737_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[14] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[14] ),
    .X(_01497_));
 sg13g2_xor2_1 _06738_ (.B(\ChiselTop.wild.cpu.decExReg_pc[14] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[14] ),
    .X(_01498_));
 sg13g2_nand2_1 _06739_ (.Y(_01499_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[13] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[13] ));
 sg13g2_and2_1 _06740_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[12] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[12] ),
    .X(_01500_));
 sg13g2_nand2_1 _06741_ (.Y(_01501_),
    .A(net1530),
    .B(\ChiselTop.wild.cpu.decExReg_pc[11] ));
 sg13g2_and2_1 _06742_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[10] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[10] ),
    .X(_01502_));
 sg13g2_xnor2_1 _06743_ (.Y(_01503_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[10] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[9] ));
 sg13g2_inv_1 _06744_ (.Y(_01504_),
    .A(_01503_));
 sg13g2_xor2_1 _06745_ (.B(\ChiselTop.wild.cpu.decExReg_pc[8] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[10] ),
    .X(_01505_));
 sg13g2_inv_1 _06746_ (.Y(_01506_),
    .A(_01505_));
 sg13g2_or2_1 _06747_ (.X(_01507_),
    .B(\ChiselTop.wild.cpu.decExReg_pc[7] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[6] ));
 sg13g2_xnor2_1 _06748_ (.Y(_01508_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[6] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[6] ));
 sg13g2_and2_1 _06749_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[5] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[5] ),
    .X(_01509_));
 sg13g2_nand2_1 _06750_ (.Y(_01510_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[4] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[4] ));
 sg13g2_xnor2_1 _06751_ (.Y(_01511_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[4] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[4] ));
 sg13g2_and2_1 _06752_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[3] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[3] ),
    .X(_01512_));
 sg13g2_nand2_1 _06753_ (.Y(_01513_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[2] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[2] ));
 sg13g2_nor2_1 _06754_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[2] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[2] ),
    .Y(_01514_));
 sg13g2_xor2_1 _06755_ (.B(\ChiselTop.wild.cpu.decExReg_pc[2] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[2] ),
    .X(_01515_));
 sg13g2_and2_1 _06756_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[1] ),
    .B(\ChiselTop.wild.cpu._wbData_T_1[1] ),
    .X(_01516_));
 sg13g2_and2_1 _06757_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[0] ),
    .B(\ChiselTop.wild.cpu._wbData_T_1[0] ),
    .X(_01517_));
 sg13g2_xor2_1 _06758_ (.B(\ChiselTop.wild.cpu._wbData_T_1[1] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[1] ),
    .X(_01518_));
 sg13g2_a21oi_1 _06759_ (.A1(_01517_),
    .A2(_01518_),
    .Y(_01519_),
    .B1(_01516_));
 sg13g2_o21ai_1 _06760_ (.B1(_01513_),
    .Y(_01520_),
    .A1(_01514_),
    .A2(_01519_));
 sg13g2_xor2_1 _06761_ (.B(\ChiselTop.wild.cpu.decExReg_pc[3] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[3] ),
    .X(_01521_));
 sg13g2_a21oi_1 _06762_ (.A1(_01520_),
    .A2(_01521_),
    .Y(_01522_),
    .B1(_01512_));
 sg13g2_o21ai_1 _06763_ (.B1(_01510_),
    .Y(_01523_),
    .A1(_01511_),
    .A2(_01522_));
 sg13g2_xor2_1 _06764_ (.B(\ChiselTop.wild.cpu.decExReg_pc[5] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[5] ),
    .X(_01524_));
 sg13g2_a21o_2 _06765_ (.A2(_01524_),
    .A1(_01523_),
    .B1(_01509_),
    .X(_01525_));
 sg13g2_nor2b_1 _06766_ (.A(_01508_),
    .B_N(_01525_),
    .Y(_01526_));
 sg13g2_a21o_1 _06767_ (.A2(\ChiselTop.wild.cpu.decExReg_pc[6] ),
    .A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[6] ),
    .B1(_01526_),
    .X(_01527_));
 sg13g2_nand3b_1 _06768_ (.B(_01525_),
    .C(_01507_),
    .Y(_01528_),
    .A_N(_01508_));
 sg13g2_o21ai_1 _06769_ (.B1(\ChiselTop.wild.cpu.decExReg_decOut_imm[6] ),
    .Y(_01529_),
    .A1(\ChiselTop.wild.cpu.decExReg_pc[7] ),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[6] ));
 sg13g2_a21oi_2 _06770_ (.B1(_01506_),
    .Y(_01530_),
    .A2(_01529_),
    .A1(_01528_));
 sg13g2_o21ai_1 _06771_ (.B1(\ChiselTop.wild.cpu.decExReg_decOut_imm[10] ),
    .Y(_01531_),
    .A1(\ChiselTop.wild.cpu.decExReg_pc[9] ),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[8] ));
 sg13g2_inv_1 _06772_ (.Y(_01532_),
    .A(_01531_));
 sg13g2_a21o_1 _06773_ (.A2(_01530_),
    .A1(_01504_),
    .B1(_01532_),
    .X(_01533_));
 sg13g2_xor2_1 _06774_ (.B(\ChiselTop.wild.cpu.decExReg_pc[10] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[10] ),
    .X(_01534_));
 sg13g2_a21oi_1 _06775_ (.A1(_01533_),
    .A2(_01534_),
    .Y(_01535_),
    .B1(_01502_));
 sg13g2_xnor2_1 _06776_ (.Y(_01536_),
    .A(net1397),
    .B(\ChiselTop.wild.cpu.decExReg_pc[11] ));
 sg13g2_o21ai_1 _06777_ (.B1(_01501_),
    .Y(_01537_),
    .A1(_01535_),
    .A2(_01536_));
 sg13g2_xor2_1 _06778_ (.B(\ChiselTop.wild.cpu.decExReg_pc[12] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[12] ),
    .X(_01538_));
 sg13g2_a21oi_2 _06779_ (.B1(_01500_),
    .Y(_01539_),
    .A2(_01538_),
    .A1(_01537_));
 sg13g2_xnor2_1 _06780_ (.Y(_01540_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[13] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[13] ));
 sg13g2_o21ai_1 _06781_ (.B1(_01499_),
    .Y(_01541_),
    .A1(_01539_),
    .A2(_01540_));
 sg13g2_a21oi_1 _06782_ (.A1(_01498_),
    .A2(_01541_),
    .Y(_01542_),
    .B1(_01497_));
 sg13g2_a221oi_1 _06783_ (.B2(_01541_),
    .C1(_01497_),
    .B1(_01498_),
    .A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[15] ),
    .Y(_01543_),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[15] ));
 sg13g2_nor3_1 _06784_ (.A(_01495_),
    .B(_01496_),
    .C(_01543_),
    .Y(_01544_));
 sg13g2_o21ai_1 _06785_ (.B1(_01495_),
    .Y(_01545_),
    .A1(_01496_),
    .A2(_01543_));
 sg13g2_nand2b_1 _06786_ (.Y(_01546_),
    .B(_01545_),
    .A_N(_01544_));
 sg13g2_nor2b_2 _06787_ (.A(net2185),
    .B_N(_00003_),
    .Y(_01547_));
 sg13g2_nand2b_1 _06788_ (.Y(_01548_),
    .B(_00003_),
    .A_N(net2185));
 sg13g2_o21ai_1 _06789_ (.B1(_01547_),
    .Y(_01549_),
    .A1(net2623),
    .A2(_01494_));
 sg13g2_a21oi_1 _06790_ (.A1(net2623),
    .A2(_01546_),
    .Y(_01550_),
    .B1(_01549_));
 sg13g2_a21o_1 _06791_ (.A2(_01243_),
    .A1(net2184),
    .B1(_01550_),
    .X(_01551_));
 sg13g2_nor2_1 _06792_ (.A(net2540),
    .B(_00987_),
    .Y(_01552_));
 sg13g2_a22oi_1 _06793_ (.Y(_01553_),
    .B1(_01552_),
    .B2(_00986_),
    .A2(_01551_),
    .A1(net2541));
 sg13g2_mux4_1 _06794_ (.S0(net2682),
    .A0(\ChiselTop.wild.cpu.regs[0][16] ),
    .A1(\ChiselTop.wild.cpu.regs[1][16] ),
    .A2(\ChiselTop.wild.cpu.regs[2][16] ),
    .A3(\ChiselTop.wild.cpu.regs[3][16] ),
    .S1(net2664),
    .X(_01554_));
 sg13g2_nor2_1 _06795_ (.A(net2651),
    .B(_01554_),
    .Y(_01555_));
 sg13g2_nor2_1 _06796_ (.A(net2703),
    .B(net2676),
    .Y(_01556_));
 sg13g2_nand2_1 _06797_ (.Y(_01557_),
    .A(net1539),
    .B(_01556_));
 sg13g2_nor2b_1 _06798_ (.A(\ChiselTop.wild.cpu.regs[5][16] ),
    .B_N(net2682),
    .Y(_01558_));
 sg13g2_nor2_1 _06799_ (.A(net2682),
    .B(\ChiselTop.wild.cpu.regs[4][16] ),
    .Y(_01559_));
 sg13g2_nor3_1 _06800_ (.A(net2664),
    .B(_01558_),
    .C(_01559_),
    .Y(_01560_));
 sg13g2_nor2b_1 _06801_ (.A(\ChiselTop.wild.cpu.regs[7][16] ),
    .B_N(net2692),
    .Y(_01561_));
 sg13g2_o21ai_1 _06802_ (.B1(net2670),
    .Y(_01562_),
    .A1(net2692),
    .A2(\ChiselTop.wild.cpu.regs[6][16] ));
 sg13g2_o21ai_1 _06803_ (.B1(net2659),
    .Y(_01563_),
    .A1(_01561_),
    .A2(_01562_));
 sg13g2_o21ai_1 _06804_ (.B1(net2466),
    .Y(_01564_),
    .A1(_01560_),
    .A2(_01563_));
 sg13g2_nor2_1 _06805_ (.A(_01555_),
    .B(_01564_),
    .Y(_01565_));
 sg13g2_nor2_1 _06806_ (.A(net2439),
    .B(_01565_),
    .Y(_01566_));
 sg13g2_a21oi_2 _06807_ (.B1(_01566_),
    .Y(_01567_),
    .A2(net2113),
    .A1(net2440));
 sg13g2_xor2_1 _06808_ (.B(_01567_),
    .A(_00965_),
    .X(_01568_));
 sg13g2_and2_2 _06809_ (.A(\ChiselTop.wild.cpu._GEN_176[6] ),
    .B(net2523),
    .X(_01569_));
 sg13g2_nor2_1 _06810_ (.A(_00117_),
    .B(_00978_),
    .Y(_01570_));
 sg13g2_xnor2_1 _06811_ (.Y(_01571_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[7] ),
    .B(_01570_));
 sg13g2_nand2_1 _06812_ (.Y(_01572_),
    .A(net2614),
    .B(_01571_));
 sg13g2_nand2_1 _06813_ (.Y(_01573_),
    .A(_00037_),
    .B(net2637));
 sg13g2_nand3_1 _06814_ (.B(_01304_),
    .C(_01365_),
    .A(_01302_),
    .Y(_01574_));
 sg13g2_nand3b_1 _06815_ (.B(net2499),
    .C(_01574_),
    .Y(_01575_),
    .A_N(_01366_));
 sg13g2_nor2_2 _06816_ (.A(_01054_),
    .B(net2385),
    .Y(_01576_));
 sg13g2_nand2_1 _06817_ (.Y(_01577_),
    .A(net2432),
    .B(net2384));
 sg13g2_nor2_1 _06818_ (.A(_00999_),
    .B(net2335),
    .Y(_01578_));
 sg13g2_nand2_1 _06819_ (.Y(_01579_),
    .A(_01112_),
    .B(net2335));
 sg13g2_mux2_1 _06820_ (.A0(_00999_),
    .A1(_01113_),
    .S(net2329),
    .X(_01580_));
 sg13g2_mux4_1 _06821_ (.S0(net2342),
    .A0(_00999_),
    .A1(_01064_),
    .A2(_01113_),
    .A3(net2424),
    .S1(net2328),
    .X(_01581_));
 sg13g2_mux2_1 _06822_ (.A0(net2414),
    .A1(net2416),
    .S(net2332),
    .X(_01582_));
 sg13g2_mux2_1 _06823_ (.A0(net2419),
    .A1(_01141_),
    .S(net2329),
    .X(_01583_));
 sg13g2_mux4_1 _06824_ (.S0(net2328),
    .A0(net2419),
    .A1(_01141_),
    .A2(net2414),
    .A3(net2416),
    .S1(net2352),
    .X(_01584_));
 sg13g2_mux2_1 _06825_ (.A0(_01581_),
    .A1(_01584_),
    .S(net2356),
    .X(_01585_));
 sg13g2_nor2_1 _06826_ (.A(net2377),
    .B(_01585_),
    .Y(_01586_));
 sg13g2_nor2_1 _06827_ (.A(_01576_),
    .B(_01586_),
    .Y(_01587_));
 sg13g2_o21ai_1 _06828_ (.B1(net2319),
    .Y(_01588_),
    .A1(net2480),
    .A2(_01587_));
 sg13g2_nand2_1 _06829_ (.Y(_01589_),
    .A(net2431),
    .B(net2332));
 sg13g2_nand3_1 _06830_ (.B(net2343),
    .C(net2332),
    .A(net2431),
    .Y(_01590_));
 sg13g2_nor2_1 _06831_ (.A(net2357),
    .B(_01590_),
    .Y(_01591_));
 sg13g2_a21oi_1 _06832_ (.A1(net2377),
    .A2(_01591_),
    .Y(_01592_),
    .B1(_01586_));
 sg13g2_mux2_1 _06833_ (.A0(_01104_),
    .A1(_01047_),
    .S(net2330),
    .X(_01593_));
 sg13g2_mux2_1 _06834_ (.A0(net2429),
    .A1(_01093_),
    .S(net2330),
    .X(_01594_));
 sg13g2_mux2_1 _06835_ (.A0(_01593_),
    .A1(_01594_),
    .S(net2342),
    .X(_01595_));
 sg13g2_nor2_1 _06836_ (.A(net2365),
    .B(_01595_),
    .Y(_01596_));
 sg13g2_nand2_1 _06837_ (.Y(_01597_),
    .A(net2420),
    .B(net2334));
 sg13g2_mux2_1 _06838_ (.A0(net2434),
    .A1(net2420),
    .S(net2330),
    .X(_01598_));
 sg13g2_mux2_1 _06839_ (.A0(_01172_),
    .A1(net2436),
    .S(net2330),
    .X(_01599_));
 sg13g2_mux2_1 _06840_ (.A0(_01598_),
    .A1(_01599_),
    .S(net2342),
    .X(_01600_));
 sg13g2_o21ai_1 _06841_ (.B1(net2386),
    .Y(_01601_),
    .A1(net2357),
    .A2(_01600_));
 sg13g2_nand2_1 _06842_ (.Y(_01602_),
    .A(_01131_),
    .B(net2335));
 sg13g2_mux2_1 _06843_ (.A0(net2422),
    .A1(_01131_),
    .S(net2328),
    .X(_01603_));
 sg13g2_mux4_1 _06844_ (.S0(net2350),
    .A0(net2422),
    .A1(net2415),
    .A2(_01131_),
    .A3(net2430),
    .S1(net2332),
    .X(_01604_));
 sg13g2_nand2_1 _06845_ (.Y(_01605_),
    .A(net2418),
    .B(net2334));
 sg13g2_nand2_1 _06846_ (.Y(_01606_),
    .A(net2426),
    .B(net2334));
 sg13g2_mux4_1 _06847_ (.S0(net2328),
    .A0(net2437),
    .A1(net2426),
    .A2(net2421),
    .A3(net2417),
    .S1(net2350),
    .X(_01607_));
 sg13g2_mux2_1 _06848_ (.A0(_01604_),
    .A1(_01607_),
    .S(net2357),
    .X(_01608_));
 sg13g2_nand2_1 _06849_ (.Y(_01609_),
    .A(net2376),
    .B(_01608_));
 sg13g2_o21ai_1 _06850_ (.B1(_01609_),
    .Y(_01610_),
    .A1(_01596_),
    .A2(_01601_));
 sg13g2_a22oi_1 _06851_ (.Y(_01611_),
    .B1(_01610_),
    .B2(net2397),
    .A2(_01592_),
    .A1(net2318));
 sg13g2_nand3_1 _06852_ (.B(_01588_),
    .C(_01611_),
    .A(net2481),
    .Y(_01612_));
 sg13g2_o21ai_1 _06853_ (.B1(net2489),
    .Y(_01613_),
    .A1(_01302_),
    .A2(net2472));
 sg13g2_nor2b_1 _06854_ (.A(net2333),
    .B_N(_01078_),
    .Y(_01614_));
 sg13g2_a21oi_1 _06855_ (.A1(net2435),
    .A2(net2333),
    .Y(_01615_),
    .B1(_01614_));
 sg13g2_nor2_1 _06856_ (.A(_01036_),
    .B(net2335),
    .Y(_01616_));
 sg13g2_a21oi_1 _06857_ (.A1(net2436),
    .A2(net2333),
    .Y(_01617_),
    .B1(_01616_));
 sg13g2_mux2_1 _06858_ (.A0(_01615_),
    .A1(_01617_),
    .S(net2344),
    .X(_01618_));
 sg13g2_mux2_1 _06859_ (.A0(_01024_),
    .A1(_01120_),
    .S(net2333),
    .X(_01619_));
 sg13g2_nand3_1 _06860_ (.B(_01352_),
    .C(_01354_),
    .A(net2427),
    .Y(_01620_));
 sg13g2_nand2_2 _06861_ (.Y(_01621_),
    .A(_01394_),
    .B(_01620_));
 sg13g2_mux2_1 _06862_ (.A0(_01619_),
    .A1(_01621_),
    .S(net2351),
    .X(_01622_));
 sg13g2_nand2_1 _06863_ (.Y(_01623_),
    .A(net2360),
    .B(_01622_));
 sg13g2_o21ai_1 _06864_ (.B1(_01623_),
    .Y(_01624_),
    .A1(net2360),
    .A2(_01618_));
 sg13g2_nor2_1 _06865_ (.A(net2380),
    .B(_01624_),
    .Y(_01625_));
 sg13g2_a21oi_1 _06866_ (.A1(net2317),
    .A2(_01625_),
    .Y(_01626_),
    .B1(_01613_));
 sg13g2_nand2_1 _06867_ (.Y(_01627_),
    .A(_01612_),
    .B(_01626_));
 sg13g2_nand2b_1 _06868_ (.Y(_01628_),
    .B(_01398_),
    .A_N(_01403_));
 sg13g2_o21ai_1 _06869_ (.B1(_01324_),
    .Y(_01629_),
    .A1(_01397_),
    .A2(_01403_));
 sg13g2_nand2_1 _06870_ (.Y(_01630_),
    .A(_01323_),
    .B(_01629_));
 sg13g2_and3_1 _06871_ (.X(_01631_),
    .A(_01313_),
    .B(_01323_),
    .C(_01629_));
 sg13g2_or3_1 _06872_ (.A(_01307_),
    .B(_01314_),
    .C(_01631_),
    .X(_01632_));
 sg13g2_nor2b_1 _06873_ (.A(_01306_),
    .B_N(_01632_),
    .Y(_01633_));
 sg13g2_xnor2_1 _06874_ (.Y(_01634_),
    .A(_01302_),
    .B(_01633_));
 sg13g2_o21ai_1 _06875_ (.B1(_01627_),
    .Y(_01635_),
    .A1(net2489),
    .A2(_01634_));
 sg13g2_nand3_1 _06876_ (.B(_01575_),
    .C(_01635_),
    .A(net2530),
    .Y(_01636_));
 sg13g2_a21oi_1 _06877_ (.A1(_01573_),
    .A2(_01636_),
    .Y(_01637_),
    .B1(net2626));
 sg13g2_xor2_1 _06878_ (.B(\ChiselTop.wild.cpu.decExReg_pc[7] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[6] ),
    .X(_01638_));
 sg13g2_xnor2_1 _06879_ (.Y(_01639_),
    .A(_01527_),
    .B(_01638_));
 sg13g2_a21o_1 _06880_ (.A2(_01639_),
    .A1(net2625),
    .B1(net2171),
    .X(_01640_));
 sg13g2_nand2_1 _06881_ (.Y(_01641_),
    .A(net2185),
    .B(_01238_));
 sg13g2_nor2_2 _06882_ (.A(net2611),
    .B(_01234_),
    .Y(_01642_));
 sg13g2_nor2_2 _06883_ (.A(_01178_),
    .B(_01234_),
    .Y(_01643_));
 sg13g2_nand2_2 _06884_ (.Y(_01644_),
    .A(_01177_),
    .B(_01233_));
 sg13g2_nor2_2 _06885_ (.A(net2525),
    .B(_01643_),
    .Y(_01645_));
 sg13g2_inv_1 _06886_ (.Y(_01646_),
    .A(_01645_));
 sg13g2_nand3_1 _06887_ (.B(_01176_),
    .C(net2501),
    .A(\ChiselTop.wild.dmem.MEM_2[0][7] ),
    .Y(_01647_));
 sg13g2_a22oi_1 _06888_ (.Y(_01648_),
    .B1(_01646_),
    .B2(_01647_),
    .A2(_01644_),
    .A1(_01227_));
 sg13g2_o21ai_1 _06889_ (.B1(net2183),
    .Y(_01649_),
    .A1(net2322),
    .A2(_01648_));
 sg13g2_o21ai_1 _06890_ (.B1(_01649_),
    .Y(_01650_),
    .A1(_01637_),
    .A2(_01640_));
 sg13g2_o21ai_1 _06891_ (.B1(_01572_),
    .Y(_01651_),
    .A1(net2613),
    .A2(_01650_));
 sg13g2_mux4_1 _06892_ (.S0(net2689),
    .A0(\ChiselTop.wild.cpu.regs[0][7] ),
    .A1(\ChiselTop.wild.cpu.regs[1][7] ),
    .A2(\ChiselTop.wild.cpu.regs[2][7] ),
    .A3(\ChiselTop.wild.cpu.regs[3][7] ),
    .S1(net2668),
    .X(_01652_));
 sg13g2_nor2_1 _06893_ (.A(net2655),
    .B(_01652_),
    .Y(_01653_));
 sg13g2_nor2b_1 _06894_ (.A(\ChiselTop.wild.cpu.regs[5][7] ),
    .B_N(net2689),
    .Y(_01654_));
 sg13g2_nor2_1 _06895_ (.A(net2689),
    .B(\ChiselTop.wild.cpu.regs[4][7] ),
    .Y(_01655_));
 sg13g2_nor3_1 _06896_ (.A(net2669),
    .B(_01654_),
    .C(_01655_),
    .Y(_01656_));
 sg13g2_nor2b_1 _06897_ (.A(\ChiselTop.wild.cpu.regs[7][7] ),
    .B_N(net2689),
    .Y(_01657_));
 sg13g2_o21ai_1 _06898_ (.B1(net2669),
    .Y(_01658_),
    .A1(net2689),
    .A2(\ChiselTop.wild.cpu.regs[6][7] ));
 sg13g2_o21ai_1 _06899_ (.B1(net2655),
    .Y(_01659_),
    .A1(_01657_),
    .A2(_01658_));
 sg13g2_o21ai_1 _06900_ (.B1(net2470),
    .Y(_01660_),
    .A1(_01656_),
    .A2(_01659_));
 sg13g2_nor2_1 _06901_ (.A(_01653_),
    .B(_01660_),
    .Y(_01661_));
 sg13g2_nor2_1 _06902_ (.A(net2440),
    .B(_01661_),
    .Y(_01662_));
 sg13g2_a21oi_1 _06903_ (.A1(net2441),
    .A2(net2146),
    .Y(_01663_),
    .B1(_01662_));
 sg13g2_mux4_1 _06904_ (.S0(net2350),
    .A0(net2424),
    .A1(_01113_),
    .A2(net2421),
    .A3(_01064_),
    .S1(net2328),
    .X(_01664_));
 sg13g2_mux4_1 _06905_ (.S0(net2342),
    .A0(net2416),
    .A1(_01141_),
    .A2(net2419),
    .A3(_00999_),
    .S1(net2328),
    .X(_01665_));
 sg13g2_mux2_1 _06906_ (.A0(_01664_),
    .A1(_01665_),
    .S(net2358),
    .X(_01666_));
 sg13g2_nand2_1 _06907_ (.Y(_01667_),
    .A(net2391),
    .B(_01666_));
 sg13g2_inv_1 _06908_ (.Y(_01668_),
    .A(_01667_));
 sg13g2_nand3_1 _06909_ (.B(_01434_),
    .C(_01435_),
    .A(net2348),
    .Y(_01669_));
 sg13g2_or2_1 _06910_ (.X(_01670_),
    .B(_01669_),
    .A(net2358));
 sg13g2_and2_1 _06911_ (.A(net2381),
    .B(_01670_),
    .X(_01671_));
 sg13g2_nor2_1 _06912_ (.A(_01668_),
    .B(_01671_),
    .Y(_01672_));
 sg13g2_nand2_1 _06913_ (.Y(_01673_),
    .A(net2431),
    .B(net2354));
 sg13g2_o21ai_1 _06914_ (.B1(net2431),
    .Y(_01674_),
    .A1(net2358),
    .A2(net2354));
 sg13g2_nand2_1 _06915_ (.Y(_01675_),
    .A(_01670_),
    .B(_01674_));
 sg13g2_o21ai_1 _06916_ (.B1(_01667_),
    .Y(_01676_),
    .A1(net2391),
    .A2(_01675_));
 sg13g2_o21ai_1 _06917_ (.B1(net2320),
    .Y(_01677_),
    .A1(_01450_),
    .A2(_01676_));
 sg13g2_o21ai_1 _06918_ (.B1(net2318),
    .Y(_01678_),
    .A1(_01668_),
    .A2(_01671_));
 sg13g2_mux4_1 _06919_ (.S0(net2338),
    .A0(_01023_),
    .A1(_01037_),
    .A2(_01108_),
    .A3(_01172_),
    .S1(net2354),
    .X(_01679_));
 sg13g2_inv_1 _06920_ (.Y(_01680_),
    .A(_01679_));
 sg13g2_mux4_1 _06921_ (.S0(net2341),
    .A0(_01047_),
    .A1(net2428),
    .A2(_01093_),
    .A3(net2433),
    .S1(net2349),
    .X(_01681_));
 sg13g2_o21ai_1 _06922_ (.B1(net2392),
    .Y(_01682_),
    .A1(net2371),
    .A2(_01681_));
 sg13g2_a21oi_1 _06923_ (.A1(net2370),
    .A2(_01680_),
    .Y(_01683_),
    .B1(_01682_));
 sg13g2_mux4_1 _06924_ (.S0(net2338),
    .A0(net2430),
    .A1(net2422),
    .A2(_01131_),
    .A3(_01104_),
    .S1(net2349),
    .X(_01684_));
 sg13g2_and2_1 _06925_ (.A(net2370),
    .B(_01684_),
    .X(_01685_));
 sg13g2_mux4_1 _06926_ (.S0(net2328),
    .A0(net2426),
    .A1(net2415),
    .A2(net2417),
    .A3(net2437),
    .S1(net2350),
    .X(_01686_));
 sg13g2_a21oi_1 _06927_ (.A1(net2358),
    .A2(_01686_),
    .Y(_01687_),
    .B1(_01685_));
 sg13g2_nor2_1 _06928_ (.A(net2391),
    .B(_01687_),
    .Y(_01688_));
 sg13g2_o21ai_1 _06929_ (.B1(net2398),
    .Y(_01689_),
    .A1(_01683_),
    .A2(_01688_));
 sg13g2_nand4_1 _06930_ (.B(_01677_),
    .C(_01678_),
    .A(net2483),
    .Y(_01690_),
    .D(_01689_));
 sg13g2_a21oi_1 _06931_ (.A1(_01465_),
    .A2(_01466_),
    .Y(_01691_),
    .B1(net2355));
 sg13g2_a21oi_1 _06932_ (.A1(net2355),
    .A2(_01463_),
    .Y(_01692_),
    .B1(_01691_));
 sg13g2_nand2_1 _06933_ (.Y(_01693_),
    .A(net2353),
    .B(_01395_));
 sg13g2_o21ai_1 _06934_ (.B1(_01693_),
    .Y(_01694_),
    .A1(net2353),
    .A2(_01461_));
 sg13g2_mux2_1 _06935_ (.A0(_01692_),
    .A1(_01694_),
    .S(net2363),
    .X(_01695_));
 sg13g2_nand2_1 _06936_ (.Y(_01696_),
    .A(net2395),
    .B(_01695_));
 sg13g2_nand3_1 _06937_ (.B(net2317),
    .C(_01695_),
    .A(net2395),
    .Y(_01697_));
 sg13g2_a21oi_1 _06938_ (.A1(_01307_),
    .A2(net2476),
    .Y(_01698_),
    .B1(net2491));
 sg13g2_nand3_1 _06939_ (.B(_01697_),
    .C(_01698_),
    .A(_01690_),
    .Y(_01699_));
 sg13g2_o21ai_1 _06940_ (.B1(_01307_),
    .Y(_01700_),
    .A1(_01314_),
    .A2(_01631_));
 sg13g2_and2_1 _06941_ (.A(_01632_),
    .B(_01700_),
    .X(_01701_));
 sg13g2_o21ai_1 _06942_ (.B1(_01699_),
    .Y(_01702_),
    .A1(net2489),
    .A2(_01701_));
 sg13g2_nor3_1 _06943_ (.A(_01307_),
    .B(_01311_),
    .C(_01364_),
    .Y(_01703_));
 sg13g2_nor2_1 _06944_ (.A(net2496),
    .B(_01703_),
    .Y(_01704_));
 sg13g2_a21oi_1 _06945_ (.A1(_01365_),
    .A2(_01704_),
    .Y(_01705_),
    .B1(net2635));
 sg13g2_a22oi_1 _06946_ (.Y(_01706_),
    .B1(_01702_),
    .B2(_01705_),
    .A2(net2635),
    .A1(_00037_));
 sg13g2_xor2_1 _06947_ (.B(_01525_),
    .A(_01508_),
    .X(_01707_));
 sg13g2_a21oi_1 _06948_ (.A1(net2625),
    .A2(_01707_),
    .Y(_01708_),
    .B1(net2171));
 sg13g2_o21ai_1 _06949_ (.B1(_01708_),
    .Y(_01709_),
    .A1(net2625),
    .A2(_01706_));
 sg13g2_nand3_1 _06950_ (.B(net2501),
    .C(_01229_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][6] ),
    .Y(_01710_));
 sg13g2_nand3_1 _06951_ (.B(net2501),
    .C(_01231_),
    .A(\ChiselTop.wild.dmem.MEM_3[0][6] ),
    .Y(_01711_));
 sg13g2_a21oi_1 _06952_ (.A1(_01710_),
    .A2(_01711_),
    .Y(_01712_),
    .B1(_01176_));
 sg13g2_nor2_2 _06953_ (.A(_01223_),
    .B(_01225_),
    .Y(_01713_));
 sg13g2_a22oi_1 _06954_ (.Y(_01714_),
    .B1(net2448),
    .B2(\ChiselTop.wild.rx._shiftReg_T_1[5] ),
    .A2(net2506),
    .A1(\ChiselTop.wild.dmem.MEM[0][6] ));
 sg13g2_nand3_1 _06955_ (.B(net2502),
    .C(_01642_),
    .A(\ChiselTop.wild.dmem.MEM_2[0][6] ),
    .Y(_01715_));
 sg13g2_o21ai_1 _06956_ (.B1(_01715_),
    .Y(_01716_),
    .A1(_01713_),
    .A2(_01714_));
 sg13g2_o21ai_1 _06957_ (.B1(net2183),
    .Y(_01717_),
    .A1(_01712_),
    .A2(_01716_));
 sg13g2_nand2_1 _06958_ (.Y(_01718_),
    .A(_01709_),
    .B(_01717_));
 sg13g2_nand2_1 _06959_ (.Y(_01719_),
    .A(_00117_),
    .B(_00978_));
 sg13g2_nor2_1 _06960_ (.A(net2543),
    .B(_01570_),
    .Y(_01720_));
 sg13g2_a22oi_1 _06961_ (.Y(_01721_),
    .B1(_01719_),
    .B2(_01720_),
    .A2(_01718_),
    .A1(net2543));
 sg13g2_mux4_1 _06962_ (.S0(net2689),
    .A0(\ChiselTop.wild.cpu.regs[0][6] ),
    .A1(\ChiselTop.wild.cpu.regs[1][6] ),
    .A2(\ChiselTop.wild.cpu.regs[2][6] ),
    .A3(\ChiselTop.wild.cpu.regs[3][6] ),
    .S1(net2668),
    .X(_01722_));
 sg13g2_nor2_1 _06963_ (.A(net2655),
    .B(_01722_),
    .Y(_01723_));
 sg13g2_nor2b_1 _06964_ (.A(\ChiselTop.wild.cpu.regs[5][6] ),
    .B_N(net2690),
    .Y(_01724_));
 sg13g2_nor2_1 _06965_ (.A(net2689),
    .B(\ChiselTop.wild.cpu.regs[4][6] ),
    .Y(_01725_));
 sg13g2_nor3_1 _06966_ (.A(net2668),
    .B(_01724_),
    .C(_01725_),
    .Y(_01726_));
 sg13g2_nor2b_1 _06967_ (.A(\ChiselTop.wild.cpu.regs[7][6] ),
    .B_N(net2690),
    .Y(_01727_));
 sg13g2_o21ai_1 _06968_ (.B1(net2668),
    .Y(_01728_),
    .A1(net2690),
    .A2(\ChiselTop.wild.cpu.regs[6][6] ));
 sg13g2_o21ai_1 _06969_ (.B1(net2655),
    .Y(_01729_),
    .A1(_01727_),
    .A2(_01728_));
 sg13g2_o21ai_1 _06970_ (.B1(net2467),
    .Y(_01730_),
    .A1(_01726_),
    .A2(_01729_));
 sg13g2_nor2_1 _06971_ (.A(_01723_),
    .B(_01730_),
    .Y(_01731_));
 sg13g2_nor2_1 _06972_ (.A(net2442),
    .B(_01731_),
    .Y(_01732_));
 sg13g2_a21oi_1 _06973_ (.A1(net2441),
    .A2(net2144),
    .Y(_01733_),
    .B1(_01732_));
 sg13g2_o21ai_1 _06974_ (.B1(_01569_),
    .Y(_01734_),
    .A1(_01663_),
    .A2(_01733_));
 sg13g2_inv_1 _06975_ (.Y(_01735_),
    .A(_01734_));
 sg13g2_a21oi_2 _06976_ (.B1(_01569_),
    .Y(_01736_),
    .A2(_01733_),
    .A1(_01663_));
 sg13g2_inv_1 _06977_ (.Y(_01737_),
    .A(_01736_));
 sg13g2_nand2_2 _06978_ (.Y(_01738_),
    .A(net1528),
    .B(net2523));
 sg13g2_xor2_1 _06979_ (.B(_00977_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[5] ),
    .X(_01739_));
 sg13g2_nand2_1 _06980_ (.Y(_01740_),
    .A(_01316_),
    .B(net2475));
 sg13g2_mux4_1 _06981_ (.S0(net2329),
    .A0(_01064_),
    .A1(net2424),
    .A2(net2421),
    .A3(net2417),
    .S1(net2343),
    .X(_01741_));
 sg13g2_mux2_1 _06982_ (.A0(_01580_),
    .A1(_01583_),
    .S(net2350),
    .X(_01742_));
 sg13g2_mux2_1 _06983_ (.A0(_01741_),
    .A1(_01742_),
    .S(net2356),
    .X(_01743_));
 sg13g2_o21ai_1 _06984_ (.B1(_01673_),
    .Y(_01744_),
    .A1(net2354),
    .A2(_01582_));
 sg13g2_nand2_1 _06985_ (.Y(_01745_),
    .A(net2366),
    .B(_01744_));
 sg13g2_a21oi_2 _06986_ (.B1(net2390),
    .Y(_01746_),
    .A2(net2358),
    .A1(net2431));
 sg13g2_inv_1 _06987_ (.Y(_01747_),
    .A(_01746_));
 sg13g2_a22oi_1 _06988_ (.Y(_01748_),
    .B1(_01745_),
    .B2(_01746_),
    .A2(_01743_),
    .A1(net2385));
 sg13g2_nand2_1 _06989_ (.Y(_01749_),
    .A(_01449_),
    .B(_01748_));
 sg13g2_mux2_1 _06990_ (.A0(_01594_),
    .A1(_01598_),
    .S(net2342),
    .X(_01750_));
 sg13g2_a21oi_1 _06991_ (.A1(net2435),
    .A2(net2333),
    .Y(_01751_),
    .B1(_01616_));
 sg13g2_mux4_1 _06992_ (.S0(net2345),
    .A0(_01172_),
    .A1(_01037_),
    .A2(net2436),
    .A3(net2435),
    .S1(net2330),
    .X(_01752_));
 sg13g2_mux2_1 _06993_ (.A0(_01593_),
    .A1(_01603_),
    .S(net2350),
    .X(_01753_));
 sg13g2_and2_1 _06994_ (.A(net2365),
    .B(_01753_),
    .X(_01754_));
 sg13g2_mux4_1 _06995_ (.S0(net2329),
    .A0(net2437),
    .A1(net2426),
    .A2(net2415),
    .A3(net2430),
    .S1(net2343),
    .X(_01755_));
 sg13g2_a21oi_1 _06996_ (.A1(net2356),
    .A2(_01755_),
    .Y(_01756_),
    .B1(_01754_));
 sg13g2_mux4_1 _06997_ (.S0(net2365),
    .A0(_01750_),
    .A1(_01752_),
    .A2(_01755_),
    .A3(_01753_),
    .S1(net2375),
    .X(_01757_));
 sg13g2_nand3_1 _06998_ (.B(net2354),
    .C(net2338),
    .A(net2431),
    .Y(_01758_));
 sg13g2_o21ai_1 _06999_ (.B1(_01758_),
    .Y(_01759_),
    .A1(net2352),
    .A2(_01582_));
 sg13g2_a21oi_1 _07000_ (.A1(net2366),
    .A2(_01759_),
    .Y(_01760_),
    .B1(net2385));
 sg13g2_a21oi_1 _07001_ (.A1(net2385),
    .A2(_01743_),
    .Y(_01761_),
    .B1(_01760_));
 sg13g2_o21ai_1 _07002_ (.B1(net2481),
    .Y(_01762_),
    .A1(_01457_),
    .A2(_01761_));
 sg13g2_a221oi_1 _07003_ (.B2(net2397),
    .C1(_01762_),
    .B1(_01757_),
    .A1(net2319),
    .Y(_01763_),
    .A2(_01749_));
 sg13g2_nand3b_1 _07004_ (.B(net2346),
    .C(net2360),
    .Y(_01764_),
    .A_N(_01621_));
 sg13g2_nor2_1 _07005_ (.A(net2346),
    .B(_01619_),
    .Y(_01765_));
 sg13g2_a21oi_1 _07006_ (.A1(net2346),
    .A2(_01615_),
    .Y(_01766_),
    .B1(_01765_));
 sg13g2_o21ai_1 _07007_ (.B1(_01764_),
    .Y(_01767_),
    .A1(net2360),
    .A2(_01766_));
 sg13g2_nand2_1 _07008_ (.Y(_01768_),
    .A(net2388),
    .B(_01767_));
 sg13g2_o21ai_1 _07009_ (.B1(net2471),
    .Y(_01769_),
    .A1(net2314),
    .A2(_01768_));
 sg13g2_o21ai_1 _07010_ (.B1(_01740_),
    .Y(_01770_),
    .A1(_01763_),
    .A2(_01769_));
 sg13g2_nand3_1 _07011_ (.B(_01321_),
    .C(_01363_),
    .A(_01316_),
    .Y(_01771_));
 sg13g2_nand2b_1 _07012_ (.Y(_01772_),
    .B(_01771_),
    .A_N(_01364_));
 sg13g2_xor2_1 _07013_ (.B(_01630_),
    .A(_01316_),
    .X(_01773_));
 sg13g2_o21ai_1 _07014_ (.B1(net2530),
    .Y(_01774_),
    .A1(net2488),
    .A2(_01773_));
 sg13g2_a221oi_1 _07015_ (.B2(net2498),
    .C1(_01774_),
    .B1(_01772_),
    .A1(_01386_),
    .Y(_01775_),
    .A2(_01770_));
 sg13g2_a21oi_1 _07016_ (.A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[5] ),
    .A2(net2638),
    .Y(_01776_),
    .B1(net2628));
 sg13g2_nand2b_1 _07017_ (.Y(_01777_),
    .B(_01776_),
    .A_N(_01775_));
 sg13g2_xnor2_1 _07018_ (.Y(_01778_),
    .A(_01523_),
    .B(_01524_));
 sg13g2_a21oi_1 _07019_ (.A1(net2627),
    .A2(_01778_),
    .Y(_01779_),
    .B1(net2622));
 sg13g2_a221oi_1 _07020_ (.B2(_01779_),
    .C1(net2186),
    .B1(_01777_),
    .A1(net2622),
    .Y(_01780_),
    .A2(\ChiselTop.wild.cpu.decExReg_csrVal[3] ));
 sg13g2_nand3_1 _07021_ (.B(net2502),
    .C(_01229_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][5] ),
    .Y(_01781_));
 sg13g2_nand2_2 _07022_ (.Y(_01782_),
    .A(\ChiselTop.wild.dmem.MEM_3[0][5] ),
    .B(net2505));
 sg13g2_o21ai_1 _07023_ (.B1(_01781_),
    .Y(_01783_),
    .A1(_01232_),
    .A2(_01782_));
 sg13g2_nand3_1 _07024_ (.B(net2505),
    .C(_01642_),
    .A(\ChiselTop.wild.dmem.MEM_2[0][5] ),
    .Y(_01784_));
 sg13g2_a22oi_1 _07025_ (.Y(_01785_),
    .B1(net2448),
    .B2(\ChiselTop.wild.rx._shiftReg_T_1[4] ),
    .A2(net2507),
    .A1(\ChiselTop.wild.dmem.MEM[0][5] ));
 sg13g2_o21ai_1 _07026_ (.B1(_01784_),
    .Y(_01786_),
    .A1(_01713_),
    .A2(_01785_));
 sg13g2_a21oi_1 _07027_ (.A1(net2525),
    .A2(_01783_),
    .Y(_01787_),
    .B1(_01786_));
 sg13g2_a21o_1 _07028_ (.A2(_01787_),
    .A1(net2186),
    .B1(_01780_),
    .X(_01788_));
 sg13g2_mux2_2 _07029_ (.A0(_01739_),
    .A1(_01788_),
    .S(net2547),
    .X(_01789_));
 sg13g2_nand2_1 _07030_ (.Y(_01790_),
    .A(net2445),
    .B(_01789_));
 sg13g2_mux4_1 _07031_ (.S0(net2694),
    .A0(\ChiselTop.wild.cpu.regs[0][5] ),
    .A1(\ChiselTop.wild.cpu.regs[1][5] ),
    .A2(\ChiselTop.wild.cpu.regs[2][5] ),
    .A3(\ChiselTop.wild.cpu.regs[3][5] ),
    .S1(net2671),
    .X(_01791_));
 sg13g2_nor2_1 _07032_ (.A(net2659),
    .B(_01791_),
    .Y(_01792_));
 sg13g2_nor2b_1 _07033_ (.A(\ChiselTop.wild.cpu.regs[5][5] ),
    .B_N(net2694),
    .Y(_01793_));
 sg13g2_nor2_1 _07034_ (.A(net2694),
    .B(\ChiselTop.wild.cpu.regs[4][5] ),
    .Y(_01794_));
 sg13g2_nor3_1 _07035_ (.A(net2670),
    .B(_01793_),
    .C(_01794_),
    .Y(_01795_));
 sg13g2_nor2b_1 _07036_ (.A(\ChiselTop.wild.cpu.regs[7][5] ),
    .B_N(net2697),
    .Y(_01796_));
 sg13g2_o21ai_1 _07037_ (.B1(net2673),
    .Y(_01797_),
    .A1(net2697),
    .A2(\ChiselTop.wild.cpu.regs[6][5] ));
 sg13g2_o21ai_1 _07038_ (.B1(net2657),
    .Y(_01798_),
    .A1(_01796_),
    .A2(_01797_));
 sg13g2_o21ai_1 _07039_ (.B1(net2469),
    .Y(_01799_),
    .A1(_01795_),
    .A2(_01798_));
 sg13g2_nor2_1 _07040_ (.A(_01792_),
    .B(_01799_),
    .Y(_01800_));
 sg13g2_o21ai_1 _07041_ (.B1(_01790_),
    .Y(_01801_),
    .A1(net2445),
    .A2(_01800_));
 sg13g2_nand2_1 _07042_ (.Y(_01802_),
    .A(_01738_),
    .B(_01801_));
 sg13g2_a21o_1 _07043_ (.A2(_01801_),
    .A1(_01738_),
    .B1(_01736_),
    .X(_01803_));
 sg13g2_nand2_1 _07044_ (.Y(_01804_),
    .A(\ChiselTop.wild.cpu.decOut_opcode[5] ),
    .B(net2551));
 sg13g2_nor2_1 _07045_ (.A(\ChiselTop.wild.cpu.decOut_opcode[4] ),
    .B(_01804_),
    .Y(_01805_));
 sg13g2_nor2b_2 _07046_ (.A(\ChiselTop.wild.cpu.decOut_opcode[2] ),
    .B_N(\ChiselTop.wild.cpu.decOut_opcode[4] ),
    .Y(_01806_));
 sg13g2_nor2_1 _07047_ (.A(\ChiselTop.wild.cpu.decOut_opcode[5] ),
    .B(net2551),
    .Y(_01807_));
 sg13g2_a22oi_1 _07048_ (.Y(_01808_),
    .B1(_01806_),
    .B2(_01807_),
    .A2(_01805_),
    .A1(net1534));
 sg13g2_nor2b_1 _07049_ (.A(_01804_),
    .B_N(_01806_),
    .Y(_01809_));
 sg13g2_nor2_1 _07050_ (.A(\ChiselTop.wild.cpu.decOut_opcode[4] ),
    .B(\ChiselTop.wild.cpu.decOut_opcode[2] ),
    .Y(_01810_));
 sg13g2_and2_1 _07051_ (.A(_01807_),
    .B(_01810_),
    .X(_01811_));
 sg13g2_nor2_1 _07052_ (.A(_01809_),
    .B(_01811_),
    .Y(_01812_));
 sg13g2_nand2_2 _07053_ (.Y(_01813_),
    .A(_01808_),
    .B(_01812_));
 sg13g2_nand2_1 _07054_ (.Y(_01814_),
    .A(net1518),
    .B(_01813_));
 sg13g2_and2_1 _07055_ (.A(\ChiselTop.wild.cpu.decOut_opcode[5] ),
    .B(_01810_),
    .X(_01815_));
 sg13g2_nand2_2 _07056_ (.Y(_01816_),
    .A(\ChiselTop.wild.cpu.decOut_opcode[5] ),
    .B(_01810_));
 sg13g2_a21oi_1 _07057_ (.A1(\ChiselTop.wild.cpu._GEN_176[2] ),
    .A2(net2523),
    .Y(_01817_),
    .B1(net2465));
 sg13g2_a21oi_1 _07058_ (.A1(_00114_),
    .A2(net2465),
    .Y(_01818_),
    .B1(_01817_));
 sg13g2_o21ai_1 _07059_ (.B1(_01814_),
    .Y(_01819_),
    .A1(_01813_),
    .A2(_01818_));
 sg13g2_inv_1 _07060_ (.Y(_01820_),
    .A(_01819_));
 sg13g2_a21o_1 _07061_ (.A2(\ChiselTop.wild.cpu.decExReg_pc[2] ),
    .A1(\ChiselTop.wild.cpu.decExReg_pc[3] ),
    .B1(\ChiselTop.wild.cpu.decExReg_pc[4] ),
    .X(_01821_));
 sg13g2_nand3_1 _07062_ (.B(net2502),
    .C(_01229_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][4] ),
    .Y(_01822_));
 sg13g2_nand2_2 _07063_ (.Y(_01823_),
    .A(\ChiselTop.wild.dmem.MEM_3[0][4] ),
    .B(net2504));
 sg13g2_o21ai_1 _07064_ (.B1(_01822_),
    .Y(_01824_),
    .A1(_01232_),
    .A2(_01823_));
 sg13g2_nand3_1 _07065_ (.B(net2505),
    .C(_01642_),
    .A(\ChiselTop.wild.dmem.MEM_2[0][4] ),
    .Y(_01825_));
 sg13g2_a22oi_1 _07066_ (.Y(_01826_),
    .B1(_01226_),
    .B2(\ChiselTop.wild.rx._shiftReg_T_1[3] ),
    .A2(net2507),
    .A1(\ChiselTop.wild.dmem.MEM[0][4] ));
 sg13g2_o21ai_1 _07067_ (.B1(_01825_),
    .Y(_01827_),
    .A1(_01713_),
    .A2(_01826_));
 sg13g2_a21oi_1 _07068_ (.A1(net2525),
    .A2(_01824_),
    .Y(_01828_),
    .B1(_01827_));
 sg13g2_nand2b_1 _07069_ (.Y(_01829_),
    .B(net2186),
    .A_N(_01828_));
 sg13g2_nor3_1 _07070_ (.A(net2640),
    .B(_01361_),
    .C(_01362_),
    .Y(_01830_));
 sg13g2_a21oi_1 _07071_ (.A1(net2640),
    .A2(_01628_),
    .Y(_01831_),
    .B1(_01830_));
 sg13g2_o21ai_1 _07072_ (.B1(_01385_),
    .Y(_01832_),
    .A1(_01324_),
    .A2(_01831_));
 sg13g2_a21oi_1 _07073_ (.A1(_01324_),
    .A2(_01831_),
    .Y(_01833_),
    .B1(_01832_));
 sg13g2_mux2_1 _07074_ (.A0(_01430_),
    .A1(_01442_),
    .S(net2370),
    .X(_01834_));
 sg13g2_nand2_1 _07075_ (.Y(_01835_),
    .A(net2392),
    .B(_01834_));
 sg13g2_and2_1 _07076_ (.A(net2370),
    .B(_01437_),
    .X(_01836_));
 sg13g2_o21ai_1 _07077_ (.B1(_01835_),
    .Y(_01837_),
    .A1(net2391),
    .A2(_01836_));
 sg13g2_inv_1 _07078_ (.Y(_01838_),
    .A(_01837_));
 sg13g2_o21ai_1 _07079_ (.B1(_01835_),
    .Y(_01839_),
    .A1(_01747_),
    .A2(_01836_));
 sg13g2_o21ai_1 _07080_ (.B1(net2320),
    .Y(_01840_),
    .A1(net2480),
    .A2(_01839_));
 sg13g2_mux4_1 _07081_ (.S0(net2349),
    .A0(_01093_),
    .A1(net2420),
    .A2(net2433),
    .A3(_01172_),
    .S1(net2338),
    .X(_01841_));
 sg13g2_nor2_1 _07082_ (.A(net2371),
    .B(_01841_),
    .Y(_01842_));
 sg13g2_nand3_1 _07083_ (.B(_01466_),
    .C(_01467_),
    .A(net2353),
    .Y(_01843_));
 sg13g2_nand3_1 _07084_ (.B(_01462_),
    .C(_01465_),
    .A(net2348),
    .Y(_01844_));
 sg13g2_and2_1 _07085_ (.A(_01843_),
    .B(_01844_),
    .X(_01845_));
 sg13g2_o21ai_1 _07086_ (.B1(net2393),
    .Y(_01846_),
    .A1(net2359),
    .A2(_01845_));
 sg13g2_mux4_1 _07087_ (.S0(net2338),
    .A0(_01047_),
    .A1(net2428),
    .A2(_01131_),
    .A3(_01104_),
    .S1(net2354),
    .X(_01847_));
 sg13g2_mux2_1 _07088_ (.A0(_01440_),
    .A1(_01847_),
    .S(net2370),
    .X(_01848_));
 sg13g2_nand2_1 _07089_ (.Y(_01849_),
    .A(net2381),
    .B(_01848_));
 sg13g2_o21ai_1 _07090_ (.B1(_01849_),
    .Y(_01850_),
    .A1(_01842_),
    .A2(_01846_));
 sg13g2_a221oi_1 _07091_ (.B2(net2399),
    .C1(net2485),
    .B1(_01850_),
    .A1(net2318),
    .Y(_01851_),
    .A2(_01837_));
 sg13g2_a21oi_1 _07092_ (.A1(_01325_),
    .A2(net2476),
    .Y(_01852_),
    .B1(_01385_));
 sg13g2_mux2_1 _07093_ (.A0(_01464_),
    .A1(_01487_),
    .S(net2363),
    .X(_01853_));
 sg13g2_nand2b_1 _07094_ (.Y(_01854_),
    .B(net2395),
    .A_N(_01853_));
 sg13g2_o21ai_1 _07095_ (.B1(_01852_),
    .Y(_01855_),
    .A1(net2315),
    .A2(_01854_));
 sg13g2_a21oi_2 _07096_ (.B1(_01855_),
    .Y(_01856_),
    .A2(_01851_),
    .A1(_01840_));
 sg13g2_nor3_2 _07097_ (.A(net2635),
    .B(_01833_),
    .C(_01856_),
    .Y(_01857_));
 sg13g2_o21ai_1 _07098_ (.B1(net2529),
    .Y(_01858_),
    .A1(net2531),
    .A2(_00118_));
 sg13g2_xnor2_1 _07099_ (.Y(_01859_),
    .A(_01511_),
    .B(_01522_));
 sg13g2_and2_1 _07100_ (.A(net2628),
    .B(_01859_),
    .X(_01860_));
 sg13g2_o21ai_1 _07101_ (.B1(_01547_),
    .Y(_01861_),
    .A1(_01857_),
    .A2(_01858_));
 sg13g2_o21ai_1 _07102_ (.B1(_01829_),
    .Y(_01862_),
    .A1(_01860_),
    .A2(_01861_));
 sg13g2_and2_1 _07103_ (.A(net2616),
    .B(_00977_),
    .X(_01863_));
 sg13g2_a22oi_1 _07104_ (.Y(_01864_),
    .B1(_01863_),
    .B2(_01821_),
    .A2(_01862_),
    .A1(net2548));
 sg13g2_mux4_1 _07105_ (.S0(net2697),
    .A0(\ChiselTop.wild.cpu.regs[0][4] ),
    .A1(\ChiselTop.wild.cpu.regs[1][4] ),
    .A2(\ChiselTop.wild.cpu.regs[2][4] ),
    .A3(\ChiselTop.wild.cpu.regs[3][4] ),
    .S1(net2673),
    .X(_01865_));
 sg13g2_nor2_2 _07106_ (.A(net2658),
    .B(_01865_),
    .Y(_01866_));
 sg13g2_nor2b_1 _07107_ (.A(\ChiselTop.wild.cpu.regs[5][4] ),
    .B_N(net2695),
    .Y(_01867_));
 sg13g2_nor2_1 _07108_ (.A(net2696),
    .B(\ChiselTop.wild.cpu.regs[4][4] ),
    .Y(_01868_));
 sg13g2_nor3_1 _07109_ (.A(net2672),
    .B(_01867_),
    .C(_01868_),
    .Y(_01869_));
 sg13g2_nor2b_1 _07110_ (.A(\ChiselTop.wild.cpu.regs[7][4] ),
    .B_N(net2695),
    .Y(_01870_));
 sg13g2_o21ai_1 _07111_ (.B1(net2672),
    .Y(_01871_),
    .A1(net2695),
    .A2(\ChiselTop.wild.cpu.regs[6][4] ));
 sg13g2_o21ai_1 _07112_ (.B1(net2657),
    .Y(_01872_),
    .A1(_01870_),
    .A2(_01871_));
 sg13g2_o21ai_1 _07113_ (.B1(net2468),
    .Y(_01873_),
    .A1(_01869_),
    .A2(_01872_));
 sg13g2_nor2_1 _07114_ (.A(_01866_),
    .B(_01873_),
    .Y(_01874_));
 sg13g2_nor2_1 _07115_ (.A(net2445),
    .B(_01874_),
    .Y(_01875_));
 sg13g2_a21oi_1 _07116_ (.A1(net2445),
    .A2(net2152),
    .Y(_01876_),
    .B1(_01875_));
 sg13g2_nand2_1 _07117_ (.Y(_01877_),
    .A(_01820_),
    .B(_01876_));
 sg13g2_o21ai_1 _07118_ (.B1(_01877_),
    .Y(_01878_),
    .A1(_01738_),
    .A2(_01801_));
 sg13g2_a21oi_1 _07119_ (.A1(_00122_),
    .A2(net2465),
    .Y(_01879_),
    .B1(_01817_));
 sg13g2_o21ai_1 _07120_ (.B1(_01814_),
    .Y(_01880_),
    .A1(_01813_),
    .A2(_01879_));
 sg13g2_nand2b_1 _07121_ (.Y(_01881_),
    .B(net2638),
    .A_N(\ChiselTop.wild.cpu.decExReg_decOut_imm[2] ));
 sg13g2_mux2_1 _07122_ (.A0(_01664_),
    .A1(_01686_),
    .S(net2371),
    .X(_01882_));
 sg13g2_nand2_1 _07123_ (.Y(_01883_),
    .A(net2390),
    .B(_01882_));
 sg13g2_inv_1 _07124_ (.Y(_01884_),
    .A(_01883_));
 sg13g2_and2_1 _07125_ (.A(net2371),
    .B(_01665_),
    .X(_01885_));
 sg13g2_a21o_1 _07126_ (.A2(_01669_),
    .A1(net2358),
    .B1(_01885_),
    .X(_01886_));
 sg13g2_inv_1 _07127_ (.Y(_01887_),
    .A(_01886_));
 sg13g2_a21oi_1 _07128_ (.A1(net2381),
    .A2(_01886_),
    .Y(_01888_),
    .B1(_01884_));
 sg13g2_o21ai_1 _07129_ (.B1(_01883_),
    .Y(_01889_),
    .A1(net2390),
    .A2(_01887_));
 sg13g2_o21ai_1 _07130_ (.B1(_01886_),
    .Y(_01890_),
    .A1(_01673_),
    .A2(_01885_));
 sg13g2_o21ai_1 _07131_ (.B1(_01883_),
    .Y(_01891_),
    .A1(net2390),
    .A2(_01890_));
 sg13g2_o21ai_1 _07132_ (.B1(net2319),
    .Y(_01892_),
    .A1(net2480),
    .A2(_01891_));
 sg13g2_a21oi_1 _07133_ (.A1(_01462_),
    .A2(_01465_),
    .Y(_01893_),
    .B1(net2348));
 sg13g2_mux2_1 _07134_ (.A0(_01119_),
    .A1(_01025_),
    .S(net2339),
    .X(_01894_));
 sg13g2_nor2_1 _07135_ (.A(net2353),
    .B(_01894_),
    .Y(_01895_));
 sg13g2_nand2_1 _07136_ (.Y(_01896_),
    .A(net2359),
    .B(_01679_));
 sg13g2_or2_1 _07137_ (.X(_01897_),
    .B(_01895_),
    .A(_01893_));
 sg13g2_a21oi_1 _07138_ (.A1(net2371),
    .A2(_01897_),
    .Y(_01898_),
    .B1(net2381));
 sg13g2_and2_1 _07139_ (.A(net2370),
    .B(_01681_),
    .X(_01899_));
 sg13g2_a21oi_1 _07140_ (.A1(net2358),
    .A2(_01684_),
    .Y(_01900_),
    .B1(_01899_));
 sg13g2_a22oi_1 _07141_ (.Y(_01901_),
    .B1(_01900_),
    .B2(net2381),
    .A2(_01898_),
    .A1(_01896_));
 sg13g2_a221oi_1 _07142_ (.B2(net2399),
    .C1(net2485),
    .B1(_01901_),
    .A1(net2318),
    .Y(_01902_),
    .A2(_01889_));
 sg13g2_nand2_1 _07143_ (.Y(_01903_),
    .A(net2372),
    .B(_01694_));
 sg13g2_nor2_1 _07144_ (.A(net2382),
    .B(_01903_),
    .Y(_01904_));
 sg13g2_a221oi_1 _07145_ (.B2(net2316),
    .C1(net2474),
    .B1(_01904_),
    .A1(_01892_),
    .Y(_01905_),
    .A2(_01902_));
 sg13g2_o21ai_1 _07146_ (.B1(net2488),
    .Y(_01906_),
    .A1(_01339_),
    .A2(net2472));
 sg13g2_a21oi_1 _07147_ (.A1(_01338_),
    .A2(_01358_),
    .Y(_01907_),
    .B1(net2495));
 sg13g2_a21oi_1 _07148_ (.A1(_01349_),
    .A2(_01394_),
    .Y(_01908_),
    .B1(_01347_));
 sg13g2_nor2_1 _07149_ (.A(_01339_),
    .B(_01908_),
    .Y(_01909_));
 sg13g2_xnor2_1 _07150_ (.Y(_01910_),
    .A(_01338_),
    .B(_01908_));
 sg13g2_a221oi_1 _07151_ (.B2(net2490),
    .C1(net2634),
    .B1(_01910_),
    .A1(_01359_),
    .Y(_01911_),
    .A2(_01907_));
 sg13g2_o21ai_1 _07152_ (.B1(_01911_),
    .Y(_01912_),
    .A1(_01905_),
    .A2(_01906_));
 sg13g2_xnor2_1 _07153_ (.Y(_01913_),
    .A(_01515_),
    .B(_01519_));
 sg13g2_nand3_1 _07154_ (.B(_01881_),
    .C(_01912_),
    .A(_00925_),
    .Y(_01914_));
 sg13g2_nand2_1 _07155_ (.Y(_01915_),
    .A(net2628),
    .B(_01913_));
 sg13g2_a21o_1 _07156_ (.A2(_01915_),
    .A1(_01914_),
    .B1(\ChiselTop.wild.cpu.decExReg_decOut_isCssrw ),
    .X(_01916_));
 sg13g2_a21oi_1 _07157_ (.A1(net2622),
    .A2(\ChiselTop.wild.cpu.decExReg_csrVal[2] ),
    .Y(_01917_),
    .B1(net2187));
 sg13g2_a22oi_1 _07158_ (.Y(_01918_),
    .B1(net2448),
    .B2(\ChiselTop.wild.rx._shiftReg_T_1[1] ),
    .A2(net2506),
    .A1(\ChiselTop.wild.dmem.MEM[0][2] ));
 sg13g2_nor2_1 _07159_ (.A(_01713_),
    .B(_01918_),
    .Y(_01919_));
 sg13g2_and2_1 _07160_ (.A(\ChiselTop.wild.dmem.MEM_2[0][2] ),
    .B(net2500),
    .X(_01920_));
 sg13g2_nand3_1 _07161_ (.B(net2504),
    .C(_01229_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][2] ),
    .Y(_01921_));
 sg13g2_nand2_2 _07162_ (.Y(_01922_),
    .A(\ChiselTop.wild.dmem.MEM_3[0][2] ),
    .B(net2505));
 sg13g2_o21ai_1 _07163_ (.B1(_01921_),
    .Y(_01923_),
    .A1(_01232_),
    .A2(_01922_));
 sg13g2_a221oi_1 _07164_ (.B2(net2526),
    .C1(_01919_),
    .B1(_01923_),
    .A1(_01642_),
    .Y(_01924_),
    .A2(_01920_));
 sg13g2_a22oi_1 _07165_ (.Y(_01925_),
    .B1(_01924_),
    .B2(net2187),
    .A2(_01917_),
    .A1(_01916_));
 sg13g2_nand2b_1 _07166_ (.Y(_01926_),
    .B(net2619),
    .A_N(net1538));
 sg13g2_o21ai_1 _07167_ (.B1(_01926_),
    .Y(_01927_),
    .A1(net2617),
    .A2(_01925_));
 sg13g2_mux4_1 _07168_ (.S0(net2697),
    .A0(\ChiselTop.wild.cpu.regs[0][2] ),
    .A1(\ChiselTop.wild.cpu.regs[1][2] ),
    .A2(\ChiselTop.wild.cpu.regs[2][2] ),
    .A3(\ChiselTop.wild.cpu.regs[3][2] ),
    .S1(net2673),
    .X(_01928_));
 sg13g2_nor2_1 _07169_ (.A(net2658),
    .B(_01928_),
    .Y(_01929_));
 sg13g2_nor2b_1 _07170_ (.A(\ChiselTop.wild.cpu.regs[5][2] ),
    .B_N(net2701),
    .Y(_01930_));
 sg13g2_nor2_1 _07171_ (.A(net2701),
    .B(\ChiselTop.wild.cpu.regs[4][2] ),
    .Y(_01931_));
 sg13g2_nor3_1 _07172_ (.A(net2673),
    .B(_01930_),
    .C(_01931_),
    .Y(_01932_));
 sg13g2_nor2b_1 _07173_ (.A(\ChiselTop.wild.cpu.regs[7][2] ),
    .B_N(net2701),
    .Y(_01933_));
 sg13g2_o21ai_1 _07174_ (.B1(net2676),
    .Y(_01934_),
    .A1(net2701),
    .A2(\ChiselTop.wild.cpu.regs[6][2] ));
 sg13g2_o21ai_1 _07175_ (.B1(net2661),
    .Y(_01935_),
    .A1(_01933_),
    .A2(_01934_));
 sg13g2_o21ai_1 _07176_ (.B1(net2468),
    .Y(_01936_),
    .A1(_01932_),
    .A2(_01935_));
 sg13g2_nor2_1 _07177_ (.A(_01929_),
    .B(_01936_),
    .Y(_01937_));
 sg13g2_nor2_1 _07178_ (.A(net2444),
    .B(_01937_),
    .Y(_01938_));
 sg13g2_a21oi_1 _07179_ (.A1(net2446),
    .A2(net2140),
    .Y(_01939_),
    .B1(_01938_));
 sg13g2_nand2b_1 _07180_ (.Y(_01940_),
    .B(_01939_),
    .A_N(_01880_));
 sg13g2_xnor2_1 _07181_ (.Y(_01941_),
    .A(_01880_),
    .B(_01939_));
 sg13g2_mux2_1 _07182_ (.A0(_01741_),
    .A1(_01755_),
    .S(net2365),
    .X(_01942_));
 sg13g2_mux4_1 _07183_ (.S0(net2343),
    .A0(_01054_),
    .A1(_01582_),
    .A2(_01583_),
    .A3(_01580_),
    .S1(net2365),
    .X(_01943_));
 sg13g2_mux2_1 _07184_ (.A0(_01942_),
    .A1(_01943_),
    .S(net2375),
    .X(_01944_));
 sg13g2_o21ai_1 _07185_ (.B1(net2319),
    .Y(_01945_),
    .A1(net2480),
    .A2(_01944_));
 sg13g2_mux2_1 _07186_ (.A0(_01750_),
    .A1(_01753_),
    .S(net2356),
    .X(_01946_));
 sg13g2_nand2_1 _07187_ (.Y(_01947_),
    .A(net2356),
    .B(_01752_));
 sg13g2_a21oi_1 _07188_ (.A1(_01120_),
    .A2(net2333),
    .Y(_01948_),
    .B1(_01614_));
 sg13g2_mux4_1 _07189_ (.S0(net2335),
    .A0(_01024_),
    .A1(net2427),
    .A2(_01078_),
    .A3(_01120_),
    .S1(net2351),
    .X(_01949_));
 sg13g2_a21oi_1 _07190_ (.A1(net2365),
    .A2(_01949_),
    .Y(_01950_),
    .B1(net2376));
 sg13g2_a21oi_1 _07191_ (.A1(_01947_),
    .A2(_01950_),
    .Y(_01951_),
    .B1(net2402));
 sg13g2_o21ai_1 _07192_ (.B1(_01951_),
    .Y(_01952_),
    .A1(net2386),
    .A2(_01946_));
 sg13g2_mux4_1 _07193_ (.S0(net2356),
    .A0(_01580_),
    .A1(_01582_),
    .A2(_01583_),
    .A3(_01589_),
    .S1(net2350),
    .X(_01953_));
 sg13g2_mux2_1 _07194_ (.A0(_01942_),
    .A1(_01953_),
    .S(net2375),
    .X(_01954_));
 sg13g2_inv_1 _07195_ (.Y(_01955_),
    .A(_01954_));
 sg13g2_a21oi_1 _07196_ (.A1(net2318),
    .A2(_01954_),
    .Y(_01956_),
    .B1(net2484));
 sg13g2_nand3_1 _07197_ (.B(_01952_),
    .C(_01956_),
    .A(_01945_),
    .Y(_01957_));
 sg13g2_nor3_1 _07198_ (.A(net2360),
    .B(net2351),
    .C(_01621_),
    .Y(_01958_));
 sg13g2_nand2_1 _07199_ (.Y(_01959_),
    .A(net2388),
    .B(_01958_));
 sg13g2_nor2_1 _07200_ (.A(net2314),
    .B(_01959_),
    .Y(_01960_));
 sg13g2_nor2_1 _07201_ (.A(net2475),
    .B(_01960_),
    .Y(_01961_));
 sg13g2_a221oi_1 _07202_ (.B2(_01961_),
    .C1(net2491),
    .B1(_01957_),
    .A1(_01350_),
    .Y(_01962_),
    .A2(net2475));
 sg13g2_xor2_1 _07203_ (.B(_01394_),
    .A(_01350_),
    .X(_01963_));
 sg13g2_xnor2_1 _07204_ (.Y(_01964_),
    .A(_01350_),
    .B(_01356_));
 sg13g2_a22oi_1 _07205_ (.Y(_01965_),
    .B1(_01964_),
    .B2(net2498),
    .A2(_01963_),
    .A1(net2490));
 sg13g2_nand2_1 _07206_ (.Y(_01966_),
    .A(net2530),
    .B(_01965_));
 sg13g2_a21oi_1 _07207_ (.A1(_00058_),
    .A2(net2634),
    .Y(_01967_),
    .B1(net2626));
 sg13g2_o21ai_1 _07208_ (.B1(_01967_),
    .Y(_01968_),
    .A1(_01962_),
    .A2(_01966_));
 sg13g2_xor2_1 _07209_ (.B(_01518_),
    .A(_01517_),
    .X(_01969_));
 sg13g2_a21oi_1 _07210_ (.A1(net2628),
    .A2(_01969_),
    .Y(_01970_),
    .B1(net2622));
 sg13g2_a221oi_1 _07211_ (.B2(_01970_),
    .C1(net2186),
    .B1(_01968_),
    .A1(net2622),
    .Y(_01971_),
    .A2(net1125));
 sg13g2_nor3_1 _07212_ (.A(\ChiselTop.wild.memAddressReg[2] ),
    .B(\ChiselTop.wild.uartStatusReg[1] ),
    .C(net2506),
    .Y(_01972_));
 sg13g2_a221oi_1 _07213_ (.B2(_00900_),
    .C1(_01972_),
    .B1(net2448),
    .A1(_00932_),
    .Y(_01973_),
    .A2(net2506));
 sg13g2_nand2_2 _07214_ (.Y(_01974_),
    .A(\ChiselTop.wild.dmem.MEM_3[0][1] ),
    .B(net2500));
 sg13g2_nand2_1 _07215_ (.Y(_01975_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][1] ),
    .B(net2500));
 sg13g2_a22oi_1 _07216_ (.Y(_01976_),
    .B1(_01975_),
    .B2(_01229_),
    .A2(_01974_),
    .A1(_01231_));
 sg13g2_inv_1 _07217_ (.Y(_01977_),
    .A(_01976_));
 sg13g2_nand2_2 _07218_ (.Y(_01978_),
    .A(\ChiselTop.wild.dmem.MEM_2[0][1] ),
    .B(net2500));
 sg13g2_nand2_1 _07219_ (.Y(_01979_),
    .A(_01642_),
    .B(_01978_));
 sg13g2_o21ai_1 _07220_ (.B1(_01979_),
    .Y(_01980_),
    .A1(_01713_),
    .A2(_01973_));
 sg13g2_a21oi_1 _07221_ (.A1(net2525),
    .A2(_01977_),
    .Y(_01981_),
    .B1(_01980_));
 sg13g2_a21oi_1 _07222_ (.A1(net2186),
    .A2(_01981_),
    .Y(_01982_),
    .B1(_01971_));
 sg13g2_nor2_1 _07223_ (.A(net2617),
    .B(_01982_),
    .Y(_01983_));
 sg13g2_a21oi_1 _07224_ (.A1(net2617),
    .A2(net1542),
    .Y(_01984_),
    .B1(_01983_));
 sg13g2_mux4_1 _07225_ (.S0(net2703),
    .A0(\ChiselTop.wild.cpu.regs[0][1] ),
    .A1(\ChiselTop.wild.cpu.regs[1][1] ),
    .A2(\ChiselTop.wild.cpu.regs[2][1] ),
    .A3(\ChiselTop.wild.cpu.regs[3][1] ),
    .S1(net2676),
    .X(_01985_));
 sg13g2_nor2_1 _07226_ (.A(net2660),
    .B(_01985_),
    .Y(_01986_));
 sg13g2_nor2b_1 _07227_ (.A(\ChiselTop.wild.cpu.regs[5][1] ),
    .B_N(net2701),
    .Y(_01987_));
 sg13g2_nor2_1 _07228_ (.A(net2703),
    .B(\ChiselTop.wild.cpu.regs[4][1] ),
    .Y(_01988_));
 sg13g2_nor3_1 _07229_ (.A(net2675),
    .B(_01987_),
    .C(_01988_),
    .Y(_01989_));
 sg13g2_nor2b_1 _07230_ (.A(\ChiselTop.wild.cpu.regs[7][1] ),
    .B_N(net2703),
    .Y(_01990_));
 sg13g2_o21ai_1 _07231_ (.B1(net2675),
    .Y(_01991_),
    .A1(net2703),
    .A2(\ChiselTop.wild.cpu.regs[6][1] ));
 sg13g2_o21ai_1 _07232_ (.B1(net2660),
    .Y(_01992_),
    .A1(_01990_),
    .A2(_01991_));
 sg13g2_o21ai_1 _07233_ (.B1(net2469),
    .Y(_01993_),
    .A1(_01989_),
    .A2(_01992_));
 sg13g2_nor2_1 _07234_ (.A(_01986_),
    .B(_01993_),
    .Y(_01994_));
 sg13g2_nor2_1 _07235_ (.A(net2445),
    .B(_01994_),
    .Y(_01995_));
 sg13g2_a21oi_1 _07236_ (.A1(net2445),
    .A2(net2149),
    .Y(_01996_),
    .B1(_01995_));
 sg13g2_nand3_1 _07237_ (.B(net2523),
    .C(_01816_),
    .A(\ChiselTop.wild.cpu._GEN_176[1] ),
    .Y(_01997_));
 sg13g2_o21ai_1 _07238_ (.B1(_01997_),
    .Y(_01998_),
    .A1(_00933_),
    .A2(_01816_));
 sg13g2_and2_1 _07239_ (.A(_01996_),
    .B(_01998_),
    .X(_01999_));
 sg13g2_xor2_1 _07240_ (.B(_01998_),
    .A(_01996_),
    .X(_02000_));
 sg13g2_nor2_2 _07241_ (.A(net2551),
    .B(_01816_),
    .Y(_02001_));
 sg13g2_and2_1 _07242_ (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_1[0] ),
    .B(net2522),
    .X(_02002_));
 sg13g2_a22oi_1 _07243_ (.Y(_02003_),
    .B1(_02002_),
    .B2(_01816_),
    .A2(_02001_),
    .A1(net1214));
 sg13g2_inv_1 _07244_ (.Y(_02004_),
    .A(_02003_));
 sg13g2_mux2_1 _07245_ (.A0(_01841_),
    .A1(_01847_),
    .S(net2359),
    .X(_02005_));
 sg13g2_nand2b_1 _07246_ (.Y(_02006_),
    .B(net2383),
    .A_N(_02005_));
 sg13g2_nand2_1 _07247_ (.Y(_02007_),
    .A(net2359),
    .B(_01845_));
 sg13g2_o21ai_1 _07248_ (.B1(_01487_),
    .Y(_02008_),
    .A1(_01348_),
    .A2(net2340));
 sg13g2_a21oi_1 _07249_ (.A1(net2353),
    .A2(_01894_),
    .Y(_02009_),
    .B1(_02008_));
 sg13g2_a21oi_1 _07250_ (.A1(net2373),
    .A2(_02009_),
    .Y(_02010_),
    .B1(net2382));
 sg13g2_a21oi_1 _07251_ (.A1(_02007_),
    .A2(_02010_),
    .Y(_02011_),
    .B1(net2403));
 sg13g2_nand2_2 _07252_ (.Y(_02012_),
    .A(net2480),
    .B(_01452_));
 sg13g2_a22oi_1 _07253_ (.Y(_02013_),
    .B1(_02006_),
    .B2(_02011_),
    .A2(_01444_),
    .A1(_01319_));
 sg13g2_nand2_1 _07254_ (.Y(_02014_),
    .A(_02012_),
    .B(_02013_));
 sg13g2_nand2_1 _07255_ (.Y(_02015_),
    .A(net2643),
    .B(_00132_));
 sg13g2_o21ai_1 _07256_ (.B1(_02015_),
    .Y(_02016_),
    .A1(net2641),
    .A2(_01017_));
 sg13g2_nand2_1 _07257_ (.Y(_02017_),
    .A(_01015_),
    .B(_02016_));
 sg13g2_xnor2_1 _07258_ (.Y(_02018_),
    .A(net2437),
    .B(_02016_));
 sg13g2_nand2_1 _07259_ (.Y(_02019_),
    .A(net2644),
    .B(_00131_));
 sg13g2_o21ai_1 _07260_ (.B1(_02019_),
    .Y(_02020_),
    .A1(net2642),
    .A2(_01136_));
 sg13g2_nand2b_1 _07261_ (.Y(_02021_),
    .B(_02020_),
    .A_N(net2418));
 sg13g2_nand2b_2 _07262_ (.Y(_02022_),
    .B(net2418),
    .A_N(_02020_));
 sg13g2_xnor2_1 _07263_ (.Y(_02023_),
    .A(net2417),
    .B(_02020_));
 sg13g2_and2_1 _07264_ (.A(net2312),
    .B(net2311),
    .X(_02024_));
 sg13g2_nand2_1 _07265_ (.Y(_02025_),
    .A(_02018_),
    .B(_02023_));
 sg13g2_and2_1 _07266_ (.A(net2643),
    .B(_00130_),
    .X(_02026_));
 sg13g2_nand2_1 _07267_ (.Y(_02027_),
    .A(net2643),
    .B(_00130_));
 sg13g2_a21oi_2 _07268_ (.B1(_02026_),
    .Y(_02028_),
    .A2(_01106_),
    .A1(net2533));
 sg13g2_and2_1 _07269_ (.A(net2421),
    .B(_02028_),
    .X(_02029_));
 sg13g2_nor2_1 _07270_ (.A(_01105_),
    .B(_02028_),
    .Y(_02030_));
 sg13g2_xnor2_1 _07271_ (.Y(_02031_),
    .A(net2421),
    .B(_02028_));
 sg13g2_inv_1 _07272_ (.Y(_02032_),
    .A(_02031_));
 sg13g2_o21ai_1 _07273_ (.B1(_02027_),
    .Y(_02033_),
    .A1(net2641),
    .A2(_01087_));
 sg13g2_nor2b_1 _07274_ (.A(_02033_),
    .B_N(net2424),
    .Y(_02034_));
 sg13g2_nand2b_1 _07275_ (.Y(_02035_),
    .B(_02033_),
    .A_N(net2424));
 sg13g2_xnor2_1 _07276_ (.Y(_02036_),
    .A(net2425),
    .B(_02033_));
 sg13g2_inv_1 _07277_ (.Y(_02037_),
    .A(_02036_));
 sg13g2_nand2b_1 _07278_ (.Y(_02038_),
    .B(_02036_),
    .A_N(_02031_));
 sg13g2_nor3_2 _07279_ (.A(net2642),
    .B(_01161_),
    .C(_01162_),
    .Y(_02039_));
 sg13g2_nor2_2 _07280_ (.A(_01253_),
    .B(_02039_),
    .Y(_02040_));
 sg13g2_nor2_1 _07281_ (.A(net2415),
    .B(_02040_),
    .Y(_02041_));
 sg13g2_o21ai_1 _07282_ (.B1(_01159_),
    .Y(_02042_),
    .A1(_01253_),
    .A2(_02039_));
 sg13g2_xnor2_1 _07283_ (.Y(_02043_),
    .A(_01159_),
    .B(_02040_));
 sg13g2_xnor2_1 _07284_ (.Y(_02044_),
    .A(net2415),
    .B(_02040_));
 sg13g2_a21oi_2 _07285_ (.B1(_01253_),
    .Y(_02045_),
    .A2(_01083_),
    .A1(net2533));
 sg13g2_and2_1 _07286_ (.A(net2426),
    .B(_02045_),
    .X(_02046_));
 sg13g2_or2_2 _07287_ (.X(_02047_),
    .B(_02045_),
    .A(net2426));
 sg13g2_nand2b_2 _07288_ (.Y(_02048_),
    .B(_02047_),
    .A_N(_02046_));
 sg13g2_inv_1 _07289_ (.Y(_02049_),
    .A(_02048_));
 sg13g2_nor4_1 _07290_ (.A(_02025_),
    .B(_02038_),
    .C(_02044_),
    .D(_02048_),
    .Y(_02050_));
 sg13g2_or4_1 _07291_ (.A(_02025_),
    .B(_02038_),
    .C(_02044_),
    .D(_02048_),
    .X(_02051_));
 sg13g2_o21ai_1 _07292_ (.B1(_02027_),
    .Y(_02052_),
    .A1(net2643),
    .A2(_01066_));
 sg13g2_a221oi_1 _07293_ (.B2(net2533),
    .C1(_02026_),
    .B1(_01067_),
    .A1(_01061_),
    .Y(_02053_),
    .A2(_01062_));
 sg13g2_nand2_1 _07294_ (.Y(_02054_),
    .A(_01063_),
    .B(_02052_));
 sg13g2_nor2b_1 _07295_ (.A(_02053_),
    .B_N(_02054_),
    .Y(_02055_));
 sg13g2_xnor2_1 _07296_ (.Y(_02056_),
    .A(_01063_),
    .B(_02052_));
 sg13g2_and2_2 _07297_ (.A(net2644),
    .B(_00127_),
    .X(_02057_));
 sg13g2_nand2_1 _07298_ (.Y(_02058_),
    .A(net2644),
    .B(_00127_));
 sg13g2_o21ai_1 _07299_ (.B1(_02058_),
    .Y(_02059_),
    .A1(net2643),
    .A2(_01156_));
 sg13g2_inv_1 _07300_ (.Y(_02060_),
    .A(_02059_));
 sg13g2_nor2_2 _07301_ (.A(_01153_),
    .B(_02059_),
    .Y(_02061_));
 sg13g2_and2_1 _07302_ (.A(_01153_),
    .B(_02059_),
    .X(_02062_));
 sg13g2_nor2_2 _07303_ (.A(_02061_),
    .B(_02062_),
    .Y(_02063_));
 sg13g2_or2_1 _07304_ (.X(_02064_),
    .B(_02062_),
    .A(_02061_));
 sg13g2_and2_1 _07305_ (.A(net2646),
    .B(_00129_),
    .X(_02065_));
 sg13g2_nor3_2 _07306_ (.A(net2642),
    .B(_01114_),
    .C(_01115_),
    .Y(_02066_));
 sg13g2_or2_1 _07307_ (.X(_02067_),
    .B(_02066_),
    .A(_02065_));
 sg13g2_inv_1 _07308_ (.Y(_02068_),
    .A(_02067_));
 sg13g2_nor2_1 _07309_ (.A(_01113_),
    .B(_02068_),
    .Y(_02069_));
 sg13g2_o21ai_1 _07310_ (.B1(_01112_),
    .Y(_02070_),
    .A1(_02065_),
    .A2(_02066_));
 sg13g2_nor3_1 _07311_ (.A(_01112_),
    .B(_02065_),
    .C(_02066_),
    .Y(_02071_));
 sg13g2_nand2_1 _07312_ (.Y(_02072_),
    .A(_01113_),
    .B(_02068_));
 sg13g2_xnor2_1 _07313_ (.Y(_02073_),
    .A(_01112_),
    .B(_02067_));
 sg13g2_a21oi_2 _07314_ (.B1(_02057_),
    .Y(_02074_),
    .A2(_01127_),
    .A1(net2533));
 sg13g2_a21o_1 _07315_ (.A2(_01127_),
    .A1(net2532),
    .B1(_02057_),
    .X(_02075_));
 sg13g2_nand2_1 _07316_ (.Y(_02076_),
    .A(_01126_),
    .B(_02075_));
 sg13g2_xnor2_1 _07317_ (.Y(_02077_),
    .A(_01126_),
    .B(_02074_));
 sg13g2_xnor2_1 _07318_ (.Y(_02078_),
    .A(_01125_),
    .B(_02074_));
 sg13g2_and2_2 _07319_ (.A(net2644),
    .B(_00128_),
    .X(_02079_));
 sg13g2_nor3_2 _07320_ (.A(net2643),
    .B(_01010_),
    .C(_01011_),
    .Y(_02080_));
 sg13g2_nor3_1 _07321_ (.A(_00998_),
    .B(_02079_),
    .C(_02080_),
    .Y(_02081_));
 sg13g2_or3_1 _07322_ (.A(_00998_),
    .B(_02079_),
    .C(_02080_),
    .X(_02082_));
 sg13g2_o21ai_1 _07323_ (.B1(_00998_),
    .Y(_02083_),
    .A1(_02079_),
    .A2(_02080_));
 sg13g2_and2_1 _07324_ (.A(_02082_),
    .B(_02083_),
    .X(_02084_));
 sg13g2_inv_1 _07325_ (.Y(_02085_),
    .A(_02084_));
 sg13g2_nor3_2 _07326_ (.A(net2643),
    .B(_01142_),
    .C(_01143_),
    .Y(_02086_));
 sg13g2_nor3_1 _07327_ (.A(_01140_),
    .B(_02079_),
    .C(_02086_),
    .Y(_02087_));
 sg13g2_or3_1 _07328_ (.A(_01140_),
    .B(_02079_),
    .C(_02086_),
    .X(_02088_));
 sg13g2_o21ai_1 _07329_ (.B1(_01140_),
    .Y(_02089_),
    .A1(_02079_),
    .A2(_02086_));
 sg13g2_and2_2 _07330_ (.A(_02088_),
    .B(_02089_),
    .X(_02090_));
 sg13g2_nand4_1 _07331_ (.B(_02083_),
    .C(_02088_),
    .A(_02082_),
    .Y(_02091_),
    .D(_02089_));
 sg13g2_a21oi_2 _07332_ (.B1(_02057_),
    .Y(_02092_),
    .A2(_01168_),
    .A1(net2534));
 sg13g2_a21o_1 _07333_ (.A2(_01168_),
    .A1(net2535),
    .B1(_02057_),
    .X(_02093_));
 sg13g2_nor2_1 _07334_ (.A(net2414),
    .B(_02092_),
    .Y(_02094_));
 sg13g2_xnor2_1 _07335_ (.Y(_02095_),
    .A(net2414),
    .B(_02092_));
 sg13g2_mux2_1 _07336_ (.A0(_00126_),
    .A1(_01056_),
    .S(net2534),
    .X(_02096_));
 sg13g2_nand2_1 _07337_ (.Y(_02097_),
    .A(net2432),
    .B(_02096_));
 sg13g2_nor2_1 _07338_ (.A(net2432),
    .B(_02096_),
    .Y(_02098_));
 sg13g2_xnor2_1 _07339_ (.Y(_02099_),
    .A(net2432),
    .B(_02096_));
 sg13g2_or4_1 _07340_ (.A(_02056_),
    .B(_02073_),
    .C(_02095_),
    .D(_02099_),
    .X(_02100_));
 sg13g2_nor4_2 _07341_ (.A(_02064_),
    .B(_02078_),
    .C(_02091_),
    .Y(_02101_),
    .D(_02100_));
 sg13g2_nand2_1 _07342_ (.Y(_02102_),
    .A(net2646),
    .B(_00937_));
 sg13g2_o21ai_1 _07343_ (.B1(_02102_),
    .Y(_02103_),
    .A1(net2641),
    .A2(_01060_));
 sg13g2_or2_1 _07344_ (.X(_02104_),
    .B(_02103_),
    .A(_01059_));
 sg13g2_inv_1 _07345_ (.Y(_02105_),
    .A(_02104_));
 sg13g2_nand2_1 _07346_ (.Y(_02106_),
    .A(net2430),
    .B(_02103_));
 sg13g2_inv_1 _07347_ (.Y(_02107_),
    .A(_02106_));
 sg13g2_nor2_2 _07348_ (.A(_02105_),
    .B(_02107_),
    .Y(_02108_));
 sg13g2_nand4_1 _07349_ (.B(_02050_),
    .C(_02101_),
    .A(_01246_),
    .Y(_02109_),
    .D(_02108_));
 sg13g2_nand2_1 _07350_ (.Y(_02110_),
    .A(_01257_),
    .B(_01262_));
 sg13g2_nand2b_1 _07351_ (.Y(_02111_),
    .B(_01271_),
    .A_N(_01252_));
 sg13g2_nor2_1 _07352_ (.A(_02110_),
    .B(_02111_),
    .Y(_02112_));
 sg13g2_nor4_1 _07353_ (.A(_01391_),
    .B(_01409_),
    .C(_02110_),
    .D(_02111_),
    .Y(_02113_));
 sg13g2_nor2b_1 _07354_ (.A(_02109_),
    .B_N(_02113_),
    .Y(_02114_));
 sg13g2_a21oi_1 _07355_ (.A1(_01399_),
    .A2(_02114_),
    .Y(_02115_),
    .B1(_02012_));
 sg13g2_nor2b_1 _07356_ (.A(_02062_),
    .B_N(_02076_),
    .Y(_02116_));
 sg13g2_o21ai_1 _07357_ (.B1(_02070_),
    .Y(_02117_),
    .A1(_02053_),
    .A2(_02071_));
 sg13g2_a221oi_1 _07358_ (.B2(_02089_),
    .C1(_02087_),
    .B1(_02081_),
    .A1(_01125_),
    .Y(_02118_),
    .A2(_02074_));
 sg13g2_o21ai_1 _07359_ (.B1(_02118_),
    .Y(_02119_),
    .A1(_02091_),
    .A2(_02117_));
 sg13g2_a21oi_1 _07360_ (.A1(_02116_),
    .A2(_02119_),
    .Y(_02120_),
    .B1(_02061_));
 sg13g2_a21oi_1 _07361_ (.A1(net2414),
    .A2(_02092_),
    .Y(_02121_),
    .B1(_02098_));
 sg13g2_o21ai_1 _07362_ (.B1(_02121_),
    .Y(_02122_),
    .A1(_02094_),
    .A2(_02120_));
 sg13g2_a22oi_1 _07363_ (.Y(_02123_),
    .B1(_02103_),
    .B2(net2430),
    .A2(_01244_),
    .A1(net2423));
 sg13g2_o21ai_1 _07364_ (.B1(_02042_),
    .Y(_02124_),
    .A1(net2430),
    .A2(_02103_));
 sg13g2_a22oi_1 _07365_ (.Y(_02125_),
    .B1(_02045_),
    .B2(net2426),
    .A2(_02040_),
    .A1(net2415));
 sg13g2_o21ai_1 _07366_ (.B1(_02125_),
    .Y(_02126_),
    .A1(_02123_),
    .A2(_02124_));
 sg13g2_and3_1 _07367_ (.X(_02127_),
    .A(net2312),
    .B(net2311),
    .C(_02047_));
 sg13g2_o21ai_1 _07368_ (.B1(_02022_),
    .Y(_02128_),
    .A1(_01015_),
    .A2(_02016_));
 sg13g2_a22oi_1 _07369_ (.Y(_02129_),
    .B1(_02128_),
    .B2(_02021_),
    .A2(_02127_),
    .A1(_02126_));
 sg13g2_a21oi_1 _07370_ (.A1(_02029_),
    .A2(_02035_),
    .Y(_02130_),
    .B1(_02034_));
 sg13g2_o21ai_1 _07371_ (.B1(_02130_),
    .Y(_02131_),
    .A1(_02038_),
    .A2(_02129_));
 sg13g2_a22oi_1 _07372_ (.Y(_02132_),
    .B1(_02131_),
    .B2(_02101_),
    .A2(_02122_),
    .A1(_02097_));
 sg13g2_o21ai_1 _07373_ (.B1(_01251_),
    .Y(_02133_),
    .A1(_01250_),
    .A2(_01270_));
 sg13g2_a21oi_1 _07374_ (.A1(_01256_),
    .A2(_01261_),
    .Y(_02134_),
    .B1(_01260_));
 sg13g2_o21ai_1 _07375_ (.B1(_02134_),
    .Y(_02135_),
    .A1(_02110_),
    .A2(_02133_));
 sg13g2_o21ai_1 _07376_ (.B1(_01290_),
    .Y(_02136_),
    .A1(_01289_),
    .A2(_01294_));
 sg13g2_o21ai_1 _07377_ (.B1(_01276_),
    .Y(_02137_),
    .A1(_01275_),
    .A2(_01284_));
 sg13g2_a21o_1 _07378_ (.A2(_02136_),
    .A1(_01390_),
    .B1(_02137_),
    .X(_02138_));
 sg13g2_a221oi_1 _07379_ (.B2(_02112_),
    .C1(_02135_),
    .B1(_02138_),
    .A1(_01406_),
    .Y(_02139_),
    .A2(_02113_));
 sg13g2_or2_1 _07380_ (.X(_02140_),
    .B(_02139_),
    .A(_02109_));
 sg13g2_nand4_1 _07381_ (.B(net2640),
    .C(_00066_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[1] ),
    .Y(_02141_),
    .D(_02099_));
 sg13g2_nand3_1 _07382_ (.B(_02140_),
    .C(_02141_),
    .A(_02132_),
    .Y(_02142_));
 sg13g2_a21o_1 _07383_ (.A2(_02140_),
    .A1(_02132_),
    .B1(_02141_),
    .X(_02143_));
 sg13g2_nand3_1 _07384_ (.B(_02142_),
    .C(_02143_),
    .A(_02115_),
    .Y(_02144_));
 sg13g2_a21oi_1 _07385_ (.A1(_02014_),
    .A2(_02144_),
    .Y(_02145_),
    .B1(net2486));
 sg13g2_nand2_1 _07386_ (.Y(_02146_),
    .A(_01386_),
    .B(net2472));
 sg13g2_a21o_1 _07387_ (.A2(_01489_),
    .A1(net2317),
    .B1(_02146_),
    .X(_02147_));
 sg13g2_nand2_1 _07388_ (.Y(_02148_),
    .A(_01396_),
    .B(_02146_));
 sg13g2_o21ai_1 _07389_ (.B1(_02148_),
    .Y(_02149_),
    .A1(_02145_),
    .A2(_02147_));
 sg13g2_a21o_1 _07390_ (.A2(net2633),
    .A1(_00062_),
    .B1(net2623),
    .X(_02150_));
 sg13g2_a21oi_2 _07391_ (.B1(_02150_),
    .Y(_02151_),
    .A2(_02149_),
    .A1(net2531));
 sg13g2_xor2_1 _07392_ (.B(\ChiselTop.wild.cpu._wbData_T_1[0] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[0] ),
    .X(_02152_));
 sg13g2_a21o_1 _07393_ (.A2(_02152_),
    .A1(net2628),
    .B1(net2622),
    .X(_02153_));
 sg13g2_a21oi_1 _07394_ (.A1(\ChiselTop.wild.cpu.decExReg_decOut_isCssrw ),
    .A2(_00125_),
    .Y(_02154_),
    .B1(net2186));
 sg13g2_o21ai_1 _07395_ (.B1(_02154_),
    .Y(_02155_),
    .A1(_02151_),
    .A2(_02153_));
 sg13g2_nor3_1 _07396_ (.A(\ChiselTop.wild.memAddressReg[2] ),
    .B(\ChiselTop.wild.uartStatusReg[0] ),
    .C(net2506),
    .Y(_02156_));
 sg13g2_a221oi_1 _07397_ (.B2(_00901_),
    .C1(_02156_),
    .B1(net2448),
    .A1(_00938_),
    .Y(_02157_),
    .A2(net2506));
 sg13g2_or2_1 _07398_ (.X(_02158_),
    .B(_02157_),
    .A(_01713_));
 sg13g2_nand2_2 _07399_ (.Y(_02159_),
    .A(\ChiselTop.wild.dmem.MEM_3[0][0] ),
    .B(net2500));
 sg13g2_nand2_1 _07400_ (.Y(_02160_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][0] ),
    .B(net2500));
 sg13g2_a22oi_1 _07401_ (.Y(_02161_),
    .B1(_02160_),
    .B2(_01229_),
    .A2(_02159_),
    .A1(_01231_));
 sg13g2_inv_1 _07402_ (.Y(_02162_),
    .A(_02161_));
 sg13g2_a22oi_1 _07403_ (.Y(_02163_),
    .B1(_02162_),
    .B2(net2525),
    .A2(_01642_),
    .A1(_01220_));
 sg13g2_nand3_1 _07404_ (.B(_02158_),
    .C(_02163_),
    .A(net2187),
    .Y(_02164_));
 sg13g2_and2_1 _07405_ (.A(_02155_),
    .B(_02164_),
    .X(_02165_));
 sg13g2_nand2_2 _07406_ (.Y(_02166_),
    .A(net2620),
    .B(net1524));
 sg13g2_nand3_1 _07407_ (.B(_02155_),
    .C(_02164_),
    .A(net2548),
    .Y(_02167_));
 sg13g2_nand2_2 _07408_ (.Y(_02168_),
    .A(_02166_),
    .B(_02167_));
 sg13g2_mux4_1 _07409_ (.S0(net2695),
    .A0(\ChiselTop.wild.cpu.regs[0][0] ),
    .A1(\ChiselTop.wild.cpu.regs[1][0] ),
    .A2(\ChiselTop.wild.cpu.regs[2][0] ),
    .A3(\ChiselTop.wild.cpu.regs[3][0] ),
    .S1(net2672),
    .X(_02169_));
 sg13g2_nor2_1 _07410_ (.A(net2657),
    .B(_02169_),
    .Y(_02170_));
 sg13g2_nor2b_1 _07411_ (.A(\ChiselTop.wild.cpu.regs[5][0] ),
    .B_N(net2695),
    .Y(_02171_));
 sg13g2_nor2_1 _07412_ (.A(net2695),
    .B(\ChiselTop.wild.cpu.regs[4][0] ),
    .Y(_02172_));
 sg13g2_nor3_1 _07413_ (.A(net2672),
    .B(_02171_),
    .C(_02172_),
    .Y(_02173_));
 sg13g2_nor2b_1 _07414_ (.A(\ChiselTop.wild.cpu.regs[7][0] ),
    .B_N(net2695),
    .Y(_02174_));
 sg13g2_o21ai_1 _07415_ (.B1(net2672),
    .Y(_02175_),
    .A1(net2695),
    .A2(\ChiselTop.wild.cpu.regs[6][0] ));
 sg13g2_o21ai_1 _07416_ (.B1(net2657),
    .Y(_02176_),
    .A1(_02174_),
    .A2(_02175_));
 sg13g2_o21ai_1 _07417_ (.B1(net2468),
    .Y(_02177_),
    .A1(_02173_),
    .A2(_02176_));
 sg13g2_nor2_2 _07418_ (.A(_02170_),
    .B(_02177_),
    .Y(_02178_));
 sg13g2_a21o_1 _07419_ (.A2(_02167_),
    .A1(_02166_),
    .B1(_00976_),
    .X(_02179_));
 sg13g2_nor2_1 _07420_ (.A(net2444),
    .B(_02178_),
    .Y(_02180_));
 sg13g2_inv_1 _07421_ (.Y(_02181_),
    .A(_02180_));
 sg13g2_and2_1 _07422_ (.A(_02179_),
    .B(_02181_),
    .X(_02182_));
 sg13g2_nand2_1 _07423_ (.Y(_02183_),
    .A(_02004_),
    .B(_02182_));
 sg13g2_and4_1 _07424_ (.A(_02000_),
    .B(_02004_),
    .C(_02179_),
    .D(_02181_),
    .X(_02184_));
 sg13g2_o21ai_1 _07425_ (.B1(_01941_),
    .Y(_02185_),
    .A1(_01999_),
    .A2(_02184_));
 sg13g2_nand2_1 _07426_ (.Y(_02186_),
    .A(_01940_),
    .B(_02185_));
 sg13g2_a21oi_1 _07427_ (.A1(_00120_),
    .A2(net2464),
    .Y(_02187_),
    .B1(_01817_));
 sg13g2_o21ai_1 _07428_ (.B1(_01814_),
    .Y(_02188_),
    .A1(_01813_),
    .A2(_02187_));
 sg13g2_inv_1 _07429_ (.Y(_02189_),
    .A(_02188_));
 sg13g2_xnor2_1 _07430_ (.Y(_02190_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[3] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[2] ));
 sg13g2_nand2_1 _07431_ (.Y(_02191_),
    .A(net2616),
    .B(_02190_));
 sg13g2_and2_1 _07432_ (.A(net2365),
    .B(_01607_),
    .X(_02192_));
 sg13g2_a21oi_1 _07433_ (.A1(net2356),
    .A2(_01581_),
    .Y(_02193_),
    .B1(_02192_));
 sg13g2_nor2_1 _07434_ (.A(net2375),
    .B(_02193_),
    .Y(_02194_));
 sg13g2_nand2b_1 _07435_ (.Y(_02195_),
    .B(net2366),
    .A_N(_01584_));
 sg13g2_a21oi_1 _07436_ (.A1(_01746_),
    .A2(_02195_),
    .Y(_02196_),
    .B1(_02194_));
 sg13g2_a21oi_1 _07437_ (.A1(_01449_),
    .A2(_02196_),
    .Y(_02197_),
    .B1(_01454_));
 sg13g2_mux2_1 _07438_ (.A0(_01584_),
    .A1(_01590_),
    .S(net2356),
    .X(_02198_));
 sg13g2_a21oi_2 _07439_ (.B1(_02194_),
    .Y(_02199_),
    .A2(_02198_),
    .A1(net2377));
 sg13g2_or2_1 _07440_ (.X(_02200_),
    .B(_01600_),
    .A(net2365));
 sg13g2_nor2_1 _07441_ (.A(net2344),
    .B(_01751_),
    .Y(_02201_));
 sg13g2_o21ai_1 _07442_ (.B1(net2367),
    .Y(_02202_),
    .A1(net2351),
    .A2(_01948_));
 sg13g2_o21ai_1 _07443_ (.B1(_02200_),
    .Y(_02203_),
    .A1(_02201_),
    .A2(_02202_));
 sg13g2_mux2_1 _07444_ (.A0(_01595_),
    .A1(_01604_),
    .S(net2357),
    .X(_02204_));
 sg13g2_o21ai_1 _07445_ (.B1(net2401),
    .Y(_02205_),
    .A1(net2386),
    .A2(_02204_));
 sg13g2_a21oi_1 _07446_ (.A1(net2386),
    .A2(_02203_),
    .Y(_02206_),
    .B1(_02205_));
 sg13g2_nor2_1 _07447_ (.A(net2486),
    .B(_02206_),
    .Y(_02207_));
 sg13g2_o21ai_1 _07448_ (.B1(_02207_),
    .Y(_02208_),
    .A1(_01457_),
    .A2(_02199_));
 sg13g2_nand2b_1 _07449_ (.Y(_02209_),
    .B(net2369),
    .A_N(_01622_));
 sg13g2_nor2_1 _07450_ (.A(net2380),
    .B(_02209_),
    .Y(_02210_));
 sg13g2_a21oi_1 _07451_ (.A1(net2316),
    .A2(_02210_),
    .Y(_02211_),
    .B1(net2474));
 sg13g2_o21ai_1 _07452_ (.B1(_02211_),
    .Y(_02212_),
    .A1(_02197_),
    .A2(_02208_));
 sg13g2_a21oi_1 _07453_ (.A1(_01332_),
    .A2(net2478),
    .Y(_02213_),
    .B1(net2490));
 sg13g2_o21ai_1 _07454_ (.B1(_01332_),
    .Y(_02214_),
    .A1(_01337_),
    .A2(_01909_));
 sg13g2_nor3_1 _07455_ (.A(_01332_),
    .B(_01337_),
    .C(_01909_),
    .Y(_02215_));
 sg13g2_nor2_1 _07456_ (.A(net2488),
    .B(_02215_),
    .Y(_02216_));
 sg13g2_a221oi_1 _07457_ (.B2(_02216_),
    .C1(net2498),
    .B1(_02214_),
    .A1(_02212_),
    .Y(_02217_),
    .A2(_02213_));
 sg13g2_xnor2_1 _07458_ (.Y(_02218_),
    .A(_01332_),
    .B(_01360_));
 sg13g2_o21ai_1 _07459_ (.B1(net2531),
    .Y(_02219_),
    .A1(net2495),
    .A2(_02218_));
 sg13g2_a21oi_1 _07460_ (.A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[3] ),
    .A2(net2633),
    .Y(_02220_),
    .B1(net2623));
 sg13g2_o21ai_1 _07461_ (.B1(_02220_),
    .Y(_02221_),
    .A1(_02217_),
    .A2(_02219_));
 sg13g2_xnor2_1 _07462_ (.Y(_02222_),
    .A(_01520_),
    .B(_01521_));
 sg13g2_a21oi_1 _07463_ (.A1(net2627),
    .A2(_02222_),
    .Y(_02223_),
    .B1(net2622));
 sg13g2_a221oi_1 _07464_ (.B2(_02223_),
    .C1(net2186),
    .B1(_02221_),
    .A1(net2622),
    .Y(_02224_),
    .A2(\ChiselTop.wild.cpu.decExReg_csrVal[3] ));
 sg13g2_nand3_1 _07465_ (.B(net2502),
    .C(_01229_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][3] ),
    .Y(_02225_));
 sg13g2_nand2_1 _07466_ (.Y(_02226_),
    .A(\ChiselTop.wild.dmem.MEM_2[0][3] ),
    .B(net2500));
 sg13g2_nor2_1 _07467_ (.A(_01234_),
    .B(_02226_),
    .Y(_02227_));
 sg13g2_nand2_1 _07468_ (.Y(_02228_),
    .A(\ChiselTop.wild.dmem.MEM_3[0][3] ),
    .B(net2504));
 sg13g2_nor2_1 _07469_ (.A(_01233_),
    .B(_02228_),
    .Y(_02229_));
 sg13g2_o21ai_1 _07470_ (.B1(\ChiselTop.wild.cpu.decExReg_memLow[1] ),
    .Y(_02230_),
    .A1(_02227_),
    .A2(_02229_));
 sg13g2_nand2_1 _07471_ (.Y(_02231_),
    .A(_02225_),
    .B(_02230_));
 sg13g2_a22oi_1 _07472_ (.Y(_02232_),
    .B1(net2448),
    .B2(\ChiselTop.wild.rx._shiftReg_T_1[2] ),
    .A2(net2507),
    .A1(\ChiselTop.wild.dmem.MEM[0][3] ));
 sg13g2_nor2_1 _07473_ (.A(_01713_),
    .B(_02232_),
    .Y(_02233_));
 sg13g2_a221oi_1 _07474_ (.B2(net2526),
    .C1(_02233_),
    .B1(_02231_),
    .A1(_01177_),
    .Y(_02234_),
    .A2(_02227_));
 sg13g2_a21oi_1 _07475_ (.A1(net2186),
    .A2(_02234_),
    .Y(_02235_),
    .B1(_02224_));
 sg13g2_o21ai_1 _07476_ (.B1(_02191_),
    .Y(_02236_),
    .A1(net2616),
    .A2(_02235_));
 sg13g2_mux4_1 _07477_ (.S0(net2696),
    .A0(\ChiselTop.wild.cpu.regs[0][3] ),
    .A1(\ChiselTop.wild.cpu.regs[1][3] ),
    .A2(\ChiselTop.wild.cpu.regs[2][3] ),
    .A3(\ChiselTop.wild.cpu.regs[3][3] ),
    .S1(net2672),
    .X(_02237_));
 sg13g2_nor2_1 _07478_ (.A(net2657),
    .B(_02237_),
    .Y(_02238_));
 sg13g2_nor2b_1 _07479_ (.A(\ChiselTop.wild.cpu.regs[5][3] ),
    .B_N(net2696),
    .Y(_02239_));
 sg13g2_nor2_1 _07480_ (.A(net2696),
    .B(\ChiselTop.wild.cpu.regs[4][3] ),
    .Y(_02240_));
 sg13g2_nor3_1 _07481_ (.A(net2672),
    .B(_02239_),
    .C(_02240_),
    .Y(_02241_));
 sg13g2_nor2b_1 _07482_ (.A(\ChiselTop.wild.cpu.regs[7][3] ),
    .B_N(net2696),
    .Y(_02242_));
 sg13g2_o21ai_1 _07483_ (.B1(net2672),
    .Y(_02243_),
    .A1(net2696),
    .A2(\ChiselTop.wild.cpu.regs[6][3] ));
 sg13g2_o21ai_1 _07484_ (.B1(net2657),
    .Y(_02244_),
    .A1(_02242_),
    .A2(_02243_));
 sg13g2_o21ai_1 _07485_ (.B1(net2468),
    .Y(_02245_),
    .A1(_02241_),
    .A2(_02244_));
 sg13g2_nor2_2 _07486_ (.A(_02238_),
    .B(_02245_),
    .Y(_02246_));
 sg13g2_nor2_1 _07487_ (.A(net2446),
    .B(_02246_),
    .Y(_02247_));
 sg13g2_a21oi_2 _07488_ (.B1(_02247_),
    .Y(_02248_),
    .A2(_02236_),
    .A1(net2446));
 sg13g2_nand2_1 _07489_ (.Y(_02249_),
    .A(_02189_),
    .B(_02248_));
 sg13g2_nand3_1 _07490_ (.B(_02185_),
    .C(_02249_),
    .A(_01940_),
    .Y(_02250_));
 sg13g2_nor2_1 _07491_ (.A(_02189_),
    .B(_02248_),
    .Y(_02251_));
 sg13g2_nor2_1 _07492_ (.A(_01820_),
    .B(_01876_),
    .Y(_02252_));
 sg13g2_and2_1 _07493_ (.A(_01802_),
    .B(_01878_),
    .X(_02253_));
 sg13g2_nor4_1 _07494_ (.A(_01803_),
    .B(_01878_),
    .C(_02251_),
    .D(_02252_),
    .Y(_02254_));
 sg13g2_a221oi_1 _07495_ (.B2(_02250_),
    .C1(_01735_),
    .B1(_02254_),
    .A1(_01737_),
    .Y(_02255_),
    .A2(_02253_));
 sg13g2_and2_2 _07496_ (.A(net1453),
    .B(net2523),
    .X(_02256_));
 sg13g2_nand2_1 _07497_ (.Y(_02257_),
    .A(_00924_),
    .B(_00981_));
 sg13g2_nand2_1 _07498_ (.Y(_02258_),
    .A(_00027_),
    .B(net2635));
 sg13g2_nand3_1 _07499_ (.B(_01369_),
    .C(_01372_),
    .A(_01285_),
    .Y(_02259_));
 sg13g2_a21oi_1 _07500_ (.A1(_01369_),
    .A2(_01372_),
    .Y(_02260_),
    .B1(_01285_));
 sg13g2_nand3b_1 _07501_ (.B(net2499),
    .C(_02259_),
    .Y(_02261_),
    .A_N(_02260_));
 sg13g2_xnor2_1 _07502_ (.Y(_02262_),
    .A(_01286_),
    .B(_01412_));
 sg13g2_a21o_1 _07503_ (.A2(_01890_),
    .A1(net2390),
    .B1(_01576_),
    .X(_02263_));
 sg13g2_a21oi_1 _07504_ (.A1(_01449_),
    .A2(_02263_),
    .Y(_02264_),
    .B1(_01454_));
 sg13g2_o21ai_1 _07505_ (.B1(net2399),
    .Y(_02265_),
    .A1(net2393),
    .A2(_01882_));
 sg13g2_a21oi_1 _07506_ (.A1(net2390),
    .A2(_01900_),
    .Y(_02266_),
    .B1(_02265_));
 sg13g2_a21oi_1 _07507_ (.A1(net2390),
    .A2(_01887_),
    .Y(_02267_),
    .B1(_01457_));
 sg13g2_nor4_2 _07508_ (.A(net2485),
    .B(_02264_),
    .C(_02266_),
    .Y(_02268_),
    .D(_02267_));
 sg13g2_a21oi_1 _07509_ (.A1(_01286_),
    .A2(net2476),
    .Y(_02269_),
    .B1(_01425_));
 sg13g2_nor2_1 _07510_ (.A(net2394),
    .B(_01903_),
    .Y(_02270_));
 sg13g2_mux4_1 _07511_ (.S0(net2349),
    .A0(net2436),
    .A1(net2420),
    .A2(_01172_),
    .A3(net2433),
    .S1(net2338),
    .X(_02271_));
 sg13g2_nor2_1 _07512_ (.A(net2372),
    .B(_01692_),
    .Y(_02272_));
 sg13g2_a21oi_1 _07513_ (.A1(net2372),
    .A2(_02271_),
    .Y(_02273_),
    .B1(_02272_));
 sg13g2_a21oi_1 _07514_ (.A1(net2394),
    .A2(_02273_),
    .Y(_02274_),
    .B1(_02270_));
 sg13g2_nor2_1 _07515_ (.A(net2315),
    .B(_02274_),
    .Y(_02275_));
 sg13g2_nor2_1 _07516_ (.A(_02268_),
    .B(_02275_),
    .Y(_02276_));
 sg13g2_a22oi_1 _07517_ (.Y(_02277_),
    .B1(_02269_),
    .B2(_02276_),
    .A2(_02262_),
    .A1(net2491));
 sg13g2_nor2_1 _07518_ (.A(net2636),
    .B(_02277_),
    .Y(_02278_));
 sg13g2_a22oi_1 _07519_ (.Y(_02279_),
    .B1(_02261_),
    .B2(_02278_),
    .A2(net2635),
    .A1(_00027_));
 sg13g2_xnor2_1 _07520_ (.Y(_02280_),
    .A(_01533_),
    .B(_01534_));
 sg13g2_a21oi_1 _07521_ (.A1(net2624),
    .A2(_02280_),
    .Y(_02281_),
    .B1(net2170));
 sg13g2_o21ai_1 _07522_ (.B1(_02281_),
    .Y(_02282_),
    .A1(net2624),
    .A2(_02279_));
 sg13g2_nand3_1 _07523_ (.B(net2501),
    .C(_01645_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][2] ),
    .Y(_02283_));
 sg13g2_o21ai_1 _07524_ (.B1(_02283_),
    .Y(_02284_),
    .A1(_01644_),
    .A2(_01922_));
 sg13g2_o21ai_1 _07525_ (.B1(net2184),
    .Y(_02285_),
    .A1(net2322),
    .A2(_02284_));
 sg13g2_nand2_1 _07526_ (.Y(_02286_),
    .A(_02282_),
    .B(_02285_));
 sg13g2_nor2_1 _07527_ (.A(net2536),
    .B(_00982_),
    .Y(_02287_));
 sg13g2_a22oi_1 _07528_ (.Y(_02288_),
    .B1(_02287_),
    .B2(_02257_),
    .A2(_02286_),
    .A1(net2536));
 sg13g2_mux4_1 _07529_ (.S0(net2682),
    .A0(\ChiselTop.wild.cpu.regs[0][10] ),
    .A1(\ChiselTop.wild.cpu.regs[1][10] ),
    .A2(\ChiselTop.wild.cpu.regs[2][10] ),
    .A3(\ChiselTop.wild.cpu.regs[3][10] ),
    .S1(net2664),
    .X(_02289_));
 sg13g2_nor2_1 _07530_ (.A(net2656),
    .B(_02289_),
    .Y(_02290_));
 sg13g2_nor2b_1 _07531_ (.A(\ChiselTop.wild.cpu.regs[5][10] ),
    .B_N(net2699),
    .Y(_02291_));
 sg13g2_nor2_1 _07532_ (.A(net2699),
    .B(\ChiselTop.wild.cpu.regs[4][10] ),
    .Y(_02292_));
 sg13g2_nor3_1 _07533_ (.A(net2664),
    .B(_02291_),
    .C(_02292_),
    .Y(_02293_));
 sg13g2_nor2b_1 _07534_ (.A(\ChiselTop.wild.cpu.regs[7][10] ),
    .B_N(net2682),
    .Y(_02294_));
 sg13g2_o21ai_1 _07535_ (.B1(net2664),
    .Y(_02295_),
    .A1(net2682),
    .A2(\ChiselTop.wild.cpu.regs[6][10] ));
 sg13g2_o21ai_1 _07536_ (.B1(net2651),
    .Y(_02296_),
    .A1(_02294_),
    .A2(_02295_));
 sg13g2_o21ai_1 _07537_ (.B1(net2466),
    .Y(_02297_),
    .A1(_02293_),
    .A2(_02296_));
 sg13g2_nor2_1 _07538_ (.A(_02290_),
    .B(_02297_),
    .Y(_02298_));
 sg13g2_nor2_1 _07539_ (.A(net2439),
    .B(_02298_),
    .Y(_02299_));
 sg13g2_a21oi_1 _07540_ (.A1(net2439),
    .A2(net2133),
    .Y(_02300_),
    .B1(_02299_));
 sg13g2_o21ai_1 _07541_ (.B1(net2185),
    .Y(_02301_),
    .A1(_01176_),
    .A2(_01237_));
 sg13g2_mux2_1 _07542_ (.A0(_02159_),
    .A1(_02160_),
    .S(_01644_),
    .X(_02302_));
 sg13g2_a21o_1 _07543_ (.A2(_02302_),
    .A1(_01176_),
    .B1(_02301_),
    .X(_02303_));
 sg13g2_or3_1 _07544_ (.A(_01296_),
    .B(_01299_),
    .C(_01366_),
    .X(_02304_));
 sg13g2_a21oi_1 _07545_ (.A1(_01367_),
    .A2(_02304_),
    .Y(_02305_),
    .B1(net2496));
 sg13g2_nor2_1 _07546_ (.A(net2383),
    .B(_01438_),
    .Y(_02306_));
 sg13g2_nor2_1 _07547_ (.A(_01576_),
    .B(_02306_),
    .Y(_02307_));
 sg13g2_o21ai_1 _07548_ (.B1(net2319),
    .Y(_02308_),
    .A1(_01450_),
    .A2(_02307_));
 sg13g2_mux2_1 _07549_ (.A0(_01443_),
    .A1(_02005_),
    .S(net2392),
    .X(_02309_));
 sg13g2_o21ai_1 _07550_ (.B1(net2483),
    .Y(_02310_),
    .A1(_01457_),
    .A2(_02306_));
 sg13g2_a21oi_1 _07551_ (.A1(net2399),
    .A2(_02309_),
    .Y(_02311_),
    .B1(_02310_));
 sg13g2_nor2_1 _07552_ (.A(net2382),
    .B(_01470_),
    .Y(_02312_));
 sg13g2_a21oi_1 _07553_ (.A1(net2382),
    .A2(_01488_),
    .Y(_02313_),
    .B1(_02312_));
 sg13g2_a221oi_1 _07554_ (.B2(_01478_),
    .C1(net2476),
    .B1(_02313_),
    .A1(_02308_),
    .Y(_02314_),
    .A2(_02311_));
 sg13g2_a21oi_1 _07555_ (.A1(_01295_),
    .A2(net2476),
    .Y(_02315_),
    .B1(_02314_));
 sg13g2_and3_1 _07556_ (.X(_02316_),
    .A(_01296_),
    .B(_01400_),
    .C(_01406_));
 sg13g2_o21ai_1 _07557_ (.B1(net2491),
    .Y(_02317_),
    .A1(_01407_),
    .A2(_02316_));
 sg13g2_o21ai_1 _07558_ (.B1(_02317_),
    .Y(_02318_),
    .A1(_01385_),
    .A2(_02315_));
 sg13g2_o21ai_1 _07559_ (.B1(net2530),
    .Y(_02319_),
    .A1(_02305_),
    .A2(_02318_));
 sg13g2_a21oi_1 _07560_ (.A1(_02258_),
    .A2(_02319_),
    .Y(_02320_),
    .B1(net2624));
 sg13g2_nand3_1 _07561_ (.B(_01528_),
    .C(_01529_),
    .A(_01506_),
    .Y(_02321_));
 sg13g2_nand2b_1 _07562_ (.Y(_02322_),
    .B(_02321_),
    .A_N(_01530_));
 sg13g2_a21o_1 _07563_ (.A2(_02322_),
    .A1(net2625),
    .B1(net2170),
    .X(_02323_));
 sg13g2_o21ai_1 _07564_ (.B1(_02303_),
    .Y(_02324_),
    .A1(_02320_),
    .A2(_02323_));
 sg13g2_nor2b_1 _07565_ (.A(_00980_),
    .B_N(net1547),
    .Y(_02325_));
 sg13g2_nor3_1 _07566_ (.A(_00116_),
    .B(_00978_),
    .C(_00979_),
    .Y(_02326_));
 sg13g2_nor3_1 _07567_ (.A(net2539),
    .B(_02325_),
    .C(_02326_),
    .Y(_02327_));
 sg13g2_a21oi_2 _07568_ (.B1(_02327_),
    .Y(_02328_),
    .A2(_02324_),
    .A1(net2539));
 sg13g2_mux4_1 _07569_ (.S0(net2682),
    .A0(\ChiselTop.wild.cpu.regs[0][8] ),
    .A1(\ChiselTop.wild.cpu.regs[1][8] ),
    .A2(\ChiselTop.wild.cpu.regs[2][8] ),
    .A3(\ChiselTop.wild.cpu.regs[3][8] ),
    .S1(net2664),
    .X(_02329_));
 sg13g2_nor2_1 _07570_ (.A(net2656),
    .B(_02329_),
    .Y(_02330_));
 sg13g2_nor2b_1 _07571_ (.A(net1540),
    .B_N(net2683),
    .Y(_02331_));
 sg13g2_nor2_1 _07572_ (.A(net2683),
    .B(net1012),
    .Y(_02332_));
 sg13g2_nor3_1 _07573_ (.A(net2665),
    .B(_02331_),
    .C(_02332_),
    .Y(_02333_));
 sg13g2_nor2b_1 _07574_ (.A(\ChiselTop.wild.cpu.regs[7][8] ),
    .B_N(net2683),
    .Y(_02334_));
 sg13g2_o21ai_1 _07575_ (.B1(net2665),
    .Y(_02335_),
    .A1(net2683),
    .A2(\ChiselTop.wild.cpu.regs[6][8] ));
 sg13g2_o21ai_1 _07576_ (.B1(net2652),
    .Y(_02336_),
    .A1(_02334_),
    .A2(_02335_));
 sg13g2_o21ai_1 _07577_ (.B1(net2466),
    .Y(_02337_),
    .A1(_02333_),
    .A2(_02336_));
 sg13g2_nor2_1 _07578_ (.A(_02330_),
    .B(_02337_),
    .Y(_02338_));
 sg13g2_nor2_1 _07579_ (.A(net2438),
    .B(_02338_),
    .Y(_02339_));
 sg13g2_a21oi_1 _07580_ (.A1(net2438),
    .A2(net2131),
    .Y(_02340_),
    .B1(_02339_));
 sg13g2_xnor2_1 _07581_ (.Y(_02341_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[9] ),
    .B(_02326_));
 sg13g2_nand2_1 _07582_ (.Y(_02342_),
    .A(net2613),
    .B(_02341_));
 sg13g2_nand3_1 _07583_ (.B(_01367_),
    .C(_01370_),
    .A(_01291_),
    .Y(_02343_));
 sg13g2_nor2_1 _07584_ (.A(_01371_),
    .B(net2496),
    .Y(_02344_));
 sg13g2_nand3_1 _07585_ (.B(_02343_),
    .C(_02344_),
    .A(_01369_),
    .Y(_02345_));
 sg13g2_o21ai_1 _07586_ (.B1(net2491),
    .Y(_02346_),
    .A1(_01291_),
    .A2(_01408_));
 sg13g2_a21oi_1 _07587_ (.A1(_01291_),
    .A2(_01408_),
    .Y(_02347_),
    .B1(_02346_));
 sg13g2_o21ai_1 _07588_ (.B1(_01577_),
    .Y(_02348_),
    .A1(net2375),
    .A2(_01943_));
 sg13g2_a21oi_1 _07589_ (.A1(_01449_),
    .A2(_02348_),
    .Y(_02349_),
    .B1(_01454_));
 sg13g2_nor2_1 _07590_ (.A(net2375),
    .B(_01946_),
    .Y(_02350_));
 sg13g2_o21ai_1 _07591_ (.B1(net2397),
    .Y(_02351_),
    .A1(net2386),
    .A2(_01942_));
 sg13g2_nor2_1 _07592_ (.A(_02350_),
    .B(_02351_),
    .Y(_02352_));
 sg13g2_nor2_1 _07593_ (.A(net2375),
    .B(_01953_),
    .Y(_02353_));
 sg13g2_nor2_1 _07594_ (.A(_01457_),
    .B(_02353_),
    .Y(_02354_));
 sg13g2_or4_2 _07595_ (.A(net2484),
    .B(_02349_),
    .C(_02352_),
    .D(_02354_),
    .X(_02355_));
 sg13g2_nand2_1 _07596_ (.Y(_02356_),
    .A(net2378),
    .B(_01958_));
 sg13g2_o21ai_1 _07597_ (.B1(_01597_),
    .Y(_02357_),
    .A1(_01171_),
    .A2(net2334));
 sg13g2_nor2_1 _07598_ (.A(net2351),
    .B(_02357_),
    .Y(_02358_));
 sg13g2_a21oi_1 _07599_ (.A1(net2351),
    .A2(_01617_),
    .Y(_02359_),
    .B1(_02358_));
 sg13g2_mux2_1 _07600_ (.A0(_01766_),
    .A1(_02359_),
    .S(net2367),
    .X(_02360_));
 sg13g2_o21ai_1 _07601_ (.B1(_02356_),
    .Y(_02361_),
    .A1(net2378),
    .A2(_02360_));
 sg13g2_a21oi_1 _07602_ (.A1(net2317),
    .A2(_02361_),
    .Y(_02362_),
    .B1(net2476));
 sg13g2_a221oi_1 _07603_ (.B2(_02362_),
    .C1(net2491),
    .B1(_02355_),
    .A1(_01291_),
    .Y(_02363_),
    .A2(net2476));
 sg13g2_nor3_1 _07604_ (.A(net2636),
    .B(_02347_),
    .C(_02363_),
    .Y(_02364_));
 sg13g2_a22oi_1 _07605_ (.Y(_02365_),
    .B1(_02345_),
    .B2(_02364_),
    .A2(net2636),
    .A1(_00027_));
 sg13g2_or2_1 _07606_ (.X(_02366_),
    .B(_02365_),
    .A(net2625));
 sg13g2_a21oi_1 _07607_ (.A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[10] ),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[8] ),
    .Y(_02367_),
    .B1(_01530_));
 sg13g2_xnor2_1 _07608_ (.Y(_02368_),
    .A(_01503_),
    .B(_02367_));
 sg13g2_a21oi_1 _07609_ (.A1(net2624),
    .A2(_02368_),
    .Y(_02369_),
    .B1(net2170));
 sg13g2_a221oi_1 _07610_ (.B2(_01645_),
    .C1(_02301_),
    .B1(_01975_),
    .A1(_01643_),
    .Y(_02370_),
    .A2(_01974_));
 sg13g2_a21o_1 _07611_ (.A2(_02369_),
    .A1(_02366_),
    .B1(_02370_),
    .X(_02371_));
 sg13g2_o21ai_1 _07612_ (.B1(_02342_),
    .Y(_02372_),
    .A1(net2613),
    .A2(_02371_));
 sg13g2_mux4_1 _07613_ (.S0(net2679),
    .A0(\ChiselTop.wild.cpu.regs[0][9] ),
    .A1(\ChiselTop.wild.cpu.regs[1][9] ),
    .A2(\ChiselTop.wild.cpu.regs[2][9] ),
    .A3(\ChiselTop.wild.cpu.regs[3][9] ),
    .S1(net2662),
    .X(_02373_));
 sg13g2_nor2_1 _07614_ (.A(net2652),
    .B(_02373_),
    .Y(_02374_));
 sg13g2_nor2b_1 _07615_ (.A(\ChiselTop.wild.cpu.regs[5][9] ),
    .B_N(net2679),
    .Y(_02375_));
 sg13g2_nor2_1 _07616_ (.A(net2679),
    .B(\ChiselTop.wild.cpu.regs[4][9] ),
    .Y(_02376_));
 sg13g2_nor3_1 _07617_ (.A(net2662),
    .B(_02375_),
    .C(_02376_),
    .Y(_02377_));
 sg13g2_nor2b_1 _07618_ (.A(\ChiselTop.wild.cpu.regs[7][9] ),
    .B_N(net2678),
    .Y(_02378_));
 sg13g2_o21ai_1 _07619_ (.B1(net2662),
    .Y(_02379_),
    .A1(net2678),
    .A2(\ChiselTop.wild.cpu.regs[6][9] ));
 sg13g2_o21ai_1 _07620_ (.B1(net2652),
    .Y(_02380_),
    .A1(_02378_),
    .A2(_02379_));
 sg13g2_o21ai_1 _07621_ (.B1(net2466),
    .Y(_02381_),
    .A1(_02377_),
    .A2(_02380_));
 sg13g2_nor2_1 _07622_ (.A(_02374_),
    .B(_02381_),
    .Y(_02382_));
 sg13g2_nor2_1 _07623_ (.A(net2438),
    .B(_02382_),
    .Y(_02383_));
 sg13g2_a21oi_2 _07624_ (.B1(_02383_),
    .Y(_02384_),
    .A2(net2129),
    .A1(net2438));
 sg13g2_nand3_1 _07625_ (.B(_02340_),
    .C(_02384_),
    .A(_02300_),
    .Y(_02385_));
 sg13g2_nor2b_1 _07626_ (.A(_02256_),
    .B_N(_02385_),
    .Y(_02386_));
 sg13g2_nor2_1 _07627_ (.A(\ChiselTop.wild.cpu.decExReg_pc[11] ),
    .B(_00982_),
    .Y(_02387_));
 sg13g2_nor2_1 _07628_ (.A(_01281_),
    .B(_02260_),
    .Y(_02388_));
 sg13g2_o21ai_1 _07629_ (.B1(net2499),
    .Y(_02389_),
    .A1(net2321),
    .A2(_02388_));
 sg13g2_a21oi_1 _07630_ (.A1(net2321),
    .A2(_02388_),
    .Y(_02390_),
    .B1(_02389_));
 sg13g2_o21ai_1 _07631_ (.B1(_01283_),
    .Y(_02391_),
    .A1(_01286_),
    .A2(_01412_));
 sg13g2_a21oi_1 _07632_ (.A1(_01277_),
    .A2(_02391_),
    .Y(_02392_),
    .B1(net2489));
 sg13g2_o21ai_1 _07633_ (.B1(_02392_),
    .Y(_02393_),
    .A1(net2321),
    .A2(_02391_));
 sg13g2_a21oi_1 _07634_ (.A1(net2375),
    .A2(_02193_),
    .Y(_02394_),
    .B1(net2402));
 sg13g2_o21ai_1 _07635_ (.B1(_02394_),
    .Y(_02395_),
    .A1(net2376),
    .A2(_02204_));
 sg13g2_o21ai_1 _07636_ (.B1(net2431),
    .Y(_02396_),
    .A1(net2377),
    .A2(net2358));
 sg13g2_o21ai_1 _07637_ (.B1(_02396_),
    .Y(_02397_),
    .A1(net2377),
    .A2(_02195_));
 sg13g2_nand2_1 _07638_ (.Y(_02398_),
    .A(_01449_),
    .B(_02397_));
 sg13g2_nand2b_1 _07639_ (.Y(_02399_),
    .B(net2385),
    .A_N(_02198_));
 sg13g2_a221oi_1 _07640_ (.B2(net2318),
    .C1(net2484),
    .B1(_02399_),
    .A1(net2319),
    .Y(_02400_),
    .A2(_02398_));
 sg13g2_mux2_1 _07641_ (.A0(net2434),
    .A1(_01093_),
    .S(net2330),
    .X(_02401_));
 sg13g2_mux2_1 _07642_ (.A0(_02357_),
    .A1(_02401_),
    .S(net2344),
    .X(_02402_));
 sg13g2_nor2_1 _07643_ (.A(net2368),
    .B(_01618_),
    .Y(_02403_));
 sg13g2_a21oi_1 _07644_ (.A1(net2368),
    .A2(_02402_),
    .Y(_02404_),
    .B1(_02403_));
 sg13g2_nand2_1 _07645_ (.Y(_02405_),
    .A(net2387),
    .B(_02404_));
 sg13g2_o21ai_1 _07646_ (.B1(_02405_),
    .Y(_02406_),
    .A1(net2387),
    .A2(_02209_));
 sg13g2_a221oi_1 _07647_ (.B2(net2316),
    .C1(net2474),
    .B1(_02406_),
    .A1(_02395_),
    .Y(_02407_),
    .A2(_02400_));
 sg13g2_nor2_1 _07648_ (.A(net2321),
    .B(net2472),
    .Y(_02408_));
 sg13g2_o21ai_1 _07649_ (.B1(_01386_),
    .Y(_02409_),
    .A1(_02407_),
    .A2(_02408_));
 sg13g2_nand3_1 _07650_ (.B(_02393_),
    .C(_02409_),
    .A(net2531),
    .Y(_02410_));
 sg13g2_a21oi_1 _07651_ (.A1(_00911_),
    .A2(net2635),
    .Y(_02411_),
    .B1(net2624));
 sg13g2_o21ai_1 _07652_ (.B1(_02411_),
    .Y(_02412_),
    .A1(_02390_),
    .A2(_02410_));
 sg13g2_xnor2_1 _07653_ (.Y(_02413_),
    .A(_01535_),
    .B(_01536_));
 sg13g2_a21oi_1 _07654_ (.A1(net2624),
    .A2(_02413_),
    .Y(_02414_),
    .B1(net2170));
 sg13g2_nand3_1 _07655_ (.B(net2502),
    .C(_01645_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][3] ),
    .Y(_02415_));
 sg13g2_o21ai_1 _07656_ (.B1(_02415_),
    .Y(_02416_),
    .A1(_01644_),
    .A2(_02228_));
 sg13g2_nand2_1 _07657_ (.Y(_02417_),
    .A(net2185),
    .B(_02416_));
 sg13g2_nand2_2 _07658_ (.Y(_02418_),
    .A(_01641_),
    .B(_02417_));
 sg13g2_a21o_1 _07659_ (.A2(_02414_),
    .A1(_02412_),
    .B1(_02418_),
    .X(_02419_));
 sg13g2_nor3_1 _07660_ (.A(net2536),
    .B(_00983_),
    .C(_02387_),
    .Y(_02420_));
 sg13g2_a21o_1 _07661_ (.A2(_02419_),
    .A1(net2536),
    .B1(_02420_),
    .X(_02421_));
 sg13g2_mux4_1 _07662_ (.S0(net2687),
    .A0(\ChiselTop.wild.cpu.regs[0][11] ),
    .A1(\ChiselTop.wild.cpu.regs[1][11] ),
    .A2(\ChiselTop.wild.cpu.regs[2][11] ),
    .A3(\ChiselTop.wild.cpu.regs[3][11] ),
    .S1(net2668),
    .X(_02422_));
 sg13g2_nor2_1 _07663_ (.A(net2654),
    .B(_02422_),
    .Y(_02423_));
 sg13g2_nor2b_1 _07664_ (.A(net1087),
    .B_N(net2687),
    .Y(_02424_));
 sg13g2_nor2_1 _07665_ (.A(net2687),
    .B(\ChiselTop.wild.cpu.regs[4][11] ),
    .Y(_02425_));
 sg13g2_nor3_1 _07666_ (.A(net2667),
    .B(_02424_),
    .C(_02425_),
    .Y(_02426_));
 sg13g2_nor2b_1 _07667_ (.A(\ChiselTop.wild.cpu.regs[7][11] ),
    .B_N(net2687),
    .Y(_02427_));
 sg13g2_o21ai_1 _07668_ (.B1(net2667),
    .Y(_02428_),
    .A1(net2687),
    .A2(\ChiselTop.wild.cpu.regs[6][11] ));
 sg13g2_o21ai_1 _07669_ (.B1(net2654),
    .Y(_02429_),
    .A1(_02427_),
    .A2(_02428_));
 sg13g2_o21ai_1 _07670_ (.B1(net2467),
    .Y(_02430_),
    .A1(_02426_),
    .A2(_02429_));
 sg13g2_nor2_2 _07671_ (.A(_02423_),
    .B(_02430_),
    .Y(_02431_));
 sg13g2_mux2_1 _07672_ (.A0(net2124),
    .A1(_02431_),
    .S(_00976_),
    .X(_02432_));
 sg13g2_nor2_1 _07673_ (.A(_01813_),
    .B(_02001_),
    .Y(_02433_));
 sg13g2_nand2_2 _07674_ (.Y(_02434_),
    .A(net2550),
    .B(net2465));
 sg13g2_mux2_1 _07675_ (.A0(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[0] ),
    .A1(_00963_),
    .S(_02434_),
    .X(_02435_));
 sg13g2_mux2_2 _07676_ (.A0(\ChiselTop.wild.cpu._GEN_176[20] ),
    .A1(_02435_),
    .S(_02433_),
    .X(_02436_));
 sg13g2_or3_1 _07677_ (.A(_02300_),
    .B(_02340_),
    .C(_02384_),
    .X(_02437_));
 sg13g2_a22oi_1 _07678_ (.Y(_02438_),
    .B1(_02437_),
    .B2(_02256_),
    .A2(_02436_),
    .A1(_02432_));
 sg13g2_o21ai_1 _07679_ (.B1(_02438_),
    .Y(_02439_),
    .A1(_02255_),
    .A2(_02386_));
 sg13g2_and2_2 _07680_ (.A(\ChiselTop.wild.cpu._GEN_176[20] ),
    .B(net2523),
    .X(_02440_));
 sg13g2_nand2_2 _07681_ (.Y(_02441_),
    .A(net1525),
    .B(net2523));
 sg13g2_a21oi_1 _07682_ (.A1(\ChiselTop.wild.cpu.decExReg_pc[13] ),
    .A2(_00984_),
    .Y(_02442_),
    .B1(\ChiselTop.wild.cpu.decExReg_pc[14] ));
 sg13g2_o21ai_1 _07683_ (.B1(net2613),
    .Y(_02443_),
    .A1(_00985_),
    .A2(_02442_));
 sg13g2_inv_1 _07684_ (.Y(_02444_),
    .A(_02443_));
 sg13g2_and2_1 _07685_ (.A(_00011_),
    .B(net2632),
    .X(_02445_));
 sg13g2_o21ai_1 _07686_ (.B1(_01252_),
    .Y(_02446_),
    .A1(_01375_),
    .A2(_01376_));
 sg13g2_a21oi_1 _07687_ (.A1(_01266_),
    .A2(_02446_),
    .Y(_02447_),
    .B1(_01257_));
 sg13g2_and3_1 _07688_ (.X(_02448_),
    .A(_01257_),
    .B(_01266_),
    .C(_02446_));
 sg13g2_o21ai_1 _07689_ (.B1(net2499),
    .Y(_02449_),
    .A1(_02447_),
    .A2(_02448_));
 sg13g2_a21oi_1 _07690_ (.A1(net2391),
    .A2(_01675_),
    .Y(_02450_),
    .B1(_01576_));
 sg13g2_o21ai_1 _07691_ (.B1(net2320),
    .Y(_02451_),
    .A1(net2480),
    .A2(_02450_));
 sg13g2_a21oi_1 _07692_ (.A1(net2391),
    .A2(_01687_),
    .Y(_02452_),
    .B1(net2403));
 sg13g2_o21ai_1 _07693_ (.B1(_02452_),
    .Y(_02453_),
    .A1(net2391),
    .A2(_01666_));
 sg13g2_nor2_1 _07694_ (.A(net2381),
    .B(_01670_),
    .Y(_02454_));
 sg13g2_o21ai_1 _07695_ (.B1(net2318),
    .Y(_02455_),
    .A1(net2381),
    .A2(_01670_));
 sg13g2_nand4_1 _07696_ (.B(_02451_),
    .C(_02453_),
    .A(net2483),
    .Y(_02456_),
    .D(_02455_));
 sg13g2_o21ai_1 _07697_ (.B1(_01386_),
    .Y(_02457_),
    .A1(_01257_),
    .A2(net2473));
 sg13g2_mux4_1 _07698_ (.S0(net2354),
    .A0(_01047_),
    .A1(_01093_),
    .A2(_01104_),
    .A3(net2428),
    .S1(net2338),
    .X(_02458_));
 sg13g2_mux2_1 _07699_ (.A0(_02271_),
    .A1(_02458_),
    .S(net2372),
    .X(_02459_));
 sg13g2_nor2_1 _07700_ (.A(net2383),
    .B(_02459_),
    .Y(_02460_));
 sg13g2_a21oi_1 _07701_ (.A1(net2383),
    .A2(_01695_),
    .Y(_02461_),
    .B1(_02460_));
 sg13g2_nor2_1 _07702_ (.A(net2315),
    .B(_02461_),
    .Y(_02462_));
 sg13g2_nor2_1 _07703_ (.A(_02457_),
    .B(_02462_),
    .Y(_02463_));
 sg13g2_xnor2_1 _07704_ (.Y(_02464_),
    .A(_01257_),
    .B(_01420_));
 sg13g2_a22oi_1 _07705_ (.Y(_02465_),
    .B1(_02464_),
    .B2(net2494),
    .A2(_02463_),
    .A1(_02456_));
 sg13g2_a21oi_1 _07706_ (.A1(_02449_),
    .A2(_02465_),
    .Y(_02466_),
    .B1(net2635));
 sg13g2_o21ai_1 _07707_ (.B1(net2529),
    .Y(_02467_),
    .A1(_02445_),
    .A2(_02466_));
 sg13g2_xnor2_1 _07708_ (.Y(_02468_),
    .A(_01498_),
    .B(_01541_));
 sg13g2_a21oi_1 _07709_ (.A1(net2625),
    .A2(_02468_),
    .Y(_02469_),
    .B1(net2170));
 sg13g2_nand3_1 _07710_ (.B(net2501),
    .C(_01645_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][6] ),
    .Y(_02470_));
 sg13g2_nand3_1 _07711_ (.B(net2501),
    .C(_01643_),
    .A(\ChiselTop.wild.dmem.MEM_3[0][6] ),
    .Y(_02471_));
 sg13g2_nand3_1 _07712_ (.B(_02470_),
    .C(_02471_),
    .A(_01239_),
    .Y(_02472_));
 sg13g2_a221oi_1 _07713_ (.B2(net2184),
    .C1(net2613),
    .B1(_02472_),
    .A1(_02467_),
    .Y(_02473_),
    .A2(_02469_));
 sg13g2_or2_1 _07714_ (.X(_02474_),
    .B(_02473_),
    .A(_02444_));
 sg13g2_mux4_1 _07715_ (.S0(net2688),
    .A0(\ChiselTop.wild.cpu.regs[0][14] ),
    .A1(\ChiselTop.wild.cpu.regs[1][14] ),
    .A2(\ChiselTop.wild.cpu.regs[2][14] ),
    .A3(\ChiselTop.wild.cpu.regs[3][14] ),
    .S1(net2667),
    .X(_02475_));
 sg13g2_nor2_1 _07716_ (.A(net2653),
    .B(_02475_),
    .Y(_02476_));
 sg13g2_nor2b_1 _07717_ (.A(\ChiselTop.wild.cpu.regs[5][14] ),
    .B_N(net2684),
    .Y(_02477_));
 sg13g2_nor2_1 _07718_ (.A(net2684),
    .B(\ChiselTop.wild.cpu.regs[4][14] ),
    .Y(_02478_));
 sg13g2_nor3_1 _07719_ (.A(net2666),
    .B(_02477_),
    .C(_02478_),
    .Y(_02479_));
 sg13g2_nor2b_1 _07720_ (.A(\ChiselTop.wild.cpu.regs[7][14] ),
    .B_N(net2684),
    .Y(_02480_));
 sg13g2_o21ai_1 _07721_ (.B1(net2666),
    .Y(_02481_),
    .A1(net2684),
    .A2(\ChiselTop.wild.cpu.regs[6][14] ));
 sg13g2_o21ai_1 _07722_ (.B1(net2653),
    .Y(_02482_),
    .A1(_02480_),
    .A2(_02481_));
 sg13g2_o21ai_1 _07723_ (.B1(net2470),
    .Y(_02483_),
    .A1(_02479_),
    .A2(_02482_));
 sg13g2_nand3b_1 _07724_ (.B(net2441),
    .C(_02443_),
    .Y(_02484_),
    .A_N(_02473_));
 sg13g2_or3_2 _07725_ (.A(net2438),
    .B(_02476_),
    .C(_02483_),
    .X(_02485_));
 sg13g2_a21o_1 _07726_ (.A2(_02485_),
    .A1(_02484_),
    .B1(_02441_),
    .X(_02486_));
 sg13g2_o21ai_1 _07727_ (.B1(_00964_),
    .Y(_02487_),
    .A1(net1541),
    .A2(net2522));
 sg13g2_inv_2 _07728_ (.Y(_02488_),
    .A(_02487_));
 sg13g2_xnor2_1 _07729_ (.Y(_02489_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[15] ),
    .B(_00985_));
 sg13g2_nand2_1 _07730_ (.Y(_02490_),
    .A(net2615),
    .B(_02489_));
 sg13g2_nor2_1 _07731_ (.A(_01230_),
    .B(_01644_),
    .Y(_02491_));
 sg13g2_nor2_1 _07732_ (.A(net2322),
    .B(_02491_),
    .Y(_02492_));
 sg13g2_o21ai_1 _07733_ (.B1(_02492_),
    .Y(_02493_),
    .A1(_01228_),
    .A2(_01646_));
 sg13g2_o21ai_1 _07734_ (.B1(_01262_),
    .Y(_02494_),
    .A1(_01265_),
    .A2(_02447_));
 sg13g2_nor3_1 _07735_ (.A(_01262_),
    .B(_01265_),
    .C(_02447_),
    .Y(_02495_));
 sg13g2_nand3b_1 _07736_ (.B(net2499),
    .C(_02494_),
    .Y(_02496_),
    .A_N(_02495_));
 sg13g2_nor2_1 _07737_ (.A(net2385),
    .B(_01585_),
    .Y(_02497_));
 sg13g2_o21ai_1 _07738_ (.B1(net2397),
    .Y(_02498_),
    .A1(net2376),
    .A2(_01608_));
 sg13g2_a21oi_1 _07739_ (.A1(net2389),
    .A2(_01591_),
    .Y(_02499_),
    .B1(_01457_));
 sg13g2_o21ai_1 _07740_ (.B1(_01455_),
    .Y(_02500_),
    .A1(_02497_),
    .A2(_02498_));
 sg13g2_nor2_1 _07741_ (.A(net2388),
    .B(_01624_),
    .Y(_02501_));
 sg13g2_mux2_1 _07742_ (.A0(net2429),
    .A1(_01047_),
    .S(net2330),
    .X(_02502_));
 sg13g2_o21ai_1 _07743_ (.B1(_01602_),
    .Y(_02503_),
    .A1(_01103_),
    .A2(net2335));
 sg13g2_mux2_1 _07744_ (.A0(_02502_),
    .A1(_02503_),
    .S(net2344),
    .X(_02504_));
 sg13g2_and2_1 _07745_ (.A(net2367),
    .B(_02504_),
    .X(_02505_));
 sg13g2_a21oi_1 _07746_ (.A1(net2360),
    .A2(_02402_),
    .Y(_02506_),
    .B1(_02505_));
 sg13g2_a21oi_1 _07747_ (.A1(net2388),
    .A2(_02506_),
    .Y(_02507_),
    .B1(_02501_));
 sg13g2_inv_1 _07748_ (.Y(_02508_),
    .A(_02507_));
 sg13g2_a221oi_1 _07749_ (.B2(net2317),
    .C1(net2490),
    .B1(_02508_),
    .A1(_01263_),
    .Y(_02509_),
    .A2(net2474));
 sg13g2_o21ai_1 _07750_ (.B1(_02509_),
    .Y(_02510_),
    .A1(_02499_),
    .A2(_02500_));
 sg13g2_xnor2_1 _07751_ (.Y(_02511_),
    .A(_01262_),
    .B(_01422_));
 sg13g2_o21ai_1 _07752_ (.B1(_02510_),
    .Y(_02512_),
    .A1(net2489),
    .A2(_02511_));
 sg13g2_a21oi_1 _07753_ (.A1(net2496),
    .A2(_02512_),
    .Y(_02513_),
    .B1(net2635));
 sg13g2_o21ai_1 _07754_ (.B1(net2529),
    .Y(_02514_),
    .A1(_00007_),
    .A2(net2531));
 sg13g2_a21o_1 _07755_ (.A2(_02513_),
    .A1(_02496_),
    .B1(_02514_),
    .X(_02515_));
 sg13g2_xnor2_1 _07756_ (.Y(_02516_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[15] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[15] ));
 sg13g2_xnor2_1 _07757_ (.Y(_02517_),
    .A(_01542_),
    .B(_02516_));
 sg13g2_a21oi_1 _07758_ (.A1(net2625),
    .A2(_02517_),
    .Y(_02518_),
    .B1(net2170));
 sg13g2_a221oi_1 _07759_ (.B2(_02518_),
    .C1(net2613),
    .B1(_02515_),
    .A1(net2184),
    .Y(_02519_),
    .A2(_02493_));
 sg13g2_a21o_2 _07760_ (.A2(_02489_),
    .A1(net2615),
    .B1(_02519_),
    .X(_02520_));
 sg13g2_mux4_1 _07761_ (.S0(net2700),
    .A0(\ChiselTop.wild.cpu.regs[0][15] ),
    .A1(\ChiselTop.wild.cpu.regs[1][15] ),
    .A2(\ChiselTop.wild.cpu.regs[2][15] ),
    .A3(\ChiselTop.wild.cpu.regs[3][15] ),
    .S1(net2677),
    .X(_02521_));
 sg13g2_nor2_1 _07762_ (.A(net2660),
    .B(_02521_),
    .Y(_02522_));
 sg13g2_nor2b_1 _07763_ (.A(\ChiselTop.wild.cpu.regs[5][15] ),
    .B_N(net2700),
    .Y(_02523_));
 sg13g2_nor2_1 _07764_ (.A(net2700),
    .B(\ChiselTop.wild.cpu.regs[4][15] ),
    .Y(_02524_));
 sg13g2_nor3_1 _07765_ (.A(net2677),
    .B(_02523_),
    .C(_02524_),
    .Y(_02525_));
 sg13g2_nor2b_1 _07766_ (.A(\ChiselTop.wild.cpu.regs[7][15] ),
    .B_N(net2700),
    .Y(_02526_));
 sg13g2_o21ai_1 _07767_ (.B1(net2677),
    .Y(_02527_),
    .A1(net2700),
    .A2(\ChiselTop.wild.cpu.regs[6][15] ));
 sg13g2_o21ai_1 _07768_ (.B1(net2660),
    .Y(_02528_),
    .A1(_02526_),
    .A2(_02527_));
 sg13g2_o21ai_1 _07769_ (.B1(net2469),
    .Y(_02529_),
    .A1(_02525_),
    .A2(_02528_));
 sg13g2_nand3b_1 _07770_ (.B(_00975_),
    .C(_02490_),
    .Y(_02530_),
    .A_N(_02519_));
 sg13g2_or3_1 _07771_ (.A(net2440),
    .B(_02522_),
    .C(_02529_),
    .X(_02531_));
 sg13g2_a21o_1 _07772_ (.A2(_02531_),
    .A1(_02530_),
    .B1(_02488_),
    .X(_02532_));
 sg13g2_nand3_1 _07773_ (.B(_02484_),
    .C(_02485_),
    .A(_02441_),
    .Y(_02533_));
 sg13g2_and3_1 _07774_ (.X(_02534_),
    .A(_02488_),
    .B(_02530_),
    .C(_02531_));
 sg13g2_nand3_1 _07775_ (.B(_02530_),
    .C(_02531_),
    .A(_02488_),
    .Y(_02535_));
 sg13g2_and4_1 _07776_ (.A(_02486_),
    .B(_02532_),
    .C(_02533_),
    .D(_02535_),
    .X(_02536_));
 sg13g2_nand4_1 _07777_ (.B(_02532_),
    .C(_02533_),
    .A(_02486_),
    .Y(_02537_),
    .D(_02535_));
 sg13g2_o21ai_1 _07778_ (.B1(_00964_),
    .Y(_02538_),
    .A1(_00113_),
    .A2(net2522));
 sg13g2_or2_1 _07779_ (.X(_02539_),
    .B(_00984_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[13] ));
 sg13g2_o21ai_1 _07780_ (.B1(_02396_),
    .Y(_02540_),
    .A1(net2377),
    .A2(_01745_));
 sg13g2_nand2_1 _07781_ (.Y(_02541_),
    .A(_01449_),
    .B(_02540_));
 sg13g2_a21oi_1 _07782_ (.A1(net2386),
    .A2(_01756_),
    .Y(_02542_),
    .B1(net2402));
 sg13g2_o21ai_1 _07783_ (.B1(_02542_),
    .Y(_02543_),
    .A1(net2386),
    .A2(_01743_));
 sg13g2_nand3_1 _07784_ (.B(net2366),
    .C(_01759_),
    .A(net2385),
    .Y(_02544_));
 sg13g2_a22oi_1 _07785_ (.Y(_02545_),
    .B1(_02544_),
    .B2(net2318),
    .A2(_02541_),
    .A1(net2319));
 sg13g2_nand3_1 _07786_ (.B(_02543_),
    .C(_02545_),
    .A(net2481),
    .Y(_02546_));
 sg13g2_mux2_1 _07787_ (.A0(_02401_),
    .A1(_02502_),
    .S(net2344),
    .X(_02547_));
 sg13g2_mux2_1 _07788_ (.A0(_02359_),
    .A1(_02547_),
    .S(net2368),
    .X(_02548_));
 sg13g2_nor2_1 _07789_ (.A(net2379),
    .B(_02548_),
    .Y(_02549_));
 sg13g2_a21oi_2 _07790_ (.B1(_02549_),
    .Y(_02550_),
    .A2(_01767_),
    .A1(net2378));
 sg13g2_nor2_1 _07791_ (.A(net2315),
    .B(_02550_),
    .Y(_02551_));
 sg13g2_a21oi_1 _07792_ (.A1(_01252_),
    .A2(net2477),
    .Y(_02552_),
    .B1(_02551_));
 sg13g2_nand3_1 _07793_ (.B(_02546_),
    .C(_02552_),
    .A(net2489),
    .Y(_02553_));
 sg13g2_xor2_1 _07794_ (.B(_01418_),
    .A(_01252_),
    .X(_02554_));
 sg13g2_o21ai_1 _07795_ (.B1(_02553_),
    .Y(_02555_),
    .A1(net2489),
    .A2(_02554_));
 sg13g2_or3_1 _07796_ (.A(_01252_),
    .B(_01375_),
    .C(_01376_),
    .X(_02556_));
 sg13g2_nand3_1 _07797_ (.B(_02446_),
    .C(_02556_),
    .A(net2499),
    .Y(_02557_));
 sg13g2_a21oi_1 _07798_ (.A1(_02555_),
    .A2(_02557_),
    .Y(_02558_),
    .B1(net2636));
 sg13g2_o21ai_1 _07799_ (.B1(net2529),
    .Y(_02559_),
    .A1(_00015_),
    .A2(net2531));
 sg13g2_xnor2_1 _07800_ (.Y(_02560_),
    .A(_01539_),
    .B(_01540_));
 sg13g2_a21oi_1 _07801_ (.A1(net2624),
    .A2(_02560_),
    .Y(_02561_),
    .B1(net2170));
 sg13g2_o21ai_1 _07802_ (.B1(_02561_),
    .Y(_02562_),
    .A1(_02558_),
    .A2(_02559_));
 sg13g2_nand3_1 _07803_ (.B(net2501),
    .C(_01645_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][5] ),
    .Y(_02563_));
 sg13g2_o21ai_1 _07804_ (.B1(_02563_),
    .Y(_02564_),
    .A1(_01644_),
    .A2(_01782_));
 sg13g2_o21ai_1 _07805_ (.B1(net2183),
    .Y(_02565_),
    .A1(net2322),
    .A2(_02564_));
 sg13g2_nand2_1 _07806_ (.Y(_02566_),
    .A(_02562_),
    .B(_02565_));
 sg13g2_a21oi_1 _07807_ (.A1(\ChiselTop.wild.cpu.decExReg_pc[13] ),
    .A2(_00984_),
    .Y(_02567_),
    .B1(net2538));
 sg13g2_a22oi_1 _07808_ (.Y(_02568_),
    .B1(_02567_),
    .B2(_02539_),
    .A2(_02566_),
    .A1(net2538));
 sg13g2_mux4_1 _07809_ (.S0(net2689),
    .A0(\ChiselTop.wild.cpu.regs[0][13] ),
    .A1(\ChiselTop.wild.cpu.regs[1][13] ),
    .A2(\ChiselTop.wild.cpu.regs[2][13] ),
    .A3(\ChiselTop.wild.cpu.regs[3][13] ),
    .S1(net2669),
    .X(_02569_));
 sg13g2_nor2_1 _07810_ (.A(net2660),
    .B(_02569_),
    .Y(_02570_));
 sg13g2_nor2b_1 _07811_ (.A(\ChiselTop.wild.cpu.regs[5][13] ),
    .B_N(net2700),
    .Y(_02571_));
 sg13g2_nor2_1 _07812_ (.A(net2700),
    .B(\ChiselTop.wild.cpu.regs[4][13] ),
    .Y(_02572_));
 sg13g2_nor3_1 _07813_ (.A(net2677),
    .B(_02571_),
    .C(_02572_),
    .Y(_02573_));
 sg13g2_nor2b_1 _07814_ (.A(\ChiselTop.wild.cpu.regs[7][13] ),
    .B_N(net2694),
    .Y(_02574_));
 sg13g2_o21ai_1 _07815_ (.B1(net2671),
    .Y(_02575_),
    .A1(net2700),
    .A2(\ChiselTop.wild.cpu.regs[6][13] ));
 sg13g2_o21ai_1 _07816_ (.B1(net2659),
    .Y(_02576_),
    .A1(_02574_),
    .A2(_02575_));
 sg13g2_o21ai_1 _07817_ (.B1(net2468),
    .Y(_02577_),
    .A1(_02573_),
    .A2(_02576_));
 sg13g2_nor2_1 _07818_ (.A(_02570_),
    .B(_02577_),
    .Y(_02578_));
 sg13g2_nor2_1 _07819_ (.A(net2440),
    .B(_02578_),
    .Y(_02579_));
 sg13g2_a21oi_1 _07820_ (.A1(net2440),
    .A2(net2122),
    .Y(_02580_),
    .B1(_02579_));
 sg13g2_a21oi_2 _07821_ (.B1(_00963_),
    .Y(_02581_),
    .A2(_00961_),
    .A1(_00930_));
 sg13g2_nor2_1 _07822_ (.A(\ChiselTop.wild.cpu.decExReg_pc[12] ),
    .B(_00983_),
    .Y(_02582_));
 sg13g2_o21ai_1 _07823_ (.B1(net2613),
    .Y(_02583_),
    .A1(_00984_),
    .A2(_02582_));
 sg13g2_nand3_1 _07824_ (.B(net2503),
    .C(_01645_),
    .A(\ChiselTop.wild.dmem.MEM_1[0][4] ),
    .Y(_02584_));
 sg13g2_o21ai_1 _07825_ (.B1(_02584_),
    .Y(_02585_),
    .A1(_01644_),
    .A2(_01823_));
 sg13g2_o21ai_1 _07826_ (.B1(net2183),
    .Y(_02586_),
    .A1(net2322),
    .A2(_02585_));
 sg13g2_and2_1 _07827_ (.A(net2391),
    .B(_01836_),
    .X(_02587_));
 sg13g2_nor2b_1 _07828_ (.A(_02587_),
    .B_N(_02396_),
    .Y(_02588_));
 sg13g2_o21ai_1 _07829_ (.B1(net2320),
    .Y(_02589_),
    .A1(net2480),
    .A2(_02588_));
 sg13g2_nor2_1 _07830_ (.A(net2381),
    .B(_01848_),
    .Y(_02590_));
 sg13g2_o21ai_1 _07831_ (.B1(net2398),
    .Y(_02591_),
    .A1(net2392),
    .A2(_01834_));
 sg13g2_o21ai_1 _07832_ (.B1(_02589_),
    .Y(_02592_),
    .A1(_01457_),
    .A2(_02587_));
 sg13g2_o21ai_1 _07833_ (.B1(net2483),
    .Y(_02593_),
    .A1(_02590_),
    .A2(_02591_));
 sg13g2_nor2_1 _07834_ (.A(_02592_),
    .B(_02593_),
    .Y(_02594_));
 sg13g2_a21oi_1 _07835_ (.A1(_01272_),
    .A2(net2477),
    .Y(_02595_),
    .B1(net2491));
 sg13g2_nor2_1 _07836_ (.A(net2395),
    .B(_01853_),
    .Y(_02596_));
 sg13g2_nor2_1 _07837_ (.A(net2373),
    .B(_01468_),
    .Y(_02597_));
 sg13g2_a21oi_1 _07838_ (.A1(net2373),
    .A2(_01476_),
    .Y(_02598_),
    .B1(_02597_));
 sg13g2_a21oi_1 _07839_ (.A1(net2395),
    .A2(_02598_),
    .Y(_02599_),
    .B1(_02596_));
 sg13g2_o21ai_1 _07840_ (.B1(_02595_),
    .Y(_02600_),
    .A1(net2315),
    .A2(_02599_));
 sg13g2_xnor2_1 _07841_ (.Y(_02601_),
    .A(_01271_),
    .B(_01416_));
 sg13g2_nand2_1 _07842_ (.Y(_02602_),
    .A(_01385_),
    .B(_02601_));
 sg13g2_o21ai_1 _07843_ (.B1(_02602_),
    .Y(_02603_),
    .A1(_02594_),
    .A2(_02600_));
 sg13g2_nor2_1 _07844_ (.A(_01272_),
    .B(_01374_),
    .Y(_02604_));
 sg13g2_nand2b_1 _07845_ (.Y(_02605_),
    .B(net2499),
    .A_N(_01375_));
 sg13g2_o21ai_1 _07846_ (.B1(_02603_),
    .Y(_02606_),
    .A1(_02604_),
    .A2(_02605_));
 sg13g2_o21ai_1 _07847_ (.B1(net2529),
    .Y(_02607_),
    .A1(_00019_),
    .A2(net2530));
 sg13g2_a21oi_1 _07848_ (.A1(net2530),
    .A2(_02606_),
    .Y(_02608_),
    .B1(_02607_));
 sg13g2_xnor2_1 _07849_ (.Y(_02609_),
    .A(_01537_),
    .B(_01538_));
 sg13g2_a21o_1 _07850_ (.A2(_02609_),
    .A1(net2624),
    .B1(net2170),
    .X(_02610_));
 sg13g2_o21ai_1 _07851_ (.B1(_02586_),
    .Y(_02611_),
    .A1(_02608_),
    .A2(_02610_));
 sg13g2_o21ai_1 _07852_ (.B1(_02583_),
    .Y(_02612_),
    .A1(net2613),
    .A2(_02611_));
 sg13g2_mux4_1 _07853_ (.S0(net2686),
    .A0(\ChiselTop.wild.cpu.regs[0][12] ),
    .A1(\ChiselTop.wild.cpu.regs[1][12] ),
    .A2(\ChiselTop.wild.cpu.regs[2][12] ),
    .A3(\ChiselTop.wild.cpu.regs[3][12] ),
    .S1(net2667),
    .X(_02613_));
 sg13g2_nor2_1 _07854_ (.A(net2654),
    .B(_02613_),
    .Y(_02614_));
 sg13g2_nor2b_1 _07855_ (.A(\ChiselTop.wild.cpu.regs[5][12] ),
    .B_N(net2686),
    .Y(_02615_));
 sg13g2_nor2_1 _07856_ (.A(net2687),
    .B(\ChiselTop.wild.cpu.regs[4][12] ),
    .Y(_02616_));
 sg13g2_nor3_1 _07857_ (.A(net2668),
    .B(_02615_),
    .C(_02616_),
    .Y(_02617_));
 sg13g2_nor2b_1 _07858_ (.A(\ChiselTop.wild.cpu.regs[7][12] ),
    .B_N(net2686),
    .Y(_02618_));
 sg13g2_o21ai_1 _07859_ (.B1(net2668),
    .Y(_02619_),
    .A1(net2686),
    .A2(\ChiselTop.wild.cpu.regs[6][12] ));
 sg13g2_o21ai_1 _07860_ (.B1(net2653),
    .Y(_02620_),
    .A1(_02618_),
    .A2(_02619_));
 sg13g2_o21ai_1 _07861_ (.B1(net2467),
    .Y(_02621_),
    .A1(_02617_),
    .A2(_02620_));
 sg13g2_nor2_2 _07862_ (.A(_02614_),
    .B(_02621_),
    .Y(_02622_));
 sg13g2_nor2_1 _07863_ (.A(net2442),
    .B(_02622_),
    .Y(_02623_));
 sg13g2_a21oi_1 _07864_ (.A1(net2442),
    .A2(net2126),
    .Y(_02624_),
    .B1(_02623_));
 sg13g2_nor2b_1 _07865_ (.A(_02581_),
    .B_N(_02624_),
    .Y(_02625_));
 sg13g2_a21o_1 _07866_ (.A2(_02580_),
    .A1(_02538_),
    .B1(_02625_),
    .X(_02626_));
 sg13g2_nor2_1 _07867_ (.A(_02538_),
    .B(_02580_),
    .Y(_02627_));
 sg13g2_nand2b_1 _07868_ (.Y(_02628_),
    .B(_02581_),
    .A_N(_02624_));
 sg13g2_o21ai_1 _07869_ (.B1(_02628_),
    .Y(_02629_),
    .A1(_02432_),
    .A2(_02436_));
 sg13g2_nor3_1 _07870_ (.A(_02626_),
    .B(_02627_),
    .C(_02629_),
    .Y(_02630_));
 sg13g2_and3_1 _07871_ (.X(_02631_),
    .A(_02439_),
    .B(_02536_),
    .C(_02630_));
 sg13g2_o21ai_1 _07872_ (.B1(_02626_),
    .Y(_02632_),
    .A1(_02538_),
    .A2(_02580_));
 sg13g2_a21o_1 _07873_ (.A2(_02532_),
    .A1(_02486_),
    .B1(_02534_),
    .X(_02633_));
 sg13g2_o21ai_1 _07874_ (.B1(_02633_),
    .Y(_02634_),
    .A1(_02537_),
    .A2(_02632_));
 sg13g2_o21ai_1 _07875_ (.B1(_01568_),
    .Y(_02635_),
    .A1(_02631_),
    .A2(_02634_));
 sg13g2_inv_1 _07876_ (.Y(_02636_),
    .A(_02635_));
 sg13g2_nor3_2 _07877_ (.A(_01568_),
    .B(_02631_),
    .C(_02634_),
    .Y(_02637_));
 sg13g2_nor2_1 _07878_ (.A(_02636_),
    .B(_02637_),
    .Y(\ChiselTop.wild.cpu.io_dmem_rdAddress[16] ));
 sg13g2_xnor2_1 _07879_ (.Y(\ChiselTop.wild.cpu.decEx_memLow[0] ),
    .A(_02003_),
    .B(_02182_));
 sg13g2_inv_1 _07880_ (.Y(_02638_),
    .A(\ChiselTop.wild.cpu.decEx_memLow[0] ));
 sg13g2_xnor2_1 _07881_ (.Y(\ChiselTop.wild.cpu.decEx_memLow[1] ),
    .A(_02000_),
    .B(_02183_));
 sg13g2_nand2_1 _07882_ (.Y(_02639_),
    .A(_00941_),
    .B(_00961_));
 sg13g2_nand2_2 _07883_ (.Y(_02640_),
    .A(_00964_),
    .B(_02639_));
 sg13g2_nor2_2 _07884_ (.A(_00940_),
    .B(_00986_),
    .Y(_02641_));
 sg13g2_nand3_1 _07885_ (.B(\ChiselTop.wild.cpu.decExReg_pc[18] ),
    .C(_02641_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[19] ),
    .Y(_02642_));
 sg13g2_nor2_1 _07886_ (.A(_00939_),
    .B(_02642_),
    .Y(_02643_));
 sg13g2_and2_1 _07887_ (.A(\ChiselTop.wild.cpu.decExReg_pc[21] ),
    .B(_02643_),
    .X(_02644_));
 sg13g2_and3_1 _07888_ (.X(_02645_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[23] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[22] ),
    .C(_02644_));
 sg13g2_and3_1 _07889_ (.X(_02646_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[25] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[24] ),
    .C(_02645_));
 sg13g2_and2_1 _07890_ (.A(\ChiselTop.wild.cpu.decExReg_pc[26] ),
    .B(_02646_),
    .X(_02647_));
 sg13g2_and2_1 _07891_ (.A(\ChiselTop.wild.cpu.decExReg_pc[27] ),
    .B(_02647_),
    .X(_02648_));
 sg13g2_nand2_1 _07892_ (.Y(_02649_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[27] ),
    .B(_02647_));
 sg13g2_nand3_1 _07893_ (.B(\ChiselTop.wild.cpu.decExReg_pc[28] ),
    .C(_02648_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[29] ),
    .Y(_02650_));
 sg13g2_nand4_1 _07894_ (.B(\ChiselTop.wild.cpu.decExReg_pc[29] ),
    .C(\ChiselTop.wild.cpu.decExReg_pc[28] ),
    .A(\ChiselTop.wild.cpu.decExReg_pc[30] ),
    .Y(_02651_),
    .D(_02648_));
 sg13g2_xor2_1 _07895_ (.B(_02650_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[30] ),
    .X(_02652_));
 sg13g2_nand2_1 _07896_ (.Y(_02653_),
    .A(net2638),
    .B(_00127_));
 sg13g2_nor2_1 _07897_ (.A(net2416),
    .B(_02059_),
    .Y(_02654_));
 sg13g2_nor2_1 _07898_ (.A(net2419),
    .B(_02075_),
    .Y(_02655_));
 sg13g2_nand2_2 _07899_ (.Y(_02656_),
    .A(_01058_),
    .B(_02103_));
 sg13g2_nand2b_1 _07900_ (.Y(_02657_),
    .B(_01244_),
    .A_N(net2422));
 sg13g2_a21o_2 _07901_ (.A2(_02657_),
    .A1(_01384_),
    .B1(_02108_),
    .X(_02658_));
 sg13g2_a21o_1 _07902_ (.A2(_02658_),
    .A1(_02656_),
    .B1(_02043_),
    .X(_02659_));
 sg13g2_nand2_1 _07903_ (.Y(_02660_),
    .A(_02044_),
    .B(_02048_));
 sg13g2_a21oi_1 _07904_ (.A1(_02656_),
    .A2(_02658_),
    .Y(_02661_),
    .B1(_02660_));
 sg13g2_a21o_1 _07905_ (.A2(_02658_),
    .A1(_02656_),
    .B1(_02660_),
    .X(_02662_));
 sg13g2_nand2b_1 _07906_ (.Y(_02663_),
    .B(_02045_),
    .A_N(_01082_));
 sg13g2_nand2_1 _07907_ (.Y(_02664_),
    .A(_01159_),
    .B(_02040_));
 sg13g2_nor2_1 _07908_ (.A(_02049_),
    .B(_02664_),
    .Y(_02665_));
 sg13g2_o21ai_1 _07909_ (.B1(_02663_),
    .Y(_02666_),
    .A1(_02049_),
    .A2(_02664_));
 sg13g2_inv_1 _07910_ (.Y(_02667_),
    .A(_02666_));
 sg13g2_nor2_1 _07911_ (.A(_02661_),
    .B(_02666_),
    .Y(_02668_));
 sg13g2_nor4_1 _07912_ (.A(net2312),
    .B(net2311),
    .C(_02032_),
    .D(_02036_),
    .Y(_02669_));
 sg13g2_o21ai_1 _07913_ (.B1(_02669_),
    .Y(_02670_),
    .A1(_02661_),
    .A2(_02666_));
 sg13g2_nor2_1 _07914_ (.A(net2425),
    .B(_02033_),
    .Y(_02671_));
 sg13g2_nand2b_1 _07915_ (.Y(_02672_),
    .B(_02028_),
    .A_N(net2421));
 sg13g2_nor2_1 _07916_ (.A(net2437),
    .B(_02016_),
    .Y(_02673_));
 sg13g2_nand2b_1 _07917_ (.Y(_02674_),
    .B(_02673_),
    .A_N(net2311));
 sg13g2_o21ai_1 _07918_ (.B1(_02674_),
    .Y(_02675_),
    .A1(net2417),
    .A2(_02020_));
 sg13g2_nand2_1 _07919_ (.Y(_02676_),
    .A(_02031_),
    .B(_02675_));
 sg13g2_a21oi_1 _07920_ (.A1(_02672_),
    .A2(_02676_),
    .Y(_02677_),
    .B1(_02036_));
 sg13g2_nor2_2 _07921_ (.A(_02671_),
    .B(_02677_),
    .Y(_02678_));
 sg13g2_a21oi_1 _07922_ (.A1(_02670_),
    .A2(_02678_),
    .Y(_02679_),
    .B1(_02055_));
 sg13g2_a221oi_1 _07923_ (.B2(_02678_),
    .C1(_02055_),
    .B1(_02670_),
    .A1(_02070_),
    .Y(_02680_),
    .A2(_02072_));
 sg13g2_nor2_1 _07924_ (.A(_02084_),
    .B(_02090_),
    .Y(_02681_));
 sg13g2_or3_1 _07925_ (.A(_00999_),
    .B(_02079_),
    .C(_02080_),
    .X(_02682_));
 sg13g2_nor2_1 _07926_ (.A(_01064_),
    .B(_02052_),
    .Y(_02683_));
 sg13g2_and2_1 _07927_ (.A(_02073_),
    .B(_02683_),
    .X(_02684_));
 sg13g2_a21o_1 _07928_ (.A2(_02068_),
    .A1(_01112_),
    .B1(_02684_),
    .X(_02685_));
 sg13g2_nand2_1 _07929_ (.Y(_02686_),
    .A(_02085_),
    .B(_02685_));
 sg13g2_a21oi_1 _07930_ (.A1(_02682_),
    .A2(_02686_),
    .Y(_02687_),
    .B1(_02090_));
 sg13g2_nor3_1 _07931_ (.A(_01141_),
    .B(_02079_),
    .C(_02086_),
    .Y(_02688_));
 sg13g2_or2_1 _07932_ (.X(_02689_),
    .B(_02688_),
    .A(_02687_));
 sg13g2_a21o_1 _07933_ (.A2(_02681_),
    .A1(_02680_),
    .B1(_02689_),
    .X(_02690_));
 sg13g2_a21oi_1 _07934_ (.A1(_02078_),
    .A2(_02690_),
    .Y(_02691_),
    .B1(_02655_));
 sg13g2_nor2_1 _07935_ (.A(_02063_),
    .B(_02691_),
    .Y(_02692_));
 sg13g2_o21ai_1 _07936_ (.B1(_02095_),
    .Y(_02693_),
    .A1(_02654_),
    .A2(_02692_));
 sg13g2_nor3_1 _07937_ (.A(_02095_),
    .B(_02654_),
    .C(_02692_),
    .Y(_02694_));
 sg13g2_nand2_1 _07938_ (.Y(_02695_),
    .A(net2498),
    .B(_02693_));
 sg13g2_nor2_1 _07939_ (.A(_01245_),
    .B(_01427_),
    .Y(_02696_));
 sg13g2_o21ai_1 _07940_ (.B1(_02106_),
    .Y(_02697_),
    .A1(_01245_),
    .A2(_01427_));
 sg13g2_nor3_1 _07941_ (.A(_01245_),
    .B(_01427_),
    .C(_02105_),
    .Y(_02698_));
 sg13g2_a21oi_1 _07942_ (.A1(_02104_),
    .A2(_02697_),
    .Y(_02699_),
    .B1(_02051_));
 sg13g2_nor2b_1 _07943_ (.A(_02030_),
    .B_N(_02035_),
    .Y(_02700_));
 sg13g2_a21oi_2 _07944_ (.B1(_02046_),
    .Y(_02701_),
    .A2(_02047_),
    .A1(_02042_));
 sg13g2_nand2_1 _07945_ (.Y(_02702_),
    .A(_02017_),
    .B(_02021_));
 sg13g2_nand2_1 _07946_ (.Y(_02703_),
    .A(_02022_),
    .B(_02702_));
 sg13g2_a22oi_1 _07947_ (.Y(_02704_),
    .B1(_02702_),
    .B2(_02022_),
    .A2(_02701_),
    .A1(_02024_));
 sg13g2_or2_1 _07948_ (.X(_02705_),
    .B(_02704_),
    .A(_02038_));
 sg13g2_o21ai_1 _07949_ (.B1(_02705_),
    .Y(_02706_),
    .A1(_02034_),
    .A2(_02700_));
 sg13g2_nor2_1 _07950_ (.A(_02699_),
    .B(_02706_),
    .Y(_02707_));
 sg13g2_o21ai_1 _07951_ (.B1(_02055_),
    .Y(_02708_),
    .A1(_02699_),
    .A2(_02706_));
 sg13g2_nand2_1 _07952_ (.Y(_02709_),
    .A(_02054_),
    .B(_02708_));
 sg13g2_a21oi_1 _07953_ (.A1(_02054_),
    .A2(_02708_),
    .Y(_02710_),
    .B1(_02071_));
 sg13g2_nor2_1 _07954_ (.A(_02069_),
    .B(_02710_),
    .Y(_02711_));
 sg13g2_o21ai_1 _07955_ (.B1(_02084_),
    .Y(_02712_),
    .A1(_02069_),
    .A2(_02710_));
 sg13g2_nand3_1 _07956_ (.B(_02089_),
    .C(_02712_),
    .A(_02083_),
    .Y(_02713_));
 sg13g2_nand3_1 _07957_ (.B(_02088_),
    .C(_02713_),
    .A(_02077_),
    .Y(_02714_));
 sg13g2_and2_1 _07958_ (.A(_02116_),
    .B(_02714_),
    .X(_02715_));
 sg13g2_o21ai_1 _07959_ (.B1(_02095_),
    .Y(_02716_),
    .A1(_02061_),
    .A2(_02715_));
 sg13g2_a221oi_1 _07960_ (.B2(_02714_),
    .C1(_02095_),
    .B1(_02116_),
    .A1(net2416),
    .Y(_02717_),
    .A2(_02060_));
 sg13g2_nor2_1 _07961_ (.A(net2488),
    .B(_02717_),
    .Y(_02718_));
 sg13g2_nand2_1 _07962_ (.Y(_02719_),
    .A(net2478),
    .B(_02095_));
 sg13g2_nand2_1 _07963_ (.Y(_02720_),
    .A(net2399),
    .B(_02450_));
 sg13g2_a21oi_1 _07964_ (.A1(_01054_),
    .A2(net2402),
    .Y(_02721_),
    .B1(net2480));
 sg13g2_nor2_1 _07965_ (.A(net2403),
    .B(_01452_),
    .Y(_02722_));
 sg13g2_a221oi_1 _07966_ (.B2(_02454_),
    .C1(net2485),
    .B1(net2308),
    .A1(_02720_),
    .Y(_02723_),
    .A2(net2310));
 sg13g2_nand2_1 _07967_ (.Y(_02724_),
    .A(_01485_),
    .B(_02461_));
 sg13g2_a21oi_1 _07968_ (.A1(_01064_),
    .A2(net2336),
    .Y(_02725_),
    .B1(_01441_));
 sg13g2_nand2_1 _07969_ (.Y(_02726_),
    .A(net2352),
    .B(_02725_));
 sg13g2_mux2_1 _07970_ (.A0(_01112_),
    .A1(_00998_),
    .S(net2335),
    .X(_02727_));
 sg13g2_nand2_1 _07971_ (.Y(_02728_),
    .A(net2346),
    .B(_02727_));
 sg13g2_and2_1 _07972_ (.A(_02726_),
    .B(_02728_),
    .X(_02729_));
 sg13g2_o21ai_1 _07973_ (.B1(net2348),
    .Y(_02730_),
    .A1(_01153_),
    .A2(net2339));
 sg13g2_nand2b_1 _07974_ (.Y(_02731_),
    .B(_01435_),
    .A_N(_02730_));
 sg13g2_mux2_1 _07975_ (.A0(_01140_),
    .A1(_01126_),
    .S(net2337),
    .X(_02732_));
 sg13g2_a21oi_1 _07976_ (.A1(net2351),
    .A2(_02732_),
    .Y(_02733_),
    .B1(net2362));
 sg13g2_a221oi_1 _07977_ (.B2(_02733_),
    .C1(net2380),
    .B1(_02731_),
    .A1(net2362),
    .Y(_02734_),
    .A2(_02729_));
 sg13g2_mux2_1 _07978_ (.A0(_01082_),
    .A1(_01014_),
    .S(net2333),
    .X(_02735_));
 sg13g2_mux2_1 _07979_ (.A0(net2418),
    .A1(_01105_),
    .S(net2336),
    .X(_02736_));
 sg13g2_mux2_1 _07980_ (.A0(_02735_),
    .A1(_02736_),
    .S(net2347),
    .X(_02737_));
 sg13g2_o21ai_1 _07981_ (.B1(_01439_),
    .Y(_02738_),
    .A1(_01058_),
    .A2(net2337));
 sg13g2_nor2_1 _07982_ (.A(net2352),
    .B(_02738_),
    .Y(_02739_));
 sg13g2_a21oi_1 _07983_ (.A1(net2353),
    .A2(_01474_),
    .Y(_02740_),
    .B1(_02739_));
 sg13g2_mux2_1 _07984_ (.A0(_02737_),
    .A1(_02740_),
    .S(net2363),
    .X(_02741_));
 sg13g2_o21ai_1 _07985_ (.B1(net2317),
    .Y(_02742_),
    .A1(net2395),
    .A2(_02741_));
 sg13g2_o21ai_1 _07986_ (.B1(_02724_),
    .Y(_02743_),
    .A1(_02734_),
    .A2(_02742_));
 sg13g2_o21ai_1 _07987_ (.B1(_02719_),
    .Y(_02744_),
    .A1(_02723_),
    .A2(_02743_));
 sg13g2_a221oi_1 _07988_ (.B2(_01386_),
    .C1(net2633),
    .B1(_02744_),
    .A1(_02716_),
    .Y(_02745_),
    .A2(_02718_));
 sg13g2_o21ai_1 _07989_ (.B1(_02745_),
    .Y(_02746_),
    .A1(_02694_),
    .A2(_02695_));
 sg13g2_a21o_1 _07990_ (.A2(_02746_),
    .A1(_02653_),
    .B1(net2627),
    .X(_02747_));
 sg13g2_and2_1 _07991_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[28] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[29] ),
    .X(_02748_));
 sg13g2_and2_1 _07992_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[26] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[27] ),
    .X(_02749_));
 sg13g2_xnor2_1 _07993_ (.Y(_02750_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[26] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[26] ));
 sg13g2_nor2_1 _07994_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[25] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[25] ),
    .Y(_02751_));
 sg13g2_nand2_1 _07995_ (.Y(_02752_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[25] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[25] ));
 sg13g2_nand2_1 _07996_ (.Y(_02753_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[22] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[24] ));
 sg13g2_xor2_1 _07997_ (.B(\ChiselTop.wild.cpu.decExReg_pc[23] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[22] ),
    .X(_02754_));
 sg13g2_nand2_1 _07998_ (.Y(_02755_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[22] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[22] ));
 sg13g2_xor2_1 _07999_ (.B(\ChiselTop.wild.cpu.decExReg_pc[22] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[22] ),
    .X(_02756_));
 sg13g2_nand2_1 _08000_ (.Y(_02757_),
    .A(_02754_),
    .B(_02756_));
 sg13g2_nand2_1 _08001_ (.Y(_02758_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[21] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[21] ));
 sg13g2_nor2_1 _08002_ (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[21] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[21] ),
    .Y(_02759_));
 sg13g2_xnor2_1 _08003_ (.Y(_02760_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[21] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[21] ));
 sg13g2_xnor2_1 _08004_ (.Y(_02761_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[14] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[19] ));
 sg13g2_nand2_1 _08005_ (.Y(_02762_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[14] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[18] ));
 sg13g2_xnor2_1 _08006_ (.Y(_02763_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[14] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[18] ));
 sg13g2_nor2_1 _08007_ (.A(_02761_),
    .B(_02763_),
    .Y(_02764_));
 sg13g2_xnor2_1 _08008_ (.Y(_02765_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[17] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[17] ));
 sg13g2_nor4_2 _08009_ (.A(_01495_),
    .B(_01496_),
    .C(_01543_),
    .Y(_02766_),
    .D(_02765_));
 sg13g2_a22oi_1 _08010_ (.Y(_02767_),
    .B1(\ChiselTop.wild.cpu.decExReg_decOut_imm[17] ),
    .B2(\ChiselTop.wild.cpu.decExReg_pc[17] ),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[16] ),
    .A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[16] ));
 sg13g2_a21oi_1 _08011_ (.A1(_00936_),
    .A2(_00940_),
    .Y(_02768_),
    .B1(_02767_));
 sg13g2_a22oi_1 _08012_ (.Y(_02769_),
    .B1(_02764_),
    .B2(_02768_),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[19] ),
    .A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[14] ));
 sg13g2_inv_1 _08013_ (.Y(_02770_),
    .A(_02769_));
 sg13g2_a221oi_1 _08014_ (.B2(_02766_),
    .C1(_02770_),
    .B1(_02764_),
    .A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[14] ),
    .Y(_02771_),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[18] ));
 sg13g2_nand2_1 _08015_ (.Y(_02772_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[20] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[20] ));
 sg13g2_xor2_1 _08016_ (.B(\ChiselTop.wild.cpu.decExReg_pc[20] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[20] ),
    .X(_02773_));
 sg13g2_inv_1 _08017_ (.Y(_02774_),
    .A(_02773_));
 sg13g2_nand2b_1 _08018_ (.Y(_02775_),
    .B(_02773_),
    .A_N(_02771_));
 sg13g2_nor2_1 _08019_ (.A(_02760_),
    .B(_02775_),
    .Y(_02776_));
 sg13g2_nor4_2 _08020_ (.A(_02757_),
    .B(_02760_),
    .C(_02771_),
    .Y(_02777_),
    .D(_02774_));
 sg13g2_o21ai_1 _08021_ (.B1(_02758_),
    .Y(_02778_),
    .A1(_02759_),
    .A2(_02772_));
 sg13g2_nand2b_1 _08022_ (.Y(_02779_),
    .B(_02778_),
    .A_N(_02757_));
 sg13g2_o21ai_1 _08023_ (.B1(\ChiselTop.wild.cpu.decExReg_decOut_imm[22] ),
    .Y(_02780_),
    .A1(\ChiselTop.wild.cpu.decExReg_pc[23] ),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[22] ));
 sg13g2_nand2_1 _08024_ (.Y(_02781_),
    .A(_02779_),
    .B(_02780_));
 sg13g2_nor2_1 _08025_ (.A(_02777_),
    .B(_02781_),
    .Y(_02782_));
 sg13g2_xor2_1 _08026_ (.B(\ChiselTop.wild.cpu.decExReg_pc[24] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[22] ),
    .X(_02783_));
 sg13g2_o21ai_1 _08027_ (.B1(_02783_),
    .Y(_02784_),
    .A1(_02777_),
    .A2(_02781_));
 sg13g2_nand2_1 _08028_ (.Y(_02785_),
    .A(_02753_),
    .B(_02784_));
 sg13g2_and3_1 _08029_ (.X(_02786_),
    .A(_02752_),
    .B(_02753_),
    .C(_02784_));
 sg13g2_nor2b_1 _08030_ (.A(_02751_),
    .B_N(_02752_),
    .Y(_02787_));
 sg13g2_nor3_1 _08031_ (.A(_02750_),
    .B(_02751_),
    .C(_02786_),
    .Y(_02788_));
 sg13g2_xor2_1 _08032_ (.B(\ChiselTop.wild.cpu.decExReg_pc[27] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[26] ),
    .X(_02789_));
 sg13g2_a221oi_1 _08033_ (.B2(_02789_),
    .C1(_02749_),
    .B1(_02788_),
    .A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[26] ),
    .Y(_02790_),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[26] ));
 sg13g2_xnor2_1 _08034_ (.Y(_02791_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[28] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[28] ));
 sg13g2_nor2_1 _08035_ (.A(_02790_),
    .B(_02791_),
    .Y(_02792_));
 sg13g2_xor2_1 _08036_ (.B(\ChiselTop.wild.cpu.decExReg_pc[29] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[28] ),
    .X(_02793_));
 sg13g2_a221oi_1 _08037_ (.B2(_02793_),
    .C1(_02748_),
    .B1(_02792_),
    .A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[28] ),
    .Y(_02794_),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[28] ));
 sg13g2_xor2_1 _08038_ (.B(\ChiselTop.wild.cpu.decExReg_pc[30] ),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[28] ),
    .X(_02795_));
 sg13g2_nor2b_1 _08039_ (.A(_02794_),
    .B_N(_02795_),
    .Y(_02796_));
 sg13g2_xor2_1 _08040_ (.B(_02795_),
    .A(_02794_),
    .X(_02797_));
 sg13g2_a21oi_1 _08041_ (.A1(net2630),
    .A2(_02797_),
    .Y(_02798_),
    .B1(net2173));
 sg13g2_a21oi_2 _08042_ (.B1(\ChiselTop.wild.cpu.decExReg_func3[1] ),
    .Y(_02799_),
    .A2(_01240_),
    .A1(net2612));
 sg13g2_a21oi_1 _08043_ (.A1(\ChiselTop.wild.dmem.MEM_3[0][6] ),
    .A2(net2503),
    .Y(_02800_),
    .B1(_01221_));
 sg13g2_o21ai_1 _08044_ (.B1(_01239_),
    .Y(_02801_),
    .A1(_02799_),
    .A2(_02800_));
 sg13g2_a22oi_1 _08045_ (.Y(_02802_),
    .B1(_02801_),
    .B2(net2185),
    .A2(_02798_),
    .A1(_02747_));
 sg13g2_mux2_2 _08046_ (.A0(_02652_),
    .A1(_02802_),
    .S(net2547),
    .X(_02803_));
 sg13g2_mux4_1 _08047_ (.S0(net2694),
    .A0(\ChiselTop.wild.cpu.regs[0][30] ),
    .A1(\ChiselTop.wild.cpu.regs[1][30] ),
    .A2(\ChiselTop.wild.cpu.regs[2][30] ),
    .A3(\ChiselTop.wild.cpu.regs[3][30] ),
    .S1(net2671),
    .X(_02804_));
 sg13g2_nor2_1 _08048_ (.A(net2657),
    .B(_02804_),
    .Y(_02805_));
 sg13g2_nor2b_1 _08049_ (.A(\ChiselTop.wild.cpu.regs[5][30] ),
    .B_N(net2697),
    .Y(_02806_));
 sg13g2_nor2_1 _08050_ (.A(net2697),
    .B(\ChiselTop.wild.cpu.regs[4][30] ),
    .Y(_02807_));
 sg13g2_nor3_1 _08051_ (.A(net2673),
    .B(_02806_),
    .C(_02807_),
    .Y(_02808_));
 sg13g2_nor2b_1 _08052_ (.A(\ChiselTop.wild.cpu.regs[7][30] ),
    .B_N(net2697),
    .Y(_02809_));
 sg13g2_o21ai_1 _08053_ (.B1(net2673),
    .Y(_02810_),
    .A1(net2697),
    .A2(\ChiselTop.wild.cpu.regs[6][30] ));
 sg13g2_o21ai_1 _08054_ (.B1(net2658),
    .Y(_02811_),
    .A1(_02809_),
    .A2(_02810_));
 sg13g2_o21ai_1 _08055_ (.B1(net2469),
    .Y(_02812_),
    .A1(_02808_),
    .A2(_02811_));
 sg13g2_nor2_1 _08056_ (.A(_02805_),
    .B(_02812_),
    .Y(_02813_));
 sg13g2_nor2_1 _08057_ (.A(net2444),
    .B(_02813_),
    .Y(_02814_));
 sg13g2_a21oi_1 _08058_ (.A1(net2444),
    .A2(net2076),
    .Y(_02815_),
    .B1(_02814_));
 sg13g2_a21o_2 _08059_ (.A2(_00961_),
    .A1(\ChiselTop.wild.cpu._GEN_176[6] ),
    .B1(_02440_),
    .X(_02816_));
 sg13g2_and2_1 _08060_ (.A(net2639),
    .B(_00128_),
    .X(_02817_));
 sg13g2_nand2_1 _08061_ (.Y(_02818_),
    .A(net2639),
    .B(_00128_));
 sg13g2_o21ai_1 _08062_ (.B1(net2309),
    .Y(_02819_),
    .A1(net2402),
    .A2(_02397_));
 sg13g2_nand2b_1 _08063_ (.Y(_02820_),
    .B(net2307),
    .A_N(_02399_));
 sg13g2_nand3_1 _08064_ (.B(_02819_),
    .C(_02820_),
    .A(net2481),
    .Y(_02821_));
 sg13g2_mux2_1 _08065_ (.A0(net2422),
    .A1(net2430),
    .S(net2334),
    .X(_02822_));
 sg13g2_o21ai_1 _08066_ (.B1(_01606_),
    .Y(_02823_),
    .A1(_01159_),
    .A2(net2334));
 sg13g2_mux2_1 _08067_ (.A0(_02822_),
    .A1(_02823_),
    .S(net2345),
    .X(_02824_));
 sg13g2_mux2_1 _08068_ (.A0(_02504_),
    .A1(_02824_),
    .S(net2367),
    .X(_02825_));
 sg13g2_o21ai_1 _08069_ (.B1(_01605_),
    .Y(_02826_),
    .A1(_01015_),
    .A2(net2333));
 sg13g2_mux2_1 _08070_ (.A0(net2421),
    .A1(net2424),
    .S(net2334),
    .X(_02827_));
 sg13g2_mux2_1 _08071_ (.A0(_02826_),
    .A1(_02827_),
    .S(net2345),
    .X(_02828_));
 sg13g2_nand2_1 _08072_ (.Y(_02829_),
    .A(net2360),
    .B(_02828_));
 sg13g2_o21ai_1 _08073_ (.B1(_01579_),
    .Y(_02830_),
    .A1(_01064_),
    .A2(net2336));
 sg13g2_a21oi_1 _08074_ (.A1(_01140_),
    .A2(net2335),
    .Y(_02831_),
    .B1(_01578_));
 sg13g2_nand2_1 _08075_ (.Y(_02832_),
    .A(net2346),
    .B(_02831_));
 sg13g2_o21ai_1 _08076_ (.B1(_02832_),
    .Y(_02833_),
    .A1(net2346),
    .A2(_02830_));
 sg13g2_a21oi_1 _08077_ (.A1(net2367),
    .A2(_02833_),
    .Y(_02834_),
    .B1(net2379));
 sg13g2_a21oi_1 _08078_ (.A1(_02829_),
    .A2(_02834_),
    .Y(_02835_),
    .B1(net2314));
 sg13g2_o21ai_1 _08079_ (.B1(_02835_),
    .Y(_02836_),
    .A1(net2387),
    .A2(_02825_));
 sg13g2_o21ai_1 _08080_ (.B1(_02836_),
    .Y(_02837_),
    .A1(_01486_),
    .A2(_02406_));
 sg13g2_nor2_2 _08081_ (.A(net2474),
    .B(_02837_),
    .Y(_02838_));
 sg13g2_o21ai_1 _08082_ (.B1(net2487),
    .Y(_02839_),
    .A1(net2473),
    .A2(_02090_));
 sg13g2_a21oi_1 _08083_ (.A1(_02821_),
    .A2(_02838_),
    .Y(_02840_),
    .B1(_02839_));
 sg13g2_a21oi_1 _08084_ (.A1(_02083_),
    .A2(_02712_),
    .Y(_02841_),
    .B1(_02090_));
 sg13g2_and3_1 _08085_ (.X(_02842_),
    .A(_02083_),
    .B(_02090_),
    .C(_02712_));
 sg13g2_nor3_1 _08086_ (.A(net2487),
    .B(_02841_),
    .C(_02842_),
    .Y(_02843_));
 sg13g2_o21ai_1 _08087_ (.B1(net2495),
    .Y(_02844_),
    .A1(_02840_),
    .A2(_02843_));
 sg13g2_o21ai_1 _08088_ (.B1(_02085_),
    .Y(_02845_),
    .A1(_02680_),
    .A2(_02685_));
 sg13g2_and3_1 _08089_ (.X(_02846_),
    .A(_02090_),
    .B(_02682_),
    .C(_02845_));
 sg13g2_a21oi_1 _08090_ (.A1(_02682_),
    .A2(_02845_),
    .Y(_02847_),
    .B1(_02090_));
 sg13g2_o21ai_1 _08091_ (.B1(net2497),
    .Y(_02848_),
    .A1(_02846_),
    .A2(_02847_));
 sg13g2_a21oi_1 _08092_ (.A1(_02844_),
    .A2(_02848_),
    .Y(_02849_),
    .B1(net2632));
 sg13g2_o21ai_1 _08093_ (.B1(_00925_),
    .Y(_02850_),
    .A1(_02817_),
    .A2(_02849_));
 sg13g2_a21oi_1 _08094_ (.A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[26] ),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[26] ),
    .Y(_02851_),
    .B1(_02788_));
 sg13g2_xor2_1 _08095_ (.B(_02851_),
    .A(_02789_),
    .X(_02852_));
 sg13g2_a21oi_1 _08096_ (.A1(net2630),
    .A2(_02852_),
    .Y(_02853_),
    .B1(net2173));
 sg13g2_a21oi_1 _08097_ (.A1(\ChiselTop.wild.cpu.decExReg_memLow[1] ),
    .A2(_01230_),
    .Y(_02854_),
    .B1(\ChiselTop.wild.cpu.decExReg_memLow[0] ));
 sg13g2_nor3_1 _08098_ (.A(_01178_),
    .B(_02229_),
    .C(_02854_),
    .Y(_02855_));
 sg13g2_and2_1 _08099_ (.A(net2611),
    .B(_02228_),
    .X(_02856_));
 sg13g2_nand2_1 _08100_ (.Y(_02857_),
    .A(_01177_),
    .B(_01225_));
 sg13g2_a21oi_1 _08101_ (.A1(\ChiselTop.wild.dmem.MEM_1[0][7] ),
    .A2(net2503),
    .Y(_02858_),
    .B1(_02857_));
 sg13g2_nor4_1 _08102_ (.A(_02301_),
    .B(_02855_),
    .C(_02856_),
    .D(_02858_),
    .Y(_02859_));
 sg13g2_a21oi_1 _08103_ (.A1(_02850_),
    .A2(_02853_),
    .Y(_02860_),
    .B1(_02859_));
 sg13g2_xnor2_1 _08104_ (.Y(_02861_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[27] ),
    .B(_02647_));
 sg13g2_mux2_1 _08105_ (.A0(_02860_),
    .A1(_02861_),
    .S(net2618),
    .X(_02862_));
 sg13g2_mux4_1 _08106_ (.S0(net2692),
    .A0(\ChiselTop.wild.cpu.regs[0][27] ),
    .A1(\ChiselTop.wild.cpu.regs[1][27] ),
    .A2(\ChiselTop.wild.cpu.regs[2][27] ),
    .A3(\ChiselTop.wild.cpu.regs[3][27] ),
    .S1(net2670),
    .X(_02863_));
 sg13g2_nor2_1 _08107_ (.A(net2659),
    .B(_02863_),
    .Y(_02864_));
 sg13g2_nor2b_1 _08108_ (.A(\ChiselTop.wild.cpu.regs[5][27] ),
    .B_N(net2693),
    .Y(_02865_));
 sg13g2_nor2_1 _08109_ (.A(net2693),
    .B(\ChiselTop.wild.cpu.regs[4][27] ),
    .Y(_02866_));
 sg13g2_nor3_1 _08110_ (.A(net2670),
    .B(_02865_),
    .C(_02866_),
    .Y(_02867_));
 sg13g2_nor2b_1 _08111_ (.A(\ChiselTop.wild.cpu.regs[7][27] ),
    .B_N(net2693),
    .Y(_02868_));
 sg13g2_o21ai_1 _08112_ (.B1(net2670),
    .Y(_02869_),
    .A1(net2693),
    .A2(\ChiselTop.wild.cpu.regs[6][27] ));
 sg13g2_o21ai_1 _08113_ (.B1(net2659),
    .Y(_02870_),
    .A1(_02868_),
    .A2(_02869_));
 sg13g2_o21ai_1 _08114_ (.B1(net2468),
    .Y(_02871_),
    .A1(_02867_),
    .A2(_02870_));
 sg13g2_nor2_1 _08115_ (.A(_02864_),
    .B(_02871_),
    .Y(_02872_));
 sg13g2_nor2_1 _08116_ (.A(net2443),
    .B(_02872_),
    .Y(_02873_));
 sg13g2_a21oi_2 _08117_ (.B1(_02873_),
    .Y(_02874_),
    .A2(net2089),
    .A1(net2443));
 sg13g2_nand2b_1 _08118_ (.Y(_02875_),
    .B(_01922_),
    .A_N(_01241_));
 sg13g2_o21ai_1 _08119_ (.B1(_02875_),
    .Y(_02876_),
    .A1(net2611),
    .A2(_01240_));
 sg13g2_nor2_1 _08120_ (.A(_01178_),
    .B(_01240_),
    .Y(_02877_));
 sg13g2_a21oi_1 _08121_ (.A1(_01176_),
    .A2(_02876_),
    .Y(_02878_),
    .B1(_02301_));
 sg13g2_nor3_1 _08122_ (.A(_02085_),
    .B(_02680_),
    .C(_02685_),
    .Y(_02879_));
 sg13g2_nand3b_1 _08123_ (.B(net2497),
    .C(_02845_),
    .Y(_02880_),
    .A_N(_02879_));
 sg13g2_o21ai_1 _08124_ (.B1(net2310),
    .Y(_02881_),
    .A1(net2403),
    .A2(_02263_));
 sg13g2_nand3_1 _08125_ (.B(_01887_),
    .C(net2308),
    .A(net2390),
    .Y(_02882_));
 sg13g2_nand3_1 _08126_ (.B(_02881_),
    .C(_02882_),
    .A(net2482),
    .Y(_02883_));
 sg13g2_nand2_1 _08127_ (.Y(_02884_),
    .A(net2361),
    .B(_02737_));
 sg13g2_a21oi_1 _08128_ (.A1(net2369),
    .A2(_02729_),
    .Y(_02885_),
    .B1(net2380));
 sg13g2_and2_1 _08129_ (.A(net2364),
    .B(_02458_),
    .X(_02886_));
 sg13g2_a21oi_1 _08130_ (.A1(net2372),
    .A2(_02740_),
    .Y(_02887_),
    .B1(_02886_));
 sg13g2_a221oi_1 _08131_ (.B2(net2380),
    .C1(net2314),
    .B1(_02887_),
    .A1(_02884_),
    .Y(_02888_),
    .A2(_02885_));
 sg13g2_a21oi_1 _08132_ (.A1(net2313),
    .A2(_02274_),
    .Y(_02889_),
    .B1(_02888_));
 sg13g2_nand3_1 _08133_ (.B(_02883_),
    .C(_02889_),
    .A(net2471),
    .Y(_02890_));
 sg13g2_a21oi_1 _08134_ (.A1(net2479),
    .A2(_02085_),
    .Y(_02891_),
    .B1(net2493));
 sg13g2_nand2_1 _08135_ (.Y(_02892_),
    .A(_02890_),
    .B(_02891_));
 sg13g2_xnor2_1 _08136_ (.Y(_02893_),
    .A(_02084_),
    .B(_02711_));
 sg13g2_o21ai_1 _08137_ (.B1(_02892_),
    .Y(_02894_),
    .A1(net2487),
    .A2(_02893_));
 sg13g2_nand3_1 _08138_ (.B(_02880_),
    .C(_02894_),
    .A(net2531),
    .Y(_02895_));
 sg13g2_a21oi_1 _08139_ (.A1(_02818_),
    .A2(_02895_),
    .Y(_02896_),
    .B1(net2629));
 sg13g2_o21ai_1 _08140_ (.B1(_02750_),
    .Y(_02897_),
    .A1(_02751_),
    .A2(_02786_));
 sg13g2_nand2b_1 _08141_ (.Y(_02898_),
    .B(_02897_),
    .A_N(_02788_));
 sg13g2_a21oi_1 _08142_ (.A1(net2629),
    .A2(_02898_),
    .Y(_02899_),
    .B1(_02896_));
 sg13g2_a21o_1 _08143_ (.A2(_02899_),
    .A1(_01547_),
    .B1(_02878_),
    .X(_02900_));
 sg13g2_nor2_1 _08144_ (.A(\ChiselTop.wild.cpu.decExReg_pc[26] ),
    .B(_02646_),
    .Y(_02901_));
 sg13g2_nor3_1 _08145_ (.A(net2545),
    .B(_02647_),
    .C(_02901_),
    .Y(_02902_));
 sg13g2_a21oi_2 _08146_ (.B1(_02902_),
    .Y(_02903_),
    .A2(_02900_),
    .A1(net2546));
 sg13g2_mux4_1 _08147_ (.S0(net2702),
    .A0(\ChiselTop.wild.cpu.regs[0][26] ),
    .A1(\ChiselTop.wild.cpu.regs[1][26] ),
    .A2(\ChiselTop.wild.cpu.regs[2][26] ),
    .A3(\ChiselTop.wild.cpu.regs[3][26] ),
    .S1(net2675),
    .X(_02904_));
 sg13g2_nor2_1 _08148_ (.A(net2661),
    .B(_02904_),
    .Y(_02905_));
 sg13g2_nor2b_1 _08149_ (.A(\ChiselTop.wild.cpu.regs[5][26] ),
    .B_N(net2701),
    .Y(_02906_));
 sg13g2_nor2_1 _08150_ (.A(net2701),
    .B(\ChiselTop.wild.cpu.regs[4][26] ),
    .Y(_02907_));
 sg13g2_nor3_1 _08151_ (.A(net2675),
    .B(_02906_),
    .C(_02907_),
    .Y(_02908_));
 sg13g2_nor2b_1 _08152_ (.A(\ChiselTop.wild.cpu.regs[7][26] ),
    .B_N(net2702),
    .Y(_02909_));
 sg13g2_o21ai_1 _08153_ (.B1(net2675),
    .Y(_02910_),
    .A1(net2701),
    .A2(\ChiselTop.wild.cpu.regs[6][26] ));
 sg13g2_o21ai_1 _08154_ (.B1(net2661),
    .Y(_02911_),
    .A1(_02909_),
    .A2(_02910_));
 sg13g2_o21ai_1 _08155_ (.B1(net2469),
    .Y(_02912_),
    .A1(_02908_),
    .A2(_02911_));
 sg13g2_nor2_1 _08156_ (.A(_02905_),
    .B(_02912_),
    .Y(_02913_));
 sg13g2_nor2_1 _08157_ (.A(net2444),
    .B(_02913_),
    .Y(_02914_));
 sg13g2_a21oi_1 _08158_ (.A1(net2444),
    .A2(net2084),
    .Y(_02915_),
    .B1(_02914_));
 sg13g2_or2_1 _08159_ (.X(_02916_),
    .B(_02915_),
    .A(_02874_));
 sg13g2_and2_1 _08160_ (.A(_02816_),
    .B(_02916_),
    .X(_02917_));
 sg13g2_a21oi_1 _08161_ (.A1(_02874_),
    .A2(_02915_),
    .Y(_02918_),
    .B1(_02816_));
 sg13g2_a21oi_2 _08162_ (.B1(_02440_),
    .Y(_02919_),
    .A2(_00961_),
    .A1(net1528));
 sg13g2_a21o_1 _08163_ (.A2(_00961_),
    .A1(\ChiselTop.wild.cpu._GEN_176[5] ),
    .B1(_02440_),
    .X(_02920_));
 sg13g2_a21oi_1 _08164_ (.A1(\ChiselTop.wild.cpu.decExReg_pc[24] ),
    .A2(_02645_),
    .Y(_02921_),
    .B1(\ChiselTop.wild.cpu.decExReg_pc[25] ));
 sg13g2_o21ai_1 _08165_ (.B1(net2618),
    .Y(_02922_),
    .A1(_02646_),
    .A2(_02921_));
 sg13g2_o21ai_1 _08166_ (.B1(_01242_),
    .Y(_02923_),
    .A1(_01224_),
    .A2(_01974_));
 sg13g2_nand2_1 _08167_ (.Y(_02924_),
    .A(net2185),
    .B(_02923_));
 sg13g2_nand2b_1 _08168_ (.Y(_02925_),
    .B(net2397),
    .A_N(_02348_));
 sg13g2_a221oi_1 _08169_ (.B2(net2309),
    .C1(net2484),
    .B1(_02925_),
    .A1(_02353_),
    .Y(_02926_),
    .A2(net2307));
 sg13g2_mux2_1 _08170_ (.A0(_02823_),
    .A1(_02826_),
    .S(net2344),
    .X(_02927_));
 sg13g2_nor2_1 _08171_ (.A(net2345),
    .B(_02827_),
    .Y(_02928_));
 sg13g2_a21oi_1 _08172_ (.A1(net2344),
    .A2(_02830_),
    .Y(_02929_),
    .B1(_02928_));
 sg13g2_nand2_1 _08173_ (.Y(_02930_),
    .A(net2368),
    .B(_02929_));
 sg13g2_a21oi_1 _08174_ (.A1(net2361),
    .A2(_02927_),
    .Y(_02931_),
    .B1(net2378));
 sg13g2_mux2_1 _08175_ (.A0(_02503_),
    .A1(_02822_),
    .S(net2344),
    .X(_02932_));
 sg13g2_and2_1 _08176_ (.A(net2368),
    .B(_02932_),
    .X(_02933_));
 sg13g2_a21oi_1 _08177_ (.A1(net2360),
    .A2(_02547_),
    .Y(_02934_),
    .B1(_02933_));
 sg13g2_a221oi_1 _08178_ (.B2(net2378),
    .C1(net2314),
    .B1(_02934_),
    .A1(_02930_),
    .Y(_02935_),
    .A2(_02931_));
 sg13g2_o21ai_1 _08179_ (.B1(net2471),
    .Y(_02936_),
    .A1(_01486_),
    .A2(_02361_));
 sg13g2_nor3_2 _08180_ (.A(_02926_),
    .B(_02935_),
    .C(_02936_),
    .Y(_02937_));
 sg13g2_a21oi_1 _08181_ (.A1(net2478),
    .A2(_02073_),
    .Y(_02938_),
    .B1(_02937_));
 sg13g2_o21ai_1 _08182_ (.B1(net2493),
    .Y(_02939_),
    .A1(_02073_),
    .A2(_02709_));
 sg13g2_a21oi_1 _08183_ (.A1(_02073_),
    .A2(_02709_),
    .Y(_02940_),
    .B1(_02939_));
 sg13g2_a21oi_1 _08184_ (.A1(net2487),
    .A2(_02938_),
    .Y(_02941_),
    .B1(_02940_));
 sg13g2_nor3_1 _08185_ (.A(_02073_),
    .B(_02679_),
    .C(_02683_),
    .Y(_02942_));
 sg13g2_nor4_1 _08186_ (.A(net2495),
    .B(_02680_),
    .C(_02684_),
    .D(_02942_),
    .Y(_02943_));
 sg13g2_nor3_2 _08187_ (.A(net2632),
    .B(_02941_),
    .C(_02943_),
    .Y(_02944_));
 sg13g2_a21oi_1 _08188_ (.A1(net2639),
    .A2(_00129_),
    .Y(_02945_),
    .B1(_02944_));
 sg13g2_xnor2_1 _08189_ (.Y(_02946_),
    .A(_02785_),
    .B(_02787_));
 sg13g2_a21oi_1 _08190_ (.A1(net2629),
    .A2(_02946_),
    .Y(_02947_),
    .B1(net2173));
 sg13g2_o21ai_1 _08191_ (.B1(_02947_),
    .Y(_02948_),
    .A1(net2629),
    .A2(_02945_));
 sg13g2_nand2_1 _08192_ (.Y(_02949_),
    .A(_02924_),
    .B(_02948_));
 sg13g2_o21ai_1 _08193_ (.B1(_02922_),
    .Y(_02950_),
    .A1(net2619),
    .A2(_02949_));
 sg13g2_mux4_1 _08194_ (.S0(net2681),
    .A0(\ChiselTop.wild.cpu.regs[0][25] ),
    .A1(\ChiselTop.wild.cpu.regs[1][25] ),
    .A2(\ChiselTop.wild.cpu.regs[2][25] ),
    .A3(\ChiselTop.wild.cpu.regs[3][25] ),
    .S1(net2663),
    .X(_02951_));
 sg13g2_nor2_1 _08195_ (.A(net2651),
    .B(_02951_),
    .Y(_02952_));
 sg13g2_nor2b_1 _08196_ (.A(\ChiselTop.wild.cpu.regs[5][25] ),
    .B_N(net2681),
    .Y(_02953_));
 sg13g2_nor2_1 _08197_ (.A(net2681),
    .B(\ChiselTop.wild.cpu.regs[4][25] ),
    .Y(_02954_));
 sg13g2_nor3_1 _08198_ (.A(net2663),
    .B(_02953_),
    .C(_02954_),
    .Y(_02955_));
 sg13g2_nor2b_1 _08199_ (.A(\ChiselTop.wild.cpu.regs[7][25] ),
    .B_N(net2681),
    .Y(_02956_));
 sg13g2_o21ai_1 _08200_ (.B1(net2664),
    .Y(_02957_),
    .A1(net2681),
    .A2(\ChiselTop.wild.cpu.regs[6][25] ));
 sg13g2_o21ai_1 _08201_ (.B1(net2651),
    .Y(_02958_),
    .A1(_02956_),
    .A2(_02957_));
 sg13g2_o21ai_1 _08202_ (.B1(net2466),
    .Y(_02959_),
    .A1(_02955_),
    .A2(_02958_));
 sg13g2_nor2_2 _08203_ (.A(_02952_),
    .B(_02959_),
    .Y(_02960_));
 sg13g2_nor2_1 _08204_ (.A(net2443),
    .B(_02960_),
    .Y(_02961_));
 sg13g2_a21oi_2 _08205_ (.B1(_02961_),
    .Y(_02962_),
    .A2(net2083),
    .A1(net2443));
 sg13g2_inv_1 _08206_ (.Y(_02963_),
    .A(_02962_));
 sg13g2_o21ai_1 _08207_ (.B1(_00964_),
    .Y(_02964_),
    .A1(_00119_),
    .A2(net2522));
 sg13g2_nor2_2 _08208_ (.A(_02301_),
    .B(_02877_),
    .Y(_02965_));
 sg13g2_a21o_1 _08209_ (.A2(net2503),
    .A1(\ChiselTop.wild.dmem.MEM_2[0][7] ),
    .B1(_01224_),
    .X(_02966_));
 sg13g2_nand2_1 _08210_ (.Y(_02967_),
    .A(net2638),
    .B(_00130_));
 sg13g2_nand2_1 _08211_ (.Y(_02968_),
    .A(net2397),
    .B(_01587_));
 sg13g2_nor2b_1 _08212_ (.A(_01592_),
    .B_N(net2307),
    .Y(_02969_));
 sg13g2_a21oi_1 _08213_ (.A1(net2309),
    .A2(_02968_),
    .Y(_02970_),
    .B1(_02969_));
 sg13g2_mux2_1 _08214_ (.A0(_02824_),
    .A1(_02828_),
    .S(net2367),
    .X(_02971_));
 sg13g2_nor2_1 _08215_ (.A(net2379),
    .B(_02971_),
    .Y(_02972_));
 sg13g2_a21oi_1 _08216_ (.A1(net2379),
    .A2(_02506_),
    .Y(_02973_),
    .B1(_02972_));
 sg13g2_o21ai_1 _08217_ (.B1(net2471),
    .Y(_02974_),
    .A1(_01486_),
    .A2(_01625_));
 sg13g2_a221oi_1 _08218_ (.B2(net2316),
    .C1(_02974_),
    .B1(_02973_),
    .A1(net2482),
    .Y(_02975_),
    .A2(_02970_));
 sg13g2_nor2_1 _08219_ (.A(net2490),
    .B(_02975_),
    .Y(_02976_));
 sg13g2_o21ai_1 _08220_ (.B1(_02976_),
    .Y(_02977_),
    .A1(net2473),
    .A2(_02036_));
 sg13g2_a21oi_1 _08221_ (.A1(_02104_),
    .A2(_02697_),
    .Y(_02978_),
    .B1(_02044_));
 sg13g2_nor4_2 _08222_ (.A(_02044_),
    .B(_02048_),
    .C(_02107_),
    .Y(_02979_),
    .D(_02698_));
 sg13g2_o21ai_1 _08223_ (.B1(_02024_),
    .Y(_02980_),
    .A1(_02701_),
    .A2(_02979_));
 sg13g2_a21oi_1 _08224_ (.A1(_02703_),
    .A2(_02980_),
    .Y(_02981_),
    .B1(_02031_));
 sg13g2_o21ai_1 _08225_ (.B1(_02037_),
    .Y(_02982_),
    .A1(_02030_),
    .A2(_02981_));
 sg13g2_nor3_1 _08226_ (.A(_02030_),
    .B(_02037_),
    .C(_02981_),
    .Y(_02983_));
 sg13g2_nand3b_1 _08227_ (.B(net2492),
    .C(_02982_),
    .Y(_02984_),
    .A_N(_02983_));
 sg13g2_a21oi_1 _08228_ (.A1(_02977_),
    .A2(_02984_),
    .Y(_02985_),
    .B1(net2498));
 sg13g2_a221oi_1 _08229_ (.B2(_02667_),
    .C1(net2312),
    .B1(_02662_),
    .A1(_02021_),
    .Y(_02986_),
    .A2(_02022_));
 sg13g2_o21ai_1 _08230_ (.B1(_02031_),
    .Y(_02987_),
    .A1(_02675_),
    .A2(_02986_));
 sg13g2_nand3_1 _08231_ (.B(_02672_),
    .C(_02987_),
    .A(_02036_),
    .Y(_02988_));
 sg13g2_a21o_1 _08232_ (.A2(_02987_),
    .A1(_02672_),
    .B1(_02036_),
    .X(_02989_));
 sg13g2_a21oi_1 _08233_ (.A1(_02988_),
    .A2(_02989_),
    .Y(_02990_),
    .B1(net2495));
 sg13g2_o21ai_1 _08234_ (.B1(net2530),
    .Y(_02991_),
    .A1(_02985_),
    .A2(_02990_));
 sg13g2_a21o_1 _08235_ (.A2(_02991_),
    .A1(_02967_),
    .B1(net2627),
    .X(_02992_));
 sg13g2_o21ai_1 _08236_ (.B1(_02756_),
    .Y(_02993_),
    .A1(_02776_),
    .A2(_02778_));
 sg13g2_nand2_1 _08237_ (.Y(_02994_),
    .A(_02755_),
    .B(_02993_));
 sg13g2_xnor2_1 _08238_ (.Y(_02995_),
    .A(_02754_),
    .B(_02994_));
 sg13g2_a21oi_1 _08239_ (.A1(net2629),
    .A2(_02995_),
    .Y(_02996_),
    .B1(net2172));
 sg13g2_a22oi_1 _08240_ (.Y(_02997_),
    .B1(_02992_),
    .B2(_02996_),
    .A2(_02966_),
    .A1(_02965_));
 sg13g2_a21oi_1 _08241_ (.A1(\ChiselTop.wild.cpu.decExReg_pc[22] ),
    .A2(_02644_),
    .Y(_02998_),
    .B1(\ChiselTop.wild.cpu.decExReg_pc[23] ));
 sg13g2_or2_1 _08242_ (.X(_02999_),
    .B(_02998_),
    .A(_02645_));
 sg13g2_mux2_1 _08243_ (.A0(_02997_),
    .A1(_02999_),
    .S(net2614),
    .X(_03000_));
 sg13g2_inv_1 _08244_ (.Y(_03001_),
    .A(net2092));
 sg13g2_mux4_1 _08245_ (.S0(net2684),
    .A0(\ChiselTop.wild.cpu.regs[0][23] ),
    .A1(\ChiselTop.wild.cpu.regs[1][23] ),
    .A2(\ChiselTop.wild.cpu.regs[2][23] ),
    .A3(\ChiselTop.wild.cpu.regs[3][23] ),
    .S1(net2666),
    .X(_03002_));
 sg13g2_nor2_2 _08246_ (.A(net2653),
    .B(_03002_),
    .Y(_03003_));
 sg13g2_nor2b_1 _08247_ (.A(\ChiselTop.wild.cpu.regs[5][23] ),
    .B_N(net2685),
    .Y(_03004_));
 sg13g2_nor2_1 _08248_ (.A(net2684),
    .B(\ChiselTop.wild.cpu.regs[4][23] ),
    .Y(_03005_));
 sg13g2_nor3_1 _08249_ (.A(net2666),
    .B(_03004_),
    .C(_03005_),
    .Y(_03006_));
 sg13g2_nor2b_1 _08250_ (.A(\ChiselTop.wild.cpu.regs[7][23] ),
    .B_N(net2684),
    .Y(_03007_));
 sg13g2_o21ai_1 _08251_ (.B1(net2666),
    .Y(_03008_),
    .A1(net2684),
    .A2(\ChiselTop.wild.cpu.regs[6][23] ));
 sg13g2_o21ai_1 _08252_ (.B1(net2653),
    .Y(_03009_),
    .A1(_03007_),
    .A2(_03008_));
 sg13g2_o21ai_1 _08253_ (.B1(net2467),
    .Y(_03010_),
    .A1(_03006_),
    .A2(_03009_));
 sg13g2_nor2_2 _08254_ (.A(_03003_),
    .B(_03010_),
    .Y(_03011_));
 sg13g2_nor2_1 _08255_ (.A(net2439),
    .B(_03011_),
    .Y(_03012_));
 sg13g2_a21oi_2 _08256_ (.B1(_03012_),
    .Y(_03013_),
    .A2(net2092),
    .A1(net2439));
 sg13g2_or2_1 _08257_ (.X(_03014_),
    .B(_02645_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[24] ));
 sg13g2_o21ai_1 _08258_ (.B1(_01242_),
    .Y(_03015_),
    .A1(_01224_),
    .A2(_02159_));
 sg13g2_nand2_1 _08259_ (.Y(_03016_),
    .A(net2183),
    .B(_03015_));
 sg13g2_and3_1 _08260_ (.X(_03017_),
    .A(_02055_),
    .B(_02670_),
    .C(_02678_));
 sg13g2_o21ai_1 _08261_ (.B1(net2497),
    .Y(_03018_),
    .A1(_02679_),
    .A2(_03017_));
 sg13g2_nand2_1 _08262_ (.Y(_03019_),
    .A(net2399),
    .B(_02307_));
 sg13g2_a221oi_1 _08263_ (.B2(net2310),
    .C1(net2485),
    .B1(_03019_),
    .A1(_02306_),
    .Y(_03020_),
    .A2(net2308));
 sg13g2_mux2_1 _08264_ (.A0(_02735_),
    .A1(_02738_),
    .S(net2352),
    .X(_03021_));
 sg13g2_nor2_1 _08265_ (.A(net2347),
    .B(_02736_),
    .Y(_03022_));
 sg13g2_a21oi_1 _08266_ (.A1(net2347),
    .A2(_02725_),
    .Y(_03023_),
    .B1(_03022_));
 sg13g2_a21o_1 _08267_ (.A2(_03023_),
    .A1(net2369),
    .B1(net2378),
    .X(_03024_));
 sg13g2_a21oi_1 _08268_ (.A1(net2362),
    .A2(_03021_),
    .Y(_03025_),
    .B1(_03024_));
 sg13g2_o21ai_1 _08269_ (.B1(net2316),
    .Y(_03026_),
    .A1(net2394),
    .A2(_01477_));
 sg13g2_nor2_1 _08270_ (.A(_01486_),
    .B(_02313_),
    .Y(_03027_));
 sg13g2_o21ai_1 _08271_ (.B1(net2471),
    .Y(_03028_),
    .A1(_03025_),
    .A2(_03026_));
 sg13g2_nor3_2 _08272_ (.A(_03020_),
    .B(_03027_),
    .C(_03028_),
    .Y(_03029_));
 sg13g2_a21oi_1 _08273_ (.A1(net2478),
    .A2(_02056_),
    .Y(_03030_),
    .B1(_03029_));
 sg13g2_xnor2_1 _08274_ (.Y(_03031_),
    .A(_02056_),
    .B(_02707_));
 sg13g2_a22oi_1 _08275_ (.Y(_03032_),
    .B1(_03031_),
    .B2(net2493),
    .A2(_03030_),
    .A1(_01386_));
 sg13g2_a21o_1 _08276_ (.A2(_03032_),
    .A1(_03018_),
    .B1(net2632),
    .X(_03033_));
 sg13g2_a21oi_1 _08277_ (.A1(_02967_),
    .A2(_03033_),
    .Y(_03034_),
    .B1(net2627));
 sg13g2_xor2_1 _08278_ (.B(_02783_),
    .A(_02782_),
    .X(_03035_));
 sg13g2_a21o_1 _08279_ (.A2(_03035_),
    .A1(net2629),
    .B1(net2172),
    .X(_03036_));
 sg13g2_o21ai_1 _08280_ (.B1(_03016_),
    .Y(_03037_),
    .A1(_03034_),
    .A2(_03036_));
 sg13g2_a21oi_1 _08281_ (.A1(\ChiselTop.wild.cpu.decExReg_pc[24] ),
    .A2(_02645_),
    .Y(_03038_),
    .B1(net2545));
 sg13g2_a22oi_1 _08282_ (.Y(_03039_),
    .B1(_03038_),
    .B2(_03014_),
    .A2(_03037_),
    .A1(net2545));
 sg13g2_mux4_1 _08283_ (.S0(net2694),
    .A0(\ChiselTop.wild.cpu.regs[0][24] ),
    .A1(\ChiselTop.wild.cpu.regs[1][24] ),
    .A2(\ChiselTop.wild.cpu.regs[2][24] ),
    .A3(\ChiselTop.wild.cpu.regs[3][24] ),
    .S1(net2671),
    .X(_03040_));
 sg13g2_nor2_1 _08284_ (.A(net2659),
    .B(_03040_),
    .Y(_03041_));
 sg13g2_nor2b_1 _08285_ (.A(\ChiselTop.wild.cpu.regs[5][24] ),
    .B_N(net2702),
    .Y(_03042_));
 sg13g2_nor2_1 _08286_ (.A(net2702),
    .B(\ChiselTop.wild.cpu.regs[4][24] ),
    .Y(_03043_));
 sg13g2_nor3_1 _08287_ (.A(net2675),
    .B(_03042_),
    .C(_03043_),
    .Y(_03044_));
 sg13g2_nor2b_1 _08288_ (.A(\ChiselTop.wild.cpu.regs[7][24] ),
    .B_N(net2705),
    .Y(_03045_));
 sg13g2_o21ai_1 _08289_ (.B1(net2675),
    .Y(_03046_),
    .A1(net2702),
    .A2(\ChiselTop.wild.cpu.regs[6][24] ));
 sg13g2_o21ai_1 _08290_ (.B1(net2658),
    .Y(_03047_),
    .A1(_03045_),
    .A2(_03046_));
 sg13g2_o21ai_1 _08291_ (.B1(net2469),
    .Y(_03048_),
    .A1(_03044_),
    .A2(_03047_));
 sg13g2_nor2_1 _08292_ (.A(_03041_),
    .B(_03048_),
    .Y(_03049_));
 sg13g2_nor2_1 _08293_ (.A(net2443),
    .B(_03049_),
    .Y(_03050_));
 sg13g2_a21oi_1 _08294_ (.A1(net2443),
    .A2(net2096),
    .Y(_03051_),
    .B1(_03050_));
 sg13g2_or3_1 _08295_ (.A(_02031_),
    .B(_02675_),
    .C(_02986_),
    .X(_03052_));
 sg13g2_a21oi_1 _08296_ (.A1(_02987_),
    .A2(_03052_),
    .Y(_03053_),
    .B1(net2495));
 sg13g2_nand3_1 _08297_ (.B(_02703_),
    .C(_02980_),
    .A(_02031_),
    .Y(_03054_));
 sg13g2_nor2_1 _08298_ (.A(net2488),
    .B(_02981_),
    .Y(_03055_));
 sg13g2_nand2_1 _08299_ (.Y(_03056_),
    .A(net2398),
    .B(_01676_));
 sg13g2_a221oi_1 _08300_ (.B2(net2310),
    .C1(net2485),
    .B1(_03056_),
    .A1(_01672_),
    .Y(_03057_),
    .A2(net2308));
 sg13g2_mux2_1 _08301_ (.A0(_02459_),
    .A1(_02741_),
    .S(net2394),
    .X(_03058_));
 sg13g2_a221oi_1 _08302_ (.B2(_01478_),
    .C1(_03057_),
    .B1(_03058_),
    .A1(_01485_),
    .Y(_03059_),
    .A2(_01696_));
 sg13g2_nor2_1 _08303_ (.A(net2475),
    .B(_03059_),
    .Y(_03060_));
 sg13g2_a21oi_1 _08304_ (.A1(net2478),
    .A2(_02032_),
    .Y(_03061_),
    .B1(_03060_));
 sg13g2_a221oi_1 _08305_ (.B2(net2488),
    .C1(net2498),
    .B1(_03061_),
    .A1(_03054_),
    .Y(_03062_),
    .A2(_03055_));
 sg13g2_o21ai_1 _08306_ (.B1(net2530),
    .Y(_03063_),
    .A1(_03053_),
    .A2(_03062_));
 sg13g2_a21oi_1 _08307_ (.A1(_02967_),
    .A2(_03063_),
    .Y(_03064_),
    .B1(net2627));
 sg13g2_or3_1 _08308_ (.A(_02756_),
    .B(_02776_),
    .C(_02778_),
    .X(_03065_));
 sg13g2_nand2_1 _08309_ (.Y(_03066_),
    .A(_02993_),
    .B(_03065_));
 sg13g2_a21o_1 _08310_ (.A2(_03066_),
    .A1(net2629),
    .B1(net2172),
    .X(_03067_));
 sg13g2_a21o_1 _08311_ (.A2(net2503),
    .A1(\ChiselTop.wild.dmem.MEM_2[0][6] ),
    .B1(_01241_),
    .X(_03068_));
 sg13g2_a22oi_1 _08312_ (.Y(_03069_),
    .B1(_02965_),
    .B2(_03068_),
    .A2(net2322),
    .A1(net2183));
 sg13g2_o21ai_1 _08313_ (.B1(_03069_),
    .Y(_03070_),
    .A1(_03064_),
    .A2(_03067_));
 sg13g2_or2_1 _08314_ (.X(_03071_),
    .B(_02644_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[22] ));
 sg13g2_a21oi_1 _08315_ (.A1(\ChiselTop.wild.cpu.decExReg_pc[22] ),
    .A2(_02644_),
    .Y(_03072_),
    .B1(net2543));
 sg13g2_a22oi_1 _08316_ (.Y(_03073_),
    .B1(_03071_),
    .B2(_03072_),
    .A2(_03070_),
    .A1(net2543));
 sg13g2_mux4_1 _08317_ (.S0(net2679),
    .A0(\ChiselTop.wild.cpu.regs[0][22] ),
    .A1(\ChiselTop.wild.cpu.regs[1][22] ),
    .A2(\ChiselTop.wild.cpu.regs[2][22] ),
    .A3(\ChiselTop.wild.cpu.regs[3][22] ),
    .S1(net2662),
    .X(_03074_));
 sg13g2_nor2_2 _08318_ (.A(net2652),
    .B(_03074_),
    .Y(_03075_));
 sg13g2_nor2b_1 _08319_ (.A(\ChiselTop.wild.cpu.regs[5][22] ),
    .B_N(net2679),
    .Y(_03076_));
 sg13g2_nor2_1 _08320_ (.A(net2679),
    .B(\ChiselTop.wild.cpu.regs[4][22] ),
    .Y(_03077_));
 sg13g2_nor3_1 _08321_ (.A(net2662),
    .B(_03076_),
    .C(_03077_),
    .Y(_03078_));
 sg13g2_nor2b_1 _08322_ (.A(\ChiselTop.wild.cpu.regs[7][22] ),
    .B_N(net2679),
    .Y(_03079_));
 sg13g2_o21ai_1 _08323_ (.B1(net2662),
    .Y(_03080_),
    .A1(net2678),
    .A2(\ChiselTop.wild.cpu.regs[6][22] ));
 sg13g2_o21ai_1 _08324_ (.B1(net2652),
    .Y(_03081_),
    .A1(_03079_),
    .A2(_03080_));
 sg13g2_o21ai_1 _08325_ (.B1(net2466),
    .Y(_03082_),
    .A1(_03078_),
    .A2(_03081_));
 sg13g2_nor2_2 _08326_ (.A(_03075_),
    .B(_03082_),
    .Y(_03083_));
 sg13g2_nor2_1 _08327_ (.A(net2439),
    .B(_03083_),
    .Y(_03084_));
 sg13g2_a21oi_2 _08328_ (.B1(_03084_),
    .Y(_03085_),
    .A2(net2095),
    .A1(net2439));
 sg13g2_and2_1 _08329_ (.A(_03051_),
    .B(_03085_),
    .X(_03086_));
 sg13g2_a21oi_1 _08330_ (.A1(_03013_),
    .A2(_03086_),
    .Y(_03087_),
    .B1(_02964_));
 sg13g2_a21o_2 _08331_ (.A2(_00961_),
    .A1(\ChiselTop.wild.cpu._GEN_176[1] ),
    .B1(_02440_),
    .X(_03088_));
 sg13g2_xnor2_1 _08332_ (.Y(_03089_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[21] ),
    .B(_02643_));
 sg13g2_o21ai_1 _08333_ (.B1(net2309),
    .Y(_03090_),
    .A1(net2402),
    .A2(_01748_));
 sg13g2_a21oi_1 _08334_ (.A1(_01761_),
    .A2(net2307),
    .Y(_03091_),
    .B1(net2484));
 sg13g2_nand2_1 _08335_ (.Y(_03092_),
    .A(_03090_),
    .B(_03091_));
 sg13g2_and2_1 _08336_ (.A(net2368),
    .B(_02927_),
    .X(_03093_));
 sg13g2_a21oi_1 _08337_ (.A1(net2361),
    .A2(_02932_),
    .Y(_03094_),
    .B1(_03093_));
 sg13g2_nor2_1 _08338_ (.A(net2387),
    .B(_02548_),
    .Y(_03095_));
 sg13g2_a21oi_1 _08339_ (.A1(net2387),
    .A2(_03094_),
    .Y(_03096_),
    .B1(_03095_));
 sg13g2_a221oi_1 _08340_ (.B2(net2316),
    .C1(net2474),
    .B1(_03096_),
    .A1(net2313),
    .Y(_03097_),
    .A2(_01768_));
 sg13g2_a21oi_2 _08341_ (.B1(net2490),
    .Y(_03098_),
    .A2(_03097_),
    .A1(_03092_));
 sg13g2_o21ai_1 _08342_ (.B1(_03098_),
    .Y(_03099_),
    .A1(net2473),
    .A2(net2311));
 sg13g2_o21ai_1 _08343_ (.B1(_02018_),
    .Y(_03100_),
    .A1(_02701_),
    .A2(_02979_));
 sg13g2_nand3_1 _08344_ (.B(net2311),
    .C(_03100_),
    .A(_02017_),
    .Y(_03101_));
 sg13g2_a21o_1 _08345_ (.A2(_03100_),
    .A1(_02017_),
    .B1(net2311),
    .X(_03102_));
 sg13g2_nand3_1 _08346_ (.B(_03101_),
    .C(_03102_),
    .A(net2492),
    .Y(_03103_));
 sg13g2_nor2b_1 _08347_ (.A(_02673_),
    .B_N(net2311),
    .Y(_03104_));
 sg13g2_o21ai_1 _08348_ (.B1(_03104_),
    .Y(_03105_),
    .A1(net2312),
    .A2(_02668_));
 sg13g2_nand2_1 _08349_ (.Y(_03106_),
    .A(net2498),
    .B(_02674_));
 sg13g2_nor2_1 _08350_ (.A(_02986_),
    .B(_03106_),
    .Y(_03107_));
 sg13g2_and2_1 _08351_ (.A(net2638),
    .B(_00131_),
    .X(_03108_));
 sg13g2_a221oi_1 _08352_ (.B2(_03107_),
    .C1(net2634),
    .B1(_03105_),
    .A1(_03099_),
    .Y(_03109_),
    .A2(_03103_));
 sg13g2_o21ai_1 _08353_ (.B1(net2529),
    .Y(_03110_),
    .A1(_03108_),
    .A2(_03109_));
 sg13g2_nand2_1 _08354_ (.Y(_03111_),
    .A(_02772_),
    .B(_02775_));
 sg13g2_xor2_1 _08355_ (.B(_03111_),
    .A(_02760_),
    .X(_03112_));
 sg13g2_a21oi_1 _08356_ (.A1(net2629),
    .A2(_03112_),
    .Y(_03113_),
    .B1(net2172));
 sg13g2_a21oi_1 _08357_ (.A1(\ChiselTop.wild.dmem.MEM_2[0][5] ),
    .A2(net2502),
    .Y(_03114_),
    .B1(_01221_));
 sg13g2_o21ai_1 _08358_ (.B1(_01239_),
    .Y(_03115_),
    .A1(_02799_),
    .A2(_03114_));
 sg13g2_a22oi_1 _08359_ (.Y(_03116_),
    .B1(_03115_),
    .B2(net2183),
    .A2(_03113_),
    .A1(_03110_));
 sg13g2_mux2_1 _08360_ (.A0(_03089_),
    .A1(_03116_),
    .S(net2544),
    .X(_03117_));
 sg13g2_inv_1 _08361_ (.Y(_03118_),
    .A(net2104));
 sg13g2_mux4_1 _08362_ (.S0(net2687),
    .A0(\ChiselTop.wild.cpu.regs[0][21] ),
    .A1(\ChiselTop.wild.cpu.regs[1][21] ),
    .A2(\ChiselTop.wild.cpu.regs[2][21] ),
    .A3(\ChiselTop.wild.cpu.regs[3][21] ),
    .S1(net2667),
    .X(_03119_));
 sg13g2_nor2_1 _08363_ (.A(net2654),
    .B(_03119_),
    .Y(_03120_));
 sg13g2_nor2b_1 _08364_ (.A(\ChiselTop.wild.cpu.regs[5][21] ),
    .B_N(net2686),
    .Y(_03121_));
 sg13g2_nor2_1 _08365_ (.A(net2686),
    .B(\ChiselTop.wild.cpu.regs[4][21] ),
    .Y(_03122_));
 sg13g2_nor3_1 _08366_ (.A(net2667),
    .B(_03121_),
    .C(_03122_),
    .Y(_03123_));
 sg13g2_nor2b_1 _08367_ (.A(\ChiselTop.wild.cpu.regs[7][21] ),
    .B_N(net2686),
    .Y(_03124_));
 sg13g2_o21ai_1 _08368_ (.B1(net2666),
    .Y(_03125_),
    .A1(net2686),
    .A2(\ChiselTop.wild.cpu.regs[6][21] ));
 sg13g2_o21ai_1 _08369_ (.B1(net2653),
    .Y(_03126_),
    .A1(_03124_),
    .A2(_03125_));
 sg13g2_o21ai_1 _08370_ (.B1(net2467),
    .Y(_03127_),
    .A1(_03123_),
    .A2(_03126_));
 sg13g2_nor2_2 _08371_ (.A(_03120_),
    .B(_03127_),
    .Y(_03128_));
 sg13g2_nor2_1 _08372_ (.A(net2440),
    .B(_03128_),
    .Y(_03129_));
 sg13g2_a21oi_2 _08373_ (.B1(_03129_),
    .Y(_03130_),
    .A2(net2104),
    .A1(net2441));
 sg13g2_nor2_1 _08374_ (.A(_03088_),
    .B(_03130_),
    .Y(_03131_));
 sg13g2_or2_1 _08375_ (.X(_03132_),
    .B(_03130_),
    .A(_03088_));
 sg13g2_o21ai_1 _08376_ (.B1(_00964_),
    .Y(_03133_),
    .A1(net1548),
    .A2(net2522));
 sg13g2_xnor2_1 _08377_ (.Y(_03134_),
    .A(_00939_),
    .B(_02642_));
 sg13g2_nor3_1 _08378_ (.A(net2312),
    .B(_02701_),
    .C(_02979_),
    .Y(_03135_));
 sg13g2_nand3b_1 _08379_ (.B(net2492),
    .C(_03100_),
    .Y(_03136_),
    .A_N(_03135_));
 sg13g2_nand2_1 _08380_ (.Y(_03137_),
    .A(net2398),
    .B(_01839_));
 sg13g2_a221oi_1 _08381_ (.B2(net2310),
    .C1(net2485),
    .B1(_03137_),
    .A1(_01838_),
    .Y(_03138_),
    .A2(net2308));
 sg13g2_mux2_1 _08382_ (.A0(_01475_),
    .A1(_03021_),
    .S(net2369),
    .X(_03139_));
 sg13g2_nor2_1 _08383_ (.A(net2382),
    .B(_03139_),
    .Y(_03140_));
 sg13g2_a21oi_1 _08384_ (.A1(net2382),
    .A2(_02598_),
    .Y(_03141_),
    .B1(_03140_));
 sg13g2_a221oi_1 _08385_ (.B2(net2317),
    .C1(_03138_),
    .B1(_03141_),
    .A1(net2313),
    .Y(_03142_),
    .A2(_01854_));
 sg13g2_a21oi_1 _08386_ (.A1(net2478),
    .A2(net2312),
    .Y(_03143_),
    .B1(net2492));
 sg13g2_o21ai_1 _08387_ (.B1(_03143_),
    .Y(_03144_),
    .A1(net2478),
    .A2(_03142_));
 sg13g2_nand3_1 _08388_ (.B(_03136_),
    .C(_03144_),
    .A(net2495),
    .Y(_03145_));
 sg13g2_xor2_1 _08389_ (.B(_02668_),
    .A(net2312),
    .X(_03146_));
 sg13g2_o21ai_1 _08390_ (.B1(_03145_),
    .Y(_03147_),
    .A1(net2496),
    .A2(_03146_));
 sg13g2_a21oi_1 _08391_ (.A1(net2638),
    .A2(_00935_),
    .Y(_03148_),
    .B1(net2623));
 sg13g2_o21ai_1 _08392_ (.B1(_03148_),
    .Y(_03149_),
    .A1(net2638),
    .A2(_03147_));
 sg13g2_xnor2_1 _08393_ (.Y(_03150_),
    .A(_02771_),
    .B(_02773_));
 sg13g2_nor2_1 _08394_ (.A(net2529),
    .B(_03150_),
    .Y(_03151_));
 sg13g2_nor2_1 _08395_ (.A(net2172),
    .B(_03151_),
    .Y(_03152_));
 sg13g2_a22oi_1 _08396_ (.Y(_03153_),
    .B1(_02854_),
    .B2(_01177_),
    .A2(net2502),
    .A1(\ChiselTop.wild.dmem.MEM_2[0][4] ));
 sg13g2_nor3_1 _08397_ (.A(_02301_),
    .B(_02877_),
    .C(_03153_),
    .Y(_03154_));
 sg13g2_a221oi_1 _08398_ (.B2(_03152_),
    .C1(_03154_),
    .B1(_03149_),
    .A1(net2183),
    .Y(_03155_),
    .A2(net2322));
 sg13g2_mux2_1 _08399_ (.A0(_03134_),
    .A1(_03155_),
    .S(net2542),
    .X(_03156_));
 sg13g2_inv_1 _08400_ (.Y(_03157_),
    .A(net2101));
 sg13g2_mux4_1 _08401_ (.S0(net2688),
    .A0(\ChiselTop.wild.cpu.regs[0][20] ),
    .A1(\ChiselTop.wild.cpu.regs[1][20] ),
    .A2(\ChiselTop.wild.cpu.regs[2][20] ),
    .A3(\ChiselTop.wild.cpu.regs[3][20] ),
    .S1(net2667),
    .X(_03158_));
 sg13g2_nor2_1 _08402_ (.A(net2653),
    .B(_03158_),
    .Y(_03159_));
 sg13g2_nor2b_1 _08403_ (.A(\ChiselTop.wild.cpu.regs[5][20] ),
    .B_N(net2685),
    .Y(_03160_));
 sg13g2_nor2_1 _08404_ (.A(net2685),
    .B(\ChiselTop.wild.cpu.regs[4][20] ),
    .Y(_03161_));
 sg13g2_nor3_1 _08405_ (.A(net2666),
    .B(_03160_),
    .C(_03161_),
    .Y(_03162_));
 sg13g2_nor2b_1 _08406_ (.A(\ChiselTop.wild.cpu.regs[7][20] ),
    .B_N(net2685),
    .Y(_03163_));
 sg13g2_o21ai_1 _08407_ (.B1(net2666),
    .Y(_03164_),
    .A1(net2685),
    .A2(\ChiselTop.wild.cpu.regs[6][20] ));
 sg13g2_o21ai_1 _08408_ (.B1(net2653),
    .Y(_03165_),
    .A1(_03163_),
    .A2(_03164_));
 sg13g2_o21ai_1 _08409_ (.B1(net2467),
    .Y(_03166_),
    .A1(_03162_),
    .A2(_03165_));
 sg13g2_nor2_2 _08410_ (.A(_03159_),
    .B(_03166_),
    .Y(_03167_));
 sg13g2_nor2_1 _08411_ (.A(net2440),
    .B(_03167_),
    .Y(_03168_));
 sg13g2_a21oi_1 _08412_ (.A1(net2440),
    .A2(net2101),
    .Y(_03169_),
    .B1(_03168_));
 sg13g2_a22oi_1 _08413_ (.Y(_03170_),
    .B1(_03133_),
    .B2(_03169_),
    .A2(_03130_),
    .A1(_03088_));
 sg13g2_or2_1 _08414_ (.X(_03171_),
    .B(_03170_),
    .A(_03131_));
 sg13g2_a21oi_2 _08415_ (.B1(_00963_),
    .Y(_03172_),
    .A2(_00961_),
    .A1(_00942_));
 sg13g2_inv_1 _08416_ (.Y(_03173_),
    .A(_03172_));
 sg13g2_nand2_1 _08417_ (.Y(_03174_),
    .A(_00940_),
    .B(_00986_));
 sg13g2_o21ai_1 _08418_ (.B1(_01242_),
    .Y(_03175_),
    .A1(_01224_),
    .A2(_01978_));
 sg13g2_nand3_1 _08419_ (.B(_02108_),
    .C(_02657_),
    .A(_01384_),
    .Y(_03176_));
 sg13g2_nand3_1 _08420_ (.B(_02658_),
    .C(_03176_),
    .A(net2497),
    .Y(_03177_));
 sg13g2_nand2_1 _08421_ (.Y(_03178_),
    .A(net2397),
    .B(_01944_));
 sg13g2_a22oi_1 _08422_ (.Y(_03179_),
    .B1(_03178_),
    .B2(net2309),
    .A2(net2307),
    .A1(_01955_));
 sg13g2_nand2_1 _08423_ (.Y(_03180_),
    .A(net2481),
    .B(_03179_));
 sg13g2_nor2_1 _08424_ (.A(net2387),
    .B(_02360_),
    .Y(_03181_));
 sg13g2_a21oi_1 _08425_ (.A1(net2387),
    .A2(_02934_),
    .Y(_03182_),
    .B1(_03181_));
 sg13g2_a221oi_1 _08426_ (.B2(net2316),
    .C1(net2474),
    .B1(_03182_),
    .A1(net2313),
    .Y(_03183_),
    .A2(_01959_));
 sg13g2_a21oi_2 _08427_ (.B1(net2490),
    .Y(_03184_),
    .A2(_03183_),
    .A1(_03180_));
 sg13g2_o21ai_1 _08428_ (.B1(_03184_),
    .Y(_03185_),
    .A1(net2473),
    .A2(_02108_));
 sg13g2_xnor2_1 _08429_ (.Y(_03186_),
    .A(_02108_),
    .B(_02696_));
 sg13g2_o21ai_1 _08430_ (.B1(_03185_),
    .Y(_03187_),
    .A1(net2488),
    .A2(_03186_));
 sg13g2_a21o_1 _08431_ (.A2(_03187_),
    .A1(_03177_),
    .B1(net2633),
    .X(_03188_));
 sg13g2_a21oi_1 _08432_ (.A1(net2632),
    .A2(_00937_),
    .Y(_03189_),
    .B1(net2626));
 sg13g2_a21oi_1 _08433_ (.A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[16] ),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[16] ),
    .Y(_03190_),
    .B1(_01544_));
 sg13g2_xnor2_1 _08434_ (.Y(_03191_),
    .A(_02765_),
    .B(_03190_));
 sg13g2_a221oi_1 _08435_ (.B2(net2623),
    .C1(net2171),
    .B1(_03191_),
    .A1(_03188_),
    .Y(_03192_),
    .A2(_03189_));
 sg13g2_a21o_1 _08436_ (.A2(_03175_),
    .A1(net2184),
    .B1(_03192_),
    .X(_03193_));
 sg13g2_nor2_1 _08437_ (.A(net2541),
    .B(_02641_),
    .Y(_03194_));
 sg13g2_a22oi_1 _08438_ (.Y(_03195_),
    .B1(_03194_),
    .B2(_03174_),
    .A2(_03193_),
    .A1(net2541));
 sg13g2_mux4_1 _08439_ (.S0(net2680),
    .A0(\ChiselTop.wild.cpu.regs[0][17] ),
    .A1(\ChiselTop.wild.cpu.regs[1][17] ),
    .A2(\ChiselTop.wild.cpu.regs[2][17] ),
    .A3(\ChiselTop.wild.cpu.regs[3][17] ),
    .S1(net2663),
    .X(_03196_));
 sg13g2_nor2_1 _08440_ (.A(net2651),
    .B(_03196_),
    .Y(_03197_));
 sg13g2_nor2b_1 _08441_ (.A(\ChiselTop.wild.cpu.regs[5][17] ),
    .B_N(net2680),
    .Y(_03198_));
 sg13g2_nor2_1 _08442_ (.A(net2680),
    .B(\ChiselTop.wild.cpu.regs[4][17] ),
    .Y(_03199_));
 sg13g2_nor3_1 _08443_ (.A(net2663),
    .B(_03198_),
    .C(_03199_),
    .Y(_03200_));
 sg13g2_nor2b_1 _08444_ (.A(\ChiselTop.wild.cpu.regs[7][17] ),
    .B_N(net2680),
    .Y(_03201_));
 sg13g2_o21ai_1 _08445_ (.B1(net2663),
    .Y(_03202_),
    .A1(net2680),
    .A2(\ChiselTop.wild.cpu.regs[6][17] ));
 sg13g2_o21ai_1 _08446_ (.B1(net2651),
    .Y(_03203_),
    .A1(_03201_),
    .A2(_03202_));
 sg13g2_o21ai_1 _08447_ (.B1(net2466),
    .Y(_03204_),
    .A1(_03200_),
    .A2(_03203_));
 sg13g2_nor2_1 _08448_ (.A(_03197_),
    .B(_03204_),
    .Y(_03205_));
 sg13g2_nor2_1 _08449_ (.A(net2438),
    .B(_03205_),
    .Y(_03206_));
 sg13g2_a21oi_2 _08450_ (.B1(_03206_),
    .Y(_03207_),
    .A2(net2116),
    .A1(net2442));
 sg13g2_inv_1 _08451_ (.Y(_03208_),
    .A(_03207_));
 sg13g2_a22oi_1 _08452_ (.Y(_03209_),
    .B1(_03173_),
    .B2(_03207_),
    .A2(_01567_),
    .A1(_00965_));
 sg13g2_a22oi_1 _08453_ (.Y(_03210_),
    .B1(_03209_),
    .B2(_02635_),
    .A2(_03208_),
    .A1(_03172_));
 sg13g2_nand2_1 _08454_ (.Y(_03211_),
    .A(_01223_),
    .B(_02226_));
 sg13g2_o21ai_1 _08455_ (.B1(net2309),
    .Y(_03212_),
    .A1(net2402),
    .A2(_02196_));
 sg13g2_nand2_1 _08456_ (.Y(_03213_),
    .A(_02199_),
    .B(net2307));
 sg13g2_nand3_1 _08457_ (.B(_03212_),
    .C(_03213_),
    .A(net2481),
    .Y(_03214_));
 sg13g2_a21oi_1 _08458_ (.A1(net2379),
    .A2(_02404_),
    .Y(_03215_),
    .B1(net2314));
 sg13g2_o21ai_1 _08459_ (.B1(_03215_),
    .Y(_03216_),
    .A1(net2379),
    .A2(_02825_));
 sg13g2_o21ai_1 _08460_ (.B1(net2313),
    .Y(_03217_),
    .A1(net2379),
    .A2(_02209_));
 sg13g2_nand4_1 _08461_ (.B(_03214_),
    .C(_03216_),
    .A(net2471),
    .Y(_03218_),
    .D(_03217_));
 sg13g2_a21oi_1 _08462_ (.A1(net2479),
    .A2(_02048_),
    .Y(_03219_),
    .B1(net2492));
 sg13g2_nand2_1 _08463_ (.Y(_03220_),
    .A(_03218_),
    .B(_03219_));
 sg13g2_or3_1 _08464_ (.A(_02041_),
    .B(_02048_),
    .C(_02978_),
    .X(_03221_));
 sg13g2_o21ai_1 _08465_ (.B1(_02048_),
    .Y(_03222_),
    .A1(_02041_),
    .A2(_02978_));
 sg13g2_nand3_1 _08466_ (.B(_03221_),
    .C(_03222_),
    .A(net2492),
    .Y(_03223_));
 sg13g2_nand3_1 _08467_ (.B(_02659_),
    .C(_02664_),
    .A(_02049_),
    .Y(_03224_));
 sg13g2_nor3_1 _08468_ (.A(net2496),
    .B(_02661_),
    .C(_02665_),
    .Y(_03225_));
 sg13g2_a221oi_1 _08469_ (.B2(_03225_),
    .C1(net2632),
    .B1(_03224_),
    .A1(_03220_),
    .Y(_03226_),
    .A2(_03223_));
 sg13g2_o21ai_1 _08470_ (.B1(net2529),
    .Y(_03227_),
    .A1(_02445_),
    .A2(_03226_));
 sg13g2_nor2_1 _08471_ (.A(_02766_),
    .B(_02768_),
    .Y(_03228_));
 sg13g2_o21ai_1 _08472_ (.B1(_02762_),
    .Y(_03229_),
    .A1(_02763_),
    .A2(_03228_));
 sg13g2_xor2_1 _08473_ (.B(_03229_),
    .A(_02761_),
    .X(_03230_));
 sg13g2_a21oi_1 _08474_ (.A1(net2627),
    .A2(_03230_),
    .Y(_03231_),
    .B1(net2172));
 sg13g2_a22oi_1 _08475_ (.Y(_03232_),
    .B1(_03227_),
    .B2(_03231_),
    .A2(_03211_),
    .A1(_02965_));
 sg13g2_a21o_1 _08476_ (.A2(_02641_),
    .A1(\ChiselTop.wild.cpu.decExReg_pc[18] ),
    .B1(\ChiselTop.wild.cpu.decExReg_pc[19] ),
    .X(_03233_));
 sg13g2_a21oi_1 _08477_ (.A1(_02642_),
    .A2(_03233_),
    .Y(_03234_),
    .B1(net2542));
 sg13g2_a21o_1 _08478_ (.A2(_03232_),
    .A1(net2542),
    .B1(_03234_),
    .X(_03235_));
 sg13g2_mux4_1 _08479_ (.S0(net2692),
    .A0(\ChiselTop.wild.cpu.regs[0][19] ),
    .A1(\ChiselTop.wild.cpu.regs[1][19] ),
    .A2(\ChiselTop.wild.cpu.regs[2][19] ),
    .A3(\ChiselTop.wild.cpu.regs[3][19] ),
    .S1(net2670),
    .X(_03236_));
 sg13g2_nor2_1 _08480_ (.A(net2659),
    .B(_03236_),
    .Y(_03237_));
 sg13g2_nor2b_1 _08481_ (.A(\ChiselTop.wild.cpu.regs[5][19] ),
    .B_N(net2692),
    .Y(_03238_));
 sg13g2_nor2_1 _08482_ (.A(net2692),
    .B(net1552),
    .Y(_03239_));
 sg13g2_nor3_1 _08483_ (.A(net2670),
    .B(_03238_),
    .C(_03239_),
    .Y(_03240_));
 sg13g2_nor2b_1 _08484_ (.A(\ChiselTop.wild.cpu.regs[7][19] ),
    .B_N(net2692),
    .Y(_03241_));
 sg13g2_o21ai_1 _08485_ (.B1(net2670),
    .Y(_03242_),
    .A1(net2692),
    .A2(\ChiselTop.wild.cpu.regs[6][19] ));
 sg13g2_o21ai_1 _08486_ (.B1(net2659),
    .Y(_03243_),
    .A1(_03241_),
    .A2(_03242_));
 sg13g2_o21ai_1 _08487_ (.B1(net2468),
    .Y(_03244_),
    .A1(_03240_),
    .A2(_03243_));
 sg13g2_nor2_2 _08488_ (.A(_03237_),
    .B(_03244_),
    .Y(_03245_));
 sg13g2_nor2_1 _08489_ (.A(net2443),
    .B(_03245_),
    .Y(_03246_));
 sg13g2_a21oi_1 _08490_ (.A1(net2445),
    .A2(net2110),
    .Y(_03247_),
    .B1(_03246_));
 sg13g2_nand2_1 _08491_ (.Y(_03248_),
    .A(_02440_),
    .B(_03247_));
 sg13g2_xnor2_1 _08492_ (.Y(_03249_),
    .A(_02440_),
    .B(_03247_));
 sg13g2_o21ai_1 _08493_ (.B1(_02965_),
    .Y(_03250_),
    .A1(_01224_),
    .A2(_01920_));
 sg13g2_nand3_1 _08494_ (.B(_02656_),
    .C(_02658_),
    .A(_02043_),
    .Y(_03251_));
 sg13g2_nand3_1 _08495_ (.B(_02659_),
    .C(_03251_),
    .A(net2497),
    .Y(_03252_));
 sg13g2_nand3_1 _08496_ (.B(_02104_),
    .C(_02697_),
    .A(_02044_),
    .Y(_03253_));
 sg13g2_nor2_1 _08497_ (.A(net2487),
    .B(_02978_),
    .Y(_03254_));
 sg13g2_nand2_1 _08498_ (.Y(_03255_),
    .A(net2397),
    .B(_01891_));
 sg13g2_a221oi_1 _08499_ (.B2(net2309),
    .C1(net2484),
    .B1(_03255_),
    .A1(_01888_),
    .Y(_03256_),
    .A2(net2308));
 sg13g2_nand2_1 _08500_ (.Y(_03257_),
    .A(net2394),
    .B(_02887_));
 sg13g2_a21oi_1 _08501_ (.A1(net2382),
    .A2(_02273_),
    .Y(_03258_),
    .B1(net2315));
 sg13g2_nand2_1 _08502_ (.Y(_03259_),
    .A(_03257_),
    .B(_03258_));
 sg13g2_o21ai_1 _08503_ (.B1(_03259_),
    .Y(_03260_),
    .A1(_01486_),
    .A2(_01904_));
 sg13g2_o21ai_1 _08504_ (.B1(net2471),
    .Y(_03261_),
    .A1(_03256_),
    .A2(_03260_));
 sg13g2_a21oi_1 _08505_ (.A1(net2478),
    .A2(_02043_),
    .Y(_03262_),
    .B1(net2492));
 sg13g2_a221oi_1 _08506_ (.B2(_03262_),
    .C1(net2632),
    .B1(_03261_),
    .A1(_03253_),
    .Y(_03263_),
    .A2(_03254_));
 sg13g2_a21oi_1 _08507_ (.A1(_03252_),
    .A2(_03263_),
    .Y(_03264_),
    .B1(_02445_));
 sg13g2_xnor2_1 _08508_ (.Y(_03265_),
    .A(_02763_),
    .B(_03228_));
 sg13g2_a21oi_1 _08509_ (.A1(net2623),
    .A2(_03265_),
    .Y(_03266_),
    .B1(net2171));
 sg13g2_o21ai_1 _08510_ (.B1(_03266_),
    .Y(_03267_),
    .A1(net2623),
    .A2(_03264_));
 sg13g2_nand2_1 _08511_ (.Y(_03268_),
    .A(_03250_),
    .B(_03267_));
 sg13g2_or2_1 _08512_ (.X(_03269_),
    .B(_02641_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[18] ));
 sg13g2_a21oi_1 _08513_ (.A1(\ChiselTop.wild.cpu.decExReg_pc[18] ),
    .A2(_02641_),
    .Y(_03270_),
    .B1(net2541));
 sg13g2_a22oi_1 _08514_ (.Y(_03271_),
    .B1(_03269_),
    .B2(_03270_),
    .A2(_03268_),
    .A1(net2541));
 sg13g2_mux4_1 _08515_ (.S0(net2680),
    .A0(\ChiselTop.wild.cpu.regs[0][18] ),
    .A1(\ChiselTop.wild.cpu.regs[1][18] ),
    .A2(\ChiselTop.wild.cpu.regs[2][18] ),
    .A3(\ChiselTop.wild.cpu.regs[3][18] ),
    .S1(net2663),
    .X(_03272_));
 sg13g2_nor2_2 _08516_ (.A(net2651),
    .B(_03272_),
    .Y(_03273_));
 sg13g2_nor2b_1 _08517_ (.A(\ChiselTop.wild.cpu.regs[5][18] ),
    .B_N(net2681),
    .Y(_03274_));
 sg13g2_nor2_1 _08518_ (.A(net2681),
    .B(net1553),
    .Y(_03275_));
 sg13g2_nor3_1 _08519_ (.A(net2663),
    .B(_03274_),
    .C(_03275_),
    .Y(_03276_));
 sg13g2_nor2b_1 _08520_ (.A(\ChiselTop.wild.cpu.regs[7][18] ),
    .B_N(net2680),
    .Y(_03277_));
 sg13g2_o21ai_1 _08521_ (.B1(net2663),
    .Y(_03278_),
    .A1(net2680),
    .A2(\ChiselTop.wild.cpu.regs[6][18] ));
 sg13g2_o21ai_1 _08522_ (.B1(net2651),
    .Y(_03279_),
    .A1(_03277_),
    .A2(_03278_));
 sg13g2_o21ai_1 _08523_ (.B1(net2467),
    .Y(_03280_),
    .A1(_03276_),
    .A2(_03279_));
 sg13g2_nor2_1 _08524_ (.A(_03273_),
    .B(_03280_),
    .Y(_03281_));
 sg13g2_nor2_1 _08525_ (.A(net2438),
    .B(_03281_),
    .Y(_03282_));
 sg13g2_a21oi_2 _08526_ (.B1(_03282_),
    .Y(_03283_),
    .A2(net2107),
    .A1(net2438));
 sg13g2_nand2_1 _08527_ (.Y(_03284_),
    .A(_02440_),
    .B(_03283_));
 sg13g2_xnor2_1 _08528_ (.Y(_03285_),
    .A(_02441_),
    .B(_03283_));
 sg13g2_nand2b_1 _08529_ (.Y(_03286_),
    .B(_03285_),
    .A_N(_03249_));
 sg13g2_a221oi_1 _08530_ (.B2(_02635_),
    .C1(_03286_),
    .B1(_03209_),
    .A1(_03172_),
    .Y(_03287_),
    .A2(_03208_));
 sg13g2_nand2_1 _08531_ (.Y(_03288_),
    .A(_03248_),
    .B(_03284_));
 sg13g2_or2_1 _08532_ (.X(_03289_),
    .B(_03169_),
    .A(_03133_));
 sg13g2_and3_1 _08533_ (.X(_03290_),
    .A(_03132_),
    .B(_03170_),
    .C(_03289_));
 sg13g2_o21ai_1 _08534_ (.B1(_03290_),
    .Y(_03291_),
    .A1(_03287_),
    .A2(_03288_));
 sg13g2_a21o_1 _08535_ (.A2(_03291_),
    .A1(_03171_),
    .B1(_03087_),
    .X(_03292_));
 sg13g2_or3_1 _08536_ (.A(_03013_),
    .B(_03051_),
    .C(_03085_),
    .X(_03293_));
 sg13g2_a22oi_1 _08537_ (.Y(_03294_),
    .B1(_02964_),
    .B2(_03293_),
    .A2(_02962_),
    .A1(_02920_));
 sg13g2_a221oi_1 _08538_ (.B2(_03294_),
    .C1(_02918_),
    .B1(_03292_),
    .A1(_02919_),
    .Y(_03295_),
    .A2(_02963_));
 sg13g2_or2_1 _08539_ (.X(_03296_),
    .B(_03295_),
    .A(_02917_));
 sg13g2_nor2_1 _08540_ (.A(_00135_),
    .B(_02649_),
    .Y(_03297_));
 sg13g2_xnor2_1 _08541_ (.Y(_03298_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[29] ),
    .B(_03297_));
 sg13g2_and2_2 _08542_ (.A(net2618),
    .B(_03298_),
    .X(_03299_));
 sg13g2_o21ai_1 _08543_ (.B1(net2309),
    .Y(_03300_),
    .A1(net2402),
    .A2(_02540_));
 sg13g2_nand2b_1 _08544_ (.Y(_03301_),
    .B(net2307),
    .A_N(_02544_));
 sg13g2_nand3_1 _08545_ (.B(_03300_),
    .C(_03301_),
    .A(net2481),
    .Y(_03302_));
 sg13g2_mux4_1 _08546_ (.S0(net2345),
    .A0(_00999_),
    .A1(net2419),
    .A2(_01141_),
    .A3(net2416),
    .S1(net2331),
    .X(_03303_));
 sg13g2_nand2_1 _08547_ (.Y(_03304_),
    .A(net2367),
    .B(_03303_));
 sg13g2_a21oi_1 _08548_ (.A1(net2361),
    .A2(_02929_),
    .Y(_03305_),
    .B1(net2378));
 sg13g2_a221oi_1 _08549_ (.B2(_03305_),
    .C1(net2314),
    .B1(_03304_),
    .A1(net2378),
    .Y(_03306_),
    .A2(_03094_));
 sg13g2_a21oi_1 _08550_ (.A1(net2313),
    .A2(_02550_),
    .Y(_03307_),
    .B1(_03306_));
 sg13g2_nand3_1 _08551_ (.B(_03302_),
    .C(_03307_),
    .A(net2471),
    .Y(_03308_));
 sg13g2_o21ai_1 _08552_ (.B1(_03308_),
    .Y(_03309_),
    .A1(net2473),
    .A2(_02063_));
 sg13g2_nor2_1 _08553_ (.A(net2492),
    .B(_03309_),
    .Y(_03310_));
 sg13g2_a21oi_1 _08554_ (.A1(_02076_),
    .A2(_02714_),
    .Y(_03311_),
    .B1(_02063_));
 sg13g2_and3_1 _08555_ (.X(_03312_),
    .A(_02063_),
    .B(_02076_),
    .C(_02714_));
 sg13g2_nor3_1 _08556_ (.A(net2487),
    .B(_03311_),
    .C(_03312_),
    .Y(_03313_));
 sg13g2_xnor2_1 _08557_ (.Y(_03314_),
    .A(_02064_),
    .B(_02691_));
 sg13g2_a21oi_1 _08558_ (.A1(net2497),
    .A2(_03314_),
    .Y(_03315_),
    .B1(net2632));
 sg13g2_o21ai_1 _08559_ (.B1(_03315_),
    .Y(_03316_),
    .A1(_03310_),
    .A2(_03313_));
 sg13g2_a21o_1 _08560_ (.A2(_03316_),
    .A1(_02653_),
    .B1(net2627),
    .X(_03317_));
 sg13g2_a21oi_1 _08561_ (.A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[28] ),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[28] ),
    .Y(_03318_),
    .B1(_02792_));
 sg13g2_xor2_1 _08562_ (.B(_03318_),
    .A(_02793_),
    .X(_03319_));
 sg13g2_a21oi_1 _08563_ (.A1(net2630),
    .A2(_03319_),
    .Y(_03320_),
    .B1(net2172));
 sg13g2_a21oi_1 _08564_ (.A1(_01222_),
    .A2(_01782_),
    .Y(_03321_),
    .B1(_02799_));
 sg13g2_or2_1 _08565_ (.X(_03322_),
    .B(_03321_),
    .A(net2322));
 sg13g2_a22oi_1 _08566_ (.Y(_03323_),
    .B1(_03322_),
    .B2(net2188),
    .A2(_03320_),
    .A1(_03317_));
 sg13g2_a221oi_1 _08567_ (.B2(net2185),
    .C1(net2618),
    .B1(_03322_),
    .A1(_03317_),
    .Y(_03324_),
    .A2(_03320_));
 sg13g2_or2_1 _08568_ (.X(_03325_),
    .B(_03324_),
    .A(_03299_));
 sg13g2_mux4_1 _08569_ (.S0(net2703),
    .A0(\ChiselTop.wild.cpu.regs[0][29] ),
    .A1(\ChiselTop.wild.cpu.regs[1][29] ),
    .A2(\ChiselTop.wild.cpu.regs[2][29] ),
    .A3(\ChiselTop.wild.cpu.regs[3][29] ),
    .S1(net2676),
    .X(_03326_));
 sg13g2_nor2_2 _08570_ (.A(net2660),
    .B(_03326_),
    .Y(_03327_));
 sg13g2_nor2b_1 _08571_ (.A(\ChiselTop.wild.cpu.regs[5][29] ),
    .B_N(net2703),
    .Y(_03328_));
 sg13g2_nor2_1 _08572_ (.A(net2703),
    .B(\ChiselTop.wild.cpu.regs[4][29] ),
    .Y(_03329_));
 sg13g2_nor3_1 _08573_ (.A(net2676),
    .B(_03328_),
    .C(_03329_),
    .Y(_03330_));
 sg13g2_nor2b_1 _08574_ (.A(\ChiselTop.wild.cpu.regs[7][29] ),
    .B_N(net2704),
    .Y(_03331_));
 sg13g2_o21ai_1 _08575_ (.B1(net2676),
    .Y(_03332_),
    .A1(net2704),
    .A2(\ChiselTop.wild.cpu.regs[6][29] ));
 sg13g2_o21ai_1 _08576_ (.B1(net2660),
    .Y(_03333_),
    .A1(_03331_),
    .A2(_03332_));
 sg13g2_o21ai_1 _08577_ (.B1(net2469),
    .Y(_03334_),
    .A1(_03330_),
    .A2(_03333_));
 sg13g2_o21ai_1 _08578_ (.B1(net2445),
    .Y(_03335_),
    .A1(_03299_),
    .A2(_03324_));
 sg13g2_o21ai_1 _08579_ (.B1(_00976_),
    .Y(_03336_),
    .A1(_03327_),
    .A2(_03334_));
 sg13g2_and3_1 _08580_ (.X(_03337_),
    .A(_02640_),
    .B(_03335_),
    .C(_03336_));
 sg13g2_a21oi_1 _08581_ (.A1(_03335_),
    .A2(_03336_),
    .Y(_03338_),
    .B1(_02640_));
 sg13g2_or2_1 _08582_ (.X(_03339_),
    .B(_03338_),
    .A(_03337_));
 sg13g2_xnor2_1 _08583_ (.Y(_03340_),
    .A(_02078_),
    .B(_02690_));
 sg13g2_a21o_1 _08584_ (.A2(_02713_),
    .A1(_02088_),
    .B1(_02077_),
    .X(_03341_));
 sg13g2_nand3_1 _08585_ (.B(_02714_),
    .C(_03341_),
    .A(net2493),
    .Y(_03342_));
 sg13g2_nand2_1 _08586_ (.Y(_03343_),
    .A(net2398),
    .B(_02588_));
 sg13g2_a221oi_1 _08587_ (.B2(net2310),
    .C1(net2485),
    .B1(_03343_),
    .A1(_02587_),
    .Y(_03344_),
    .A2(net2308));
 sg13g2_nor2_1 _08588_ (.A(net2346),
    .B(_02727_),
    .Y(_03345_));
 sg13g2_o21ai_1 _08589_ (.B1(net2369),
    .Y(_03346_),
    .A1(net2351),
    .A2(_02732_));
 sg13g2_or2_1 _08590_ (.X(_03347_),
    .B(_03023_),
    .A(net2369));
 sg13g2_o21ai_1 _08591_ (.B1(_03347_),
    .Y(_03348_),
    .A1(_03345_),
    .A2(_03346_));
 sg13g2_a21oi_1 _08592_ (.A1(net2388),
    .A2(_03348_),
    .Y(_03349_),
    .B1(net2314));
 sg13g2_o21ai_1 _08593_ (.B1(_03349_),
    .Y(_03350_),
    .A1(net2389),
    .A2(_03139_));
 sg13g2_a21oi_2 _08594_ (.B1(_03344_),
    .Y(_03351_),
    .A2(_02599_),
    .A1(_01485_));
 sg13g2_a21oi_2 _08595_ (.B1(net2475),
    .Y(_03352_),
    .A2(_03351_),
    .A1(_03350_));
 sg13g2_a21oi_1 _08596_ (.A1(net2479),
    .A2(_02077_),
    .Y(_03353_),
    .B1(_03352_));
 sg13g2_a21oi_1 _08597_ (.A1(net2487),
    .A2(_03353_),
    .Y(_03354_),
    .B1(net2497));
 sg13g2_a22oi_1 _08598_ (.Y(_03355_),
    .B1(_03342_),
    .B2(_03354_),
    .A2(_03340_),
    .A1(net2497));
 sg13g2_o21ai_1 _08599_ (.B1(_02653_),
    .Y(_03356_),
    .A1(net2638),
    .A2(_03355_));
 sg13g2_xnor2_1 _08600_ (.Y(_03357_),
    .A(_02790_),
    .B(_02791_));
 sg13g2_a21o_1 _08601_ (.A2(_03357_),
    .A1(net2630),
    .B1(net2173),
    .X(_03358_));
 sg13g2_a21oi_1 _08602_ (.A1(_00925_),
    .A2(_03356_),
    .Y(_03359_),
    .B1(_03358_));
 sg13g2_a21oi_1 _08603_ (.A1(_01222_),
    .A2(_01823_),
    .Y(_03360_),
    .B1(_02799_));
 sg13g2_o21ai_1 _08604_ (.B1(net2188),
    .Y(_03361_),
    .A1(_01238_),
    .A2(_03360_));
 sg13g2_inv_1 _08605_ (.Y(_03362_),
    .A(_03361_));
 sg13g2_nand2b_1 _08606_ (.Y(_03363_),
    .B(_03361_),
    .A_N(_03359_));
 sg13g2_and2_1 _08607_ (.A(_00135_),
    .B(_02649_),
    .X(_03364_));
 sg13g2_o21ai_1 _08608_ (.B1(net2618),
    .Y(_03365_),
    .A1(_03297_),
    .A2(_03364_));
 sg13g2_inv_1 _08609_ (.Y(_03366_),
    .A(_03365_));
 sg13g2_nor3_2 _08610_ (.A(net2618),
    .B(_03359_),
    .C(_03362_),
    .Y(_03367_));
 sg13g2_or2_1 _08611_ (.X(_03368_),
    .B(_03367_),
    .A(_03366_));
 sg13g2_mux4_1 _08612_ (.S0(net2678),
    .A0(\ChiselTop.wild.cpu.regs[0][28] ),
    .A1(\ChiselTop.wild.cpu.regs[1][28] ),
    .A2(\ChiselTop.wild.cpu.regs[2][28] ),
    .A3(\ChiselTop.wild.cpu.regs[3][28] ),
    .S1(net2662),
    .X(_03369_));
 sg13g2_nor2_1 _08613_ (.A(net2652),
    .B(_03369_),
    .Y(_03370_));
 sg13g2_nor2b_1 _08614_ (.A(\ChiselTop.wild.cpu.regs[5][28] ),
    .B_N(net2678),
    .Y(_03371_));
 sg13g2_nor2_1 _08615_ (.A(net2678),
    .B(\ChiselTop.wild.cpu.regs[4][28] ),
    .Y(_03372_));
 sg13g2_nor3_1 _08616_ (.A(net2665),
    .B(_03371_),
    .C(_03372_),
    .Y(_03373_));
 sg13g2_nor2b_1 _08617_ (.A(\ChiselTop.wild.cpu.regs[7][28] ),
    .B_N(net2678),
    .Y(_03374_));
 sg13g2_o21ai_1 _08618_ (.B1(net2662),
    .Y(_03375_),
    .A1(net2678),
    .A2(\ChiselTop.wild.cpu.regs[6][28] ));
 sg13g2_o21ai_1 _08619_ (.B1(net2652),
    .Y(_03376_),
    .A1(_03374_),
    .A2(_03375_));
 sg13g2_o21ai_1 _08620_ (.B1(net2466),
    .Y(_03377_),
    .A1(_03373_),
    .A2(_03376_));
 sg13g2_nor2_2 _08621_ (.A(_03370_),
    .B(_03377_),
    .Y(_03378_));
 sg13g2_o21ai_1 _08622_ (.B1(_00975_),
    .Y(_03379_),
    .A1(_03366_),
    .A2(_03367_));
 sg13g2_nor2_1 _08623_ (.A(net2443),
    .B(_03378_),
    .Y(_03380_));
 sg13g2_inv_1 _08624_ (.Y(_03381_),
    .A(_03380_));
 sg13g2_and3_1 _08625_ (.X(_03382_),
    .A(_02640_),
    .B(_03379_),
    .C(_03381_));
 sg13g2_a21oi_1 _08626_ (.A1(_03379_),
    .A2(_03381_),
    .Y(_03383_),
    .B1(_02640_));
 sg13g2_nor2_1 _08627_ (.A(_03382_),
    .B(_03383_),
    .Y(_03384_));
 sg13g2_nor4_1 _08628_ (.A(_03337_),
    .B(_03338_),
    .C(_03382_),
    .D(_03383_),
    .Y(_03385_));
 sg13g2_o21ai_1 _08629_ (.B1(_03385_),
    .Y(_03386_),
    .A1(_02917_),
    .A2(_03295_));
 sg13g2_nor2_1 _08630_ (.A(_03337_),
    .B(_03382_),
    .Y(_03387_));
 sg13g2_xnor2_1 _08631_ (.Y(_03388_),
    .A(_02640_),
    .B(_02815_));
 sg13g2_a21oi_1 _08632_ (.A1(_03386_),
    .A2(_03387_),
    .Y(_03389_),
    .B1(_03388_));
 sg13g2_a21oi_1 _08633_ (.A1(_02640_),
    .A2(_02815_),
    .Y(_03390_),
    .B1(_03389_));
 sg13g2_o21ai_1 _08634_ (.B1(_02693_),
    .Y(_03391_),
    .A1(net2414),
    .A2(_02093_));
 sg13g2_or2_1 _08635_ (.X(_03392_),
    .B(_03391_),
    .A(_02099_));
 sg13g2_a21oi_1 _08636_ (.A1(_02099_),
    .A2(_03391_),
    .Y(_03393_),
    .B1(net2495));
 sg13g2_mux4_1 _08637_ (.S0(net2330),
    .A0(net2419),
    .A1(net2416),
    .A2(net2414),
    .A3(_01054_),
    .S1(net2342),
    .X(_03394_));
 sg13g2_mux4_1 _08638_ (.S0(net2367),
    .A0(_02824_),
    .A1(_02828_),
    .A2(_02833_),
    .A3(_03394_),
    .S1(net2387),
    .X(_03395_));
 sg13g2_nand3_1 _08639_ (.B(_01591_),
    .C(net2307),
    .A(net2385),
    .Y(_03396_));
 sg13g2_nand3_1 _08640_ (.B(_01451_),
    .C(_03396_),
    .A(net2481),
    .Y(_03397_));
 sg13g2_a22oi_1 _08641_ (.Y(_03398_),
    .B1(_03395_),
    .B2(net2316),
    .A2(_02507_),
    .A1(net2313));
 sg13g2_a221oi_1 _08642_ (.B2(_03398_),
    .C1(net2490),
    .B1(_03397_),
    .A1(net2474),
    .Y(_03399_),
    .A2(_02099_));
 sg13g2_nor3_1 _08643_ (.A(_02094_),
    .B(_02099_),
    .C(_02717_),
    .Y(_03400_));
 sg13g2_o21ai_1 _08644_ (.B1(_02099_),
    .Y(_03401_),
    .A1(_02094_),
    .A2(_02717_));
 sg13g2_nor2_1 _08645_ (.A(net2487),
    .B(_03400_),
    .Y(_03402_));
 sg13g2_a21oi_1 _08646_ (.A1(_03401_),
    .A2(_03402_),
    .Y(_03403_),
    .B1(_03399_));
 sg13g2_a21oi_1 _08647_ (.A1(net2639),
    .A2(_00934_),
    .Y(_03404_),
    .B1(net2628));
 sg13g2_a21oi_2 _08648_ (.B1(_03403_),
    .Y(_03405_),
    .A2(_03393_),
    .A1(_03392_));
 sg13g2_o21ai_1 _08649_ (.B1(_03404_),
    .Y(_03406_),
    .A1(net2639),
    .A2(_03405_));
 sg13g2_a21oi_1 _08650_ (.A1(\ChiselTop.wild.cpu.decExReg_decOut_imm[28] ),
    .A2(\ChiselTop.wild.cpu.decExReg_pc[30] ),
    .Y(_03407_),
    .B1(_02796_));
 sg13g2_xnor2_1 _08651_ (.Y(_03408_),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_imm[31] ),
    .B(\ChiselTop.wild.cpu.decExReg_pc[31] ));
 sg13g2_xnor2_1 _08652_ (.Y(_03409_),
    .A(_03407_),
    .B(_03408_));
 sg13g2_a21oi_1 _08653_ (.A1(net2630),
    .A2(_03409_),
    .Y(_03410_),
    .B1(net2172));
 sg13g2_a21o_1 _08654_ (.A2(_02857_),
    .A1(_01230_),
    .B1(_02858_),
    .X(_03411_));
 sg13g2_o21ai_1 _08655_ (.B1(_01641_),
    .Y(_03412_),
    .A1(_02301_),
    .A2(_03411_));
 sg13g2_a21oi_2 _08656_ (.B1(_03412_),
    .Y(_03413_),
    .A2(_03410_),
    .A1(_03406_));
 sg13g2_nor2_1 _08657_ (.A(net2619),
    .B(_03413_),
    .Y(_03414_));
 sg13g2_xnor2_1 _08658_ (.Y(_03415_),
    .A(\ChiselTop.wild.cpu.decExReg_pc[31] ),
    .B(_02651_));
 sg13g2_a21oi_1 _08659_ (.A1(net2619),
    .A2(_03415_),
    .Y(_03416_),
    .B1(_03414_));
 sg13g2_mux4_1 _08660_ (.S0(net2702),
    .A0(\ChiselTop.wild.cpu.regs[0][31] ),
    .A1(\ChiselTop.wild.cpu.regs[1][31] ),
    .A2(\ChiselTop.wild.cpu.regs[2][31] ),
    .A3(\ChiselTop.wild.cpu.regs[3][31] ),
    .S1(net2675),
    .X(_03417_));
 sg13g2_nor2_1 _08661_ (.A(net2660),
    .B(_03417_),
    .Y(_03418_));
 sg13g2_nor2b_1 _08662_ (.A(\ChiselTop.wild.cpu.regs[5][31] ),
    .B_N(net2698),
    .Y(_03419_));
 sg13g2_nor2_1 _08663_ (.A(net2698),
    .B(\ChiselTop.wild.cpu.regs[4][31] ),
    .Y(_03420_));
 sg13g2_nor3_1 _08664_ (.A(net2673),
    .B(_03419_),
    .C(_03420_),
    .Y(_03421_));
 sg13g2_nor2b_1 _08665_ (.A(\ChiselTop.wild.cpu.regs[7][31] ),
    .B_N(net2698),
    .Y(_03422_));
 sg13g2_o21ai_1 _08666_ (.B1(net2673),
    .Y(_03423_),
    .A1(net2698),
    .A2(\ChiselTop.wild.cpu.regs[6][31] ));
 sg13g2_o21ai_1 _08667_ (.B1(net2657),
    .Y(_03424_),
    .A1(_03422_),
    .A2(_03423_));
 sg13g2_o21ai_1 _08668_ (.B1(net2468),
    .Y(_03425_),
    .A1(_03421_),
    .A2(_03424_));
 sg13g2_nor2_1 _08669_ (.A(_03418_),
    .B(_03425_),
    .Y(_03426_));
 sg13g2_nor2_1 _08670_ (.A(net2444),
    .B(_03426_),
    .Y(_03427_));
 sg13g2_a21oi_1 _08671_ (.A1(net2444),
    .A2(net2074),
    .Y(_03428_),
    .B1(_03427_));
 sg13g2_xnor2_1 _08672_ (.Y(_03429_),
    .A(_00110_),
    .B(_03428_));
 sg13g2_xnor2_1 _08673_ (.Y(\ChiselTop.wild.cpu.io_dmem_rdAddress[31] ),
    .A(_03390_),
    .B(_03429_));
 sg13g2_nand3_1 _08674_ (.B(_03387_),
    .C(_03388_),
    .A(_03386_),
    .Y(_03430_));
 sg13g2_nor2b_1 _08675_ (.A(_03389_),
    .B_N(_03430_),
    .Y(\ChiselTop.wild.cpu.io_dmem_rdAddress[30] ));
 sg13g2_a21oi_1 _08676_ (.A1(_03296_),
    .A2(_03384_),
    .Y(_03431_),
    .B1(_03382_));
 sg13g2_xor2_1 _08677_ (.B(_03431_),
    .A(_03339_),
    .X(\ChiselTop.wild.cpu.io_dmem_rdAddress[29] ));
 sg13g2_xor2_1 _08678_ (.B(_03384_),
    .A(_03296_),
    .X(\ChiselTop.wild.cpu.io_dmem_rdAddress[28] ));
 sg13g2_or3_1 _08679_ (.A(_01941_),
    .B(_01999_),
    .C(_02184_),
    .X(_03432_));
 sg13g2_and2_1 _08680_ (.A(_02185_),
    .B(_03432_),
    .X(\ChiselTop.wild.cpu.io_dmem_rdAddress[2] ));
 sg13g2_xnor2_1 _08681_ (.Y(_03433_),
    .A(_03173_),
    .B(_03207_));
 sg13g2_a21oi_1 _08682_ (.A1(_00965_),
    .A2(_01567_),
    .Y(_03434_),
    .B1(_02636_));
 sg13g2_xnor2_1 _08683_ (.Y(_03435_),
    .A(_03433_),
    .B(_03434_));
 sg13g2_inv_1 _08684_ (.Y(\ChiselTop.wild.cpu.io_dmem_rdAddress[17] ),
    .A(_03435_));
 sg13g2_nand2_1 _08685_ (.Y(_03436_),
    .A(_03210_),
    .B(_03285_));
 sg13g2_xnor2_1 _08686_ (.Y(_03437_),
    .A(_03210_),
    .B(_03285_));
 sg13g2_inv_1 _08687_ (.Y(\ChiselTop.wild.cpu.io_dmem_rdAddress[18] ),
    .A(_03437_));
 sg13g2_nand2_1 _08688_ (.Y(_03438_),
    .A(_03284_),
    .B(_03436_));
 sg13g2_xor2_1 _08689_ (.B(_03438_),
    .A(_03249_),
    .X(_03439_));
 sg13g2_inv_1 _08690_ (.Y(\ChiselTop.wild.cpu.io_dmem_rdAddress[19] ),
    .A(_03439_));
 sg13g2_xnor2_1 _08691_ (.Y(_03440_),
    .A(_02189_),
    .B(_02248_));
 sg13g2_xnor2_1 _08692_ (.Y(\ChiselTop.wild.cpu.io_dmem_rdAddress[3] ),
    .A(_02186_),
    .B(_03440_));
 sg13g2_nor2_1 _08693_ (.A(\ChiselTop.dec.counter[1] ),
    .B(_00949_),
    .Y(_03441_));
 sg13g2_nor2_1 _08694_ (.A(_00949_),
    .B(net2650),
    .Y(_03442_));
 sg13g2_nand2_1 _08695_ (.Y(_03443_),
    .A(_00950_),
    .B(_03441_));
 sg13g2_nand3_1 _08696_ (.B(\ChiselTop.dec.counter[0] ),
    .C(net2650),
    .A(\ChiselTop.dec.counter[1] ),
    .Y(_03444_));
 sg13g2_nand2_1 _08697_ (.Y(_03445_),
    .A(_03443_),
    .B(_03444_));
 sg13g2_nand2_1 _08698_ (.Y(_03446_),
    .A(_00951_),
    .B(_03444_));
 sg13g2_nor3_1 _08699_ (.A(_00950_),
    .B(_00951_),
    .C(_03441_),
    .Y(_03447_));
 sg13g2_a21oi_1 _08700_ (.A1(\ChiselTop.dec.counter[2] ),
    .A2(_03442_),
    .Y(_03448_),
    .B1(_03447_));
 sg13g2_o21ai_1 _08701_ (.B1(_03448_),
    .Y(uo_out[0]),
    .A1(\ChiselTop.dec.counter[2] ),
    .A2(_03445_));
 sg13g2_nor2_1 _08702_ (.A(\ChiselTop.dec.counter[1] ),
    .B(net2650),
    .Y(_03449_));
 sg13g2_nor2_1 _08703_ (.A(\ChiselTop.dec.counter[0] ),
    .B(_03449_),
    .Y(_03450_));
 sg13g2_nand2b_2 _08704_ (.Y(_03451_),
    .B(\ChiselTop.dec.counter[2] ),
    .A_N(\ChiselTop.dec.counter[1] ));
 sg13g2_o21ai_1 _08705_ (.B1(_03446_),
    .Y(uo_out[1]),
    .A1(_03445_),
    .A2(_03450_));
 sg13g2_nand2_1 _08706_ (.Y(_03452_),
    .A(\ChiselTop.dec.counter[1] ),
    .B(_00951_));
 sg13g2_nor3_1 _08707_ (.A(\ChiselTop.dec.counter[0] ),
    .B(net2650),
    .C(_03452_),
    .Y(_03453_));
 sg13g2_nor2_1 _08708_ (.A(_03447_),
    .B(_03453_),
    .Y(uo_out[2]));
 sg13g2_nand2_1 _08709_ (.Y(_03454_),
    .A(_00949_),
    .B(_03451_));
 sg13g2_a22oi_1 _08710_ (.Y(_03455_),
    .B1(_03451_),
    .B2(_03452_),
    .A2(_00950_),
    .A1(_00949_));
 sg13g2_xnor2_1 _08711_ (.Y(uo_out[3]),
    .A(_03454_),
    .B(_03455_));
 sg13g2_o21ai_1 _08712_ (.B1(net2650),
    .Y(_03456_),
    .A1(\ChiselTop.dec.counter[1] ),
    .A2(\ChiselTop.dec.counter[2] ));
 sg13g2_nand2_1 _08713_ (.Y(uo_out[4]),
    .A(_03454_),
    .B(_03456_));
 sg13g2_a22oi_1 _08714_ (.Y(_03457_),
    .B1(_03452_),
    .B2(_00949_),
    .A2(_03451_),
    .A1(net2650));
 sg13g2_o21ai_1 _08715_ (.B1(_03457_),
    .Y(uo_out[5]),
    .A1(net2650),
    .A2(_03451_));
 sg13g2_a21oi_1 _08716_ (.A1(\ChiselTop.dec.counter[2] ),
    .A2(_03442_),
    .Y(_03458_),
    .B1(_03449_));
 sg13g2_o21ai_1 _08717_ (.B1(_03458_),
    .Y(_03459_),
    .A1(\ChiselTop.dec.counter[0] ),
    .A2(_03451_));
 sg13g2_o21ai_1 _08718_ (.B1(_03459_),
    .Y(uo_out[6]),
    .A1(net2650),
    .A2(_03451_));
 sg13g2_nor2b_2 _08719_ (.A(net2553),
    .B_N(net2552),
    .Y(_03460_));
 sg13g2_nor2b_2 _08720_ (.A(net1531),
    .B_N(\ChiselTop.wild.cpu.pcReg[2] ),
    .Y(_03461_));
 sg13g2_nand2_1 _08721_ (.Y(_03462_),
    .A(_03460_),
    .B(_03461_));
 sg13g2_nor2b_2 _08722_ (.A(net1535),
    .B_N(net1531),
    .Y(_03463_));
 sg13g2_nor2_2 _08723_ (.A(net2552),
    .B(net2553),
    .Y(_03464_));
 sg13g2_a22oi_1 _08724_ (.Y(_03465_),
    .B1(_03463_),
    .B2(_03464_),
    .A2(_03461_),
    .A1(_03460_));
 sg13g2_inv_1 _08725_ (.Y(\ChiselTop.wild.cpu.io_imem_data[13] ),
    .A(_03465_));
 sg13g2_nor2_1 _08726_ (.A(net1038),
    .B(net1260),
    .Y(_03466_));
 sg13g2_or2_1 _08727_ (.X(_03467_),
    .B(net1535),
    .A(net1038));
 sg13g2_nand2_1 _08728_ (.Y(_03468_),
    .A(net2552),
    .B(_03466_));
 sg13g2_nand2_1 _08729_ (.Y(_03469_),
    .A(_03460_),
    .B(_03466_));
 sg13g2_and2_2 _08730_ (.A(net1546),
    .B(\ChiselTop.wild.cpu.pcReg[2] ),
    .X(_03470_));
 sg13g2_nand2b_1 _08731_ (.Y(_03471_),
    .B(net2553),
    .A_N(net2552));
 sg13g2_nand2_2 _08732_ (.Y(_03472_),
    .A(net856),
    .B(_03470_));
 sg13g2_o21ai_1 _08733_ (.B1(_03469_),
    .Y(_03473_),
    .A1(net2552),
    .A2(_03472_));
 sg13g2_nand3_1 _08734_ (.B(net2553),
    .C(_03466_),
    .A(net2552),
    .Y(_03474_));
 sg13g2_nand2_1 _08735_ (.Y(_03475_),
    .A(_03460_),
    .B(_03463_));
 sg13g2_nand3b_1 _08736_ (.B(_03474_),
    .C(_03475_),
    .Y(\ChiselTop.wild.cpu.io_imem_data[15] ),
    .A_N(_03473_));
 sg13g2_nor2_2 _08737_ (.A(net2553),
    .B(net1532),
    .Y(_03476_));
 sg13g2_nand2_1 _08738_ (.Y(_03477_),
    .A(_03460_),
    .B(_03470_));
 sg13g2_or2_1 _08739_ (.X(_03478_),
    .B(_03476_),
    .A(net2552));
 sg13g2_a21oi_1 _08740_ (.A1(net2553),
    .A2(_03467_),
    .Y(_03479_),
    .B1(_03478_));
 sg13g2_a21oi_1 _08741_ (.A1(net2553),
    .A2(_03467_),
    .Y(_03480_),
    .B1(_03476_));
 sg13g2_nor2_1 _08742_ (.A(_03461_),
    .B(_03463_),
    .Y(_03481_));
 sg13g2_o21ai_1 _08743_ (.B1(_03464_),
    .Y(_03482_),
    .A1(_03461_),
    .A2(_03463_));
 sg13g2_nand2_1 _08744_ (.Y(_03483_),
    .A(_03462_),
    .B(_03482_));
 sg13g2_nor3_1 _08745_ (.A(_03473_),
    .B(_03480_),
    .C(_03483_),
    .Y(\ChiselTop.wild.cpu.io_imem_data[16] ));
 sg13g2_nor2_1 _08746_ (.A(_03463_),
    .B(_03471_),
    .Y(_03484_));
 sg13g2_a21oi_2 _08747_ (.B1(_03484_),
    .Y(_03485_),
    .A2(_03470_),
    .A1(_03464_));
 sg13g2_inv_2 _08748_ (.Y(\ChiselTop.wild.cpu.io_imem_data[22] ),
    .A(_03485_));
 sg13g2_nand2b_1 _08749_ (.Y(_03486_),
    .B(_03482_),
    .A_N(_03460_));
 sg13g2_nand2_1 _08750_ (.Y(_03487_),
    .A(_03467_),
    .B(_03486_));
 sg13g2_nand2_1 _08751_ (.Y(\ChiselTop.wild.cpu.io_imem_data[20] ),
    .A(_03485_),
    .B(_03487_));
 sg13g2_nand2_1 _08752_ (.Y(\ChiselTop.wild.cpu.io_imem_data[21] ),
    .A(_03465_),
    .B(_03485_));
 sg13g2_and2_1 _08753_ (.A(\ChiselTop.ledReg ),
    .B(net1),
    .X(\ChiselTop.led ));
 sg13g2_nor3_2 _08754_ (.A(net1464),
    .B(net937),
    .C(net1495),
    .Y(_03488_));
 sg13g2_nor2b_1 _08755_ (.A(net1342),
    .B_N(_03488_),
    .Y(_03489_));
 sg13g2_nor2b_1 _08756_ (.A(net1355),
    .B_N(_03489_),
    .Y(_03490_));
 sg13g2_nor2b_1 _08757_ (.A(net1331),
    .B_N(_03490_),
    .Y(_03491_));
 sg13g2_nor2b_1 _08758_ (.A(net1367),
    .B_N(_03491_),
    .Y(_03492_));
 sg13g2_nand2b_2 _08759_ (.Y(_03493_),
    .B(_03492_),
    .A_N(net1078));
 sg13g2_nor3_2 _08760_ (.A(net1504),
    .B(net1479),
    .C(_03493_),
    .Y(_03494_));
 sg13g2_nand2b_2 _08761_ (.Y(_03495_),
    .B(_03494_),
    .A_N(net1106));
 sg13g2_nor3_2 _08762_ (.A(net1484),
    .B(net1510),
    .C(_03495_),
    .Y(_03496_));
 sg13g2_nand2b_2 _08763_ (.Y(_03497_),
    .B(_03496_),
    .A_N(net1138));
 sg13g2_nor3_2 _08764_ (.A(net1486),
    .B(net1468),
    .C(_03497_),
    .Y(_03498_));
 sg13g2_nand2b_2 _08765_ (.Y(_03499_),
    .B(_03498_),
    .A_N(net1042));
 sg13g2_nor3_2 _08766_ (.A(net1481),
    .B(net1506),
    .C(_03499_),
    .Y(_03500_));
 sg13g2_nand2_2 _08767_ (.Y(_03501_),
    .A(_00944_),
    .B(_03500_));
 sg13g2_nand2_1 _08768_ (.Y(_03502_),
    .A(net2736),
    .B(_03501_));
 sg13g2_o21ai_1 _08769_ (.B1(net1495),
    .Y(_03503_),
    .A1(net1464),
    .A2(net937));
 sg13g2_nor2b_1 _08770_ (.A(_03488_),
    .B_N(_03503_),
    .Y(_03504_));
 sg13g2_nor2_1 _08771_ (.A(net2154),
    .B(_03504_),
    .Y(_00143_));
 sg13g2_xnor2_1 _08772_ (.Y(_03505_),
    .A(net1342),
    .B(_03488_));
 sg13g2_nor2_1 _08773_ (.A(net2154),
    .B(net1343),
    .Y(_00144_));
 sg13g2_xnor2_1 _08774_ (.Y(_03506_),
    .A(net1355),
    .B(_03489_));
 sg13g2_nor2_1 _08775_ (.A(net2154),
    .B(net1356),
    .Y(_00145_));
 sg13g2_nand2b_1 _08776_ (.Y(_03507_),
    .B(net1078),
    .A_N(_03492_));
 sg13g2_a21oi_1 _08777_ (.A1(_03493_),
    .A2(net1079),
    .Y(_00146_),
    .B1(net2153));
 sg13g2_nand2b_1 _08778_ (.Y(_03508_),
    .B(net1106),
    .A_N(_03494_));
 sg13g2_a21oi_1 _08779_ (.A1(_03495_),
    .A2(net1107),
    .Y(_00147_),
    .B1(net2153));
 sg13g2_xor2_1 _08780_ (.B(_03495_),
    .A(net1484),
    .X(_03509_));
 sg13g2_nor2_1 _08781_ (.A(net2153),
    .B(net1485),
    .Y(_00148_));
 sg13g2_o21ai_1 _08782_ (.B1(net1510),
    .Y(_03510_),
    .A1(\ChiselTop.wild.tx.tx.cntReg[11] ),
    .A2(_03495_));
 sg13g2_nor2b_1 _08783_ (.A(_03496_),
    .B_N(_03510_),
    .Y(_03511_));
 sg13g2_nor2_1 _08784_ (.A(net2153),
    .B(net1511),
    .Y(_00149_));
 sg13g2_nand2b_1 _08785_ (.Y(_03512_),
    .B(net1138),
    .A_N(_03496_));
 sg13g2_a21oi_1 _08786_ (.A1(_03497_),
    .A2(net1139),
    .Y(_00150_),
    .B1(net2153));
 sg13g2_xor2_1 _08787_ (.B(_03497_),
    .A(net1468),
    .X(_03513_));
 sg13g2_nor2_1 _08788_ (.A(net2153),
    .B(net1469),
    .Y(_00151_));
 sg13g2_o21ai_1 _08789_ (.B1(net1486),
    .Y(_03514_),
    .A1(net1468),
    .A2(_03497_));
 sg13g2_nor2b_1 _08790_ (.A(net1487),
    .B_N(_03514_),
    .Y(_03515_));
 sg13g2_nor2_1 _08791_ (.A(net2153),
    .B(_03515_),
    .Y(_00152_));
 sg13g2_nand2b_1 _08792_ (.Y(_03516_),
    .B(net1042),
    .A_N(_03498_));
 sg13g2_a21oi_1 _08793_ (.A1(_03499_),
    .A2(net1043),
    .Y(_00153_),
    .B1(net2153));
 sg13g2_xor2_1 _08794_ (.B(_03499_),
    .A(net1481),
    .X(_03517_));
 sg13g2_nor2_1 _08795_ (.A(net2154),
    .B(net1482),
    .Y(_00154_));
 sg13g2_o21ai_1 _08796_ (.B1(net1506),
    .Y(_03518_),
    .A1(net1481),
    .A2(_03499_));
 sg13g2_nor2b_1 _08797_ (.A(_03500_),
    .B_N(_03518_),
    .Y(_03519_));
 sg13g2_nor2_1 _08798_ (.A(net2154),
    .B(_03519_),
    .Y(_00155_));
 sg13g2_nor3_1 _08799_ (.A(net2721),
    .B(_00944_),
    .C(_03500_),
    .Y(_00156_));
 sg13g2_nand2b_1 _08800_ (.Y(_03520_),
    .B(net2649),
    .A_N(net2648));
 sg13g2_nor2_1 _08801_ (.A(\ChiselTop.wild.cpu.decExReg_rd[2] ),
    .B(_00970_),
    .Y(_03521_));
 sg13g2_nand2_1 _08802_ (.Y(_03522_),
    .A(net2648),
    .B(net2649));
 sg13g2_nor2_2 _08803_ (.A(_00142_),
    .B(_00970_),
    .Y(_03523_));
 sg13g2_nand2b_1 _08804_ (.Y(_03524_),
    .B(net2648),
    .A_N(net2649));
 sg13g2_nor2_1 _08805_ (.A(\ChiselTop.wild.cpu._GEN_176[6] ),
    .B(\ChiselTop.wild.cpu._GEN_176[5] ),
    .Y(_03525_));
 sg13g2_nand3_1 _08806_ (.B(net1453),
    .C(_03525_),
    .A(\ChiselTop.wild.cpu._GEN_176[20] ),
    .Y(_03526_));
 sg13g2_and2_1 _08807_ (.A(net1523),
    .B(net2730),
    .X(_00563_));
 sg13g2_nor2b_1 _08808_ (.A(net1496),
    .B_N(net1518),
    .Y(_03527_));
 sg13g2_nand3_1 _08809_ (.B(_00563_),
    .C(_03527_),
    .A(net1458),
    .Y(_03528_));
 sg13g2_nor2_1 _08810_ (.A(net1454),
    .B(_03528_),
    .Y(_00158_));
 sg13g2_and2_2 _08811_ (.A(net1496),
    .B(net2730),
    .X(_00562_));
 sg13g2_nor4_1 _08812_ (.A(net1458),
    .B(\ChiselTop.wild.cpu._GEN_176[1] ),
    .C(_00941_),
    .D(_03526_),
    .Y(_03529_));
 sg13g2_a21o_1 _08813_ (.A2(_03529_),
    .A1(_00562_),
    .B1(_00158_),
    .X(_00157_));
 sg13g2_nand2_2 _08814_ (.Y(_03530_),
    .A(_00967_),
    .B(_03521_));
 sg13g2_nor2_2 _08815_ (.A(_03520_),
    .B(_03530_),
    .Y(_03531_));
 sg13g2_nor2_1 _08816_ (.A(net1215),
    .B(net2303),
    .Y(_03532_));
 sg13g2_a21oi_1 _08817_ (.A1(net2136),
    .A2(net2303),
    .Y(_00159_),
    .B1(_03532_));
 sg13g2_nor2_1 _08818_ (.A(net1212),
    .B(net2304),
    .Y(_03533_));
 sg13g2_a21oi_1 _08819_ (.A1(net2148),
    .A2(net2304),
    .Y(_00160_),
    .B1(_03533_));
 sg13g2_nor2_1 _08820_ (.A(net1385),
    .B(net2303),
    .Y(_03534_));
 sg13g2_a21oi_1 _08821_ (.A1(net2138),
    .A2(net2303),
    .Y(_00161_),
    .B1(_03534_));
 sg13g2_nor2_1 _08822_ (.A(net1322),
    .B(net2303),
    .Y(_03535_));
 sg13g2_a21oi_1 _08823_ (.A1(net2134),
    .A2(net2303),
    .Y(_00162_),
    .B1(_03535_));
 sg13g2_nor2_1 _08824_ (.A(net1341),
    .B(net2303),
    .Y(_03536_));
 sg13g2_a21oi_1 _08825_ (.A1(net2151),
    .A2(net2303),
    .Y(_00163_),
    .B1(_03536_));
 sg13g2_nor2_1 _08826_ (.A(net1347),
    .B(net2302),
    .Y(_03537_));
 sg13g2_a21oi_1 _08827_ (.A1(net2141),
    .A2(net2302),
    .Y(_00164_),
    .B1(_03537_));
 sg13g2_nor2_1 _08828_ (.A(net1207),
    .B(net2300),
    .Y(_03538_));
 sg13g2_a21oi_1 _08829_ (.A1(net2143),
    .A2(net2300),
    .Y(_00165_),
    .B1(_03538_));
 sg13g2_nor2_1 _08830_ (.A(net1253),
    .B(net2300),
    .Y(_03539_));
 sg13g2_a21oi_1 _08831_ (.A1(net2145),
    .A2(net2300),
    .Y(_00166_),
    .B1(_03539_));
 sg13g2_nor2_1 _08832_ (.A(net1357),
    .B(net2301),
    .Y(_03540_));
 sg13g2_a21oi_1 _08833_ (.A1(net2131),
    .A2(net2301),
    .Y(_00167_),
    .B1(_03540_));
 sg13g2_nor2_1 _08834_ (.A(net1319),
    .B(net2298),
    .Y(_03541_));
 sg13g2_a21oi_1 _08835_ (.A1(net2127),
    .A2(net2298),
    .Y(_00168_),
    .B1(_03541_));
 sg13g2_nor2_1 _08836_ (.A(net1318),
    .B(net2297),
    .Y(_03542_));
 sg13g2_a21oi_1 _08837_ (.A1(net2133),
    .A2(net2297),
    .Y(_00169_),
    .B1(_03542_));
 sg13g2_mux2_1 _08838_ (.A0(net1334),
    .A1(net2123),
    .S(net2300),
    .X(_00170_));
 sg13g2_nor2_1 _08839_ (.A(net1247),
    .B(net2300),
    .Y(_03543_));
 sg13g2_a21oi_1 _08840_ (.A1(net2125),
    .A2(net2300),
    .Y(_00171_),
    .B1(_03543_));
 sg13g2_nor2_1 _08841_ (.A(net1274),
    .B(net2301),
    .Y(_03544_));
 sg13g2_a21oi_1 _08842_ (.A1(net2122),
    .A2(net2301),
    .Y(_00172_),
    .B1(_03544_));
 sg13g2_nor2_1 _08843_ (.A(net1263),
    .B(net2299),
    .Y(_03545_));
 sg13g2_a21oi_1 _08844_ (.A1(net2120),
    .A2(net2299),
    .Y(_00173_),
    .B1(_03545_));
 sg13g2_nor2_1 _08845_ (.A(net1290),
    .B(net2304),
    .Y(_03546_));
 sg13g2_a21oi_1 _08846_ (.A1(net2117),
    .A2(net2304),
    .Y(_00174_),
    .B1(_03546_));
 sg13g2_nor2_1 _08847_ (.A(net1379),
    .B(net2297),
    .Y(_03547_));
 sg13g2_a21oi_1 _08848_ (.A1(net2111),
    .A2(net2297),
    .Y(_00175_),
    .B1(_03547_));
 sg13g2_nor2_1 _08849_ (.A(net1363),
    .B(net2297),
    .Y(_03548_));
 sg13g2_a21oi_1 _08850_ (.A1(net2114),
    .A2(net2297),
    .Y(_00176_),
    .B1(_03548_));
 sg13g2_nor2_1 _08851_ (.A(net1235),
    .B(net2298),
    .Y(_03549_));
 sg13g2_a21oi_1 _08852_ (.A1(net2105),
    .A2(net2298),
    .Y(_00177_),
    .B1(_03549_));
 sg13g2_nor2_1 _08853_ (.A(net1243),
    .B(net2302),
    .Y(_03550_));
 sg13g2_a21oi_1 _08854_ (.A1(net2108),
    .A2(net2302),
    .Y(_00178_),
    .B1(_03550_));
 sg13g2_nor2_1 _08855_ (.A(net1324),
    .B(net2299),
    .Y(_03551_));
 sg13g2_a21oi_1 _08856_ (.A1(net2099),
    .A2(net2299),
    .Y(_00179_),
    .B1(_03551_));
 sg13g2_nor2_1 _08857_ (.A(net1209),
    .B(net2299),
    .Y(_03552_));
 sg13g2_a21oi_1 _08858_ (.A1(net2103),
    .A2(net2299),
    .Y(_00180_),
    .B1(_03552_));
 sg13g2_nor2_1 _08859_ (.A(net1223),
    .B(net2298),
    .Y(_03553_));
 sg13g2_a21oi_1 _08860_ (.A1(net2093),
    .A2(net2298),
    .Y(_00181_),
    .B1(_03553_));
 sg13g2_nor2_1 _08861_ (.A(net1345),
    .B(net2299),
    .Y(_03554_));
 sg13g2_a21oi_1 _08862_ (.A1(net2090),
    .A2(net2299),
    .Y(_00182_),
    .B1(_03554_));
 sg13g2_nor2_1 _08863_ (.A(net1329),
    .B(net2304),
    .Y(_03555_));
 sg13g2_a21oi_1 _08864_ (.A1(net2096),
    .A2(net2304),
    .Y(_00183_),
    .B1(_03555_));
 sg13g2_nor2_1 _08865_ (.A(net1267),
    .B(net2297),
    .Y(_03556_));
 sg13g2_a21oi_1 _08866_ (.A1(net2082),
    .A2(net2297),
    .Y(_00184_),
    .B1(_03556_));
 sg13g2_nor2_1 _08867_ (.A(net1396),
    .B(net2305),
    .Y(_03557_));
 sg13g2_a21oi_1 _08868_ (.A1(net2085),
    .A2(net2305),
    .Y(_00185_),
    .B1(_03557_));
 sg13g2_nor2_1 _08869_ (.A(net1328),
    .B(net2302),
    .Y(_03558_));
 sg13g2_a21oi_1 _08870_ (.A1(net2087),
    .A2(net2302),
    .Y(_00186_),
    .B1(_03558_));
 sg13g2_nor2_1 _08871_ (.A(net1381),
    .B(net2298),
    .Y(_03559_));
 sg13g2_a21oi_1 _08872_ (.A1(net2077),
    .A2(net2298),
    .Y(_00187_),
    .B1(_03559_));
 sg13g2_nor2_1 _08873_ (.A(net1330),
    .B(net2305),
    .Y(_03560_));
 sg13g2_a21oi_1 _08874_ (.A1(net2079),
    .A2(net2305),
    .Y(_00188_),
    .B1(_03560_));
 sg13g2_nor2_1 _08875_ (.A(net1273),
    .B(net2302),
    .Y(_03561_));
 sg13g2_a21oi_1 _08876_ (.A1(net2076),
    .A2(net2302),
    .Y(_00189_),
    .B1(_03561_));
 sg13g2_nor2_1 _08877_ (.A(net1189),
    .B(net2304),
    .Y(_03562_));
 sg13g2_a21oi_1 _08878_ (.A1(net2074),
    .A2(net2304),
    .Y(_00190_),
    .B1(_03562_));
 sg13g2_nor2_2 _08879_ (.A(net2550),
    .B(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[13] ),
    .Y(_03563_));
 sg13g2_nor2_1 _08880_ (.A(net2528),
    .B(_00929_),
    .Y(_03564_));
 sg13g2_nor3_1 _08881_ (.A(net2724),
    .B(net2524),
    .C(_03564_),
    .Y(_00191_));
 sg13g2_nor2_1 _08882_ (.A(net2528),
    .B(net2723),
    .Y(_00597_));
 sg13g2_nor3_2 _08883_ (.A(net2528),
    .B(_00929_),
    .C(net2722),
    .Y(_00192_));
 sg13g2_nand2_1 _08884_ (.Y(_03565_),
    .A(net2734),
    .B(net2192));
 sg13g2_inv_1 _08885_ (.Y(_00524_),
    .A(net2182));
 sg13g2_a21oi_1 _08886_ (.A1(_03469_),
    .A2(_03478_),
    .Y(_00194_),
    .B1(net2178));
 sg13g2_nor2_1 _08887_ (.A(_03465_),
    .B(net2178),
    .Y(_00195_));
 sg13g2_nand3_1 _08888_ (.B(_03477_),
    .C(net2169),
    .A(_03474_),
    .Y(_03566_));
 sg13g2_nor2_1 _08889_ (.A(net1038),
    .B(_03471_),
    .Y(_03567_));
 sg13g2_a21oi_1 _08890_ (.A1(_03461_),
    .A2(_03464_),
    .Y(_03568_),
    .B1(_03567_));
 sg13g2_a21oi_1 _08891_ (.A1(_03475_),
    .A2(_03568_),
    .Y(_00196_),
    .B1(_03566_));
 sg13g2_a22oi_1 _08892_ (.Y(_03569_),
    .B1(_03464_),
    .B2(net1260),
    .A2(_03460_),
    .A1(net1531));
 sg13g2_nand2b_1 _08893_ (.Y(_03570_),
    .B(_03569_),
    .A_N(_03484_));
 sg13g2_nand2_1 _08894_ (.Y(_00197_),
    .A(net2169),
    .B(_03570_));
 sg13g2_nand2_2 _08895_ (.Y(_03571_),
    .A(net2191),
    .B(_02001_));
 sg13g2_inv_1 _08896_ (.Y(_03572_),
    .A(_03571_));
 sg13g2_and3_1 _08897_ (.X(_03573_),
    .A(\ChiselTop.wild.cpu.io_dmem_rdAddress[30] ),
    .B(\ChiselTop.wild.cpu.io_dmem_rdAddress[29] ),
    .C(\ChiselTop.wild.cpu.io_dmem_rdAddress[28] ));
 sg13g2_or2_1 _08898_ (.X(_03574_),
    .B(\ChiselTop.wild.cpu.decEx_memLow[1] ),
    .A(\ChiselTop.wild.cpu.decEx_memLow[0] ));
 sg13g2_a21oi_1 _08899_ (.A1(_00929_),
    .A2(_03574_),
    .Y(_03575_),
    .B1(_03571_));
 sg13g2_nand3_1 _08900_ (.B(_03573_),
    .C(_03575_),
    .A(\ChiselTop.wild.cpu.io_dmem_rdAddress[31] ),
    .Y(_03576_));
 sg13g2_nand2_1 _08901_ (.Y(_03577_),
    .A(_02638_),
    .B(\ChiselTop.wild.cpu.decEx_memLow[1] ));
 sg13g2_nand2_1 _08902_ (.Y(_03578_),
    .A(_00929_),
    .B(_03577_));
 sg13g2_nand3_1 _08903_ (.B(_03576_),
    .C(_03578_),
    .A(_03572_),
    .Y(_03579_));
 sg13g2_and4_1 _08904_ (.A(\ChiselTop.wild.cpu.decExReg_rd[2] ),
    .B(\ChiselTop.wild.cpu.decExReg_rd[3] ),
    .C(net2612),
    .D(\ChiselTop.wild.cpu._GEN_176[2] ),
    .X(_03580_));
 sg13g2_a21oi_1 _08905_ (.A1(_00931_),
    .A2(_00968_),
    .Y(_03581_),
    .B1(_03580_));
 sg13g2_xor2_1 _08906_ (.B(\ChiselTop.wild.cpu._GEN_176[1] ),
    .A(net2648),
    .X(_03582_));
 sg13g2_xor2_1 _08907_ (.B(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_1[0] ),
    .A(net2649),
    .X(_03583_));
 sg13g2_nor4_1 _08908_ (.A(_00970_),
    .B(_03581_),
    .C(_03582_),
    .D(_03583_),
    .Y(_03584_));
 sg13g2_nand2_1 _08909_ (.Y(_03585_),
    .A(_00929_),
    .B(_03572_));
 sg13g2_mux4_1 _08910_ (.S0(net2587),
    .A0(\ChiselTop.wild.cpu.regs[0][16] ),
    .A1(\ChiselTop.wild.cpu.regs[1][16] ),
    .A2(\ChiselTop.wild.cpu.regs[2][16] ),
    .A3(\ChiselTop.wild.cpu.regs[3][16] ),
    .S1(net2567),
    .X(_03586_));
 sg13g2_nor2_1 _08911_ (.A(net2559),
    .B(_03586_),
    .Y(_03587_));
 sg13g2_nor2b_1 _08912_ (.A(\ChiselTop.wild.cpu.regs[29][16] ),
    .B_N(net2587),
    .Y(_03588_));
 sg13g2_nor2_1 _08913_ (.A(net2587),
    .B(\ChiselTop.wild.cpu.regs[28][16] ),
    .Y(_03589_));
 sg13g2_nor3_1 _08914_ (.A(net2567),
    .B(_03588_),
    .C(_03589_),
    .Y(_03590_));
 sg13g2_nor2b_1 _08915_ (.A(\ChiselTop.wild.cpu.regs[31][16] ),
    .B_N(net2587),
    .Y(_03591_));
 sg13g2_o21ai_1 _08916_ (.B1(net2567),
    .Y(_03592_),
    .A1(net2587),
    .A2(\ChiselTop.wild.cpu.regs[30][16] ));
 sg13g2_o21ai_1 _08917_ (.B1(net2559),
    .Y(_03593_),
    .A1(_03591_),
    .A2(_03592_));
 sg13g2_nor2_1 _08918_ (.A(net2608),
    .B(net2580),
    .Y(_03594_));
 sg13g2_nand2_1 _08919_ (.Y(_03595_),
    .A(_00138_),
    .B(_03594_));
 sg13g2_o21ai_1 _08920_ (.B1(net2460),
    .Y(_03596_),
    .A1(_03590_),
    .A2(_03593_));
 sg13g2_nor2_1 _08921_ (.A(_03587_),
    .B(_03596_),
    .Y(_03597_));
 sg13g2_inv_2 _08922_ (.Y(_03598_),
    .A(_03597_));
 sg13g2_mux2_1 _08923_ (.A0(_03598_),
    .A1(net2113),
    .S(net2407),
    .X(_03599_));
 sg13g2_mux4_1 _08924_ (.S0(net2602),
    .A0(\ChiselTop.wild.cpu.regs[0][0] ),
    .A1(\ChiselTop.wild.cpu.regs[1][0] ),
    .A2(\ChiselTop.wild.cpu.regs[2][0] ),
    .A3(\ChiselTop.wild.cpu.regs[3][0] ),
    .S1(net2576),
    .X(_03600_));
 sg13g2_nor2_1 _08925_ (.A(net2561),
    .B(_03600_),
    .Y(_03601_));
 sg13g2_nor2b_1 _08926_ (.A(net969),
    .B_N(net2602),
    .Y(_03602_));
 sg13g2_nor2_1 _08927_ (.A(net2602),
    .B(net970),
    .Y(_03603_));
 sg13g2_nor3_1 _08928_ (.A(net2576),
    .B(_03602_),
    .C(_03603_),
    .Y(_03604_));
 sg13g2_nor2b_1 _08929_ (.A(\ChiselTop.wild.cpu.regs[31][0] ),
    .B_N(net2602),
    .Y(_03605_));
 sg13g2_o21ai_1 _08930_ (.B1(net2576),
    .Y(_03606_),
    .A1(net2602),
    .A2(\ChiselTop.wild.cpu.regs[30][0] ));
 sg13g2_o21ai_1 _08931_ (.B1(net2561),
    .Y(_03607_),
    .A1(_03605_),
    .A2(_03606_));
 sg13g2_o21ai_1 _08932_ (.B1(net2461),
    .Y(_03608_),
    .A1(_03604_),
    .A2(_03607_));
 sg13g2_nor2_1 _08933_ (.A(_03601_),
    .B(_03608_),
    .Y(_03609_));
 sg13g2_nor2_1 _08934_ (.A(net2404),
    .B(_03609_),
    .Y(_03610_));
 sg13g2_a21oi_2 _08935_ (.B1(_03610_),
    .Y(_03611_),
    .A2(net2404),
    .A1(net2137));
 sg13g2_nor2_1 _08936_ (.A(net2164),
    .B(_03611_),
    .Y(_03612_));
 sg13g2_a21oi_1 _08937_ (.A1(net2164),
    .A2(_03599_),
    .Y(_03613_),
    .B1(_03612_));
 sg13g2_mux2_1 _08938_ (.A0(_03613_),
    .A1(net1399),
    .S(_03579_),
    .X(_00198_));
 sg13g2_mux4_1 _08939_ (.S0(net2586),
    .A0(\ChiselTop.wild.cpu.regs[0][17] ),
    .A1(\ChiselTop.wild.cpu.regs[1][17] ),
    .A2(\ChiselTop.wild.cpu.regs[2][17] ),
    .A3(\ChiselTop.wild.cpu.regs[3][17] ),
    .S1(net2567),
    .X(_03614_));
 sg13g2_nor2_1 _08940_ (.A(net2554),
    .B(_03614_),
    .Y(_03615_));
 sg13g2_nor2b_1 _08941_ (.A(\ChiselTop.wild.cpu.regs[29][17] ),
    .B_N(net2586),
    .Y(_03616_));
 sg13g2_nor2_1 _08942_ (.A(net2586),
    .B(\ChiselTop.wild.cpu.regs[28][17] ),
    .Y(_03617_));
 sg13g2_nor3_1 _08943_ (.A(net2567),
    .B(_03616_),
    .C(_03617_),
    .Y(_03618_));
 sg13g2_nor2b_1 _08944_ (.A(\ChiselTop.wild.cpu.regs[31][17] ),
    .B_N(net2586),
    .Y(_03619_));
 sg13g2_o21ai_1 _08945_ (.B1(net2567),
    .Y(_03620_),
    .A1(net2586),
    .A2(\ChiselTop.wild.cpu.regs[30][17] ));
 sg13g2_o21ai_1 _08946_ (.B1(net2554),
    .Y(_03621_),
    .A1(_03619_),
    .A2(_03620_));
 sg13g2_o21ai_1 _08947_ (.B1(net2459),
    .Y(_03622_),
    .A1(_03618_),
    .A2(_03621_));
 sg13g2_nor2_1 _08948_ (.A(_03615_),
    .B(_03622_),
    .Y(_03623_));
 sg13g2_inv_2 _08949_ (.Y(_03624_),
    .A(_03623_));
 sg13g2_mux2_1 _08950_ (.A0(_03624_),
    .A1(net2116),
    .S(net2408),
    .X(_03625_));
 sg13g2_mux4_1 _08951_ (.S0(net2607),
    .A0(\ChiselTop.wild.cpu.regs[0][1] ),
    .A1(\ChiselTop.wild.cpu.regs[1][1] ),
    .A2(\ChiselTop.wild.cpu.regs[2][1] ),
    .A3(\ChiselTop.wild.cpu.regs[3][1] ),
    .S1(net2580),
    .X(_03626_));
 sg13g2_nor2_1 _08952_ (.A(net2562),
    .B(_03626_),
    .Y(_03627_));
 sg13g2_nor2b_1 _08953_ (.A(\ChiselTop.wild.cpu.regs[29][1] ),
    .B_N(net2606),
    .Y(_03628_));
 sg13g2_nor2_1 _08954_ (.A(net2608),
    .B(\ChiselTop.wild.cpu.regs[28][1] ),
    .Y(_03629_));
 sg13g2_nor3_1 _08955_ (.A(net2579),
    .B(_03628_),
    .C(_03629_),
    .Y(_03630_));
 sg13g2_nor2b_1 _08956_ (.A(\ChiselTop.wild.cpu.regs[31][1] ),
    .B_N(net2607),
    .Y(_03631_));
 sg13g2_o21ai_1 _08957_ (.B1(net2579),
    .Y(_03632_),
    .A1(net2607),
    .A2(\ChiselTop.wild.cpu.regs[30][1] ));
 sg13g2_o21ai_1 _08958_ (.B1(net2562),
    .Y(_03633_),
    .A1(_03631_),
    .A2(_03632_));
 sg13g2_o21ai_1 _08959_ (.B1(net2462),
    .Y(_03634_),
    .A1(_03630_),
    .A2(_03633_));
 sg13g2_nor2_1 _08960_ (.A(_03627_),
    .B(_03634_),
    .Y(_03635_));
 sg13g2_nor2_1 _08961_ (.A(net2412),
    .B(_03635_),
    .Y(_03636_));
 sg13g2_a21oi_2 _08962_ (.B1(_03636_),
    .Y(_03637_),
    .A2(net2412),
    .A1(net2147));
 sg13g2_nor2_1 _08963_ (.A(net2162),
    .B(_03637_),
    .Y(_03638_));
 sg13g2_a21oi_1 _08964_ (.A1(net2162),
    .A2(_03625_),
    .Y(_03639_),
    .B1(_03638_));
 sg13g2_mux2_1 _08965_ (.A0(_03639_),
    .A1(net1424),
    .S(_03579_),
    .X(_00199_));
 sg13g2_mux4_1 _08966_ (.S0(net2583),
    .A0(\ChiselTop.wild.cpu.regs[0][18] ),
    .A1(\ChiselTop.wild.cpu.regs[1][18] ),
    .A2(\ChiselTop.wild.cpu.regs[2][18] ),
    .A3(\ChiselTop.wild.cpu.regs[3][18] ),
    .S1(net2565),
    .X(_03640_));
 sg13g2_nor2_1 _08967_ (.A(net2554),
    .B(_03640_),
    .Y(_03641_));
 sg13g2_nor2b_1 _08968_ (.A(\ChiselTop.wild.cpu.regs[29][18] ),
    .B_N(net2583),
    .Y(_03642_));
 sg13g2_nor2_1 _08969_ (.A(net2590),
    .B(\ChiselTop.wild.cpu.regs[28][18] ),
    .Y(_03643_));
 sg13g2_nor3_1 _08970_ (.A(net2565),
    .B(_03642_),
    .C(_03643_),
    .Y(_03644_));
 sg13g2_nor2b_1 _08971_ (.A(\ChiselTop.wild.cpu.regs[31][18] ),
    .B_N(net2583),
    .Y(_03645_));
 sg13g2_o21ai_1 _08972_ (.B1(net2565),
    .Y(_03646_),
    .A1(net2583),
    .A2(\ChiselTop.wild.cpu.regs[30][18] ));
 sg13g2_o21ai_1 _08973_ (.B1(net2554),
    .Y(_03647_),
    .A1(_03645_),
    .A2(_03646_));
 sg13g2_o21ai_1 _08974_ (.B1(net2459),
    .Y(_03648_),
    .A1(_03644_),
    .A2(_03647_));
 sg13g2_nor2_1 _08975_ (.A(_03641_),
    .B(_03648_),
    .Y(_03649_));
 sg13g2_inv_2 _08976_ (.Y(_03650_),
    .A(_03649_));
 sg13g2_mux2_1 _08977_ (.A0(_03650_),
    .A1(net2107),
    .S(net2406),
    .X(_03651_));
 sg13g2_mux4_1 _08978_ (.S0(net2603),
    .A0(\ChiselTop.wild.cpu.regs[0][2] ),
    .A1(\ChiselTop.wild.cpu.regs[1][2] ),
    .A2(\ChiselTop.wild.cpu.regs[2][2] ),
    .A3(\ChiselTop.wild.cpu.regs[3][2] ),
    .S1(net2579),
    .X(_03652_));
 sg13g2_nor2_1 _08979_ (.A(net2563),
    .B(_03652_),
    .Y(_03653_));
 sg13g2_nor2b_1 _08980_ (.A(\ChiselTop.wild.cpu.regs[29][2] ),
    .B_N(net2608),
    .Y(_03654_));
 sg13g2_nor2_1 _08981_ (.A(net2608),
    .B(\ChiselTop.wild.cpu.regs[28][2] ),
    .Y(_03655_));
 sg13g2_nor3_1 _08982_ (.A(net2577),
    .B(_03654_),
    .C(_03655_),
    .Y(_03656_));
 sg13g2_nor2b_1 _08983_ (.A(\ChiselTop.wild.cpu.regs[31][2] ),
    .B_N(net2608),
    .Y(_03657_));
 sg13g2_o21ai_1 _08984_ (.B1(net2577),
    .Y(_03658_),
    .A1(net2606),
    .A2(\ChiselTop.wild.cpu.regs[30][2] ));
 sg13g2_o21ai_1 _08985_ (.B1(net2561),
    .Y(_03659_),
    .A1(_03657_),
    .A2(_03658_));
 sg13g2_o21ai_1 _08986_ (.B1(net2462),
    .Y(_03660_),
    .A1(_03656_),
    .A2(_03659_));
 sg13g2_nor2_1 _08987_ (.A(_03653_),
    .B(_03660_),
    .Y(_03661_));
 sg13g2_nor2_1 _08988_ (.A(net2404),
    .B(_03661_),
    .Y(_03662_));
 sg13g2_a21oi_2 _08989_ (.B1(_03662_),
    .Y(_03663_),
    .A2(net2404),
    .A1(net2138));
 sg13g2_nor2_1 _08990_ (.A(net2160),
    .B(_03663_),
    .Y(_03664_));
 sg13g2_a21oi_1 _08991_ (.A1(net2160),
    .A2(_03651_),
    .Y(_03665_),
    .B1(_03664_));
 sg13g2_mux2_1 _08992_ (.A0(_03665_),
    .A1(net1405),
    .S(_03579_),
    .X(_00200_));
 sg13g2_mux4_1 _08993_ (.S0(net2604),
    .A0(\ChiselTop.wild.cpu.regs[0][3] ),
    .A1(\ChiselTop.wild.cpu.regs[1][3] ),
    .A2(\ChiselTop.wild.cpu.regs[2][3] ),
    .A3(\ChiselTop.wild.cpu.regs[3][3] ),
    .S1(net2576),
    .X(_03666_));
 sg13g2_nor2_1 _08994_ (.A(net2561),
    .B(_03666_),
    .Y(_03667_));
 sg13g2_nor2b_1 _08995_ (.A(net1068),
    .B_N(net2604),
    .Y(_03668_));
 sg13g2_nor2_1 _08996_ (.A(net2602),
    .B(net1191),
    .Y(_03669_));
 sg13g2_nor3_1 _08997_ (.A(net2576),
    .B(_03668_),
    .C(_03669_),
    .Y(_03670_));
 sg13g2_nor2b_1 _08998_ (.A(\ChiselTop.wild.cpu.regs[31][3] ),
    .B_N(net2602),
    .Y(_03671_));
 sg13g2_o21ai_1 _08999_ (.B1(net2576),
    .Y(_03672_),
    .A1(net2602),
    .A2(\ChiselTop.wild.cpu.regs[30][3] ));
 sg13g2_o21ai_1 _09000_ (.B1(net2561),
    .Y(_03673_),
    .A1(_03671_),
    .A2(_03672_));
 sg13g2_o21ai_1 _09001_ (.B1(net2461),
    .Y(_03674_),
    .A1(_03670_),
    .A2(_03673_));
 sg13g2_nor2_1 _09002_ (.A(_03667_),
    .B(_03674_),
    .Y(_03675_));
 sg13g2_nor2_1 _09003_ (.A(net2404),
    .B(_03675_),
    .Y(_03676_));
 sg13g2_a21oi_2 _09004_ (.B1(_03676_),
    .Y(_03677_),
    .A2(net2404),
    .A1(net2135));
 sg13g2_nor2_1 _09005_ (.A(net2162),
    .B(_03677_),
    .Y(_03678_));
 sg13g2_mux4_1 _09006_ (.S0(net2598),
    .A0(\ChiselTop.wild.cpu.regs[0][19] ),
    .A1(\ChiselTop.wild.cpu.regs[1][19] ),
    .A2(\ChiselTop.wild.cpu.regs[2][19] ),
    .A3(\ChiselTop.wild.cpu.regs[3][19] ),
    .S1(net2574),
    .X(_03679_));
 sg13g2_nor2_1 _09007_ (.A(net2560),
    .B(_03679_),
    .Y(_03680_));
 sg13g2_nor2b_1 _09008_ (.A(\ChiselTop.wild.cpu.regs[29][19] ),
    .B_N(net2598),
    .Y(_03681_));
 sg13g2_nor2_1 _09009_ (.A(net2598),
    .B(\ChiselTop.wild.cpu.regs[28][19] ),
    .Y(_03682_));
 sg13g2_nor3_1 _09010_ (.A(net2574),
    .B(_03681_),
    .C(_03682_),
    .Y(_03683_));
 sg13g2_nor2b_1 _09011_ (.A(\ChiselTop.wild.cpu.regs[31][19] ),
    .B_N(net2598),
    .Y(_03684_));
 sg13g2_o21ai_1 _09012_ (.B1(net2574),
    .Y(_03685_),
    .A1(net2598),
    .A2(\ChiselTop.wild.cpu.regs[30][19] ));
 sg13g2_o21ai_1 _09013_ (.B1(net2560),
    .Y(_03686_),
    .A1(_03684_),
    .A2(_03685_));
 sg13g2_o21ai_1 _09014_ (.B1(net2461),
    .Y(_03687_),
    .A1(_03683_),
    .A2(_03686_));
 sg13g2_nor2_1 _09015_ (.A(_03680_),
    .B(_03687_),
    .Y(_03688_));
 sg13g2_inv_2 _09016_ (.Y(_03689_),
    .A(_03688_));
 sg13g2_mux2_1 _09017_ (.A0(_03689_),
    .A1(net2110),
    .S(net2410),
    .X(_03690_));
 sg13g2_a21oi_1 _09018_ (.A1(net2162),
    .A2(_03690_),
    .Y(_03691_),
    .B1(_03678_));
 sg13g2_mux2_1 _09019_ (.A0(_03691_),
    .A1(net1346),
    .S(_03579_),
    .X(_00201_));
 sg13g2_mux4_1 _09020_ (.S0(net2594),
    .A0(\ChiselTop.wild.cpu.regs[0][20] ),
    .A1(\ChiselTop.wild.cpu.regs[1][20] ),
    .A2(\ChiselTop.wild.cpu.regs[2][20] ),
    .A3(\ChiselTop.wild.cpu.regs[3][20] ),
    .S1(net2570),
    .X(_03692_));
 sg13g2_nor2_1 _09021_ (.A(net2557),
    .B(_03692_),
    .Y(_03693_));
 sg13g2_nor2b_1 _09022_ (.A(\ChiselTop.wild.cpu.regs[29][20] ),
    .B_N(net2593),
    .Y(_03694_));
 sg13g2_nor2_1 _09023_ (.A(net2593),
    .B(\ChiselTop.wild.cpu.regs[28][20] ),
    .Y(_03695_));
 sg13g2_nor3_1 _09024_ (.A(net2570),
    .B(_03694_),
    .C(_03695_),
    .Y(_03696_));
 sg13g2_nor2b_1 _09025_ (.A(\ChiselTop.wild.cpu.regs[31][20] ),
    .B_N(net2593),
    .Y(_03697_));
 sg13g2_o21ai_1 _09026_ (.B1(net2570),
    .Y(_03698_),
    .A1(net2593),
    .A2(\ChiselTop.wild.cpu.regs[30][20] ));
 sg13g2_o21ai_1 _09027_ (.B1(net2556),
    .Y(_03699_),
    .A1(_03697_),
    .A2(_03698_));
 sg13g2_o21ai_1 _09028_ (.B1(net2463),
    .Y(_03700_),
    .A1(_03696_),
    .A2(_03699_));
 sg13g2_nor3_2 _09029_ (.A(net2406),
    .B(_03693_),
    .C(_03700_),
    .Y(_03701_));
 sg13g2_a21oi_1 _09030_ (.A1(_03157_),
    .A2(net2412),
    .Y(_03702_),
    .B1(_03701_));
 sg13g2_mux4_1 _09031_ (.S0(net2603),
    .A0(\ChiselTop.wild.cpu.regs[0][4] ),
    .A1(\ChiselTop.wild.cpu.regs[1][4] ),
    .A2(\ChiselTop.wild.cpu.regs[2][4] ),
    .A3(\ChiselTop.wild.cpu.regs[3][4] ),
    .S1(net2577),
    .X(_03703_));
 sg13g2_nor2_1 _09032_ (.A(net2561),
    .B(_03703_),
    .Y(_03704_));
 sg13g2_nor2b_1 _09033_ (.A(\ChiselTop.wild.cpu.regs[29][4] ),
    .B_N(net2604),
    .Y(_03705_));
 sg13g2_nor2_1 _09034_ (.A(net2604),
    .B(\ChiselTop.wild.cpu.regs[28][4] ),
    .Y(_03706_));
 sg13g2_nor3_1 _09035_ (.A(net2576),
    .B(_03705_),
    .C(_03706_),
    .Y(_03707_));
 sg13g2_nor2b_1 _09036_ (.A(\ChiselTop.wild.cpu.regs[31][4] ),
    .B_N(net2603),
    .Y(_03708_));
 sg13g2_o21ai_1 _09037_ (.B1(net2577),
    .Y(_03709_),
    .A1(net2603),
    .A2(\ChiselTop.wild.cpu.regs[30][4] ));
 sg13g2_o21ai_1 _09038_ (.B1(net2561),
    .Y(_03710_),
    .A1(_03708_),
    .A2(_03709_));
 sg13g2_o21ai_1 _09039_ (.B1(net2461),
    .Y(_03711_),
    .A1(_03707_),
    .A2(_03710_));
 sg13g2_nor2_1 _09040_ (.A(_03704_),
    .B(_03711_),
    .Y(_03712_));
 sg13g2_nor2_1 _09041_ (.A(net2404),
    .B(_03712_),
    .Y(_03713_));
 sg13g2_a21oi_2 _09042_ (.B1(_03713_),
    .Y(_03714_),
    .A2(net2405),
    .A1(net2152));
 sg13g2_nor2_1 _09043_ (.A(net2163),
    .B(_03714_),
    .Y(_03715_));
 sg13g2_a21oi_2 _09044_ (.B1(_03715_),
    .Y(_03716_),
    .A2(_03702_),
    .A1(net2161));
 sg13g2_mux2_1 _09045_ (.A0(_03716_),
    .A1(net1446),
    .S(_03579_),
    .X(_00202_));
 sg13g2_mux4_1 _09046_ (.S0(net2594),
    .A0(\ChiselTop.wild.cpu.regs[0][21] ),
    .A1(\ChiselTop.wild.cpu.regs[1][21] ),
    .A2(\ChiselTop.wild.cpu.regs[2][21] ),
    .A3(\ChiselTop.wild.cpu.regs[3][21] ),
    .S1(net2570),
    .X(_03717_));
 sg13g2_nor2_1 _09047_ (.A(net2557),
    .B(_03717_),
    .Y(_03718_));
 sg13g2_nor2b_1 _09048_ (.A(\ChiselTop.wild.cpu.regs[29][21] ),
    .B_N(net2592),
    .Y(_03719_));
 sg13g2_nor2_1 _09049_ (.A(net2592),
    .B(\ChiselTop.wild.cpu.regs[28][21] ),
    .Y(_03720_));
 sg13g2_nor3_1 _09050_ (.A(net2571),
    .B(_03719_),
    .C(_03720_),
    .Y(_03721_));
 sg13g2_nor2b_1 _09051_ (.A(\ChiselTop.wild.cpu.regs[31][21] ),
    .B_N(net2591),
    .Y(_03722_));
 sg13g2_o21ai_1 _09052_ (.B1(net2571),
    .Y(_03723_),
    .A1(net2591),
    .A2(\ChiselTop.wild.cpu.regs[30][21] ));
 sg13g2_o21ai_1 _09053_ (.B1(net2556),
    .Y(_03724_),
    .A1(_03722_),
    .A2(_03723_));
 sg13g2_o21ai_1 _09054_ (.B1(net2463),
    .Y(_03725_),
    .A1(_03721_),
    .A2(_03724_));
 sg13g2_nor3_2 _09055_ (.A(net2407),
    .B(_03718_),
    .C(_03725_),
    .Y(_03726_));
 sg13g2_a21oi_1 _09056_ (.A1(_03118_),
    .A2(net2410),
    .Y(_03727_),
    .B1(_03726_));
 sg13g2_mux4_1 _09057_ (.S0(net2600),
    .A0(\ChiselTop.wild.cpu.regs[0][5] ),
    .A1(\ChiselTop.wild.cpu.regs[1][5] ),
    .A2(\ChiselTop.wild.cpu.regs[2][5] ),
    .A3(\ChiselTop.wild.cpu.regs[3][5] ),
    .S1(net2575),
    .X(_03728_));
 sg13g2_nor2_1 _09058_ (.A(net2560),
    .B(_03728_),
    .Y(_03729_));
 sg13g2_nor2b_1 _09059_ (.A(\ChiselTop.wild.cpu.regs[29][5] ),
    .B_N(net2598),
    .Y(_03730_));
 sg13g2_nor2_1 _09060_ (.A(net2598),
    .B(\ChiselTop.wild.cpu.regs[28][5] ),
    .Y(_03731_));
 sg13g2_nor3_1 _09061_ (.A(net2574),
    .B(_03730_),
    .C(_03731_),
    .Y(_03732_));
 sg13g2_nor2b_1 _09062_ (.A(\ChiselTop.wild.cpu.regs[31][5] ),
    .B_N(net2599),
    .Y(_03733_));
 sg13g2_o21ai_1 _09063_ (.B1(net2574),
    .Y(_03734_),
    .A1(net2598),
    .A2(\ChiselTop.wild.cpu.regs[30][5] ));
 sg13g2_o21ai_1 _09064_ (.B1(net2560),
    .Y(_03735_),
    .A1(_03733_),
    .A2(_03734_));
 sg13g2_o21ai_1 _09065_ (.B1(net2461),
    .Y(_03736_),
    .A1(_03732_),
    .A2(_03735_));
 sg13g2_nor2_1 _09066_ (.A(_03729_),
    .B(_03736_),
    .Y(_03737_));
 sg13g2_nor2_1 _09067_ (.A(net2404),
    .B(_03737_),
    .Y(_03738_));
 sg13g2_a21oi_2 _09068_ (.B1(_03738_),
    .Y(_03739_),
    .A2(net2413),
    .A1(net2142));
 sg13g2_nor2_1 _09069_ (.A(net2160),
    .B(_03739_),
    .Y(_03740_));
 sg13g2_a21oi_1 _09070_ (.A1(net2161),
    .A2(_03727_),
    .Y(_03741_),
    .B1(_03740_));
 sg13g2_mux2_1 _09071_ (.A0(_03741_),
    .A1(net1451),
    .S(_03579_),
    .X(_00203_));
 sg13g2_mux4_1 _09072_ (.S0(net2596),
    .A0(\ChiselTop.wild.cpu.regs[0][6] ),
    .A1(\ChiselTop.wild.cpu.regs[1][6] ),
    .A2(\ChiselTop.wild.cpu.regs[2][6] ),
    .A3(\ChiselTop.wild.cpu.regs[3][6] ),
    .S1(net2572),
    .X(_03742_));
 sg13g2_nor2_1 _09073_ (.A(net2558),
    .B(_03742_),
    .Y(_03743_));
 sg13g2_nor2b_1 _09074_ (.A(\ChiselTop.wild.cpu.regs[29][6] ),
    .B_N(net2596),
    .Y(_03744_));
 sg13g2_nor2_1 _09075_ (.A(net2596),
    .B(\ChiselTop.wild.cpu.regs[28][6] ),
    .Y(_03745_));
 sg13g2_nor3_1 _09076_ (.A(net2573),
    .B(_03744_),
    .C(_03745_),
    .Y(_03746_));
 sg13g2_nor2b_1 _09077_ (.A(\ChiselTop.wild.cpu.regs[31][6] ),
    .B_N(net2596),
    .Y(_03747_));
 sg13g2_o21ai_1 _09078_ (.B1(net2572),
    .Y(_03748_),
    .A1(net2596),
    .A2(\ChiselTop.wild.cpu.regs[30][6] ));
 sg13g2_o21ai_1 _09079_ (.B1(net2558),
    .Y(_03749_),
    .A1(_03747_),
    .A2(_03748_));
 sg13g2_o21ai_1 _09080_ (.B1(net2460),
    .Y(_03750_),
    .A1(_03746_),
    .A2(_03749_));
 sg13g2_nor2_1 _09081_ (.A(_03743_),
    .B(_03750_),
    .Y(_03751_));
 sg13g2_nor2_1 _09082_ (.A(net2408),
    .B(_03751_),
    .Y(_03752_));
 sg13g2_a21oi_2 _09083_ (.B1(_03752_),
    .Y(_03753_),
    .A2(net2407),
    .A1(net2144));
 sg13g2_nor2_1 _09084_ (.A(net2163),
    .B(_03753_),
    .Y(_03754_));
 sg13g2_mux4_1 _09085_ (.S0(net2583),
    .A0(\ChiselTop.wild.cpu.regs[0][22] ),
    .A1(\ChiselTop.wild.cpu.regs[1][22] ),
    .A2(\ChiselTop.wild.cpu.regs[2][22] ),
    .A3(\ChiselTop.wild.cpu.regs[3][22] ),
    .S1(net2566),
    .X(_03755_));
 sg13g2_nor2_1 _09086_ (.A(net2555),
    .B(_03755_),
    .Y(_03756_));
 sg13g2_nor2b_1 _09087_ (.A(\ChiselTop.wild.cpu.regs[29][22] ),
    .B_N(net2583),
    .Y(_03757_));
 sg13g2_nor2_1 _09088_ (.A(net2584),
    .B(\ChiselTop.wild.cpu.regs[28][22] ),
    .Y(_03758_));
 sg13g2_nor3_1 _09089_ (.A(net2565),
    .B(_03757_),
    .C(_03758_),
    .Y(_03759_));
 sg13g2_nor2b_1 _09090_ (.A(\ChiselTop.wild.cpu.regs[31][22] ),
    .B_N(net2583),
    .Y(_03760_));
 sg13g2_o21ai_1 _09091_ (.B1(net2565),
    .Y(_03761_),
    .A1(net2583),
    .A2(\ChiselTop.wild.cpu.regs[30][22] ));
 sg13g2_o21ai_1 _09092_ (.B1(net2554),
    .Y(_03762_),
    .A1(_03760_),
    .A2(_03761_));
 sg13g2_o21ai_1 _09093_ (.B1(net2459),
    .Y(_03763_),
    .A1(_03759_),
    .A2(_03762_));
 sg13g2_nor2_1 _09094_ (.A(_03756_),
    .B(_03763_),
    .Y(_03764_));
 sg13g2_inv_2 _09095_ (.Y(_03765_),
    .A(_03764_));
 sg13g2_mux2_2 _09096_ (.A0(_03765_),
    .A1(net2095),
    .S(net2407),
    .X(_03766_));
 sg13g2_a21oi_1 _09097_ (.A1(net2162),
    .A2(_03766_),
    .Y(_03767_),
    .B1(_03754_));
 sg13g2_mux2_1 _09098_ (.A0(_03767_),
    .A1(net1474),
    .S(_03579_),
    .X(_00204_));
 sg13g2_mux4_1 _09099_ (.S0(net2592),
    .A0(\ChiselTop.wild.cpu.regs[0][23] ),
    .A1(\ChiselTop.wild.cpu.regs[1][23] ),
    .A2(\ChiselTop.wild.cpu.regs[2][23] ),
    .A3(\ChiselTop.wild.cpu.regs[3][23] ),
    .S1(net2571),
    .X(_03768_));
 sg13g2_nor2_2 _09100_ (.A(net2556),
    .B(_03768_),
    .Y(_03769_));
 sg13g2_nor2b_1 _09101_ (.A(\ChiselTop.wild.cpu.regs[29][23] ),
    .B_N(net2592),
    .Y(_03770_));
 sg13g2_nor2_1 _09102_ (.A(net2591),
    .B(\ChiselTop.wild.cpu.regs[28][23] ),
    .Y(_03771_));
 sg13g2_nor3_1 _09103_ (.A(net2571),
    .B(_03770_),
    .C(_03771_),
    .Y(_03772_));
 sg13g2_nor2b_1 _09104_ (.A(\ChiselTop.wild.cpu.regs[31][23] ),
    .B_N(net2591),
    .Y(_03773_));
 sg13g2_o21ai_1 _09105_ (.B1(net2572),
    .Y(_03774_),
    .A1(net2595),
    .A2(\ChiselTop.wild.cpu.regs[30][23] ));
 sg13g2_o21ai_1 _09106_ (.B1(net2556),
    .Y(_03775_),
    .A1(_03773_),
    .A2(_03774_));
 sg13g2_o21ai_1 _09107_ (.B1(net2463),
    .Y(_03776_),
    .A1(_03772_),
    .A2(_03775_));
 sg13g2_nor3_2 _09108_ (.A(net2406),
    .B(_03769_),
    .C(_03776_),
    .Y(_03777_));
 sg13g2_a21oi_1 _09109_ (.A1(_03001_),
    .A2(net2412),
    .Y(_03778_),
    .B1(_03777_));
 sg13g2_mux4_1 _09110_ (.S0(net2595),
    .A0(\ChiselTop.wild.cpu.regs[0][7] ),
    .A1(\ChiselTop.wild.cpu.regs[1][7] ),
    .A2(\ChiselTop.wild.cpu.regs[2][7] ),
    .A3(\ChiselTop.wild.cpu.regs[3][7] ),
    .S1(net2572),
    .X(_03779_));
 sg13g2_nor2_1 _09111_ (.A(net2558),
    .B(_03779_),
    .Y(_03780_));
 sg13g2_nor2b_1 _09112_ (.A(\ChiselTop.wild.cpu.regs[29][7] ),
    .B_N(net2595),
    .Y(_03781_));
 sg13g2_nor2_1 _09113_ (.A(net2595),
    .B(\ChiselTop.wild.cpu.regs[28][7] ),
    .Y(_03782_));
 sg13g2_nor3_1 _09114_ (.A(net2572),
    .B(_03781_),
    .C(_03782_),
    .Y(_03783_));
 sg13g2_nor2b_1 _09115_ (.A(\ChiselTop.wild.cpu.regs[31][7] ),
    .B_N(net2595),
    .Y(_03784_));
 sg13g2_o21ai_1 _09116_ (.B1(net2572),
    .Y(_03785_),
    .A1(net2595),
    .A2(\ChiselTop.wild.cpu.regs[30][7] ));
 sg13g2_o21ai_1 _09117_ (.B1(net2558),
    .Y(_03786_),
    .A1(_03784_),
    .A2(_03785_));
 sg13g2_o21ai_1 _09118_ (.B1(net2460),
    .Y(_03787_),
    .A1(_03783_),
    .A2(_03786_));
 sg13g2_nor2_1 _09119_ (.A(_03780_),
    .B(_03787_),
    .Y(_03788_));
 sg13g2_nor2_1 _09120_ (.A(net2406),
    .B(_03788_),
    .Y(_03789_));
 sg13g2_a21oi_2 _09121_ (.B1(_03789_),
    .Y(_03790_),
    .A2(net2406),
    .A1(net2146));
 sg13g2_nor2_1 _09122_ (.A(net2160),
    .B(_03790_),
    .Y(_03791_));
 sg13g2_a21oi_2 _09123_ (.B1(_03791_),
    .Y(_03792_),
    .A2(_03778_),
    .A1(net2160));
 sg13g2_mux2_1 _09124_ (.A0(_03792_),
    .A1(net1459),
    .S(_03579_),
    .X(_00205_));
 sg13g2_o21ai_1 _09125_ (.B1(net2550),
    .Y(_03793_),
    .A1(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[13] ),
    .A2(_03574_));
 sg13g2_o21ai_1 _09126_ (.B1(_03563_),
    .Y(_03794_),
    .A1(_02000_),
    .A2(_02638_));
 sg13g2_nor2_1 _09127_ (.A(net2527),
    .B(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[13] ),
    .Y(_03795_));
 sg13g2_nand4_1 _09128_ (.B(_03576_),
    .C(_03793_),
    .A(_03572_),
    .Y(_03796_),
    .D(_03794_));
 sg13g2_mux4_1 _09129_ (.S0(net2588),
    .A0(\ChiselTop.wild.cpu.regs[0][8] ),
    .A1(\ChiselTop.wild.cpu.regs[1][8] ),
    .A2(\ChiselTop.wild.cpu.regs[2][8] ),
    .A3(\ChiselTop.wild.cpu.regs[3][8] ),
    .S1(net2568),
    .X(_03797_));
 sg13g2_nor2_1 _09130_ (.A(net2554),
    .B(_03797_),
    .Y(_03798_));
 sg13g2_nor2b_1 _09131_ (.A(\ChiselTop.wild.cpu.regs[29][8] ),
    .B_N(net2588),
    .Y(_03799_));
 sg13g2_nor2_1 _09132_ (.A(net2588),
    .B(\ChiselTop.wild.cpu.regs[28][8] ),
    .Y(_03800_));
 sg13g2_nor3_1 _09133_ (.A(net2568),
    .B(_03799_),
    .C(_03800_),
    .Y(_03801_));
 sg13g2_nor2b_1 _09134_ (.A(\ChiselTop.wild.cpu.regs[31][8] ),
    .B_N(net2588),
    .Y(_03802_));
 sg13g2_o21ai_1 _09135_ (.B1(net2568),
    .Y(_03803_),
    .A1(net2588),
    .A2(\ChiselTop.wild.cpu.regs[30][8] ));
 sg13g2_o21ai_1 _09136_ (.B1(net2554),
    .Y(_03804_),
    .A1(_03802_),
    .A2(_03803_));
 sg13g2_o21ai_1 _09137_ (.B1(net2459),
    .Y(_03805_),
    .A1(_03801_),
    .A2(_03804_));
 sg13g2_nor2_1 _09138_ (.A(_03798_),
    .B(_03805_),
    .Y(_03806_));
 sg13g2_nor2_1 _09139_ (.A(net2405),
    .B(_03806_),
    .Y(_03807_));
 sg13g2_a21oi_2 _09140_ (.B1(_03807_),
    .Y(_03808_),
    .A2(net2405),
    .A1(net2131));
 sg13g2_mux2_1 _09141_ (.A0(_03611_),
    .A1(_03808_),
    .S(net2164),
    .X(_03809_));
 sg13g2_mux2_1 _09142_ (.A0(_03809_),
    .A1(net1423),
    .S(_03796_),
    .X(_00206_));
 sg13g2_mux4_1 _09143_ (.S0(net2585),
    .A0(\ChiselTop.wild.cpu.regs[0][9] ),
    .A1(\ChiselTop.wild.cpu.regs[1][9] ),
    .A2(\ChiselTop.wild.cpu.regs[2][9] ),
    .A3(\ChiselTop.wild.cpu.regs[3][9] ),
    .S1(net2565),
    .X(_03810_));
 sg13g2_nor2_1 _09144_ (.A(net2554),
    .B(_03810_),
    .Y(_03811_));
 sg13g2_nor2b_1 _09145_ (.A(net1039),
    .B_N(net2584),
    .Y(_03812_));
 sg13g2_nor2_1 _09146_ (.A(net2584),
    .B(net1549),
    .Y(_03813_));
 sg13g2_nor3_1 _09147_ (.A(net2565),
    .B(_03812_),
    .C(_03813_),
    .Y(_03814_));
 sg13g2_nor2b_1 _09148_ (.A(\ChiselTop.wild.cpu.regs[31][9] ),
    .B_N(net2584),
    .Y(_03815_));
 sg13g2_o21ai_1 _09149_ (.B1(net2566),
    .Y(_03816_),
    .A1(net2584),
    .A2(\ChiselTop.wild.cpu.regs[30][9] ));
 sg13g2_o21ai_1 _09150_ (.B1(net2555),
    .Y(_03817_),
    .A1(_03815_),
    .A2(_03816_));
 sg13g2_o21ai_1 _09151_ (.B1(net2459),
    .Y(_03818_),
    .A1(_03814_),
    .A2(_03817_));
 sg13g2_nor2_1 _09152_ (.A(_03811_),
    .B(_03818_),
    .Y(_03819_));
 sg13g2_nand2_1 _09153_ (.Y(_03820_),
    .A(net2129),
    .B(net2405));
 sg13g2_o21ai_1 _09154_ (.B1(_03820_),
    .Y(_03821_),
    .A1(net2405),
    .A2(_03819_));
 sg13g2_a21oi_1 _09155_ (.A1(net2162),
    .A2(_03821_),
    .Y(_03822_),
    .B1(_03638_));
 sg13g2_mux2_1 _09156_ (.A0(_03822_),
    .A1(net1439),
    .S(_03796_),
    .X(_00207_));
 sg13g2_mux4_1 _09157_ (.S0(net2589),
    .A0(\ChiselTop.wild.cpu.regs[0][10] ),
    .A1(\ChiselTop.wild.cpu.regs[1][10] ),
    .A2(\ChiselTop.wild.cpu.regs[2][10] ),
    .A3(\ChiselTop.wild.cpu.regs[3][10] ),
    .S1(net2568),
    .X(_03823_));
 sg13g2_nor2_1 _09158_ (.A(net2555),
    .B(_03823_),
    .Y(_03824_));
 sg13g2_nor2b_1 _09159_ (.A(net1550),
    .B_N(net2600),
    .Y(_03825_));
 sg13g2_nor2_1 _09160_ (.A(net2600),
    .B(\ChiselTop.wild.cpu.regs[28][10] ),
    .Y(_03826_));
 sg13g2_nor3_1 _09161_ (.A(net2575),
    .B(_03825_),
    .C(_03826_),
    .Y(_03827_));
 sg13g2_nor2b_1 _09162_ (.A(\ChiselTop.wild.cpu.regs[31][10] ),
    .B_N(net2589),
    .Y(_03828_));
 sg13g2_o21ai_1 _09163_ (.B1(net2575),
    .Y(_03829_),
    .A1(net2600),
    .A2(\ChiselTop.wild.cpu.regs[30][10] ));
 sg13g2_o21ai_1 _09164_ (.B1(net2555),
    .Y(_03830_),
    .A1(_03828_),
    .A2(_03829_));
 sg13g2_o21ai_1 _09165_ (.B1(net2459),
    .Y(_03831_),
    .A1(net1551),
    .A2(_03830_));
 sg13g2_nor2_1 _09166_ (.A(_03824_),
    .B(_03831_),
    .Y(_03832_));
 sg13g2_nand2_1 _09167_ (.Y(_03833_),
    .A(net2133),
    .B(net2405));
 sg13g2_o21ai_1 _09168_ (.B1(_03833_),
    .Y(_03834_),
    .A1(net2405),
    .A2(_03832_));
 sg13g2_a21oi_1 _09169_ (.A1(net2160),
    .A2(_03834_),
    .Y(_03835_),
    .B1(_03664_));
 sg13g2_mux2_1 _09170_ (.A0(_03835_),
    .A1(net1492),
    .S(_03796_),
    .X(_00208_));
 sg13g2_mux4_1 _09171_ (.S0(net2594),
    .A0(\ChiselTop.wild.cpu.regs[0][11] ),
    .A1(\ChiselTop.wild.cpu.regs[1][11] ),
    .A2(\ChiselTop.wild.cpu.regs[2][11] ),
    .A3(\ChiselTop.wild.cpu.regs[3][11] ),
    .S1(net2570),
    .X(_03836_));
 sg13g2_nor2_1 _09172_ (.A(net2557),
    .B(_03836_),
    .Y(_03837_));
 sg13g2_nor2b_1 _09173_ (.A(net1053),
    .B_N(net2597),
    .Y(_03838_));
 sg13g2_nor2_1 _09174_ (.A(net2594),
    .B(net1117),
    .Y(_03839_));
 sg13g2_nor3_1 _09175_ (.A(net2571),
    .B(_03838_),
    .C(_03839_),
    .Y(_03840_));
 sg13g2_nor2b_1 _09176_ (.A(\ChiselTop.wild.cpu.regs[31][11] ),
    .B_N(net2593),
    .Y(_03841_));
 sg13g2_o21ai_1 _09177_ (.B1(net2573),
    .Y(_03842_),
    .A1(net2593),
    .A2(\ChiselTop.wild.cpu.regs[30][11] ));
 sg13g2_o21ai_1 _09178_ (.B1(net2557),
    .Y(_03843_),
    .A1(_03841_),
    .A2(_03842_));
 sg13g2_o21ai_1 _09179_ (.B1(net2460),
    .Y(_03844_),
    .A1(_03840_),
    .A2(_03843_));
 sg13g2_nor3_1 _09180_ (.A(net2407),
    .B(_03837_),
    .C(_03844_),
    .Y(_03845_));
 sg13g2_a21oi_2 _09181_ (.B1(_03845_),
    .Y(_03846_),
    .A2(net2407),
    .A1(net2124));
 sg13g2_a21oi_1 _09182_ (.A1(net2164),
    .A2(_03846_),
    .Y(_03847_),
    .B1(_03678_));
 sg13g2_mux2_1 _09183_ (.A0(_03847_),
    .A1(net1471),
    .S(_03796_),
    .X(_00209_));
 sg13g2_mux4_1 _09184_ (.S0(net2594),
    .A0(\ChiselTop.wild.cpu.regs[0][12] ),
    .A1(\ChiselTop.wild.cpu.regs[1][12] ),
    .A2(\ChiselTop.wild.cpu.regs[2][12] ),
    .A3(\ChiselTop.wild.cpu.regs[3][12] ),
    .S1(net2570),
    .X(_03848_));
 sg13g2_nor2_1 _09185_ (.A(net2557),
    .B(_03848_),
    .Y(_03849_));
 sg13g2_nor2b_1 _09186_ (.A(net1545),
    .B_N(net2594),
    .Y(_03850_));
 sg13g2_nor2_1 _09187_ (.A(net2594),
    .B(net1179),
    .Y(_03851_));
 sg13g2_nor3_1 _09188_ (.A(net2570),
    .B(_03850_),
    .C(_03851_),
    .Y(_03852_));
 sg13g2_nor2b_1 _09189_ (.A(\ChiselTop.wild.cpu.regs[31][12] ),
    .B_N(net2593),
    .Y(_03853_));
 sg13g2_o21ai_1 _09190_ (.B1(net2570),
    .Y(_03854_),
    .A1(net2593),
    .A2(\ChiselTop.wild.cpu.regs[30][12] ));
 sg13g2_o21ai_1 _09191_ (.B1(net2556),
    .Y(_03855_),
    .A1(_03853_),
    .A2(_03854_));
 sg13g2_o21ai_1 _09192_ (.B1(net2460),
    .Y(_03856_),
    .A1(_03852_),
    .A2(_03855_));
 sg13g2_nor2_1 _09193_ (.A(_03849_),
    .B(_03856_),
    .Y(_03857_));
 sg13g2_nand2_1 _09194_ (.Y(_03858_),
    .A(net2126),
    .B(net2406));
 sg13g2_o21ai_1 _09195_ (.B1(_03858_),
    .Y(_03859_),
    .A1(net2406),
    .A2(_03857_));
 sg13g2_a21oi_1 _09196_ (.A1(net2161),
    .A2(_03859_),
    .Y(_03860_),
    .B1(_03715_));
 sg13g2_mux2_1 _09197_ (.A0(_03860_),
    .A1(net1490),
    .S(_03796_),
    .X(_00210_));
 sg13g2_mux4_1 _09198_ (.S0(net2595),
    .A0(\ChiselTop.wild.cpu.regs[0][13] ),
    .A1(\ChiselTop.wild.cpu.regs[1][13] ),
    .A2(\ChiselTop.wild.cpu.regs[2][13] ),
    .A3(\ChiselTop.wild.cpu.regs[3][13] ),
    .S1(net2572),
    .X(_03861_));
 sg13g2_nor2_1 _09199_ (.A(net2558),
    .B(_03861_),
    .Y(_03862_));
 sg13g2_nor2b_1 _09200_ (.A(\ChiselTop.wild.cpu.regs[29][13] ),
    .B_N(net2589),
    .Y(_03863_));
 sg13g2_nor2_1 _09201_ (.A(net2596),
    .B(\ChiselTop.wild.cpu.regs[28][13] ),
    .Y(_03864_));
 sg13g2_nor3_1 _09202_ (.A(net2568),
    .B(_03863_),
    .C(_03864_),
    .Y(_03865_));
 sg13g2_nor2b_1 _09203_ (.A(\ChiselTop.wild.cpu.regs[31][13] ),
    .B_N(net2588),
    .Y(_03866_));
 sg13g2_o21ai_1 _09204_ (.B1(net2568),
    .Y(_03867_),
    .A1(net2588),
    .A2(\ChiselTop.wild.cpu.regs[30][13] ));
 sg13g2_o21ai_1 _09205_ (.B1(net2555),
    .Y(_03868_),
    .A1(_03866_),
    .A2(_03867_));
 sg13g2_o21ai_1 _09206_ (.B1(net2459),
    .Y(_03869_),
    .A1(_03865_),
    .A2(_03868_));
 sg13g2_nor2_1 _09207_ (.A(_03862_),
    .B(_03869_),
    .Y(_03870_));
 sg13g2_nand2_1 _09208_ (.Y(_03871_),
    .A(net2122),
    .B(net2408));
 sg13g2_o21ai_1 _09209_ (.B1(_03871_),
    .Y(_03872_),
    .A1(net2406),
    .A2(_03870_));
 sg13g2_a21oi_1 _09210_ (.A1(net2160),
    .A2(_03872_),
    .Y(_03873_),
    .B1(_03740_));
 sg13g2_mux2_1 _09211_ (.A0(_03873_),
    .A1(net1493),
    .S(_03796_),
    .X(_00211_));
 sg13g2_mux4_1 _09212_ (.S0(net2591),
    .A0(\ChiselTop.wild.cpu.regs[0][14] ),
    .A1(\ChiselTop.wild.cpu.regs[1][14] ),
    .A2(\ChiselTop.wild.cpu.regs[2][14] ),
    .A3(\ChiselTop.wild.cpu.regs[3][14] ),
    .S1(net2571),
    .X(_03874_));
 sg13g2_nor2_1 _09213_ (.A(net2556),
    .B(_03874_),
    .Y(_03875_));
 sg13g2_nor2b_1 _09214_ (.A(net951),
    .B_N(net2591),
    .Y(_03876_));
 sg13g2_nor2_1 _09215_ (.A(net2591),
    .B(net1055),
    .Y(_03877_));
 sg13g2_nor3_1 _09216_ (.A(net2571),
    .B(_03876_),
    .C(_03877_),
    .Y(_03878_));
 sg13g2_nor2b_1 _09217_ (.A(net1543),
    .B_N(net2591),
    .Y(_03879_));
 sg13g2_o21ai_1 _09218_ (.B1(net2572),
    .Y(_03880_),
    .A1(net2595),
    .A2(\ChiselTop.wild.cpu.regs[30][14] ));
 sg13g2_o21ai_1 _09219_ (.B1(net2556),
    .Y(_03881_),
    .A1(_03879_),
    .A2(_03880_));
 sg13g2_o21ai_1 _09220_ (.B1(net2460),
    .Y(_03882_),
    .A1(_03878_),
    .A2(_03881_));
 sg13g2_nor2_1 _09221_ (.A(_03875_),
    .B(_03882_),
    .Y(_03883_));
 sg13g2_nand2_1 _09222_ (.Y(_03884_),
    .A(net2120),
    .B(net2407));
 sg13g2_o21ai_1 _09223_ (.B1(_03884_),
    .Y(_03885_),
    .A1(net2407),
    .A2(_03883_));
 sg13g2_a21oi_1 _09224_ (.A1(net2162),
    .A2(_03885_),
    .Y(_03886_),
    .B1(_03754_));
 sg13g2_mux2_1 _09225_ (.A0(_03886_),
    .A1(net1465),
    .S(_03796_),
    .X(_00212_));
 sg13g2_mux4_1 _09226_ (.S0(net2605),
    .A0(\ChiselTop.wild.cpu.regs[0][15] ),
    .A1(\ChiselTop.wild.cpu.regs[1][15] ),
    .A2(\ChiselTop.wild.cpu.regs[2][15] ),
    .A3(\ChiselTop.wild.cpu.regs[3][15] ),
    .S1(net2581),
    .X(_03887_));
 sg13g2_nor2_1 _09227_ (.A(net2562),
    .B(_03887_),
    .Y(_03888_));
 sg13g2_nor2b_1 _09228_ (.A(\ChiselTop.wild.cpu.regs[29][15] ),
    .B_N(net2605),
    .Y(_03889_));
 sg13g2_nor2_1 _09229_ (.A(net2605),
    .B(\ChiselTop.wild.cpu.regs[28][15] ),
    .Y(_03890_));
 sg13g2_nor3_1 _09230_ (.A(net2581),
    .B(_03889_),
    .C(_03890_),
    .Y(_03891_));
 sg13g2_nor2b_1 _09231_ (.A(\ChiselTop.wild.cpu.regs[31][15] ),
    .B_N(net2605),
    .Y(_03892_));
 sg13g2_o21ai_1 _09232_ (.B1(net2581),
    .Y(_03893_),
    .A1(net2605),
    .A2(\ChiselTop.wild.cpu.regs[30][15] ));
 sg13g2_o21ai_1 _09233_ (.B1(net2562),
    .Y(_03894_),
    .A1(_03892_),
    .A2(_03893_));
 sg13g2_o21ai_1 _09234_ (.B1(net2462),
    .Y(_03895_),
    .A1(_03891_),
    .A2(_03894_));
 sg13g2_nor2_1 _09235_ (.A(_03888_),
    .B(_03895_),
    .Y(_03896_));
 sg13g2_nand2_1 _09236_ (.Y(_03897_),
    .A(net2117),
    .B(net2412));
 sg13g2_o21ai_1 _09237_ (.B1(_03897_),
    .Y(_03898_),
    .A1(net2412),
    .A2(_03896_));
 sg13g2_a21oi_1 _09238_ (.A1(net2160),
    .A2(_03898_),
    .Y(_03899_),
    .B1(_03791_));
 sg13g2_mux2_1 _09239_ (.A0(_03899_),
    .A1(net1491),
    .S(_03796_),
    .X(_00213_));
 sg13g2_a221oi_1 _09240_ (.B2(_00929_),
    .C1(_03571_),
    .B1(_03574_),
    .A1(\ChiselTop.wild.cpu.io_dmem_rdAddress[31] ),
    .Y(_03900_),
    .A2(_03573_));
 sg13g2_nand2_1 _09241_ (.Y(_03901_),
    .A(_03611_),
    .B(_03900_));
 sg13g2_o21ai_1 _09242_ (.B1(_03901_),
    .Y(_00214_),
    .A1(_00938_),
    .A2(_03900_));
 sg13g2_nand2_1 _09243_ (.Y(_03902_),
    .A(_03637_),
    .B(net2072));
 sg13g2_o21ai_1 _09244_ (.B1(_03902_),
    .Y(_00215_),
    .A1(_00932_),
    .A2(net2072));
 sg13g2_mux2_1 _09245_ (.A0(net1149),
    .A1(_03663_),
    .S(net2072),
    .X(_00216_));
 sg13g2_mux2_1 _09246_ (.A0(net993),
    .A1(_03677_),
    .S(net2072),
    .X(_00217_));
 sg13g2_mux2_1 _09247_ (.A0(net1112),
    .A1(_03714_),
    .S(net2072),
    .X(_00218_));
 sg13g2_mux2_1 _09248_ (.A0(net1120),
    .A1(_03739_),
    .S(net2072),
    .X(_00219_));
 sg13g2_mux2_1 _09249_ (.A0(net1242),
    .A1(_03753_),
    .S(net2072),
    .X(_00220_));
 sg13g2_mux2_1 _09250_ (.A0(net1249),
    .A1(_03790_),
    .S(net2072),
    .X(_00221_));
 sg13g2_nor2_2 _09251_ (.A(_03522_),
    .B(_03530_),
    .Y(_03903_));
 sg13g2_nor2_1 _09252_ (.A(net1382),
    .B(net2294),
    .Y(_03904_));
 sg13g2_a21oi_1 _09253_ (.A1(net2136),
    .A2(net2294),
    .Y(_00222_),
    .B1(_03904_));
 sg13g2_nor2_1 _09254_ (.A(net1377),
    .B(net2295),
    .Y(_03905_));
 sg13g2_a21oi_1 _09255_ (.A1(net2148),
    .A2(net2295),
    .Y(_00223_),
    .B1(_03905_));
 sg13g2_nor2_1 _09256_ (.A(net1380),
    .B(net2294),
    .Y(_03906_));
 sg13g2_a21oi_1 _09257_ (.A1(net2138),
    .A2(net2294),
    .Y(_00224_),
    .B1(_03906_));
 sg13g2_nor2_1 _09258_ (.A(net1285),
    .B(net2294),
    .Y(_03907_));
 sg13g2_a21oi_1 _09259_ (.A1(net2134),
    .A2(net2294),
    .Y(_00225_),
    .B1(_03907_));
 sg13g2_nor2_1 _09260_ (.A(net1296),
    .B(net2296),
    .Y(_03908_));
 sg13g2_a21oi_1 _09261_ (.A1(net2151),
    .A2(net2296),
    .Y(_00226_),
    .B1(_03908_));
 sg13g2_nor2_1 _09262_ (.A(net1315),
    .B(net2293),
    .Y(_03909_));
 sg13g2_a21oi_1 _09263_ (.A1(net2141),
    .A2(net2293),
    .Y(_00227_),
    .B1(_03909_));
 sg13g2_nor2_1 _09264_ (.A(net1335),
    .B(net2291),
    .Y(_03910_));
 sg13g2_a21oi_1 _09265_ (.A1(net2143),
    .A2(net2291),
    .Y(_00228_),
    .B1(_03910_));
 sg13g2_nor2_1 _09266_ (.A(net1281),
    .B(net2291),
    .Y(_03911_));
 sg13g2_a21oi_1 _09267_ (.A1(net2145),
    .A2(net2291),
    .Y(_00229_),
    .B1(_03911_));
 sg13g2_nor2_1 _09268_ (.A(net1344),
    .B(net2292),
    .Y(_03912_));
 sg13g2_a21oi_1 _09269_ (.A1(net2130),
    .A2(net2292),
    .Y(_00230_),
    .B1(_03912_));
 sg13g2_nor2_1 _09270_ (.A(net1282),
    .B(net2289),
    .Y(_03913_));
 sg13g2_a21oi_1 _09271_ (.A1(net2127),
    .A2(net2289),
    .Y(_00231_),
    .B1(_03913_));
 sg13g2_nor2_1 _09272_ (.A(net1339),
    .B(net2288),
    .Y(_03914_));
 sg13g2_a21oi_1 _09273_ (.A1(net2133),
    .A2(net2288),
    .Y(_00232_),
    .B1(_03914_));
 sg13g2_mux2_1 _09274_ (.A0(net1338),
    .A1(net2123),
    .S(net2291),
    .X(_00233_));
 sg13g2_nor2_1 _09275_ (.A(net1386),
    .B(net2291),
    .Y(_03915_));
 sg13g2_a21oi_1 _09276_ (.A1(net2125),
    .A2(net2291),
    .Y(_00234_),
    .B1(_03915_));
 sg13g2_nor2_1 _09277_ (.A(net1310),
    .B(net2292),
    .Y(_03916_));
 sg13g2_a21oi_1 _09278_ (.A1(net2122),
    .A2(net2292),
    .Y(_00235_),
    .B1(_03916_));
 sg13g2_nor2_1 _09279_ (.A(net1275),
    .B(net2290),
    .Y(_03917_));
 sg13g2_a21oi_1 _09280_ (.A1(net2120),
    .A2(net2290),
    .Y(_00236_),
    .B1(_03917_));
 sg13g2_nor2_1 _09281_ (.A(net1196),
    .B(net2295),
    .Y(_03918_));
 sg13g2_a21oi_1 _09282_ (.A1(net2117),
    .A2(net2295),
    .Y(_00237_),
    .B1(_03918_));
 sg13g2_nor2_1 _09283_ (.A(net1403),
    .B(net2288),
    .Y(_03919_));
 sg13g2_a21oi_1 _09284_ (.A1(net2111),
    .A2(net2288),
    .Y(_00238_),
    .B1(_03919_));
 sg13g2_nor2_1 _09285_ (.A(net1321),
    .B(net2288),
    .Y(_03920_));
 sg13g2_a21oi_1 _09286_ (.A1(net2114),
    .A2(net2288),
    .Y(_00239_),
    .B1(_03920_));
 sg13g2_nor2_1 _09287_ (.A(net1414),
    .B(net2289),
    .Y(_03921_));
 sg13g2_a21oi_1 _09288_ (.A1(net2105),
    .A2(net2289),
    .Y(_00240_),
    .B1(_03921_));
 sg13g2_nor2_1 _09289_ (.A(net1251),
    .B(net2293),
    .Y(_03922_));
 sg13g2_a21oi_1 _09290_ (.A1(net2108),
    .A2(net2293),
    .Y(_00241_),
    .B1(_03922_));
 sg13g2_nor2_1 _09291_ (.A(net1316),
    .B(net2290),
    .Y(_03923_));
 sg13g2_a21oi_1 _09292_ (.A1(net2099),
    .A2(net2290),
    .Y(_00242_),
    .B1(_03923_));
 sg13g2_nor2_1 _09293_ (.A(net1295),
    .B(net2290),
    .Y(_03924_));
 sg13g2_a21oi_1 _09294_ (.A1(net2103),
    .A2(net2290),
    .Y(_00243_),
    .B1(_03924_));
 sg13g2_nor2_1 _09295_ (.A(net1270),
    .B(net2289),
    .Y(_03925_));
 sg13g2_a21oi_1 _09296_ (.A1(net2093),
    .A2(net2289),
    .Y(_00244_),
    .B1(_03925_));
 sg13g2_nor2_1 _09297_ (.A(net1301),
    .B(net2290),
    .Y(_03926_));
 sg13g2_a21oi_1 _09298_ (.A1(net2090),
    .A2(net2290),
    .Y(_00245_),
    .B1(_03926_));
 sg13g2_nor2_1 _09299_ (.A(net1431),
    .B(net2295),
    .Y(_03927_));
 sg13g2_a21oi_1 _09300_ (.A1(net2096),
    .A2(net2293),
    .Y(_00246_),
    .B1(_03927_));
 sg13g2_nor2_1 _09301_ (.A(net1323),
    .B(net2288),
    .Y(_03928_));
 sg13g2_a21oi_1 _09302_ (.A1(net2081),
    .A2(net2288),
    .Y(_00247_),
    .B1(_03928_));
 sg13g2_nor2_1 _09303_ (.A(net1248),
    .B(net2296),
    .Y(_03929_));
 sg13g2_a21oi_1 _09304_ (.A1(net2085),
    .A2(net2296),
    .Y(_00248_),
    .B1(_03929_));
 sg13g2_nor2_1 _09305_ (.A(net1265),
    .B(net2293),
    .Y(_03930_));
 sg13g2_a21oi_1 _09306_ (.A1(net2087),
    .A2(net2293),
    .Y(_00249_),
    .B1(_03930_));
 sg13g2_nor2_1 _09307_ (.A(net1294),
    .B(net2289),
    .Y(_03931_));
 sg13g2_a21oi_1 _09308_ (.A1(net2077),
    .A2(net2289),
    .Y(_00250_),
    .B1(_03931_));
 sg13g2_nor2_1 _09309_ (.A(net1371),
    .B(net2295),
    .Y(_03932_));
 sg13g2_a21oi_1 _09310_ (.A1(net2079),
    .A2(net2295),
    .Y(_00251_),
    .B1(_03932_));
 sg13g2_nor2_1 _09311_ (.A(net1268),
    .B(net2294),
    .Y(_03933_));
 sg13g2_a21oi_1 _09312_ (.A1(net2076),
    .A2(net2293),
    .Y(_00252_),
    .B1(_03933_));
 sg13g2_nor2_1 _09313_ (.A(net1291),
    .B(net2296),
    .Y(_03934_));
 sg13g2_a21oi_1 _09314_ (.A1(net2074),
    .A2(net2295),
    .Y(_00253_),
    .B1(_03934_));
 sg13g2_nand3_1 _09315_ (.B(net2612),
    .C(_03523_),
    .A(\ChiselTop.wild.cpu.decExReg_rd[3] ),
    .Y(_03935_));
 sg13g2_nor2_1 _09316_ (.A(_03522_),
    .B(_03935_),
    .Y(_03936_));
 sg13g2_nor2_1 _09317_ (.A(net963),
    .B(net2284),
    .Y(_03937_));
 sg13g2_a21oi_1 _09318_ (.A1(net2136),
    .A2(net2284),
    .Y(_00254_),
    .B1(_03937_));
 sg13g2_nor2_1 _09319_ (.A(net1073),
    .B(net2286),
    .Y(_03938_));
 sg13g2_a21oi_1 _09320_ (.A1(net2147),
    .A2(net2286),
    .Y(_00255_),
    .B1(_03938_));
 sg13g2_nor2_1 _09321_ (.A(net1122),
    .B(net2286),
    .Y(_03939_));
 sg13g2_a21oi_1 _09322_ (.A1(net2138),
    .A2(net2286),
    .Y(_00256_),
    .B1(_03939_));
 sg13g2_nor2_1 _09323_ (.A(net1049),
    .B(net2284),
    .Y(_03940_));
 sg13g2_a21oi_1 _09324_ (.A1(net2134),
    .A2(net2284),
    .Y(_00257_),
    .B1(_03940_));
 sg13g2_nor2_1 _09325_ (.A(net962),
    .B(net2284),
    .Y(_03941_));
 sg13g2_a21oi_1 _09326_ (.A1(net2150),
    .A2(net2284),
    .Y(_00258_),
    .B1(_03941_));
 sg13g2_nor2_1 _09327_ (.A(net1224),
    .B(net2283),
    .Y(_03942_));
 sg13g2_a21oi_1 _09328_ (.A1(net2141),
    .A2(net2283),
    .Y(_00259_),
    .B1(_03942_));
 sg13g2_nor2_1 _09329_ (.A(net1137),
    .B(net2281),
    .Y(_03943_));
 sg13g2_a21oi_1 _09330_ (.A1(net2144),
    .A2(net2281),
    .Y(_00260_),
    .B1(_03943_));
 sg13g2_nor2_1 _09331_ (.A(net1115),
    .B(net2281),
    .Y(_03944_));
 sg13g2_a21oi_1 _09332_ (.A1(net2145),
    .A2(net2281),
    .Y(_00261_),
    .B1(_03944_));
 sg13g2_nor2_1 _09333_ (.A(net1217),
    .B(net2277),
    .Y(_03945_));
 sg13g2_a21oi_1 _09334_ (.A1(net2131),
    .A2(net2277),
    .Y(_00262_),
    .B1(_03945_));
 sg13g2_nor2_1 _09335_ (.A(net1037),
    .B(net2278),
    .Y(_03946_));
 sg13g2_a21oi_1 _09336_ (.A1(net2128),
    .A2(net2278),
    .Y(_00263_),
    .B1(_03946_));
 sg13g2_nor2_1 _09337_ (.A(net1011),
    .B(net2278),
    .Y(_03947_));
 sg13g2_a21oi_1 _09338_ (.A1(net2132),
    .A2(net2278),
    .Y(_00264_),
    .B1(_03947_));
 sg13g2_mux2_1 _09339_ (.A0(net1096),
    .A1(net2124),
    .S(net2280),
    .X(_00265_));
 sg13g2_nor2_1 _09340_ (.A(net1174),
    .B(net2280),
    .Y(_03948_));
 sg13g2_a21oi_1 _09341_ (.A1(net2126),
    .A2(net2280),
    .Y(_00266_),
    .B1(_03948_));
 sg13g2_nor2_1 _09342_ (.A(net1143),
    .B(net2281),
    .Y(_03949_));
 sg13g2_a21oi_1 _09343_ (.A1(net2121),
    .A2(net2281),
    .Y(_00267_),
    .B1(_03949_));
 sg13g2_nor2_1 _09344_ (.A(net1188),
    .B(net2279),
    .Y(_03950_));
 sg13g2_a21oi_1 _09345_ (.A1(net2120),
    .A2(net2279),
    .Y(_00268_),
    .B1(_03950_));
 sg13g2_nor2_1 _09346_ (.A(net1172),
    .B(net2285),
    .Y(_03951_));
 sg13g2_a21oi_1 _09347_ (.A1(net2117),
    .A2(net2285),
    .Y(_00269_),
    .B1(_03951_));
 sg13g2_nor2_1 _09348_ (.A(net1168),
    .B(net2282),
    .Y(_03952_));
 sg13g2_a21oi_1 _09349_ (.A1(net2111),
    .A2(net2282),
    .Y(_00270_),
    .B1(_03952_));
 sg13g2_nor2_1 _09350_ (.A(net1114),
    .B(net2277),
    .Y(_03953_));
 sg13g2_a21oi_1 _09351_ (.A1(net2114),
    .A2(net2277),
    .Y(_00271_),
    .B1(_03953_));
 sg13g2_nor2_1 _09352_ (.A(net1103),
    .B(net2277),
    .Y(_03954_));
 sg13g2_a21oi_1 _09353_ (.A1(net2105),
    .A2(net2277),
    .Y(_00272_),
    .B1(_03954_));
 sg13g2_nor2_1 _09354_ (.A(net1072),
    .B(net2283),
    .Y(_03955_));
 sg13g2_a21oi_1 _09355_ (.A1(net2108),
    .A2(net2283),
    .Y(_00273_),
    .B1(_03955_));
 sg13g2_nor2_1 _09356_ (.A(net1144),
    .B(net2280),
    .Y(_03956_));
 sg13g2_a21oi_1 _09357_ (.A1(net2100),
    .A2(net2279),
    .Y(_00274_),
    .B1(_03956_));
 sg13g2_nor2_1 _09358_ (.A(net1221),
    .B(net2279),
    .Y(_03957_));
 sg13g2_a21oi_1 _09359_ (.A1(net2102),
    .A2(net2279),
    .Y(_00275_),
    .B1(_03957_));
 sg13g2_nor2_1 _09360_ (.A(net956),
    .B(net2277),
    .Y(_03958_));
 sg13g2_a21oi_1 _09361_ (.A1(net2094),
    .A2(net2277),
    .Y(_00276_),
    .B1(_03958_));
 sg13g2_nor2_1 _09362_ (.A(net954),
    .B(net2279),
    .Y(_03959_));
 sg13g2_a21oi_1 _09363_ (.A1(net2091),
    .A2(net2279),
    .Y(_00277_),
    .B1(_03959_));
 sg13g2_nor2_1 _09364_ (.A(net986),
    .B(net2285),
    .Y(_03960_));
 sg13g2_a21oi_1 _09365_ (.A1(net2097),
    .A2(net2285),
    .Y(_00278_),
    .B1(_03960_));
 sg13g2_nor2_1 _09366_ (.A(net947),
    .B(net2278),
    .Y(_03961_));
 sg13g2_a21oi_1 _09367_ (.A1(net2081),
    .A2(net2278),
    .Y(_00279_),
    .B1(_03961_));
 sg13g2_nor2_1 _09368_ (.A(net1101),
    .B(net2285),
    .Y(_03962_));
 sg13g2_a21oi_1 _09369_ (.A1(net2084),
    .A2(net2285),
    .Y(_00280_),
    .B1(_03962_));
 sg13g2_nor2_1 _09370_ (.A(net1102),
    .B(net2283),
    .Y(_03963_));
 sg13g2_a21oi_1 _09371_ (.A1(net2087),
    .A2(net2283),
    .Y(_00281_),
    .B1(_03963_));
 sg13g2_nor2_1 _09372_ (.A(net1089),
    .B(net2279),
    .Y(_03964_));
 sg13g2_a21oi_1 _09373_ (.A1(net2078),
    .A2(net2278),
    .Y(_00282_),
    .B1(_03964_));
 sg13g2_nor2_1 _09374_ (.A(net1000),
    .B(net2285),
    .Y(_03965_));
 sg13g2_a21oi_1 _09375_ (.A1(net2080),
    .A2(net2285),
    .Y(_00283_),
    .B1(_03965_));
 sg13g2_nor2_1 _09376_ (.A(net1062),
    .B(net2283),
    .Y(_03966_));
 sg13g2_a21oi_1 _09377_ (.A1(net2075),
    .A2(net2283),
    .Y(_00284_),
    .B1(_03966_));
 sg13g2_nor2_1 _09378_ (.A(net1024),
    .B(net2284),
    .Y(_03967_));
 sg13g2_a21oi_1 _09379_ (.A1(net2073),
    .A2(net2284),
    .Y(_00285_),
    .B1(_03967_));
 sg13g2_nor2_1 _09380_ (.A(_03520_),
    .B(_03935_),
    .Y(_03968_));
 sg13g2_nor2_1 _09381_ (.A(net969),
    .B(net2273),
    .Y(_03969_));
 sg13g2_a21oi_1 _09382_ (.A1(net2136),
    .A2(net2273),
    .Y(_00286_),
    .B1(_03969_));
 sg13g2_nor2_1 _09383_ (.A(net975),
    .B(net2274),
    .Y(_03970_));
 sg13g2_a21oi_1 _09384_ (.A1(net2147),
    .A2(net2274),
    .Y(_00287_),
    .B1(_03970_));
 sg13g2_nor2_1 _09385_ (.A(net983),
    .B(net2275),
    .Y(_03971_));
 sg13g2_a21oi_1 _09386_ (.A1(net2138),
    .A2(net2275),
    .Y(_00288_),
    .B1(_03971_));
 sg13g2_nor2_1 _09387_ (.A(net1068),
    .B(net2273),
    .Y(_03972_));
 sg13g2_a21oi_1 _09388_ (.A1(net2135),
    .A2(net2273),
    .Y(_00289_),
    .B1(_03972_));
 sg13g2_nor2_1 _09389_ (.A(net1074),
    .B(net2275),
    .Y(_03973_));
 sg13g2_a21oi_1 _09390_ (.A1(net2150),
    .A2(net2275),
    .Y(_00290_),
    .B1(_03973_));
 sg13g2_nor2_1 _09391_ (.A(net959),
    .B(net2272),
    .Y(_03974_));
 sg13g2_a21oi_1 _09392_ (.A1(net2141),
    .A2(net2272),
    .Y(_00291_),
    .B1(_03974_));
 sg13g2_nor2_1 _09393_ (.A(net1018),
    .B(net2271),
    .Y(_03975_));
 sg13g2_a21oi_1 _09394_ (.A1(net2144),
    .A2(net2271),
    .Y(_00292_),
    .B1(_03975_));
 sg13g2_nor2_1 _09395_ (.A(net974),
    .B(net2270),
    .Y(_03976_));
 sg13g2_a21oi_1 _09396_ (.A1(net2145),
    .A2(net2270),
    .Y(_00293_),
    .B1(_03976_));
 sg13g2_nor2_1 _09397_ (.A(net1147),
    .B(net2266),
    .Y(_03977_));
 sg13g2_a21oi_1 _09398_ (.A1(net2130),
    .A2(net2266),
    .Y(_00294_),
    .B1(_03977_));
 sg13g2_nor2_1 _09399_ (.A(net1039),
    .B(net2267),
    .Y(_03978_));
 sg13g2_a21oi_1 _09400_ (.A1(net2128),
    .A2(net2267),
    .Y(_00295_),
    .B1(_03978_));
 sg13g2_nor2_1 _09401_ (.A(net943),
    .B(net2273),
    .Y(_03979_));
 sg13g2_a21oi_1 _09402_ (.A1(net2132),
    .A2(net2273),
    .Y(_00296_),
    .B1(_03979_));
 sg13g2_mux2_1 _09403_ (.A0(net1053),
    .A1(net2124),
    .S(net2270),
    .X(_00297_));
 sg13g2_nor2_1 _09404_ (.A(net976),
    .B(net2270),
    .Y(_03980_));
 sg13g2_a21oi_1 _09405_ (.A1(net2125),
    .A2(net2270),
    .Y(_00298_),
    .B1(_03980_));
 sg13g2_nor2_1 _09406_ (.A(net1311),
    .B(net2271),
    .Y(_03981_));
 sg13g2_a21oi_1 _09407_ (.A1(net2121),
    .A2(net2271),
    .Y(_00299_),
    .B1(_03981_));
 sg13g2_nor2_1 _09408_ (.A(net951),
    .B(net2269),
    .Y(_03982_));
 sg13g2_a21oi_1 _09409_ (.A1(net2119),
    .A2(net2269),
    .Y(_00300_),
    .B1(_03982_));
 sg13g2_nor2_1 _09410_ (.A(net1292),
    .B(net2270),
    .Y(_03983_));
 sg13g2_a21oi_1 _09411_ (.A1(net2117),
    .A2(net2270),
    .Y(_00301_),
    .B1(_03983_));
 sg13g2_nor2_1 _09412_ (.A(net1166),
    .B(net2268),
    .Y(_03984_));
 sg13g2_a21oi_1 _09413_ (.A1(net2111),
    .A2(net2268),
    .Y(_00302_),
    .B1(_03984_));
 sg13g2_nor2_1 _09414_ (.A(net1045),
    .B(net2266),
    .Y(_03985_));
 sg13g2_a21oi_1 _09415_ (.A1(net2114),
    .A2(net2266),
    .Y(_00303_),
    .B1(_03985_));
 sg13g2_nor2_1 _09416_ (.A(net1153),
    .B(net2266),
    .Y(_03986_));
 sg13g2_a21oi_1 _09417_ (.A1(net2105),
    .A2(net2266),
    .Y(_00304_),
    .B1(_03986_));
 sg13g2_nor2_1 _09418_ (.A(net1129),
    .B(net2272),
    .Y(_03987_));
 sg13g2_a21oi_1 _09419_ (.A1(net2108),
    .A2(net2272),
    .Y(_00305_),
    .B1(_03987_));
 sg13g2_nor2_1 _09420_ (.A(net1031),
    .B(net2269),
    .Y(_03988_));
 sg13g2_a21oi_1 _09421_ (.A1(net2100),
    .A2(net2269),
    .Y(_00306_),
    .B1(_03988_));
 sg13g2_nor2_1 _09422_ (.A(net957),
    .B(net2269),
    .Y(_03989_));
 sg13g2_a21oi_1 _09423_ (.A1(net2102),
    .A2(net2269),
    .Y(_00307_),
    .B1(_03989_));
 sg13g2_nor2_1 _09424_ (.A(net1354),
    .B(net2266),
    .Y(_03990_));
 sg13g2_a21oi_1 _09425_ (.A1(net2093),
    .A2(net2266),
    .Y(_00308_),
    .B1(_03990_));
 sg13g2_nor2_1 _09426_ (.A(net1171),
    .B(net2269),
    .Y(_03991_));
 sg13g2_a21oi_1 _09427_ (.A1(net2091),
    .A2(net2269),
    .Y(_00309_),
    .B1(_03991_));
 sg13g2_nor2_1 _09428_ (.A(net949),
    .B(net2274),
    .Y(_03992_));
 sg13g2_a21oi_1 _09429_ (.A1(net2097),
    .A2(net2274),
    .Y(_00310_),
    .B1(_03992_));
 sg13g2_nor2_1 _09430_ (.A(net1016),
    .B(net2268),
    .Y(_03993_));
 sg13g2_a21oi_1 _09431_ (.A1(net2081),
    .A2(net2268),
    .Y(_00311_),
    .B1(_03993_));
 sg13g2_nor2_1 _09432_ (.A(net1216),
    .B(net2274),
    .Y(_03994_));
 sg13g2_a21oi_1 _09433_ (.A1(net2084),
    .A2(net2274),
    .Y(_00312_),
    .B1(_03994_));
 sg13g2_nor2_1 _09434_ (.A(net978),
    .B(net2272),
    .Y(_03995_));
 sg13g2_a21oi_1 _09435_ (.A1(net2087),
    .A2(net2272),
    .Y(_00313_),
    .B1(_03995_));
 sg13g2_nor2_1 _09436_ (.A(net1232),
    .B(net2267),
    .Y(_03996_));
 sg13g2_a21oi_1 _09437_ (.A1(net2078),
    .A2(net2267),
    .Y(_00314_),
    .B1(_03996_));
 sg13g2_nor2_1 _09438_ (.A(net999),
    .B(net2274),
    .Y(_03997_));
 sg13g2_a21oi_1 _09439_ (.A1(net2079),
    .A2(net2274),
    .Y(_00315_),
    .B1(_03997_));
 sg13g2_nor2_1 _09440_ (.A(net1056),
    .B(net2272),
    .Y(_03998_));
 sg13g2_a21oi_1 _09441_ (.A1(net2075),
    .A2(net2272),
    .Y(_00316_),
    .B1(_03998_));
 sg13g2_nor2_1 _09442_ (.A(net979),
    .B(net2275),
    .Y(_03999_));
 sg13g2_a21oi_1 _09443_ (.A1(net2073),
    .A2(net2273),
    .Y(_00317_),
    .B1(_03999_));
 sg13g2_nor2_1 _09444_ (.A(_03524_),
    .B(_03935_),
    .Y(_04000_));
 sg13g2_nor2_1 _09445_ (.A(net1009),
    .B(net2257),
    .Y(_04001_));
 sg13g2_a21oi_1 _09446_ (.A1(net2136),
    .A2(net2257),
    .Y(_00318_),
    .B1(_04001_));
 sg13g2_nor2_1 _09447_ (.A(net1213),
    .B(net2264),
    .Y(_04002_));
 sg13g2_a21oi_1 _09448_ (.A1(net2147),
    .A2(net2263),
    .Y(_00319_),
    .B1(_04002_));
 sg13g2_nor2_1 _09449_ (.A(net1027),
    .B(net2263),
    .Y(_04003_));
 sg13g2_a21oi_1 _09450_ (.A1(net2138),
    .A2(net2263),
    .Y(_00320_),
    .B1(_04003_));
 sg13g2_nor2_1 _09451_ (.A(net1041),
    .B(net2257),
    .Y(_04004_));
 sg13g2_a21oi_1 _09452_ (.A1(net2134),
    .A2(net2257),
    .Y(_00321_),
    .B1(_04004_));
 sg13g2_nor2_1 _09453_ (.A(net1257),
    .B(net2258),
    .Y(_04005_));
 sg13g2_a21oi_1 _09454_ (.A1(net2150),
    .A2(net2258),
    .Y(_00322_),
    .B1(_04005_));
 sg13g2_nor2_1 _09455_ (.A(net1181),
    .B(net2258),
    .Y(_04006_));
 sg13g2_a21oi_1 _09456_ (.A1(net2141),
    .A2(net2258),
    .Y(_00323_),
    .B1(_04006_));
 sg13g2_nor2_1 _09457_ (.A(net1029),
    .B(net2262),
    .Y(_04007_));
 sg13g2_a21oi_1 _09458_ (.A1(net2144),
    .A2(net2262),
    .Y(_00324_),
    .B1(_04007_));
 sg13g2_nor2_1 _09459_ (.A(net1148),
    .B(net2260),
    .Y(_04008_));
 sg13g2_a21oi_1 _09460_ (.A1(net2145),
    .A2(net2260),
    .Y(_00325_),
    .B1(_04008_));
 sg13g2_nor2_1 _09461_ (.A(net1252),
    .B(net2256),
    .Y(_04009_));
 sg13g2_a21oi_1 _09462_ (.A1(net2131),
    .A2(net2256),
    .Y(_00326_),
    .B1(_04009_));
 sg13g2_nor2_1 _09463_ (.A(net987),
    .B(net2256),
    .Y(_04010_));
 sg13g2_a21oi_1 _09464_ (.A1(net2128),
    .A2(net2256),
    .Y(_00327_),
    .B1(_04010_));
 sg13g2_nor2_1 _09465_ (.A(net1035),
    .B(net2256),
    .Y(_04011_));
 sg13g2_a21oi_1 _09466_ (.A1(net2132),
    .A2(net2256),
    .Y(_00328_),
    .B1(_04011_));
 sg13g2_mux2_1 _09467_ (.A0(net1158),
    .A1(net2124),
    .S(net2261),
    .X(_00329_));
 sg13g2_nor2_1 _09468_ (.A(net1020),
    .B(net2261),
    .Y(_04012_));
 sg13g2_a21oi_1 _09469_ (.A1(net2126),
    .A2(net2261),
    .Y(_00330_),
    .B1(_04012_));
 sg13g2_nor2_1 _09470_ (.A(net1110),
    .B(net2262),
    .Y(_04013_));
 sg13g2_a21oi_1 _09471_ (.A1(net2121),
    .A2(net2260),
    .Y(_00331_),
    .B1(_04013_));
 sg13g2_nor2_1 _09472_ (.A(net1026),
    .B(net2260),
    .Y(_04014_));
 sg13g2_a21oi_1 _09473_ (.A1(net2119),
    .A2(net2260),
    .Y(_00332_),
    .B1(_04014_));
 sg13g2_nor2_1 _09474_ (.A(net1141),
    .B(net2264),
    .Y(_04015_));
 sg13g2_a21oi_1 _09475_ (.A1(net2117),
    .A2(net2263),
    .Y(_00333_),
    .B1(_04015_));
 sg13g2_nor2_1 _09476_ (.A(net988),
    .B(net2256),
    .Y(_04016_));
 sg13g2_a21oi_1 _09477_ (.A1(net2111),
    .A2(net2255),
    .Y(_00334_),
    .B1(_04016_));
 sg13g2_nor2_1 _09478_ (.A(net1255),
    .B(net2255),
    .Y(_04017_));
 sg13g2_a21oi_1 _09479_ (.A1(net2114),
    .A2(net2255),
    .Y(_00335_),
    .B1(_04017_));
 sg13g2_nor2_1 _09480_ (.A(net1208),
    .B(net2255),
    .Y(_04018_));
 sg13g2_a21oi_1 _09481_ (.A1(net2105),
    .A2(net2255),
    .Y(_00336_),
    .B1(_04018_));
 sg13g2_nor2_1 _09482_ (.A(net1132),
    .B(net2257),
    .Y(_04019_));
 sg13g2_a21oi_1 _09483_ (.A1(net2108),
    .A2(net2257),
    .Y(_00337_),
    .B1(_04019_));
 sg13g2_nor2_1 _09484_ (.A(net1193),
    .B(net2261),
    .Y(_04020_));
 sg13g2_a21oi_1 _09485_ (.A1(net2100),
    .A2(net2261),
    .Y(_00338_),
    .B1(_04020_));
 sg13g2_nor2_1 _09486_ (.A(net1283),
    .B(net2261),
    .Y(_04021_));
 sg13g2_a21oi_1 _09487_ (.A1(net2102),
    .A2(net2261),
    .Y(_00339_),
    .B1(_04021_));
 sg13g2_nor2_1 _09488_ (.A(net1157),
    .B(net2259),
    .Y(_04022_));
 sg13g2_a21oi_1 _09489_ (.A1(net2094),
    .A2(net2255),
    .Y(_00340_),
    .B1(_04022_));
 sg13g2_nor2_1 _09490_ (.A(net1195),
    .B(net2261),
    .Y(_04023_));
 sg13g2_a21oi_1 _09491_ (.A1(net2092),
    .A2(net2260),
    .Y(_00341_),
    .B1(_04023_));
 sg13g2_nor2_1 _09492_ (.A(net1085),
    .B(net2263),
    .Y(_04024_));
 sg13g2_a21oi_1 _09493_ (.A1(net2097),
    .A2(net2263),
    .Y(_00342_),
    .B1(_04024_));
 sg13g2_nor2_1 _09494_ (.A(net1021),
    .B(net2255),
    .Y(_04025_));
 sg13g2_a21oi_1 _09495_ (.A1(net2081),
    .A2(net2255),
    .Y(_00343_),
    .B1(_04025_));
 sg13g2_nor2_1 _09496_ (.A(net1123),
    .B(net2264),
    .Y(_04026_));
 sg13g2_a21oi_1 _09497_ (.A1(net2084),
    .A2(net2264),
    .Y(_00344_),
    .B1(_04026_));
 sg13g2_nor2_1 _09498_ (.A(net1146),
    .B(net2257),
    .Y(_04027_));
 sg13g2_a21oi_1 _09499_ (.A1(net2087),
    .A2(net2257),
    .Y(_00345_),
    .B1(_04027_));
 sg13g2_nor2_1 _09500_ (.A(net1218),
    .B(net2260),
    .Y(_04028_));
 sg13g2_a21oi_1 _09501_ (.A1(net2078),
    .A2(net2260),
    .Y(_00346_),
    .B1(_04028_));
 sg13g2_nor2_1 _09502_ (.A(net1194),
    .B(net2263),
    .Y(_04029_));
 sg13g2_a21oi_1 _09503_ (.A1(net2080),
    .A2(net2263),
    .Y(_00347_),
    .B1(_04029_));
 sg13g2_nor2_1 _09504_ (.A(net1206),
    .B(net2258),
    .Y(_04030_));
 sg13g2_a21oi_1 _09505_ (.A1(net2076),
    .A2(net2258),
    .Y(_00348_),
    .B1(_04030_));
 sg13g2_nor2_1 _09506_ (.A(net1228),
    .B(net2258),
    .Y(_04031_));
 sg13g2_a21oi_1 _09507_ (.A1(net2073),
    .A2(net2258),
    .Y(_00349_),
    .B1(_04031_));
 sg13g2_nand2_2 _09508_ (.Y(_04032_),
    .A(_00967_),
    .B(_03523_));
 sg13g2_nor3_1 _09509_ (.A(net2648),
    .B(net2649),
    .C(_04032_),
    .Y(_04033_));
 sg13g2_nor2_1 _09510_ (.A(net968),
    .B(net2248),
    .Y(_04034_));
 sg13g2_a21oi_1 _09511_ (.A1(net2137),
    .A2(net2248),
    .Y(_00350_),
    .B1(_04034_));
 sg13g2_nor2_1 _09512_ (.A(net1317),
    .B(net2251),
    .Y(_04035_));
 sg13g2_a21oi_1 _09513_ (.A1(net2148),
    .A2(net2251),
    .Y(_00351_),
    .B1(_04035_));
 sg13g2_nor2_1 _09514_ (.A(net982),
    .B(net2249),
    .Y(_04036_));
 sg13g2_a21oi_1 _09515_ (.A1(net2139),
    .A2(net2248),
    .Y(_00352_),
    .B1(_04036_));
 sg13g2_nor2_1 _09516_ (.A(net973),
    .B(net2248),
    .Y(_04037_));
 sg13g2_a21oi_1 _09517_ (.A1(net2135),
    .A2(net2248),
    .Y(_00353_),
    .B1(_04037_));
 sg13g2_nor2_1 _09518_ (.A(net991),
    .B(net2248),
    .Y(_04038_));
 sg13g2_a21oi_1 _09519_ (.A1(net2150),
    .A2(net2248),
    .Y(_00354_),
    .B1(_04038_));
 sg13g2_nor2_1 _09520_ (.A(net1184),
    .B(net2250),
    .Y(_04039_));
 sg13g2_a21oi_1 _09521_ (.A1(net2142),
    .A2(net2250),
    .Y(_00355_),
    .B1(_04039_));
 sg13g2_nor2_1 _09522_ (.A(net1116),
    .B(net2247),
    .Y(_04040_));
 sg13g2_a21oi_1 _09523_ (.A1(net2143),
    .A2(net2247),
    .Y(_00356_),
    .B1(_04040_));
 sg13g2_nor2_1 _09524_ (.A(net1134),
    .B(net2247),
    .Y(_04041_));
 sg13g2_a21oi_1 _09525_ (.A1(net2146),
    .A2(net2247),
    .Y(_00357_),
    .B1(_04041_));
 sg13g2_nor2_1 _09526_ (.A(net1012),
    .B(net2245),
    .Y(_04042_));
 sg13g2_a21oi_1 _09527_ (.A1(net2130),
    .A2(net2245),
    .Y(_00358_),
    .B1(_04042_));
 sg13g2_nor2_1 _09528_ (.A(net996),
    .B(net2244),
    .Y(_04043_));
 sg13g2_a21oi_1 _09529_ (.A1(net2127),
    .A2(net2244),
    .Y(_00359_),
    .B1(_04043_));
 sg13g2_nor2_1 _09530_ (.A(net1142),
    .B(net2250),
    .Y(_04044_));
 sg13g2_a21oi_1 _09531_ (.A1(net2132),
    .A2(net2250),
    .Y(_00360_),
    .B1(_04044_));
 sg13g2_mux2_1 _09532_ (.A0(net1151),
    .A1(net2123),
    .S(net2247),
    .X(_00361_));
 sg13g2_nor2_1 _09533_ (.A(net1182),
    .B(net2247),
    .Y(_04045_));
 sg13g2_a21oi_1 _09534_ (.A1(net2125),
    .A2(net2247),
    .Y(_00362_),
    .B1(_04045_));
 sg13g2_nor2_1 _09535_ (.A(net1010),
    .B(net2251),
    .Y(_04046_));
 sg13g2_a21oi_1 _09536_ (.A1(net2121),
    .A2(net2251),
    .Y(_00363_),
    .B1(_04046_));
 sg13g2_nor2_1 _09537_ (.A(net1048),
    .B(net2246),
    .Y(_04047_));
 sg13g2_a21oi_1 _09538_ (.A1(net2119),
    .A2(net2246),
    .Y(_00364_),
    .B1(_04047_));
 sg13g2_nor2_1 _09539_ (.A(net1052),
    .B(net2251),
    .Y(_04048_));
 sg13g2_a21oi_1 _09540_ (.A1(net2118),
    .A2(net2251),
    .Y(_00365_),
    .B1(_04048_));
 sg13g2_nor2_1 _09541_ (.A(net1007),
    .B(net2245),
    .Y(_04049_));
 sg13g2_a21oi_1 _09542_ (.A1(net2111),
    .A2(net2245),
    .Y(_00366_),
    .B1(_04049_));
 sg13g2_nor2_1 _09543_ (.A(net1040),
    .B(net2245),
    .Y(_04050_));
 sg13g2_a21oi_1 _09544_ (.A1(net2115),
    .A2(net2245),
    .Y(_00367_),
    .B1(_04050_));
 sg13g2_nor2_1 _09545_ (.A(net1004),
    .B(net2244),
    .Y(_04051_));
 sg13g2_a21oi_1 _09546_ (.A1(net2106),
    .A2(net2244),
    .Y(_00368_),
    .B1(_04051_));
 sg13g2_nor2_1 _09547_ (.A(net1075),
    .B(net2250),
    .Y(_04052_));
 sg13g2_a21oi_1 _09548_ (.A1(net2109),
    .A2(net2250),
    .Y(_00369_),
    .B1(_04052_));
 sg13g2_nor2_1 _09549_ (.A(net1240),
    .B(net2246),
    .Y(_04053_));
 sg13g2_a21oi_1 _09550_ (.A1(net2099),
    .A2(net2246),
    .Y(_00370_),
    .B1(_04053_));
 sg13g2_nor2_1 _09551_ (.A(net1033),
    .B(net2246),
    .Y(_04054_));
 sg13g2_a21oi_1 _09552_ (.A1(net2102),
    .A2(net2246),
    .Y(_00371_),
    .B1(_04054_));
 sg13g2_nor2_1 _09553_ (.A(net1086),
    .B(net2244),
    .Y(_04055_));
 sg13g2_a21oi_1 _09554_ (.A1(net2093),
    .A2(net2244),
    .Y(_00372_),
    .B1(_04055_));
 sg13g2_nor2_1 _09555_ (.A(net1028),
    .B(net2246),
    .Y(_04056_));
 sg13g2_a21oi_1 _09556_ (.A1(net2090),
    .A2(net2246),
    .Y(_00373_),
    .B1(_04056_));
 sg13g2_nor2_1 _09557_ (.A(net1083),
    .B(net2252),
    .Y(_04057_));
 sg13g2_a21oi_1 _09558_ (.A1(net2097),
    .A2(net2252),
    .Y(_00374_),
    .B1(_04057_));
 sg13g2_nor2_1 _09559_ (.A(net1210),
    .B(net2245),
    .Y(_04058_));
 sg13g2_a21oi_1 _09560_ (.A1(net2081),
    .A2(net2245),
    .Y(_00375_),
    .B1(_04058_));
 sg13g2_nor2_1 _09561_ (.A(net1006),
    .B(net2252),
    .Y(_04059_));
 sg13g2_a21oi_1 _09562_ (.A1(net2085),
    .A2(net2252),
    .Y(_00376_),
    .B1(_04059_));
 sg13g2_nor2_1 _09563_ (.A(net1118),
    .B(net2250),
    .Y(_04060_));
 sg13g2_a21oi_1 _09564_ (.A1(net2088),
    .A2(net2250),
    .Y(_00377_),
    .B1(_04060_));
 sg13g2_nor2_1 _09565_ (.A(net1200),
    .B(net2244),
    .Y(_04061_));
 sg13g2_a21oi_1 _09566_ (.A1(net2077),
    .A2(net2244),
    .Y(_00378_),
    .B1(_04061_));
 sg13g2_nor2_1 _09567_ (.A(net1302),
    .B(net2251),
    .Y(_04062_));
 sg13g2_a21oi_1 _09568_ (.A1(net2079),
    .A2(net2251),
    .Y(_00379_),
    .B1(_04062_));
 sg13g2_nor2_1 _09569_ (.A(net1237),
    .B(net2249),
    .Y(_04063_));
 sg13g2_a21oi_1 _09570_ (.A1(net2075),
    .A2(net2249),
    .Y(_00380_),
    .B1(_04063_));
 sg13g2_nor2_1 _09571_ (.A(net1192),
    .B(net2249),
    .Y(_04064_));
 sg13g2_a21oi_1 _09572_ (.A1(net2073),
    .A2(net2248),
    .Y(_00381_),
    .B1(_04064_));
 sg13g2_nor2_2 _09573_ (.A(_03524_),
    .B(_03530_),
    .Y(_04065_));
 sg13g2_nor2_1 _09574_ (.A(net1306),
    .B(net2240),
    .Y(_04066_));
 sg13g2_a21oi_1 _09575_ (.A1(net2136),
    .A2(net2240),
    .Y(_00382_),
    .B1(_04066_));
 sg13g2_nor2_1 _09576_ (.A(net1238),
    .B(net2241),
    .Y(_04067_));
 sg13g2_a21oi_1 _09577_ (.A1(net2147),
    .A2(net2241),
    .Y(_00383_),
    .B1(_04067_));
 sg13g2_nor2_1 _09578_ (.A(net1336),
    .B(net2240),
    .Y(_04068_));
 sg13g2_a21oi_1 _09579_ (.A1(net2138),
    .A2(net2240),
    .Y(_00384_),
    .B1(_04068_));
 sg13g2_nor2_1 _09580_ (.A(net1340),
    .B(net2240),
    .Y(_04069_));
 sg13g2_a21oi_1 _09581_ (.A1(net2134),
    .A2(net2240),
    .Y(_00385_),
    .B1(_04069_));
 sg13g2_nor2_1 _09582_ (.A(net1378),
    .B(net2240),
    .Y(_04070_));
 sg13g2_a21oi_1 _09583_ (.A1(net2151),
    .A2(net2240),
    .Y(_00386_),
    .B1(_04070_));
 sg13g2_nor2_1 _09584_ (.A(net1300),
    .B(net2239),
    .Y(_04071_));
 sg13g2_a21oi_1 _09585_ (.A1(net2141),
    .A2(net2239),
    .Y(_00387_),
    .B1(_04071_));
 sg13g2_nor2_1 _09586_ (.A(net1314),
    .B(net2237),
    .Y(_04072_));
 sg13g2_a21oi_1 _09587_ (.A1(net2143),
    .A2(net2237),
    .Y(_00388_),
    .B1(_04072_));
 sg13g2_nor2_1 _09588_ (.A(net1350),
    .B(net2237),
    .Y(_04073_));
 sg13g2_a21oi_1 _09589_ (.A1(net2146),
    .A2(net2237),
    .Y(_00389_),
    .B1(_04073_));
 sg13g2_nor2_1 _09590_ (.A(net1197),
    .B(net2238),
    .Y(_04074_));
 sg13g2_a21oi_1 _09591_ (.A1(net2130),
    .A2(net2238),
    .Y(_00390_),
    .B1(_04074_));
 sg13g2_nor2_1 _09592_ (.A(net1370),
    .B(net2235),
    .Y(_04075_));
 sg13g2_a21oi_1 _09593_ (.A1(net2127),
    .A2(net2235),
    .Y(_00391_),
    .B1(_04075_));
 sg13g2_nor2_1 _09594_ (.A(net1313),
    .B(net2234),
    .Y(_04076_));
 sg13g2_a21oi_1 _09595_ (.A1(net2133),
    .A2(net2234),
    .Y(_00392_),
    .B1(_04076_));
 sg13g2_mux2_1 _09596_ (.A0(net1366),
    .A1(net2123),
    .S(net2237),
    .X(_00393_));
 sg13g2_nor2_1 _09597_ (.A(net1299),
    .B(net2237),
    .Y(_04077_));
 sg13g2_a21oi_1 _09598_ (.A1(net2126),
    .A2(net2237),
    .Y(_00394_),
    .B1(_04077_));
 sg13g2_nor2_1 _09599_ (.A(net1280),
    .B(net2238),
    .Y(_04078_));
 sg13g2_a21oi_1 _09600_ (.A1(net2122),
    .A2(net2238),
    .Y(_00395_),
    .B1(_04078_));
 sg13g2_nor2_1 _09601_ (.A(net1298),
    .B(net2236),
    .Y(_04079_));
 sg13g2_a21oi_1 _09602_ (.A1(net2119),
    .A2(net2236),
    .Y(_00396_),
    .B1(_04079_));
 sg13g2_nor2_1 _09603_ (.A(net1320),
    .B(net2241),
    .Y(_04080_));
 sg13g2_a21oi_1 _09604_ (.A1(net2117),
    .A2(net2241),
    .Y(_00397_),
    .B1(_04080_));
 sg13g2_nor2_1 _09605_ (.A(net1272),
    .B(net2234),
    .Y(_04081_));
 sg13g2_a21oi_1 _09606_ (.A1(net2111),
    .A2(net2234),
    .Y(_00398_),
    .B1(_04081_));
 sg13g2_nor2_1 _09607_ (.A(net1327),
    .B(net2234),
    .Y(_04082_));
 sg13g2_a21oi_1 _09608_ (.A1(net2114),
    .A2(net2234),
    .Y(_00399_),
    .B1(_04082_));
 sg13g2_nor2_1 _09609_ (.A(net1262),
    .B(net2235),
    .Y(_04083_));
 sg13g2_a21oi_1 _09610_ (.A1(net2105),
    .A2(net2235),
    .Y(_00400_),
    .B1(_04083_));
 sg13g2_nor2_1 _09611_ (.A(net1352),
    .B(net2239),
    .Y(_04084_));
 sg13g2_a21oi_1 _09612_ (.A1(net2108),
    .A2(net2239),
    .Y(_00401_),
    .B1(_04084_));
 sg13g2_nor2_1 _09613_ (.A(net1258),
    .B(net2236),
    .Y(_04085_));
 sg13g2_a21oi_1 _09614_ (.A1(net2099),
    .A2(net2236),
    .Y(_00402_),
    .B1(_04085_));
 sg13g2_nor2_1 _09615_ (.A(net1289),
    .B(net2236),
    .Y(_04086_));
 sg13g2_a21oi_1 _09616_ (.A1(net2103),
    .A2(net2236),
    .Y(_00403_),
    .B1(_04086_));
 sg13g2_nor2_1 _09617_ (.A(net1229),
    .B(net2235),
    .Y(_04087_));
 sg13g2_a21oi_1 _09618_ (.A1(net2094),
    .A2(net2235),
    .Y(_00404_),
    .B1(_04087_));
 sg13g2_nor2_1 _09619_ (.A(net1333),
    .B(net2236),
    .Y(_04088_));
 sg13g2_a21oi_1 _09620_ (.A1(net2090),
    .A2(net2236),
    .Y(_00405_),
    .B1(_04088_));
 sg13g2_nor2_1 _09621_ (.A(net1271),
    .B(net2241),
    .Y(_04089_));
 sg13g2_a21oi_1 _09622_ (.A1(net2096),
    .A2(net2241),
    .Y(_00406_),
    .B1(_04089_));
 sg13g2_nor2_1 _09623_ (.A(net1190),
    .B(net2234),
    .Y(_04090_));
 sg13g2_a21oi_1 _09624_ (.A1(net2082),
    .A2(net2234),
    .Y(_00407_),
    .B1(_04090_));
 sg13g2_nor2_1 _09625_ (.A(net1376),
    .B(net2242),
    .Y(_04091_));
 sg13g2_a21oi_1 _09626_ (.A1(net2084),
    .A2(net2242),
    .Y(_00408_),
    .B1(_04091_));
 sg13g2_nor2_1 _09627_ (.A(net1293),
    .B(net2239),
    .Y(_04092_));
 sg13g2_a21oi_1 _09628_ (.A1(net2087),
    .A2(net2239),
    .Y(_00409_),
    .B1(_04092_));
 sg13g2_nor2_1 _09629_ (.A(net1254),
    .B(net2235),
    .Y(_04093_));
 sg13g2_a21oi_1 _09630_ (.A1(net2077),
    .A2(net2235),
    .Y(_00410_),
    .B1(_04093_));
 sg13g2_nor2_1 _09631_ (.A(net1241),
    .B(net2242),
    .Y(_04094_));
 sg13g2_a21oi_1 _09632_ (.A1(net2079),
    .A2(net2242),
    .Y(_00411_),
    .B1(_04094_));
 sg13g2_nor2_1 _09633_ (.A(net1286),
    .B(net2239),
    .Y(_04095_));
 sg13g2_a21oi_1 _09634_ (.A1(net2075),
    .A2(net2239),
    .Y(_00412_),
    .B1(_04095_));
 sg13g2_nor2_1 _09635_ (.A(net1266),
    .B(net2241),
    .Y(_04096_));
 sg13g2_a21oi_1 _09636_ (.A1(net2074),
    .A2(net2241),
    .Y(_00413_),
    .B1(_04096_));
 sg13g2_nor3_1 _09637_ (.A(net2648),
    .B(net2649),
    .C(_03935_),
    .Y(_04097_));
 sg13g2_nor2_1 _09638_ (.A(net970),
    .B(net2230),
    .Y(_04098_));
 sg13g2_a21oi_1 _09639_ (.A1(net2136),
    .A2(net2230),
    .Y(_00414_),
    .B1(_04098_));
 sg13g2_nor2_1 _09640_ (.A(net989),
    .B(net2231),
    .Y(_04099_));
 sg13g2_a21oi_1 _09641_ (.A1(net2147),
    .A2(net2231),
    .Y(_00415_),
    .B1(_04099_));
 sg13g2_nor2_1 _09642_ (.A(net1180),
    .B(net2232),
    .Y(_04100_));
 sg13g2_a21oi_1 _09643_ (.A1(net2138),
    .A2(net2232),
    .Y(_00416_),
    .B1(_04100_));
 sg13g2_nor2_1 _09644_ (.A(net1191),
    .B(net2230),
    .Y(_04101_));
 sg13g2_a21oi_1 _09645_ (.A1(net2134),
    .A2(net2230),
    .Y(_00417_),
    .B1(_04101_));
 sg13g2_nor2_1 _09646_ (.A(net944),
    .B(net2230),
    .Y(_04102_));
 sg13g2_a21oi_1 _09647_ (.A1(net2150),
    .A2(net2230),
    .Y(_00418_),
    .B1(_04102_));
 sg13g2_nor2_1 _09648_ (.A(net1017),
    .B(net2229),
    .Y(_04103_));
 sg13g2_a21oi_1 _09649_ (.A1(net2141),
    .A2(net2229),
    .Y(_00419_),
    .B1(_04103_));
 sg13g2_nor2_1 _09650_ (.A(net1152),
    .B(net2228),
    .Y(_04104_));
 sg13g2_a21oi_1 _09651_ (.A1(net2144),
    .A2(net2228),
    .Y(_00420_),
    .B1(_04104_));
 sg13g2_nor2_1 _09652_ (.A(net1066),
    .B(net2227),
    .Y(_04105_));
 sg13g2_a21oi_1 _09653_ (.A1(net2145),
    .A2(net2227),
    .Y(_00421_),
    .B1(_04105_));
 sg13g2_nor2_1 _09654_ (.A(net1135),
    .B(net2223),
    .Y(_04106_));
 sg13g2_a21oi_1 _09655_ (.A1(net2130),
    .A2(net2223),
    .Y(_00422_),
    .B1(_04106_));
 sg13g2_nor2_1 _09656_ (.A(net1051),
    .B(net2224),
    .Y(_04107_));
 sg13g2_a21oi_1 _09657_ (.A1(net2127),
    .A2(net2224),
    .Y(_00423_),
    .B1(_04107_));
 sg13g2_nor2_1 _09658_ (.A(net985),
    .B(net2225),
    .Y(_04108_));
 sg13g2_a21oi_1 _09659_ (.A1(net2132),
    .A2(net2225),
    .Y(_00424_),
    .B1(_04108_));
 sg13g2_mux2_1 _09660_ (.A0(net1117),
    .A1(net2123),
    .S(net2227),
    .X(_00425_));
 sg13g2_nor2_1 _09661_ (.A(net1179),
    .B(net2227),
    .Y(_04109_));
 sg13g2_a21oi_1 _09662_ (.A1(net2126),
    .A2(net2227),
    .Y(_00426_),
    .B1(_04109_));
 sg13g2_nor2_1 _09663_ (.A(net1109),
    .B(net2228),
    .Y(_04110_));
 sg13g2_a21oi_1 _09664_ (.A1(net2121),
    .A2(net2228),
    .Y(_00427_),
    .B1(_04110_));
 sg13g2_nor2_1 _09665_ (.A(net1055),
    .B(net2226),
    .Y(_04111_));
 sg13g2_a21oi_1 _09666_ (.A1(net2119),
    .A2(net2226),
    .Y(_00428_),
    .B1(_04111_));
 sg13g2_nor2_1 _09667_ (.A(net1297),
    .B(net2227),
    .Y(_04112_));
 sg13g2_a21oi_1 _09668_ (.A1(net2117),
    .A2(net2227),
    .Y(_00429_),
    .B1(_04112_));
 sg13g2_nor2_1 _09669_ (.A(net1244),
    .B(net2225),
    .Y(_04113_));
 sg13g2_a21oi_1 _09670_ (.A1(net2111),
    .A2(net2225),
    .Y(_00430_),
    .B1(_04113_));
 sg13g2_nor2_1 _09671_ (.A(net1133),
    .B(net2223),
    .Y(_04114_));
 sg13g2_a21oi_1 _09672_ (.A1(net2114),
    .A2(net2223),
    .Y(_00431_),
    .B1(_04114_));
 sg13g2_nor2_1 _09673_ (.A(net955),
    .B(net2223),
    .Y(_04115_));
 sg13g2_a21oi_1 _09674_ (.A1(net2105),
    .A2(net2223),
    .Y(_00432_),
    .B1(_04115_));
 sg13g2_nor2_1 _09675_ (.A(net1002),
    .B(net2229),
    .Y(_04116_));
 sg13g2_a21oi_1 _09676_ (.A1(net2108),
    .A2(net2229),
    .Y(_00433_),
    .B1(_04116_));
 sg13g2_nor2_1 _09677_ (.A(net1094),
    .B(net2226),
    .Y(_04117_));
 sg13g2_a21oi_1 _09678_ (.A1(net2099),
    .A2(net2226),
    .Y(_00434_),
    .B1(_04117_));
 sg13g2_nor2_1 _09679_ (.A(net1167),
    .B(net2226),
    .Y(_04118_));
 sg13g2_a21oi_1 _09680_ (.A1(net2102),
    .A2(net2226),
    .Y(_00435_),
    .B1(_04118_));
 sg13g2_nor2_1 _09681_ (.A(net1076),
    .B(net2224),
    .Y(_04119_));
 sg13g2_a21oi_1 _09682_ (.A1(net2093),
    .A2(net2224),
    .Y(_00436_),
    .B1(_04119_));
 sg13g2_nor2_1 _09683_ (.A(net965),
    .B(net2226),
    .Y(_04120_));
 sg13g2_a21oi_1 _09684_ (.A1(net2090),
    .A2(net2226),
    .Y(_00437_),
    .B1(_04120_));
 sg13g2_nor2_1 _09685_ (.A(net1264),
    .B(net2231),
    .Y(_04121_));
 sg13g2_a21oi_1 _09686_ (.A1(net2096),
    .A2(net2231),
    .Y(_00438_),
    .B1(_04121_));
 sg13g2_nor2_1 _09687_ (.A(net1013),
    .B(net2225),
    .Y(_04122_));
 sg13g2_a21oi_1 _09688_ (.A1(net2081),
    .A2(net2225),
    .Y(_00439_),
    .B1(_04122_));
 sg13g2_nor2_1 _09689_ (.A(net1236),
    .B(net2231),
    .Y(_04123_));
 sg13g2_a21oi_1 _09690_ (.A1(net2084),
    .A2(net2231),
    .Y(_00440_),
    .B1(_04123_));
 sg13g2_nor2_1 _09691_ (.A(net1060),
    .B(net2229),
    .Y(_04124_));
 sg13g2_a21oi_1 _09692_ (.A1(net2087),
    .A2(net2229),
    .Y(_00441_),
    .B1(_04124_));
 sg13g2_nor2_1 _09693_ (.A(net960),
    .B(net2223),
    .Y(_04125_));
 sg13g2_a21oi_1 _09694_ (.A1(net2077),
    .A2(net2223),
    .Y(_00442_),
    .B1(_04125_));
 sg13g2_nor2_1 _09695_ (.A(net1233),
    .B(net2231),
    .Y(_04126_));
 sg13g2_a21oi_1 _09696_ (.A1(net2079),
    .A2(net2231),
    .Y(_00443_),
    .B1(_04126_));
 sg13g2_nor2_1 _09697_ (.A(net997),
    .B(net2229),
    .Y(_04127_));
 sg13g2_a21oi_1 _09698_ (.A1(net2075),
    .A2(net2229),
    .Y(_00444_),
    .B1(_04127_));
 sg13g2_nor2_1 _09699_ (.A(net946),
    .B(net2230),
    .Y(_04128_));
 sg13g2_a21oi_1 _09700_ (.A1(net2073),
    .A2(net2230),
    .Y(_00445_),
    .B1(_04128_));
 sg13g2_nor2_1 _09701_ (.A(net2721),
    .B(net937),
    .Y(_00446_));
 sg13g2_xor2_1 _09702_ (.B(net937),
    .A(net1464),
    .X(_04129_));
 sg13g2_nor2_1 _09703_ (.A(net2721),
    .B(_04129_),
    .Y(_00447_));
 sg13g2_xnor2_1 _09704_ (.Y(_04130_),
    .A(net1331),
    .B(_03490_));
 sg13g2_nor2_1 _09705_ (.A(net2720),
    .B(net1332),
    .Y(_00448_));
 sg13g2_xnor2_1 _09706_ (.Y(_04131_),
    .A(net1367),
    .B(_03491_));
 sg13g2_nor2_1 _09707_ (.A(net2720),
    .B(_04131_),
    .Y(_00449_));
 sg13g2_xor2_1 _09708_ (.B(_03493_),
    .A(net1479),
    .X(_04132_));
 sg13g2_nor2_1 _09709_ (.A(net2720),
    .B(_04132_),
    .Y(_00450_));
 sg13g2_o21ai_1 _09710_ (.B1(net1504),
    .Y(_04133_),
    .A1(net1479),
    .A2(_03493_));
 sg13g2_nor2b_1 _09711_ (.A(_03494_),
    .B_N(_04133_),
    .Y(_04134_));
 sg13g2_nor2_1 _09712_ (.A(net2720),
    .B(_04134_),
    .Y(_00451_));
 sg13g2_nand3_1 _09713_ (.B(_03437_),
    .C(_03439_),
    .A(_03435_),
    .Y(_04135_));
 sg13g2_nor3_1 _09714_ (.A(_02636_),
    .B(_02637_),
    .C(_04135_),
    .Y(_04136_));
 sg13g2_nand4_1 _09715_ (.B(_03573_),
    .C(_03575_),
    .A(\ChiselTop.wild.cpu.io_dmem_rdAddress[31] ),
    .Y(_04137_),
    .D(_04136_));
 sg13g2_o21ai_1 _09716_ (.B1(net2729),
    .Y(_04138_),
    .A1(_03611_),
    .A2(_04137_));
 sg13g2_a21oi_1 _09717_ (.A1(_00906_),
    .A2(_04137_),
    .Y(_00452_),
    .B1(_04138_));
 sg13g2_o21ai_1 _09718_ (.B1(net2729),
    .Y(_04139_),
    .A1(_03637_),
    .A2(_04137_));
 sg13g2_a21oi_1 _09719_ (.A1(_00905_),
    .A2(_04137_),
    .Y(_00453_),
    .B1(_04139_));
 sg13g2_o21ai_1 _09720_ (.B1(net2729),
    .Y(_04140_),
    .A1(_03663_),
    .A2(_04137_));
 sg13g2_a21oi_1 _09721_ (.A1(_00904_),
    .A2(_04137_),
    .Y(_00454_),
    .B1(_04140_));
 sg13g2_o21ai_1 _09722_ (.B1(net2729),
    .Y(_04141_),
    .A1(_03677_),
    .A2(_04137_));
 sg13g2_a21oi_1 _09723_ (.A1(_00903_),
    .A2(_04137_),
    .Y(_00455_),
    .B1(_04141_));
 sg13g2_and2_1 _09724_ (.A(net1214),
    .B(net2730),
    .X(_00456_));
 sg13g2_nor2_1 _09725_ (.A(_00933_),
    .B(net2718),
    .Y(_00457_));
 sg13g2_and2_1 _09726_ (.A(net902),
    .B(net2745),
    .X(_00458_));
 sg13g2_and2_1 _09727_ (.A(net894),
    .B(net2732),
    .X(_00459_));
 sg13g2_nand4_1 _09728_ (.B(_03477_),
    .C(_03478_),
    .A(_03468_),
    .Y(_04142_),
    .D(net2169));
 sg13g2_a21oi_1 _09729_ (.A1(_03467_),
    .A2(_03476_),
    .Y(_00460_),
    .B1(_04142_));
 sg13g2_nor2_1 _09730_ (.A(net2723),
    .B(_02434_),
    .Y(_00529_));
 sg13g2_a21oi_2 _09731_ (.B1(net2723),
    .Y(_00461_),
    .A2(_02434_),
    .A1(_01808_));
 sg13g2_nor2_1 _09732_ (.A(\ChiselTop.wild.cpu._GEN_176[20] ),
    .B(\ChiselTop.wild.cpu._GEN_176[10] ),
    .Y(_04143_));
 sg13g2_a22oi_1 _09733_ (.Y(_04144_),
    .B1(_03525_),
    .B2(_04143_),
    .A2(_01807_),
    .A1(_01806_));
 sg13g2_o21ai_1 _09734_ (.B1(net2731),
    .Y(_04145_),
    .A1(net1521),
    .A2(_04144_));
 sg13g2_nor2_2 _09735_ (.A(net2550),
    .B(_04145_),
    .Y(_00462_));
 sg13g2_nand3_1 _09736_ (.B(net1472),
    .C(net2732),
    .A(net1497),
    .Y(_04146_));
 sg13g2_nor3_1 _09737_ (.A(_00927_),
    .B(net2551),
    .C(_04146_),
    .Y(_00463_));
 sg13g2_nor2_1 _09738_ (.A(net2724),
    .B(_02003_),
    .Y(_00464_));
 sg13g2_and2_1 _09739_ (.A(net2733),
    .B(_01998_),
    .X(_00465_));
 sg13g2_nor2_1 _09740_ (.A(net2724),
    .B(_01880_),
    .Y(_00466_));
 sg13g2_nor2_1 _09741_ (.A(net2722),
    .B(_02188_),
    .Y(_00467_));
 sg13g2_nor2_1 _09742_ (.A(net2722),
    .B(_01819_),
    .Y(_00468_));
 sg13g2_nor2_1 _09743_ (.A(net2725),
    .B(_01738_),
    .Y(_00469_));
 sg13g2_and2_1 _09744_ (.A(net2739),
    .B(_01569_),
    .X(_00470_));
 sg13g2_and2_1 _09745_ (.A(net2739),
    .B(_02256_),
    .X(_00471_));
 sg13g2_and2_1 _09746_ (.A(net2739),
    .B(_02436_),
    .X(_00472_));
 sg13g2_nor2_1 _09747_ (.A(net2721),
    .B(_02581_),
    .Y(_00473_));
 sg13g2_and2_1 _09748_ (.A(net2739),
    .B(_02538_),
    .X(_00474_));
 sg13g2_nor2_1 _09749_ (.A(net2725),
    .B(_02488_),
    .Y(_00475_));
 sg13g2_and2_1 _09750_ (.A(net2735),
    .B(_00965_),
    .X(_00476_));
 sg13g2_nor2_1 _09751_ (.A(net2725),
    .B(_03172_),
    .Y(_00477_));
 sg13g2_and2_1 _09752_ (.A(net1525),
    .B(net2734),
    .X(_00485_));
 sg13g2_nor2_1 _09753_ (.A(net2722),
    .B(_02441_),
    .Y(_00478_));
 sg13g2_and2_1 _09754_ (.A(net2735),
    .B(_03133_),
    .X(_00479_));
 sg13g2_and2_1 _09755_ (.A(net2735),
    .B(_03088_),
    .X(_00480_));
 sg13g2_and2_1 _09756_ (.A(net2735),
    .B(_02964_),
    .X(_00481_));
 sg13g2_nor2_1 _09757_ (.A(net2726),
    .B(_02919_),
    .Y(_00482_));
 sg13g2_and2_1 _09758_ (.A(net2742),
    .B(_02816_),
    .X(_00483_));
 sg13g2_a21oi_1 _09759_ (.A1(_00964_),
    .A2(_02639_),
    .Y(_00484_),
    .B1(net2723));
 sg13g2_and2_1 _09760_ (.A(net2742),
    .B(net895),
    .X(_00486_));
 sg13g2_and2_1 _09761_ (.A(net2741),
    .B(net887),
    .X(_00487_));
 sg13g2_and2_1 _09762_ (.A(net2740),
    .B(net898),
    .X(_00488_));
 sg13g2_and2_1 _09763_ (.A(net2733),
    .B(net882),
    .X(_00489_));
 sg13g2_and2_1 _09764_ (.A(net2733),
    .B(net889),
    .X(_00490_));
 sg13g2_and2_1 _09765_ (.A(net2740),
    .B(net881),
    .X(_00491_));
 sg13g2_and2_1 _09766_ (.A(net2737),
    .B(net900),
    .X(_00492_));
 sg13g2_and2_1 _09767_ (.A(net2737),
    .B(net875),
    .X(_00493_));
 sg13g2_and2_1 _09768_ (.A(net2736),
    .B(net888),
    .X(_00494_));
 sg13g2_and2_1 _09769_ (.A(net2738),
    .B(net871),
    .X(_00495_));
 sg13g2_and2_1 _09770_ (.A(net2736),
    .B(net867),
    .X(_00496_));
 sg13g2_and2_1 _09771_ (.A(net2736),
    .B(net878),
    .X(_00497_));
 sg13g2_and2_1 _09772_ (.A(net2736),
    .B(net890),
    .X(_00498_));
 sg13g2_and2_1 _09773_ (.A(net2736),
    .B(net876),
    .X(_00499_));
 sg13g2_and2_1 _09774_ (.A(net2736),
    .B(net877),
    .X(_00500_));
 sg13g2_and2_1 _09775_ (.A(net2736),
    .B(net903),
    .X(_00501_));
 sg13g2_and2_1 _09776_ (.A(net2737),
    .B(net879),
    .X(_00502_));
 sg13g2_and2_1 _09777_ (.A(net2737),
    .B(net872),
    .X(_00503_));
 sg13g2_and2_1 _09778_ (.A(net2737),
    .B(net873),
    .X(_00504_));
 sg13g2_and2_1 _09779_ (.A(net2737),
    .B(net899),
    .X(_00505_));
 sg13g2_and2_1 _09780_ (.A(net2738),
    .B(net880),
    .X(_00506_));
 sg13g2_and2_1 _09781_ (.A(net2738),
    .B(net896),
    .X(_00507_));
 sg13g2_and2_1 _09782_ (.A(net2738),
    .B(net886),
    .X(_00508_));
 sg13g2_and2_1 _09783_ (.A(net2737),
    .B(net883),
    .X(_00509_));
 sg13g2_and2_1 _09784_ (.A(net2737),
    .B(net901),
    .X(_00510_));
 sg13g2_and2_1 _09785_ (.A(net2743),
    .B(net891),
    .X(_00511_));
 sg13g2_and2_1 _09786_ (.A(net2743),
    .B(net892),
    .X(_00512_));
 sg13g2_and2_1 _09787_ (.A(net2743),
    .B(net885),
    .X(_00513_));
 sg13g2_and2_1 _09788_ (.A(net2743),
    .B(net874),
    .X(_00514_));
 sg13g2_and2_1 _09789_ (.A(net2743),
    .B(net893),
    .X(_00515_));
 sg13g2_and2_1 _09790_ (.A(net2743),
    .B(net868),
    .X(_00516_));
 sg13g2_and2_1 _09791_ (.A(net2743),
    .B(net884),
    .X(_00517_));
 sg13g2_nor3_1 _09792_ (.A(net1499),
    .B(net2551),
    .C(_04146_),
    .Y(_00518_));
 sg13g2_nand3_1 _09793_ (.B(_03527_),
    .C(_03529_),
    .A(net2731),
    .Y(_04147_));
 sg13g2_nand2b_1 _09794_ (.Y(_00519_),
    .B(_04147_),
    .A_N(_00157_));
 sg13g2_and2_1 _09795_ (.A(net2733),
    .B(_01809_),
    .X(_00520_));
 sg13g2_nor2_1 _09796_ (.A(net2723),
    .B(_02638_),
    .Y(_00521_));
 sg13g2_and2_1 _09797_ (.A(net2734),
    .B(\ChiselTop.wild.cpu.decEx_memLow[1] ),
    .X(_00522_));
 sg13g2_and2_1 _09798_ (.A(net2733),
    .B(_01811_),
    .X(_00523_));
 sg13g2_and3_1 _09799_ (.X(_00525_),
    .A(net1472),
    .B(net2733),
    .C(_01805_));
 sg13g2_and2_1 _09800_ (.A(net1312),
    .B(net2730),
    .X(_00526_));
 sg13g2_and2_1 _09801_ (.A(net952),
    .B(net2730),
    .X(_00527_));
 sg13g2_and2_1 _09802_ (.A(net1351),
    .B(net2730),
    .X(_00528_));
 sg13g2_nor3_1 _09803_ (.A(net2715),
    .B(_03601_),
    .C(_03608_),
    .Y(_00530_));
 sg13g2_nor3_2 _09804_ (.A(net2718),
    .B(_03627_),
    .C(_03634_),
    .Y(_00531_));
 sg13g2_nor3_2 _09805_ (.A(net2715),
    .B(_03653_),
    .C(_03660_),
    .Y(_00532_));
 sg13g2_nor3_1 _09806_ (.A(net2715),
    .B(_03667_),
    .C(_03674_),
    .Y(_00533_));
 sg13g2_nor3_1 _09807_ (.A(net2716),
    .B(_03704_),
    .C(_03711_),
    .Y(_00534_));
 sg13g2_nor3_1 _09808_ (.A(net2714),
    .B(_03729_),
    .C(_03736_),
    .Y(_00535_));
 sg13g2_nor3_1 _09809_ (.A(net2711),
    .B(_03743_),
    .C(_03750_),
    .Y(_00536_));
 sg13g2_nor3_1 _09810_ (.A(net2712),
    .B(_03780_),
    .C(_03787_),
    .Y(_00537_));
 sg13g2_nor3_1 _09811_ (.A(net2707),
    .B(_03798_),
    .C(_03805_),
    .Y(_00538_));
 sg13g2_nor3_1 _09812_ (.A(net2706),
    .B(_03811_),
    .C(_03818_),
    .Y(_00539_));
 sg13g2_nor3_1 _09813_ (.A(net2716),
    .B(_03824_),
    .C(_03831_),
    .Y(_00540_));
 sg13g2_nor3_1 _09814_ (.A(net2708),
    .B(_03837_),
    .C(_03844_),
    .Y(_00541_));
 sg13g2_nor3_1 _09815_ (.A(net2709),
    .B(_03849_),
    .C(_03856_),
    .Y(_00542_));
 sg13g2_nor3_1 _09816_ (.A(net2717),
    .B(_03862_),
    .C(_03869_),
    .Y(_00543_));
 sg13g2_nor3_1 _09817_ (.A(net2712),
    .B(_03875_),
    .C(_03882_),
    .Y(_00544_));
 sg13g2_nor3_1 _09818_ (.A(net2717),
    .B(_03888_),
    .C(_03895_),
    .Y(_00545_));
 sg13g2_nor2_1 _09819_ (.A(net2711),
    .B(_03598_),
    .Y(_00546_));
 sg13g2_nor2_1 _09820_ (.A(net2711),
    .B(_03624_),
    .Y(_00547_));
 sg13g2_nor2_1 _09821_ (.A(net2710),
    .B(_03650_),
    .Y(_00548_));
 sg13g2_nor2_1 _09822_ (.A(net2717),
    .B(_03689_),
    .Y(_00549_));
 sg13g2_nor3_1 _09823_ (.A(net2710),
    .B(_03693_),
    .C(_03700_),
    .Y(_00550_));
 sg13g2_nor3_1 _09824_ (.A(net2708),
    .B(_03718_),
    .C(_03725_),
    .Y(_00551_));
 sg13g2_nor2_1 _09825_ (.A(net2709),
    .B(_03765_),
    .Y(_00552_));
 sg13g2_nor3_1 _09826_ (.A(net2712),
    .B(_03769_),
    .C(_03776_),
    .Y(_00553_));
 sg13g2_mux4_1 _09827_ (.S0(net2605),
    .A0(\ChiselTop.wild.cpu.regs[0][24] ),
    .A1(\ChiselTop.wild.cpu.regs[1][24] ),
    .A2(\ChiselTop.wild.cpu.regs[2][24] ),
    .A3(\ChiselTop.wild.cpu.regs[3][24] ),
    .S1(net2581),
    .X(_04148_));
 sg13g2_nor2_1 _09828_ (.A(net2562),
    .B(_04148_),
    .Y(_04149_));
 sg13g2_nor2b_1 _09829_ (.A(\ChiselTop.wild.cpu.regs[29][24] ),
    .B_N(net2609),
    .Y(_04150_));
 sg13g2_nor2_1 _09830_ (.A(net2609),
    .B(\ChiselTop.wild.cpu.regs[28][24] ),
    .Y(_04151_));
 sg13g2_nor3_1 _09831_ (.A(net2581),
    .B(_04150_),
    .C(_04151_),
    .Y(_04152_));
 sg13g2_nor2b_1 _09832_ (.A(\ChiselTop.wild.cpu.regs[31][24] ),
    .B_N(net2605),
    .Y(_04153_));
 sg13g2_o21ai_1 _09833_ (.B1(net2581),
    .Y(_04154_),
    .A1(net2605),
    .A2(\ChiselTop.wild.cpu.regs[30][24] ));
 sg13g2_o21ai_1 _09834_ (.B1(net2562),
    .Y(_04155_),
    .A1(_04153_),
    .A2(_04154_));
 sg13g2_o21ai_1 _09835_ (.B1(net2462),
    .Y(_04156_),
    .A1(_04152_),
    .A2(_04155_));
 sg13g2_nor2_2 _09836_ (.A(_04149_),
    .B(_04156_),
    .Y(_04157_));
 sg13g2_nor3_1 _09837_ (.A(net2714),
    .B(_04149_),
    .C(_04156_),
    .Y(_00554_));
 sg13g2_mux4_1 _09838_ (.S0(net2588),
    .A0(\ChiselTop.wild.cpu.regs[0][25] ),
    .A1(\ChiselTop.wild.cpu.regs[1][25] ),
    .A2(\ChiselTop.wild.cpu.regs[2][25] ),
    .A3(\ChiselTop.wild.cpu.regs[3][25] ),
    .S1(net2568),
    .X(_04158_));
 sg13g2_nor2_1 _09839_ (.A(net2555),
    .B(_04158_),
    .Y(_04159_));
 sg13g2_nor2b_1 _09840_ (.A(\ChiselTop.wild.cpu.regs[29][25] ),
    .B_N(net2586),
    .Y(_04160_));
 sg13g2_nor2_1 _09841_ (.A(net2586),
    .B(\ChiselTop.wild.cpu.regs[28][25] ),
    .Y(_04161_));
 sg13g2_nor3_1 _09842_ (.A(net2567),
    .B(_04160_),
    .C(_04161_),
    .Y(_04162_));
 sg13g2_nor2b_1 _09843_ (.A(\ChiselTop.wild.cpu.regs[31][25] ),
    .B_N(net2587),
    .Y(_04163_));
 sg13g2_o21ai_1 _09844_ (.B1(net2567),
    .Y(_04164_),
    .A1(net2586),
    .A2(\ChiselTop.wild.cpu.regs[30][25] ));
 sg13g2_o21ai_1 _09845_ (.B1(net2559),
    .Y(_04165_),
    .A1(_04163_),
    .A2(_04164_));
 sg13g2_o21ai_1 _09846_ (.B1(net2460),
    .Y(_04166_),
    .A1(_04162_),
    .A2(_04165_));
 sg13g2_nor2_2 _09847_ (.A(_04159_),
    .B(_04166_),
    .Y(_04167_));
 sg13g2_nor3_1 _09848_ (.A(net2707),
    .B(_04159_),
    .C(_04166_),
    .Y(_00555_));
 sg13g2_mux4_1 _09849_ (.S0(net2606),
    .A0(\ChiselTop.wild.cpu.regs[0][26] ),
    .A1(\ChiselTop.wild.cpu.regs[1][26] ),
    .A2(\ChiselTop.wild.cpu.regs[2][26] ),
    .A3(\ChiselTop.wild.cpu.regs[3][26] ),
    .S1(net2579),
    .X(_04168_));
 sg13g2_nor2_1 _09850_ (.A(net2563),
    .B(_04168_),
    .Y(_04169_));
 sg13g2_nor2b_1 _09851_ (.A(\ChiselTop.wild.cpu.regs[29][26] ),
    .B_N(net2606),
    .Y(_04170_));
 sg13g2_nor2_1 _09852_ (.A(net2606),
    .B(\ChiselTop.wild.cpu.regs[28][26] ),
    .Y(_04171_));
 sg13g2_nor3_1 _09853_ (.A(net2579),
    .B(_04170_),
    .C(_04171_),
    .Y(_04172_));
 sg13g2_nor2b_1 _09854_ (.A(\ChiselTop.wild.cpu.regs[31][26] ),
    .B_N(net2606),
    .Y(_04173_));
 sg13g2_o21ai_1 _09855_ (.B1(net2579),
    .Y(_04174_),
    .A1(net2606),
    .A2(\ChiselTop.wild.cpu.regs[30][26] ));
 sg13g2_o21ai_1 _09856_ (.B1(net2563),
    .Y(_04175_),
    .A1(_04173_),
    .A2(_04174_));
 sg13g2_o21ai_1 _09857_ (.B1(net2462),
    .Y(_04176_),
    .A1(_04172_),
    .A2(_04175_));
 sg13g2_nor2_1 _09858_ (.A(_04169_),
    .B(_04176_),
    .Y(_04177_));
 sg13g2_nor3_2 _09859_ (.A(net2718),
    .B(_04169_),
    .C(_04176_),
    .Y(_00556_));
 sg13g2_mux4_1 _09860_ (.S0(net2599),
    .A0(\ChiselTop.wild.cpu.regs[0][27] ),
    .A1(\ChiselTop.wild.cpu.regs[1][27] ),
    .A2(\ChiselTop.wild.cpu.regs[2][27] ),
    .A3(\ChiselTop.wild.cpu.regs[3][27] ),
    .S1(net2574),
    .X(_04178_));
 sg13g2_nor2_1 _09861_ (.A(net2560),
    .B(_04178_),
    .Y(_04179_));
 sg13g2_nor2b_1 _09862_ (.A(\ChiselTop.wild.cpu.regs[29][27] ),
    .B_N(net2599),
    .Y(_04180_));
 sg13g2_nor2_1 _09863_ (.A(net2599),
    .B(\ChiselTop.wild.cpu.regs[28][27] ),
    .Y(_04181_));
 sg13g2_nor3_1 _09864_ (.A(net2574),
    .B(_04180_),
    .C(_04181_),
    .Y(_04182_));
 sg13g2_nor2b_1 _09865_ (.A(\ChiselTop.wild.cpu.regs[31][27] ),
    .B_N(net2599),
    .Y(_04183_));
 sg13g2_o21ai_1 _09866_ (.B1(net2574),
    .Y(_04184_),
    .A1(net2599),
    .A2(\ChiselTop.wild.cpu.regs[30][27] ));
 sg13g2_o21ai_1 _09867_ (.B1(net2560),
    .Y(_04185_),
    .A1(_04183_),
    .A2(_04184_));
 sg13g2_o21ai_1 _09868_ (.B1(net2461),
    .Y(_04186_),
    .A1(_04182_),
    .A2(_04185_));
 sg13g2_nor2_2 _09869_ (.A(_04179_),
    .B(_04186_),
    .Y(_04187_));
 sg13g2_nor3_1 _09870_ (.A(net2714),
    .B(_04179_),
    .C(_04186_),
    .Y(_00557_));
 sg13g2_mux4_1 _09871_ (.S0(net2585),
    .A0(\ChiselTop.wild.cpu.regs[0][28] ),
    .A1(\ChiselTop.wild.cpu.regs[1][28] ),
    .A2(\ChiselTop.wild.cpu.regs[2][28] ),
    .A3(\ChiselTop.wild.cpu.regs[3][28] ),
    .S1(net2565),
    .X(_04188_));
 sg13g2_nor2_1 _09872_ (.A(net2556),
    .B(_04188_),
    .Y(_04189_));
 sg13g2_nor2b_1 _09873_ (.A(\ChiselTop.wild.cpu.regs[29][28] ),
    .B_N(net2585),
    .Y(_04190_));
 sg13g2_nor2_1 _09874_ (.A(net2584),
    .B(net1554),
    .Y(_04191_));
 sg13g2_nor3_1 _09875_ (.A(net2566),
    .B(_04190_),
    .C(_04191_),
    .Y(_04192_));
 sg13g2_nor2b_1 _09876_ (.A(\ChiselTop.wild.cpu.regs[31][28] ),
    .B_N(net2584),
    .Y(_04193_));
 sg13g2_o21ai_1 _09877_ (.B1(net2566),
    .Y(_04194_),
    .A1(net2584),
    .A2(\ChiselTop.wild.cpu.regs[30][28] ));
 sg13g2_o21ai_1 _09878_ (.B1(net2555),
    .Y(_04195_),
    .A1(_04193_),
    .A2(_04194_));
 sg13g2_o21ai_1 _09879_ (.B1(net2459),
    .Y(_04196_),
    .A1(net1555),
    .A2(_04195_));
 sg13g2_nor2_2 _09880_ (.A(_04189_),
    .B(_04196_),
    .Y(_04197_));
 sg13g2_nor3_1 _09881_ (.A(net2706),
    .B(_04189_),
    .C(_04196_),
    .Y(_00558_));
 sg13g2_mux4_1 _09882_ (.S0(net2607),
    .A0(\ChiselTop.wild.cpu.regs[0][29] ),
    .A1(\ChiselTop.wild.cpu.regs[1][29] ),
    .A2(\ChiselTop.wild.cpu.regs[2][29] ),
    .A3(\ChiselTop.wild.cpu.regs[3][29] ),
    .S1(net2580),
    .X(_04198_));
 sg13g2_nor2_1 _09883_ (.A(net2562),
    .B(_04198_),
    .Y(_04199_));
 sg13g2_nor2b_1 _09884_ (.A(\ChiselTop.wild.cpu.regs[29][29] ),
    .B_N(net2607),
    .Y(_04200_));
 sg13g2_nor2_1 _09885_ (.A(net2607),
    .B(\ChiselTop.wild.cpu.regs[28][29] ),
    .Y(_04201_));
 sg13g2_nor3_1 _09886_ (.A(net2579),
    .B(_04200_),
    .C(_04201_),
    .Y(_04202_));
 sg13g2_nor2b_1 _09887_ (.A(\ChiselTop.wild.cpu.regs[31][29] ),
    .B_N(net2607),
    .Y(_04203_));
 sg13g2_o21ai_1 _09888_ (.B1(net2580),
    .Y(_04204_),
    .A1(net2607),
    .A2(\ChiselTop.wild.cpu.regs[30][29] ));
 sg13g2_o21ai_1 _09889_ (.B1(net2562),
    .Y(_04205_),
    .A1(_04203_),
    .A2(_04204_));
 sg13g2_o21ai_1 _09890_ (.B1(net2462),
    .Y(_04206_),
    .A1(_04202_),
    .A2(_04205_));
 sg13g2_nor2_1 _09891_ (.A(_04199_),
    .B(_04206_),
    .Y(_04207_));
 sg13g2_nor3_2 _09892_ (.A(net2719),
    .B(_04199_),
    .C(_04206_),
    .Y(_00559_));
 sg13g2_mux4_1 _09893_ (.S0(net2600),
    .A0(\ChiselTop.wild.cpu.regs[0][30] ),
    .A1(\ChiselTop.wild.cpu.regs[1][30] ),
    .A2(\ChiselTop.wild.cpu.regs[2][30] ),
    .A3(\ChiselTop.wild.cpu.regs[3][30] ),
    .S1(net2575),
    .X(_04208_));
 sg13g2_nor2_1 _09894_ (.A(net2560),
    .B(_04208_),
    .Y(_04209_));
 sg13g2_nor2b_1 _09895_ (.A(\ChiselTop.wild.cpu.regs[29][30] ),
    .B_N(net2601),
    .Y(_04210_));
 sg13g2_nor2_1 _09896_ (.A(net2600),
    .B(\ChiselTop.wild.cpu.regs[28][30] ),
    .Y(_04211_));
 sg13g2_nor3_1 _09897_ (.A(net2575),
    .B(_04210_),
    .C(_04211_),
    .Y(_04212_));
 sg13g2_nor2b_1 _09898_ (.A(\ChiselTop.wild.cpu.regs[31][30] ),
    .B_N(net2600),
    .Y(_04213_));
 sg13g2_o21ai_1 _09899_ (.B1(net2575),
    .Y(_04214_),
    .A1(net2600),
    .A2(\ChiselTop.wild.cpu.regs[30][30] ));
 sg13g2_o21ai_1 _09900_ (.B1(net2560),
    .Y(_04215_),
    .A1(_04213_),
    .A2(_04214_));
 sg13g2_o21ai_1 _09901_ (.B1(net2461),
    .Y(_04216_),
    .A1(_04212_),
    .A2(_04215_));
 sg13g2_nor2_2 _09902_ (.A(_04209_),
    .B(_04216_),
    .Y(_04217_));
 sg13g2_nor3_1 _09903_ (.A(net2714),
    .B(_04209_),
    .C(_04216_),
    .Y(_00560_));
 sg13g2_mux4_1 _09904_ (.S0(net2606),
    .A0(\ChiselTop.wild.cpu.regs[0][31] ),
    .A1(\ChiselTop.wild.cpu.regs[1][31] ),
    .A2(\ChiselTop.wild.cpu.regs[2][31] ),
    .A3(\ChiselTop.wild.cpu.regs[3][31] ),
    .S1(net2579),
    .X(_04218_));
 sg13g2_nor2_1 _09905_ (.A(net2563),
    .B(_04218_),
    .Y(_04219_));
 sg13g2_nor2b_1 _09906_ (.A(\ChiselTop.wild.cpu.regs[29][31] ),
    .B_N(net2603),
    .Y(_04220_));
 sg13g2_nor2_1 _09907_ (.A(net2603),
    .B(\ChiselTop.wild.cpu.regs[28][31] ),
    .Y(_04221_));
 sg13g2_nor3_1 _09908_ (.A(net2577),
    .B(_04220_),
    .C(_04221_),
    .Y(_04222_));
 sg13g2_nor2b_1 _09909_ (.A(\ChiselTop.wild.cpu.regs[31][31] ),
    .B_N(net2603),
    .Y(_04223_));
 sg13g2_o21ai_1 _09910_ (.B1(net2576),
    .Y(_04224_),
    .A1(net2603),
    .A2(\ChiselTop.wild.cpu.regs[30][31] ));
 sg13g2_o21ai_1 _09911_ (.B1(net2561),
    .Y(_04225_),
    .A1(_04223_),
    .A2(_04224_));
 sg13g2_o21ai_1 _09912_ (.B1(net2461),
    .Y(_04226_),
    .A1(_04222_),
    .A2(_04225_));
 sg13g2_nor2_2 _09913_ (.A(_04219_),
    .B(_04226_),
    .Y(_04227_));
 sg13g2_nor3_2 _09914_ (.A(net2715),
    .B(_04219_),
    .C(_04226_),
    .Y(_00561_));
 sg13g2_nor2_1 _09915_ (.A(_00931_),
    .B(net2718),
    .Y(_00564_));
 sg13g2_nor3_2 _09916_ (.A(net2715),
    .B(_02170_),
    .C(_02177_),
    .Y(_00565_));
 sg13g2_nor3_2 _09917_ (.A(net2718),
    .B(_01986_),
    .C(_01993_),
    .Y(_00566_));
 sg13g2_nor3_2 _09918_ (.A(net2715),
    .B(_01929_),
    .C(_01936_),
    .Y(_00567_));
 sg13g2_nor3_1 _09919_ (.A(net2715),
    .B(_02238_),
    .C(_02245_),
    .Y(_00568_));
 sg13g2_nor3_2 _09920_ (.A(net2716),
    .B(_01866_),
    .C(_01873_),
    .Y(_00569_));
 sg13g2_nor3_1 _09921_ (.A(net2714),
    .B(_01792_),
    .C(_01799_),
    .Y(_00570_));
 sg13g2_nor3_1 _09922_ (.A(net2710),
    .B(_01723_),
    .C(_01730_),
    .Y(_00571_));
 sg13g2_nor3_1 _09923_ (.A(net2712),
    .B(_01653_),
    .C(_01660_),
    .Y(_00572_));
 sg13g2_nor3_1 _09924_ (.A(net2707),
    .B(_02330_),
    .C(_02337_),
    .Y(_00573_));
 sg13g2_nor3_2 _09925_ (.A(net2706),
    .B(_02374_),
    .C(_02381_),
    .Y(_00574_));
 sg13g2_nor3_1 _09926_ (.A(net2706),
    .B(_02290_),
    .C(_02297_),
    .Y(_00575_));
 sg13g2_nor3_1 _09927_ (.A(net2708),
    .B(_02423_),
    .C(_02430_),
    .Y(_00576_));
 sg13g2_nor3_1 _09928_ (.A(net2708),
    .B(_02614_),
    .C(_02621_),
    .Y(_00577_));
 sg13g2_nor3_1 _09929_ (.A(net2717),
    .B(_02570_),
    .C(_02577_),
    .Y(_00578_));
 sg13g2_nor3_1 _09930_ (.A(net2712),
    .B(_02476_),
    .C(_02483_),
    .Y(_00579_));
 sg13g2_nor3_1 _09931_ (.A(net2717),
    .B(_02522_),
    .C(_02529_),
    .Y(_00580_));
 sg13g2_nor3_1 _09932_ (.A(net2706),
    .B(_01555_),
    .C(_01564_),
    .Y(_00581_));
 sg13g2_nor3_1 _09933_ (.A(net2707),
    .B(_03197_),
    .C(_03204_),
    .Y(_00582_));
 sg13g2_nor3_1 _09934_ (.A(net2707),
    .B(_03273_),
    .C(_03280_),
    .Y(_00583_));
 sg13g2_nor3_1 _09935_ (.A(net2714),
    .B(_03237_),
    .C(_03244_),
    .Y(_00584_));
 sg13g2_nor3_1 _09936_ (.A(net2709),
    .B(_03159_),
    .C(_03166_),
    .Y(_00585_));
 sg13g2_nor3_1 _09937_ (.A(net2708),
    .B(_03120_),
    .C(_03127_),
    .Y(_00586_));
 sg13g2_nor3_2 _09938_ (.A(net2706),
    .B(_03075_),
    .C(_03082_),
    .Y(_00587_));
 sg13g2_nor3_2 _09939_ (.A(net2709),
    .B(_03003_),
    .C(_03010_),
    .Y(_00588_));
 sg13g2_nor3_1 _09940_ (.A(net2714),
    .B(_03041_),
    .C(_03048_),
    .Y(_00589_));
 sg13g2_nor3_1 _09941_ (.A(net2706),
    .B(_02952_),
    .C(_02959_),
    .Y(_00590_));
 sg13g2_nor3_2 _09942_ (.A(net2718),
    .B(_02905_),
    .C(_02912_),
    .Y(_00591_));
 sg13g2_nor3_2 _09943_ (.A(net2714),
    .B(_02864_),
    .C(_02871_),
    .Y(_00592_));
 sg13g2_nor3_2 _09944_ (.A(net2706),
    .B(_03370_),
    .C(_03377_),
    .Y(_00593_));
 sg13g2_nor3_2 _09945_ (.A(net2719),
    .B(_03327_),
    .C(_03334_),
    .Y(_00594_));
 sg13g2_nor3_2 _09946_ (.A(net2715),
    .B(_02805_),
    .C(_02812_),
    .Y(_00595_));
 sg13g2_nor3_2 _09947_ (.A(net2718),
    .B(_03418_),
    .C(_03425_),
    .Y(_00596_));
 sg13g2_nor2_1 _09948_ (.A(_00929_),
    .B(net2724),
    .Y(_00598_));
 sg13g2_nor2_1 _09949_ (.A(net2717),
    .B(_02168_),
    .Y(_00599_));
 sg13g2_nor2_1 _09950_ (.A(net2723),
    .B(net2149),
    .Y(_00600_));
 sg13g2_nor2_2 _09951_ (.A(net2718),
    .B(net2140),
    .Y(_00601_));
 sg13g2_nor2_2 _09952_ (.A(net2723),
    .B(_02236_),
    .Y(_00602_));
 sg13g2_nor2_1 _09953_ (.A(net2717),
    .B(net2152),
    .Y(_00603_));
 sg13g2_nor2_1 _09954_ (.A(net2719),
    .B(_01789_),
    .Y(_00604_));
 sg13g2_nor2_1 _09955_ (.A(net2710),
    .B(net2143),
    .Y(_00605_));
 sg13g2_nor2_1 _09956_ (.A(net2710),
    .B(net2146),
    .Y(_00606_));
 sg13g2_nor2_1 _09957_ (.A(net2710),
    .B(_02328_),
    .Y(_00607_));
 sg13g2_nor2_1 _09958_ (.A(net2708),
    .B(net2129),
    .Y(_00608_));
 sg13g2_nor2_1 _09959_ (.A(net2711),
    .B(_02288_),
    .Y(_00609_));
 sg13g2_and2_1 _09960_ (.A(net2735),
    .B(net2124),
    .X(_00610_));
 sg13g2_nor2_1 _09961_ (.A(net2708),
    .B(net2125),
    .Y(_00611_));
 sg13g2_nor2_1 _09962_ (.A(net2711),
    .B(net2122),
    .Y(_00612_));
 sg13g2_nor2_1 _09963_ (.A(net2710),
    .B(net2120),
    .Y(_00613_));
 sg13g2_nor2_1 _09964_ (.A(net2722),
    .B(_02520_),
    .Y(_00614_));
 sg13g2_nor2_1 _09965_ (.A(net2710),
    .B(net2113),
    .Y(_00615_));
 sg13g2_nor2_1 _09966_ (.A(net2711),
    .B(net2116),
    .Y(_00616_));
 sg13g2_nor2_1 _09967_ (.A(net2720),
    .B(net2107),
    .Y(_00617_));
 sg13g2_nor2_1 _09968_ (.A(net2719),
    .B(net2110),
    .Y(_00618_));
 sg13g2_nor2_1 _09969_ (.A(net2709),
    .B(net2101),
    .Y(_00619_));
 sg13g2_nor2_1 _09970_ (.A(net2720),
    .B(net2103),
    .Y(_00620_));
 sg13g2_nor2_1 _09971_ (.A(net2720),
    .B(net2095),
    .Y(_00621_));
 sg13g2_nor2_1 _09972_ (.A(net2708),
    .B(net2091),
    .Y(_00622_));
 sg13g2_nor2_1 _09973_ (.A(net2722),
    .B(net2098),
    .Y(_00623_));
 sg13g2_nor2_1 _09974_ (.A(net2711),
    .B(net2083),
    .Y(_00624_));
 sg13g2_nor2_1 _09975_ (.A(net2722),
    .B(net2086),
    .Y(_00625_));
 sg13g2_nor2_1 _09976_ (.A(net2722),
    .B(net2089),
    .Y(_00626_));
 sg13g2_nor2_1 _09977_ (.A(net2720),
    .B(net2078),
    .Y(_00627_));
 sg13g2_nor2_1 _09978_ (.A(net2717),
    .B(net2080),
    .Y(_00628_));
 sg13g2_nor2_1 _09979_ (.A(net2719),
    .B(_02803_),
    .Y(_00629_));
 sg13g2_nor2_2 _09980_ (.A(net2723),
    .B(net2074),
    .Y(_00630_));
 sg13g2_and2_1 _09981_ (.A(net2649),
    .B(net2731),
    .X(_00631_));
 sg13g2_and2_1 _09982_ (.A(net2648),
    .B(net2730),
    .X(_00632_));
 sg13g2_and2_1 _09983_ (.A(net1450),
    .B(net2730),
    .X(_00633_));
 sg13g2_and2_1 _09984_ (.A(net1475),
    .B(net2745),
    .X(_00634_));
 sg13g2_and2_1 _09985_ (.A(net2612),
    .B(net2729),
    .X(_00635_));
 sg13g2_nor2_1 _09986_ (.A(net2719),
    .B(_00970_),
    .Y(_00636_));
 sg13g2_nor4_1 _09987_ (.A(\ChiselTop.cntReg[25] ),
    .B(_00948_),
    .C(\ChiselTop.cntReg[27] ),
    .D(\ChiselTop.cntReg[26] ),
    .Y(_04228_));
 sg13g2_nor4_1 _09988_ (.A(\ChiselTop.cntReg[14] ),
    .B(_00946_),
    .C(\ChiselTop.cntReg[19] ),
    .D(_00947_),
    .Y(_04229_));
 sg13g2_nor4_2 _09989_ (.A(\ChiselTop.cntReg[29] ),
    .B(\ChiselTop.cntReg[28] ),
    .C(\ChiselTop.cntReg[31] ),
    .Y(_04230_),
    .D(\ChiselTop.cntReg[30] ));
 sg13g2_and4_1 _09990_ (.A(\ChiselTop.cntReg[20] ),
    .B(\ChiselTop.cntReg[21] ),
    .C(\ChiselTop.cntReg[22] ),
    .D(\ChiselTop.cntReg[23] ),
    .X(_04231_));
 sg13g2_nand4_1 _09991_ (.B(_04229_),
    .C(_04230_),
    .A(_04228_),
    .Y(_04232_),
    .D(_04231_));
 sg13g2_nor4_1 _09992_ (.A(\ChiselTop.cntReg[10] ),
    .B(_00945_),
    .C(\ChiselTop.cntReg[13] ),
    .D(\ChiselTop.cntReg[12] ),
    .Y(_04233_));
 sg13g2_nor2_1 _09993_ (.A(\ChiselTop.cntReg[7] ),
    .B(\ChiselTop.cntReg[8] ),
    .Y(_04234_));
 sg13g2_nand4_1 _09994_ (.B(\ChiselTop.cntReg[9] ),
    .C(_04233_),
    .A(\ChiselTop.cntReg[6] ),
    .Y(_04235_),
    .D(_04234_));
 sg13g2_nor4_1 _09995_ (.A(\ChiselTop.cntReg[3] ),
    .B(\ChiselTop.cntReg[2] ),
    .C(\ChiselTop.cntReg[5] ),
    .D(\ChiselTop.cntReg[4] ),
    .Y(_04236_));
 sg13g2_nor2_1 _09996_ (.A(\ChiselTop.cntReg[1] ),
    .B(net1460),
    .Y(_04237_));
 sg13g2_nand4_1 _09997_ (.B(\ChiselTop.cntReg[17] ),
    .C(_04236_),
    .A(\ChiselTop.cntReg[16] ),
    .Y(_04238_),
    .D(_04237_));
 sg13g2_nor3_1 _09998_ (.A(_04232_),
    .B(_04235_),
    .C(_04238_),
    .Y(_04239_));
 sg13g2_nand2b_1 _09999_ (.Y(_04240_),
    .B(net2729),
    .A_N(_04239_));
 sg13g2_nor2_1 _10000_ (.A(_00959_),
    .B(net2324),
    .Y(_00637_));
 sg13g2_and2_1 _10001_ (.A(\ChiselTop.cntReg[1] ),
    .B(net1460),
    .X(_04241_));
 sg13g2_nor3_1 _10002_ (.A(net1461),
    .B(net2324),
    .C(_04241_),
    .Y(_00638_));
 sg13g2_and2_1 _10003_ (.A(net1400),
    .B(_04241_),
    .X(_04242_));
 sg13g2_nor2_1 _10004_ (.A(net1400),
    .B(_04241_),
    .Y(_04243_));
 sg13g2_nor3_1 _10005_ (.A(net2324),
    .B(_04242_),
    .C(net1401),
    .Y(_00639_));
 sg13g2_and2_1 _10006_ (.A(net1442),
    .B(_04242_),
    .X(_04244_));
 sg13g2_nor2_1 _10007_ (.A(net1442),
    .B(_04242_),
    .Y(_04245_));
 sg13g2_nor3_1 _10008_ (.A(net2327),
    .B(_04244_),
    .C(_04245_),
    .Y(_00640_));
 sg13g2_and2_1 _10009_ (.A(net1348),
    .B(_04244_),
    .X(_04246_));
 sg13g2_nor2_1 _10010_ (.A(net1348),
    .B(_04244_),
    .Y(_04247_));
 sg13g2_nor3_1 _10011_ (.A(net2324),
    .B(_04246_),
    .C(net1349),
    .Y(_00641_));
 sg13g2_xnor2_1 _10012_ (.Y(_04248_),
    .A(net1457),
    .B(_04246_));
 sg13g2_nor2_1 _10013_ (.A(net2324),
    .B(_04248_),
    .Y(_00642_));
 sg13g2_a21oi_1 _10014_ (.A1(\ChiselTop.cntReg[5] ),
    .A2(_04246_),
    .Y(_04249_),
    .B1(net1162));
 sg13g2_and3_1 _10015_ (.X(_04250_),
    .A(\ChiselTop.cntReg[5] ),
    .B(net1162),
    .C(_04246_));
 sg13g2_nor3_1 _10016_ (.A(net2325),
    .B(net1163),
    .C(_04250_),
    .Y(_00643_));
 sg13g2_nor2_1 _10017_ (.A(net1433),
    .B(_04250_),
    .Y(_04251_));
 sg13g2_and2_1 _10018_ (.A(net1433),
    .B(_04250_),
    .X(_04252_));
 sg13g2_nor3_1 _10019_ (.A(net2325),
    .B(net1434),
    .C(_04252_),
    .Y(_00644_));
 sg13g2_nor2_1 _10020_ (.A(net1444),
    .B(_04252_),
    .Y(_04253_));
 sg13g2_and2_1 _10021_ (.A(net1444),
    .B(_04252_),
    .X(_04254_));
 sg13g2_nor3_1 _10022_ (.A(net2325),
    .B(_04253_),
    .C(_04254_),
    .Y(_00645_));
 sg13g2_nor2_1 _10023_ (.A(net1435),
    .B(_04254_),
    .Y(_04255_));
 sg13g2_and2_1 _10024_ (.A(net1435),
    .B(_04254_),
    .X(_04256_));
 sg13g2_nor3_1 _10025_ (.A(net2325),
    .B(net1436),
    .C(_04256_),
    .Y(_00646_));
 sg13g2_nor2_1 _10026_ (.A(net1364),
    .B(_04256_),
    .Y(_04257_));
 sg13g2_and2_1 _10027_ (.A(net1364),
    .B(_04256_),
    .X(_04258_));
 sg13g2_nor3_1 _10028_ (.A(net2327),
    .B(net1365),
    .C(_04258_),
    .Y(_00647_));
 sg13g2_nor2_1 _10029_ (.A(net1360),
    .B(_04258_),
    .Y(_04259_));
 sg13g2_and2_1 _10030_ (.A(net1360),
    .B(_04258_),
    .X(_04260_));
 sg13g2_nor3_1 _10031_ (.A(net2325),
    .B(net1361),
    .C(_04260_),
    .Y(_00648_));
 sg13g2_nor2_1 _10032_ (.A(net1362),
    .B(_04260_),
    .Y(_04261_));
 sg13g2_and2_1 _10033_ (.A(net1362),
    .B(_04260_),
    .X(_04262_));
 sg13g2_nor3_1 _10034_ (.A(net2325),
    .B(_04261_),
    .C(_04262_),
    .Y(_00649_));
 sg13g2_nor2_1 _10035_ (.A(net1404),
    .B(_04262_),
    .Y(_04263_));
 sg13g2_and2_1 _10036_ (.A(net1404),
    .B(_04262_),
    .X(_04264_));
 sg13g2_nor3_1 _10037_ (.A(net2325),
    .B(_04263_),
    .C(_04264_),
    .Y(_00650_));
 sg13g2_nor2_1 _10038_ (.A(net1421),
    .B(_04264_),
    .Y(_04265_));
 sg13g2_and2_1 _10039_ (.A(net1421),
    .B(_04264_),
    .X(_04266_));
 sg13g2_nor3_1 _10040_ (.A(net2326),
    .B(_04265_),
    .C(_04266_),
    .Y(_00651_));
 sg13g2_nor2_1 _10041_ (.A(net1390),
    .B(_04266_),
    .Y(_04267_));
 sg13g2_and2_1 _10042_ (.A(net1390),
    .B(_04266_),
    .X(_04268_));
 sg13g2_nor3_1 _10043_ (.A(net2326),
    .B(net1391),
    .C(_04268_),
    .Y(_00652_));
 sg13g2_nor2_1 _10044_ (.A(net1422),
    .B(_04268_),
    .Y(_04269_));
 sg13g2_and2_1 _10045_ (.A(net1422),
    .B(_04268_),
    .X(_04270_));
 sg13g2_nor3_1 _10046_ (.A(net2325),
    .B(_04269_),
    .C(_04270_),
    .Y(_00653_));
 sg13g2_nor2_1 _10047_ (.A(net1393),
    .B(_04270_),
    .Y(_04271_));
 sg13g2_and2_1 _10048_ (.A(net1393),
    .B(_04270_),
    .X(_04272_));
 sg13g2_nor3_1 _10049_ (.A(net2326),
    .B(net1394),
    .C(_04272_),
    .Y(_00654_));
 sg13g2_nor2_1 _10050_ (.A(net1372),
    .B(_04272_),
    .Y(_04273_));
 sg13g2_and2_1 _10051_ (.A(net1372),
    .B(_04272_),
    .X(_04274_));
 sg13g2_nor3_1 _10052_ (.A(net2326),
    .B(net1373),
    .C(_04274_),
    .Y(_00655_));
 sg13g2_nor2_1 _10053_ (.A(net1395),
    .B(_04274_),
    .Y(_04275_));
 sg13g2_and2_1 _10054_ (.A(net1395),
    .B(_04274_),
    .X(_04276_));
 sg13g2_nor3_1 _10055_ (.A(net2326),
    .B(_04275_),
    .C(_04276_),
    .Y(_00656_));
 sg13g2_nor2_1 _10056_ (.A(net1430),
    .B(_04276_),
    .Y(_04277_));
 sg13g2_and2_1 _10057_ (.A(net1430),
    .B(_04276_),
    .X(_04278_));
 sg13g2_nor3_1 _10058_ (.A(net2326),
    .B(_04277_),
    .C(_04278_),
    .Y(_00657_));
 sg13g2_nor2_1 _10059_ (.A(net1416),
    .B(_04278_),
    .Y(_04279_));
 sg13g2_and3_1 _10060_ (.X(_04280_),
    .A(\ChiselTop.cntReg[20] ),
    .B(net1416),
    .C(_04276_));
 sg13g2_nor3_1 _10061_ (.A(net2326),
    .B(net1417),
    .C(_04280_),
    .Y(_00658_));
 sg13g2_nor2_1 _10062_ (.A(net1409),
    .B(_04280_),
    .Y(_04281_));
 sg13g2_and2_1 _10063_ (.A(net1409),
    .B(_04280_),
    .X(_04282_));
 sg13g2_nor3_1 _10064_ (.A(net2323),
    .B(net1410),
    .C(_04282_),
    .Y(_00659_));
 sg13g2_xnor2_1 _10065_ (.Y(_04283_),
    .A(net1447),
    .B(_04282_));
 sg13g2_nor2_1 _10066_ (.A(net2324),
    .B(_04283_),
    .Y(_00660_));
 sg13g2_a21oi_1 _10067_ (.A1(\ChiselTop.cntReg[23] ),
    .A2(_04282_),
    .Y(_04284_),
    .B1(net1097));
 sg13g2_and3_1 _10068_ (.X(_04285_),
    .A(\ChiselTop.cntReg[23] ),
    .B(net1097),
    .C(_04282_));
 sg13g2_nor3_1 _10069_ (.A(net2324),
    .B(net1098),
    .C(_04285_),
    .Y(_00661_));
 sg13g2_nor2_1 _10070_ (.A(net1419),
    .B(_04285_),
    .Y(_04286_));
 sg13g2_and2_1 _10071_ (.A(net1419),
    .B(_04285_),
    .X(_04287_));
 sg13g2_nor3_1 _10072_ (.A(net2323),
    .B(net1420),
    .C(_04287_),
    .Y(_00662_));
 sg13g2_xnor2_1 _10073_ (.Y(_04288_),
    .A(net1452),
    .B(_04287_));
 sg13g2_nor2_1 _10074_ (.A(net2323),
    .B(_04288_),
    .Y(_00663_));
 sg13g2_a21oi_1 _10075_ (.A1(\ChiselTop.cntReg[26] ),
    .A2(_04287_),
    .Y(_04289_),
    .B1(net1154));
 sg13g2_and3_1 _10076_ (.X(_04290_),
    .A(net1154),
    .B(net1452),
    .C(_04287_));
 sg13g2_nor3_1 _10077_ (.A(net2323),
    .B(net1155),
    .C(_04290_),
    .Y(_00664_));
 sg13g2_nor2_1 _10078_ (.A(net1456),
    .B(_04290_),
    .Y(_04291_));
 sg13g2_and2_1 _10079_ (.A(net1456),
    .B(_04290_),
    .X(_04292_));
 sg13g2_nor3_1 _10080_ (.A(net2323),
    .B(_04291_),
    .C(_04292_),
    .Y(_00665_));
 sg13g2_xnor2_1 _10081_ (.Y(_04293_),
    .A(net1463),
    .B(_04292_));
 sg13g2_nor2_1 _10082_ (.A(net2323),
    .B(_04293_),
    .Y(_00666_));
 sg13g2_a21oi_1 _10083_ (.A1(\ChiselTop.cntReg[29] ),
    .A2(_04292_),
    .Y(_04294_),
    .B1(net1303));
 sg13g2_and3_1 _10084_ (.X(_04295_),
    .A(\ChiselTop.cntReg[29] ),
    .B(net1303),
    .C(_04292_));
 sg13g2_nor3_1 _10085_ (.A(net2323),
    .B(net1304),
    .C(_04295_),
    .Y(_00667_));
 sg13g2_xnor2_1 _10086_ (.Y(_04296_),
    .A(net1425),
    .B(_04295_));
 sg13g2_nor2_1 _10087_ (.A(net2323),
    .B(net1426),
    .Y(_00668_));
 sg13g2_nor2_1 _10088_ (.A(_03522_),
    .B(_04032_),
    .Y(_04297_));
 sg13g2_nor2_1 _10089_ (.A(net984),
    .B(net2218),
    .Y(_04298_));
 sg13g2_a21oi_1 _10090_ (.A1(net2137),
    .A2(net2217),
    .Y(_00669_),
    .B1(_04298_));
 sg13g2_nor2_1 _10091_ (.A(net1136),
    .B(net2221),
    .Y(_04299_));
 sg13g2_a21oi_1 _10092_ (.A1(net2147),
    .A2(net2220),
    .Y(_00670_),
    .B1(_04299_));
 sg13g2_nor2_1 _10093_ (.A(net1061),
    .B(net2220),
    .Y(_04300_));
 sg13g2_a21oi_1 _10094_ (.A1(net2139),
    .A2(net2220),
    .Y(_00671_),
    .B1(_04300_));
 sg13g2_nor2_1 _10095_ (.A(net1003),
    .B(net2217),
    .Y(_04301_));
 sg13g2_a21oi_1 _10096_ (.A1(net2135),
    .A2(net2217),
    .Y(_00672_),
    .B1(_04301_));
 sg13g2_nor2_1 _10097_ (.A(net967),
    .B(net2217),
    .Y(_04302_));
 sg13g2_a21oi_1 _10098_ (.A1(net2150),
    .A2(net2217),
    .Y(_00673_),
    .B1(_04302_));
 sg13g2_nor2_1 _10099_ (.A(net1222),
    .B(net2218),
    .Y(_04303_));
 sg13g2_a21oi_1 _10100_ (.A1(net2142),
    .A2(net2217),
    .Y(_00674_),
    .B1(_04303_));
 sg13g2_nor2_1 _10101_ (.A(net1084),
    .B(net2216),
    .Y(_04304_));
 sg13g2_a21oi_1 _10102_ (.A1(net2143),
    .A2(net2216),
    .Y(_00675_),
    .B1(_04304_));
 sg13g2_nor2_1 _10103_ (.A(net1050),
    .B(net2216),
    .Y(_04305_));
 sg13g2_a21oi_1 _10104_ (.A1(net2145),
    .A2(net2216),
    .Y(_00676_),
    .B1(_04305_));
 sg13g2_nor2_1 _10105_ (.A(net1067),
    .B(net2222),
    .Y(_04306_));
 sg13g2_a21oi_1 _10106_ (.A1(net2130),
    .A2(net2214),
    .Y(_00677_),
    .B1(_04306_));
 sg13g2_nor2_1 _10107_ (.A(net1005),
    .B(net2214),
    .Y(_04307_));
 sg13g2_a21oi_1 _10108_ (.A1(net2127),
    .A2(net2214),
    .Y(_00678_),
    .B1(_04307_));
 sg13g2_nor2_1 _10109_ (.A(net1231),
    .B(net2213),
    .Y(_04308_));
 sg13g2_a21oi_1 _10110_ (.A1(net2132),
    .A2(net2213),
    .Y(_00679_),
    .B1(_04308_));
 sg13g2_mux2_1 _10111_ (.A0(net1131),
    .A1(net2123),
    .S(net2216),
    .X(_00680_));
 sg13g2_nor2_1 _10112_ (.A(net1014),
    .B(net2215),
    .Y(_04309_));
 sg13g2_a21oi_1 _10113_ (.A1(net2125),
    .A2(net2215),
    .Y(_00681_),
    .B1(_04309_));
 sg13g2_nor2_1 _10114_ (.A(net1069),
    .B(net2219),
    .Y(_04310_));
 sg13g2_a21oi_1 _10115_ (.A1(net2121),
    .A2(net2219),
    .Y(_00682_),
    .B1(_04310_));
 sg13g2_nor2_1 _10116_ (.A(net980),
    .B(net2215),
    .Y(_04311_));
 sg13g2_a21oi_1 _10117_ (.A1(net2119),
    .A2(net2215),
    .Y(_00683_),
    .B1(_04311_));
 sg13g2_nor2_1 _10118_ (.A(net1211),
    .B(net2220),
    .Y(_04312_));
 sg13g2_a21oi_1 _10119_ (.A1(net2118),
    .A2(net2220),
    .Y(_00684_),
    .B1(_04312_));
 sg13g2_nor2_1 _10120_ (.A(net1019),
    .B(net2219),
    .Y(_04313_));
 sg13g2_a21oi_1 _10121_ (.A1(net2112),
    .A2(net2219),
    .Y(_00685_),
    .B1(_04313_));
 sg13g2_nor2_1 _10122_ (.A(net1090),
    .B(net2213),
    .Y(_04314_));
 sg13g2_a21oi_1 _10123_ (.A1(net2115),
    .A2(net2213),
    .Y(_00686_),
    .B1(_04314_));
 sg13g2_nor2_1 _10124_ (.A(net1111),
    .B(net2213),
    .Y(_04315_));
 sg13g2_a21oi_1 _10125_ (.A1(net2105),
    .A2(net2213),
    .Y(_00687_),
    .B1(_04315_));
 sg13g2_nor2_1 _10126_ (.A(net1036),
    .B(net2219),
    .Y(_04316_));
 sg13g2_a21oi_1 _10127_ (.A1(net2108),
    .A2(net2219),
    .Y(_00688_),
    .B1(_04316_));
 sg13g2_nor2_1 _10128_ (.A(net966),
    .B(net2216),
    .Y(_04317_));
 sg13g2_a21oi_1 _10129_ (.A1(net2099),
    .A2(net2216),
    .Y(_00689_),
    .B1(_04317_));
 sg13g2_nor2_1 _10130_ (.A(net1219),
    .B(net2215),
    .Y(_04318_));
 sg13g2_a21oi_1 _10131_ (.A1(net2102),
    .A2(net2215),
    .Y(_00690_),
    .B1(_04318_));
 sg13g2_nor2_1 _10132_ (.A(net1124),
    .B(net2214),
    .Y(_04319_));
 sg13g2_a21oi_1 _10133_ (.A1(net2093),
    .A2(net2214),
    .Y(_00691_),
    .B1(_04319_));
 sg13g2_nor2_1 _10134_ (.A(net1091),
    .B(net2215),
    .Y(_04320_));
 sg13g2_a21oi_1 _10135_ (.A1(net2090),
    .A2(net2215),
    .Y(_00692_),
    .B1(_04320_));
 sg13g2_nor2_1 _10136_ (.A(net1269),
    .B(net2220),
    .Y(_04321_));
 sg13g2_a21oi_1 _10137_ (.A1(net2096),
    .A2(net2218),
    .Y(_00693_),
    .B1(_04321_));
 sg13g2_nor2_1 _10138_ (.A(net977),
    .B(net2213),
    .Y(_04322_));
 sg13g2_a21oi_1 _10139_ (.A1(net2082),
    .A2(net2213),
    .Y(_00694_),
    .B1(_04322_));
 sg13g2_nor2_1 _10140_ (.A(net1128),
    .B(net2220),
    .Y(_04323_));
 sg13g2_a21oi_1 _10141_ (.A1(net2084),
    .A2(net2220),
    .Y(_00695_),
    .B1(_04323_));
 sg13g2_nor2_1 _10142_ (.A(net1130),
    .B(net2219),
    .Y(_04324_));
 sg13g2_a21oi_1 _10143_ (.A1(net2088),
    .A2(net2219),
    .Y(_00696_),
    .B1(_04324_));
 sg13g2_nor2_1 _10144_ (.A(net953),
    .B(net2214),
    .Y(_04325_));
 sg13g2_a21oi_1 _10145_ (.A1(net2077),
    .A2(net2214),
    .Y(_00697_),
    .B1(_04325_));
 sg13g2_nor2_1 _10146_ (.A(net961),
    .B(net2221),
    .Y(_04326_));
 sg13g2_a21oi_1 _10147_ (.A1(net2079),
    .A2(net2221),
    .Y(_00698_),
    .B1(_04326_));
 sg13g2_nor2_1 _10148_ (.A(net1250),
    .B(net2218),
    .Y(_04327_));
 sg13g2_a21oi_1 _10149_ (.A1(net2075),
    .A2(net2218),
    .Y(_00699_),
    .B1(_04327_));
 sg13g2_nor2_1 _10150_ (.A(net1198),
    .B(net2217),
    .Y(_04328_));
 sg13g2_a21oi_1 _10151_ (.A1(net2073),
    .A2(net2217),
    .Y(_00700_),
    .B1(_04328_));
 sg13g2_nand2_1 _10152_ (.Y(_04329_),
    .A(_02000_),
    .B(\ChiselTop.wild.cpu.decEx_memLow[0] ));
 sg13g2_a22oi_1 _10153_ (.Y(_04330_),
    .B1(_04329_),
    .B2(_03563_),
    .A2(_03577_),
    .A1(net2550));
 sg13g2_nand3_1 _10154_ (.B(_03576_),
    .C(_04330_),
    .A(_03572_),
    .Y(_04331_));
 sg13g2_o21ai_1 _10155_ (.B1(net2164),
    .Y(_04332_),
    .A1(net2409),
    .A2(_04157_));
 sg13g2_a21o_1 _10156_ (.A2(net2409),
    .A1(net2098),
    .B1(_04332_),
    .X(_04333_));
 sg13g2_a22oi_1 _10157_ (.Y(_04334_),
    .B1(_03795_),
    .B2(_03808_),
    .A2(_03611_),
    .A1(net2524));
 sg13g2_o21ai_1 _10158_ (.B1(_04333_),
    .Y(_04335_),
    .A1(_03571_),
    .A2(_04334_));
 sg13g2_mux2_1 _10159_ (.A0(_04335_),
    .A1(net1432),
    .S(_04331_),
    .X(_00701_));
 sg13g2_o21ai_1 _10160_ (.B1(net2164),
    .Y(_04336_),
    .A1(net2410),
    .A2(_04167_));
 sg13g2_a21oi_1 _10161_ (.A1(net2083),
    .A2(net2409),
    .Y(_04337_),
    .B1(_04336_));
 sg13g2_and2_1 _10162_ (.A(net2524),
    .B(_03637_),
    .X(_04338_));
 sg13g2_nand4_1 _10163_ (.B(net2191),
    .C(net2464),
    .A(net2527),
    .Y(_04339_),
    .D(_04338_));
 sg13g2_nand2b_1 _10164_ (.Y(_04340_),
    .B(_04339_),
    .A_N(_04337_));
 sg13g2_mux2_1 _10165_ (.A0(_04340_),
    .A1(net1445),
    .S(_04331_),
    .X(_00702_));
 sg13g2_and2_1 _10166_ (.A(net2524),
    .B(_03663_),
    .X(_04341_));
 sg13g2_nand4_1 _10167_ (.B(net2191),
    .C(net2464),
    .A(net2527),
    .Y(_04342_),
    .D(_04341_));
 sg13g2_and2_1 _10168_ (.A(net2086),
    .B(net2411),
    .X(_04343_));
 sg13g2_o21ai_1 _10169_ (.B1(net2165),
    .Y(_04344_),
    .A1(net2411),
    .A2(_04177_));
 sg13g2_o21ai_1 _10170_ (.B1(_04342_),
    .Y(_04345_),
    .A1(_04343_),
    .A2(_04344_));
 sg13g2_mux2_1 _10171_ (.A0(_04345_),
    .A1(net1438),
    .S(_04331_),
    .X(_00703_));
 sg13g2_and2_1 _10172_ (.A(net2524),
    .B(_03677_),
    .X(_04346_));
 sg13g2_nand4_1 _10173_ (.B(net2191),
    .C(net2464),
    .A(net2527),
    .Y(_04347_),
    .D(_04346_));
 sg13g2_and2_1 _10174_ (.A(net2089),
    .B(net2409),
    .X(_04348_));
 sg13g2_o21ai_1 _10175_ (.B1(net2165),
    .Y(_04349_),
    .A1(net2409),
    .A2(_04187_));
 sg13g2_o21ai_1 _10176_ (.B1(_04347_),
    .Y(_04350_),
    .A1(_04348_),
    .A2(_04349_));
 sg13g2_mux2_1 _10177_ (.A0(_04350_),
    .A1(net1392),
    .S(_04331_),
    .X(_00704_));
 sg13g2_o21ai_1 _10178_ (.B1(net2164),
    .Y(_04351_),
    .A1(net2409),
    .A2(_04197_));
 sg13g2_a21oi_1 _10179_ (.A1(_03368_),
    .A2(net2409),
    .Y(_04352_),
    .B1(_04351_));
 sg13g2_and2_1 _10180_ (.A(net2524),
    .B(_03714_),
    .X(_04353_));
 sg13g2_nand4_1 _10181_ (.B(net2191),
    .C(net2464),
    .A(net2527),
    .Y(_04354_),
    .D(_04353_));
 sg13g2_nand2b_1 _10182_ (.Y(_04355_),
    .B(_04354_),
    .A_N(_04352_));
 sg13g2_mux2_1 _10183_ (.A0(_04355_),
    .A1(net1437),
    .S(_04331_),
    .X(_00705_));
 sg13g2_o21ai_1 _10184_ (.B1(net2163),
    .Y(_04356_),
    .A1(net2411),
    .A2(_04207_));
 sg13g2_a21oi_1 _10185_ (.A1(net2080),
    .A2(net2411),
    .Y(_04357_),
    .B1(_04356_));
 sg13g2_and2_1 _10186_ (.A(net2524),
    .B(_03739_),
    .X(_04358_));
 sg13g2_nand4_1 _10187_ (.B(net2191),
    .C(net2464),
    .A(net2527),
    .Y(_04359_),
    .D(_04358_));
 sg13g2_nand2b_1 _10188_ (.Y(_04360_),
    .B(_04359_),
    .A_N(_04357_));
 sg13g2_mux2_1 _10189_ (.A0(_04360_),
    .A1(net1443),
    .S(_04331_),
    .X(_00706_));
 sg13g2_o21ai_1 _10190_ (.B1(net2164),
    .Y(_04361_),
    .A1(net2409),
    .A2(_04217_));
 sg13g2_a21oi_1 _10191_ (.A1(_02803_),
    .A2(net2410),
    .Y(_04362_),
    .B1(_04361_));
 sg13g2_and2_1 _10192_ (.A(net2524),
    .B(_03753_),
    .X(_04363_));
 sg13g2_nand4_1 _10193_ (.B(net2191),
    .C(net2464),
    .A(net2527),
    .Y(_04364_),
    .D(_04363_));
 sg13g2_nand2b_1 _10194_ (.Y(_04365_),
    .B(_04364_),
    .A_N(_04362_));
 sg13g2_mux2_1 _10195_ (.A0(_04365_),
    .A1(net1483),
    .S(_04331_),
    .X(_00707_));
 sg13g2_o21ai_1 _10196_ (.B1(net2165),
    .Y(_04366_),
    .A1(net2411),
    .A2(_04227_));
 sg13g2_a21oi_1 _10197_ (.A1(net2074),
    .A2(net2411),
    .Y(_04367_),
    .B1(_04366_));
 sg13g2_and2_1 _10198_ (.A(_03563_),
    .B(_03790_),
    .X(_04368_));
 sg13g2_nand4_1 _10199_ (.B(net2191),
    .C(net2464),
    .A(net2527),
    .Y(_04369_),
    .D(_04368_));
 sg13g2_nand2b_1 _10200_ (.Y(_04370_),
    .B(_04369_),
    .A_N(_04367_));
 sg13g2_mux2_1 _10201_ (.A0(_04370_),
    .A1(net1440),
    .S(_04331_),
    .X(_00708_));
 sg13g2_nor2_1 _10202_ (.A(_03524_),
    .B(_04032_),
    .Y(_04371_));
 sg13g2_nor2_1 _10203_ (.A(net1259),
    .B(net2208),
    .Y(_04372_));
 sg13g2_a21oi_1 _10204_ (.A1(net2136),
    .A2(net2207),
    .Y(_00709_),
    .B1(_04372_));
 sg13g2_nor2_1 _10205_ (.A(net958),
    .B(net2210),
    .Y(_04373_));
 sg13g2_a21oi_1 _10206_ (.A1(net2147),
    .A2(net2210),
    .Y(_00710_),
    .B1(_04373_));
 sg13g2_nor2_1 _10207_ (.A(net1126),
    .B(net2210),
    .Y(_04374_));
 sg13g2_a21oi_1 _10208_ (.A1(net2139),
    .A2(net2210),
    .Y(_00711_),
    .B1(_04374_));
 sg13g2_nor2_1 _10209_ (.A(net972),
    .B(net2207),
    .Y(_04375_));
 sg13g2_a21oi_1 _10210_ (.A1(net2134),
    .A2(net2207),
    .Y(_00712_),
    .B1(_04375_));
 sg13g2_nor2_1 _10211_ (.A(net1127),
    .B(net2207),
    .Y(_04376_));
 sg13g2_a21oi_1 _10212_ (.A1(net2150),
    .A2(net2207),
    .Y(_00713_),
    .B1(_04376_));
 sg13g2_nor2_1 _10213_ (.A(net1104),
    .B(net2208),
    .Y(_04377_));
 sg13g2_a21oi_1 _10214_ (.A1(net2142),
    .A2(net2207),
    .Y(_00714_),
    .B1(_04377_));
 sg13g2_nor2_1 _10215_ (.A(net1170),
    .B(net2206),
    .Y(_04378_));
 sg13g2_a21oi_1 _10216_ (.A1(net2143),
    .A2(net2206),
    .Y(_00715_),
    .B1(_04378_));
 sg13g2_nor2_1 _10217_ (.A(net1239),
    .B(net2206),
    .Y(_04379_));
 sg13g2_a21oi_1 _10218_ (.A1(net2145),
    .A2(net2206),
    .Y(_00716_),
    .B1(_04379_));
 sg13g2_nor2_1 _10219_ (.A(net1113),
    .B(net2212),
    .Y(_04380_));
 sg13g2_a21oi_1 _10220_ (.A1(net2130),
    .A2(net2204),
    .Y(_00717_),
    .B1(_04380_));
 sg13g2_nor2_1 _10221_ (.A(net1230),
    .B(net2204),
    .Y(_04381_));
 sg13g2_a21oi_1 _10222_ (.A1(net2127),
    .A2(net2204),
    .Y(_00718_),
    .B1(_04381_));
 sg13g2_nor2_1 _10223_ (.A(net1092),
    .B(net2203),
    .Y(_04382_));
 sg13g2_a21oi_1 _10224_ (.A1(net2132),
    .A2(net2203),
    .Y(_00719_),
    .B1(_04382_));
 sg13g2_mux2_1 _10225_ (.A0(net1187),
    .A1(net2123),
    .S(net2206),
    .X(_00720_));
 sg13g2_nor2_1 _10226_ (.A(net1047),
    .B(net2205),
    .Y(_04383_));
 sg13g2_a21oi_1 _10227_ (.A1(net2125),
    .A2(net2205),
    .Y(_00721_),
    .B1(_04383_));
 sg13g2_nor2_1 _10228_ (.A(net1093),
    .B(net2209),
    .Y(_04384_));
 sg13g2_a21oi_1 _10229_ (.A1(net2121),
    .A2(net2209),
    .Y(_00722_),
    .B1(_04384_));
 sg13g2_nor2_1 _10230_ (.A(net1030),
    .B(net2205),
    .Y(_04385_));
 sg13g2_a21oi_1 _10231_ (.A1(net2119),
    .A2(net2205),
    .Y(_00723_),
    .B1(_04385_));
 sg13g2_nor2_1 _10232_ (.A(net1082),
    .B(net2211),
    .Y(_04386_));
 sg13g2_a21oi_1 _10233_ (.A1(net2118),
    .A2(net2211),
    .Y(_00724_),
    .B1(_04386_));
 sg13g2_nor2_1 _10234_ (.A(net1205),
    .B(net2209),
    .Y(_04387_));
 sg13g2_a21oi_1 _10235_ (.A1(net2112),
    .A2(net2209),
    .Y(_00725_),
    .B1(_04387_));
 sg13g2_nor2_1 _10236_ (.A(net1246),
    .B(net2203),
    .Y(_04388_));
 sg13g2_a21oi_1 _10237_ (.A1(net2114),
    .A2(net2203),
    .Y(_00726_),
    .B1(_04388_));
 sg13g2_nor2_1 _10238_ (.A(net998),
    .B(net2203),
    .Y(_04389_));
 sg13g2_a21oi_1 _10239_ (.A1(net2106),
    .A2(net2203),
    .Y(_00727_),
    .B1(_04389_));
 sg13g2_nor2_1 _10240_ (.A(net1063),
    .B(net2209),
    .Y(_04390_));
 sg13g2_a21oi_1 _10241_ (.A1(net2109),
    .A2(net2209),
    .Y(_00728_),
    .B1(_04390_));
 sg13g2_nor2_1 _10242_ (.A(net1284),
    .B(net2206),
    .Y(_04391_));
 sg13g2_a21oi_1 _10243_ (.A1(net2099),
    .A2(net2206),
    .Y(_00729_),
    .B1(_04391_));
 sg13g2_nor2_1 _10244_ (.A(net1201),
    .B(net2205),
    .Y(_04392_));
 sg13g2_a21oi_1 _10245_ (.A1(net2102),
    .A2(net2205),
    .Y(_00730_),
    .B1(_04392_));
 sg13g2_nor2_1 _10246_ (.A(net1278),
    .B(net2204),
    .Y(_04393_));
 sg13g2_a21oi_1 _10247_ (.A1(net2093),
    .A2(net2204),
    .Y(_00731_),
    .B1(_04393_));
 sg13g2_nor2_1 _10248_ (.A(net1081),
    .B(net2205),
    .Y(_04394_));
 sg13g2_a21oi_1 _10249_ (.A1(net2090),
    .A2(net2205),
    .Y(_00732_),
    .B1(_04394_));
 sg13g2_nor2_1 _10250_ (.A(net992),
    .B(net2210),
    .Y(_04395_));
 sg13g2_a21oi_1 _10251_ (.A1(net2096),
    .A2(net2210),
    .Y(_00733_),
    .B1(_04395_));
 sg13g2_nor2_1 _10252_ (.A(net1105),
    .B(net2203),
    .Y(_04396_));
 sg13g2_a21oi_1 _10253_ (.A1(net2081),
    .A2(net2203),
    .Y(_00734_),
    .B1(_04396_));
 sg13g2_nor2_1 _10254_ (.A(net1234),
    .B(net2210),
    .Y(_04397_));
 sg13g2_a21oi_1 _10255_ (.A1(net2084),
    .A2(net2210),
    .Y(_00735_),
    .B1(_04397_));
 sg13g2_nor2_1 _10256_ (.A(net1261),
    .B(net2209),
    .Y(_04398_));
 sg13g2_a21oi_1 _10257_ (.A1(net2088),
    .A2(net2209),
    .Y(_00736_),
    .B1(_04398_));
 sg13g2_nor2_1 _10258_ (.A(net1119),
    .B(net2204),
    .Y(_04399_));
 sg13g2_a21oi_1 _10259_ (.A1(net2077),
    .A2(net2204),
    .Y(_00737_),
    .B1(_04399_));
 sg13g2_nor2_1 _10260_ (.A(net1034),
    .B(net2211),
    .Y(_04400_));
 sg13g2_a21oi_1 _10261_ (.A1(net2080),
    .A2(net2211),
    .Y(_00738_),
    .B1(_04400_));
 sg13g2_nor2_1 _10262_ (.A(net981),
    .B(net2208),
    .Y(_04401_));
 sg13g2_a21oi_1 _10263_ (.A1(net2075),
    .A2(net2208),
    .Y(_00739_),
    .B1(_04401_));
 sg13g2_nor2_1 _10264_ (.A(net1183),
    .B(net2207),
    .Y(_04402_));
 sg13g2_a21oi_1 _10265_ (.A1(net2073),
    .A2(net2207),
    .Y(_00740_),
    .B1(_04402_));
 sg13g2_nor2_1 _10266_ (.A(_03520_),
    .B(_04032_),
    .Y(_04403_));
 sg13g2_nor2_1 _10267_ (.A(net990),
    .B(net2197),
    .Y(_04404_));
 sg13g2_a21oi_1 _10268_ (.A1(net2137),
    .A2(net2197),
    .Y(_00741_),
    .B1(_04404_));
 sg13g2_nor2_1 _10269_ (.A(net1070),
    .B(net2199),
    .Y(_04405_));
 sg13g2_a21oi_1 _10270_ (.A1(net2148),
    .A2(net2199),
    .Y(_00742_),
    .B1(_04405_));
 sg13g2_nor2_1 _10271_ (.A(net1100),
    .B(net2199),
    .Y(_04406_));
 sg13g2_a21oi_1 _10272_ (.A1(net2139),
    .A2(net2199),
    .Y(_00743_),
    .B1(_04406_));
 sg13g2_nor2_1 _10273_ (.A(net1245),
    .B(net2197),
    .Y(_04407_));
 sg13g2_a21oi_1 _10274_ (.A1(net2134),
    .A2(net2197),
    .Y(_00744_),
    .B1(_04407_));
 sg13g2_nor2_1 _10275_ (.A(net1025),
    .B(net2197),
    .Y(_04408_));
 sg13g2_a21oi_1 _10276_ (.A1(net2150),
    .A2(net2197),
    .Y(_00745_),
    .B1(_04408_));
 sg13g2_nor2_1 _10277_ (.A(net1077),
    .B(net2198),
    .Y(_04409_));
 sg13g2_a21oi_1 _10278_ (.A1(net2141),
    .A2(net2198),
    .Y(_00746_),
    .B1(_04409_));
 sg13g2_nor2_1 _10279_ (.A(net995),
    .B(net2196),
    .Y(_04410_));
 sg13g2_a21oi_1 _10280_ (.A1(net2143),
    .A2(net2196),
    .Y(_00747_),
    .B1(_04410_));
 sg13g2_nor2_1 _10281_ (.A(net1256),
    .B(net2196),
    .Y(_04411_));
 sg13g2_a21oi_1 _10282_ (.A1(net2146),
    .A2(net2196),
    .Y(_00748_),
    .B1(_04411_));
 sg13g2_nor2_1 _10283_ (.A(net1088),
    .B(net2194),
    .Y(_04412_));
 sg13g2_a21oi_1 _10284_ (.A1(net2130),
    .A2(net2202),
    .Y(_00749_),
    .B1(_04412_));
 sg13g2_nor2_1 _10285_ (.A(net1173),
    .B(net2194),
    .Y(_04413_));
 sg13g2_a21oi_1 _10286_ (.A1(net2127),
    .A2(net2194),
    .Y(_00750_),
    .B1(_04413_));
 sg13g2_nor2_1 _10287_ (.A(net945),
    .B(net2198),
    .Y(_04414_));
 sg13g2_a21oi_1 _10288_ (.A1(net2132),
    .A2(net2198),
    .Y(_00751_),
    .B1(_04414_));
 sg13g2_mux2_1 _10289_ (.A0(net1087),
    .A1(net2123),
    .S(net2196),
    .X(_00752_));
 sg13g2_nor2_1 _10290_ (.A(net1008),
    .B(net2196),
    .Y(_04415_));
 sg13g2_a21oi_1 _10291_ (.A1(net2125),
    .A2(net2196),
    .Y(_00753_),
    .B1(_04415_));
 sg13g2_nor2_1 _10292_ (.A(net1001),
    .B(net2200),
    .Y(_04416_));
 sg13g2_a21oi_1 _10293_ (.A1(net2121),
    .A2(net2200),
    .Y(_00754_),
    .B1(_04416_));
 sg13g2_nor2_1 _10294_ (.A(net1326),
    .B(net2195),
    .Y(_04417_));
 sg13g2_a21oi_1 _10295_ (.A1(net2119),
    .A2(net2195),
    .Y(_00755_),
    .B1(_04417_));
 sg13g2_nor2_1 _10296_ (.A(net1199),
    .B(net2200),
    .Y(_04418_));
 sg13g2_a21oi_1 _10297_ (.A1(net2118),
    .A2(net2200),
    .Y(_00756_),
    .B1(_04418_));
 sg13g2_nor2_1 _10298_ (.A(net1071),
    .B(net2193),
    .Y(_04419_));
 sg13g2_a21oi_1 _10299_ (.A1(net2112),
    .A2(net2193),
    .Y(_00757_),
    .B1(_04419_));
 sg13g2_nor2_1 _10300_ (.A(net964),
    .B(net2193),
    .Y(_04420_));
 sg13g2_a21oi_1 _10301_ (.A1(net2115),
    .A2(net2193),
    .Y(_00758_),
    .B1(_04420_));
 sg13g2_nor2_1 _10302_ (.A(net1150),
    .B(net2193),
    .Y(_04421_));
 sg13g2_a21oi_1 _10303_ (.A1(net2106),
    .A2(net2193),
    .Y(_00759_),
    .B1(_04421_));
 sg13g2_nor2_1 _10304_ (.A(net1169),
    .B(net2198),
    .Y(_04422_));
 sg13g2_a21oi_1 _10305_ (.A1(net2109),
    .A2(net2198),
    .Y(_00760_),
    .B1(_04422_));
 sg13g2_nor2_1 _10306_ (.A(net1178),
    .B(net2195),
    .Y(_04423_));
 sg13g2_a21oi_1 _10307_ (.A1(net2099),
    .A2(net2195),
    .Y(_00761_),
    .B1(_04423_));
 sg13g2_nor2_1 _10308_ (.A(net1095),
    .B(net2195),
    .Y(_04424_));
 sg13g2_a21oi_1 _10309_ (.A1(net2102),
    .A2(net2195),
    .Y(_00762_),
    .B1(_04424_));
 sg13g2_nor2_1 _10310_ (.A(net948),
    .B(net2194),
    .Y(_04425_));
 sg13g2_a21oi_1 _10311_ (.A1(net2093),
    .A2(net2194),
    .Y(_00763_),
    .B1(_04425_));
 sg13g2_nor2_1 _10312_ (.A(net1054),
    .B(net2195),
    .Y(_04426_));
 sg13g2_a21oi_1 _10313_ (.A1(net2090),
    .A2(net2195),
    .Y(_00764_),
    .B1(_04426_));
 sg13g2_nor2_1 _10314_ (.A(net950),
    .B(net2199),
    .Y(_04427_));
 sg13g2_a21oi_1 _10315_ (.A1(net2096),
    .A2(net2199),
    .Y(_00765_),
    .B1(_04427_));
 sg13g2_nor2_1 _10316_ (.A(net1015),
    .B(net2193),
    .Y(_04428_));
 sg13g2_a21oi_1 _10317_ (.A1(net2081),
    .A2(net2193),
    .Y(_00766_),
    .B1(_04428_));
 sg13g2_nor2_1 _10318_ (.A(net1165),
    .B(net2199),
    .Y(_04429_));
 sg13g2_a21oi_1 _10319_ (.A1(net2085),
    .A2(net2199),
    .Y(_00767_),
    .B1(_04429_));
 sg13g2_nor2_1 _10320_ (.A(net994),
    .B(net2198),
    .Y(_04430_));
 sg13g2_a21oi_1 _10321_ (.A1(net2087),
    .A2(net2198),
    .Y(_00768_),
    .B1(_04430_));
 sg13g2_nor2_1 _10322_ (.A(net1145),
    .B(net2194),
    .Y(_04431_));
 sg13g2_a21oi_1 _10323_ (.A1(net2077),
    .A2(net2194),
    .Y(_00769_),
    .B1(_04431_));
 sg13g2_nor2_1 _10324_ (.A(net1032),
    .B(net2200),
    .Y(_04432_));
 sg13g2_a21oi_1 _10325_ (.A1(net2079),
    .A2(net2200),
    .Y(_00770_),
    .B1(_04432_));
 sg13g2_nor2_1 _10326_ (.A(net971),
    .B(net2201),
    .Y(_04433_));
 sg13g2_a21oi_1 _10327_ (.A1(net2075),
    .A2(net2201),
    .Y(_00771_),
    .B1(_04433_));
 sg13g2_nor2_1 _10328_ (.A(net1121),
    .B(net2197),
    .Y(_04434_));
 sg13g2_a21oi_1 _10329_ (.A1(net2073),
    .A2(net2197),
    .Y(_00772_),
    .B1(_04434_));
 sg13g2_nand2_1 _10330_ (.Y(_04435_),
    .A(net859),
    .B(net2168));
 sg13g2_nor2_2 _10331_ (.A(net2724),
    .B(net2192),
    .Y(_04436_));
 sg13g2_nand3_1 _10332_ (.B(net2734),
    .C(_01213_),
    .A(net1488),
    .Y(_04437_));
 sg13g2_nor2_1 _10333_ (.A(net2547),
    .B(_01925_),
    .Y(_04438_));
 sg13g2_o21ai_1 _10334_ (.B1(_04436_),
    .Y(_04439_),
    .A1(net2616),
    .A2(_01913_));
 sg13g2_o21ai_1 _10335_ (.B1(_04435_),
    .Y(_00773_),
    .A1(_04438_),
    .A2(_04439_));
 sg13g2_o21ai_1 _10336_ (.B1(_04436_),
    .Y(_04440_),
    .A1(net2547),
    .A2(_02235_));
 sg13g2_a21o_1 _10337_ (.A2(_02222_),
    .A1(net2547),
    .B1(_04440_),
    .X(_04441_));
 sg13g2_o21ai_1 _10338_ (.B1(_04441_),
    .Y(_00774_),
    .A1(_03481_),
    .A2(net2179));
 sg13g2_o21ai_1 _10339_ (.B1(_04436_),
    .Y(_04442_),
    .A1(net2547),
    .A2(_01862_));
 sg13g2_a21o_1 _10340_ (.A2(_01859_),
    .A1(net2547),
    .B1(_04442_),
    .X(_04443_));
 sg13g2_nand2_1 _10341_ (.Y(_04444_),
    .A(_03472_),
    .B(net2169));
 sg13g2_o21ai_1 _10342_ (.B1(_04443_),
    .Y(_00775_),
    .A1(_03476_),
    .A2(_04444_));
 sg13g2_nand2_1 _10343_ (.Y(_04445_),
    .A(net2547),
    .B(_01778_));
 sg13g2_a21oi_1 _10344_ (.A1(net2616),
    .A2(_01788_),
    .Y(_04446_),
    .B1(net2190));
 sg13g2_nand2_1 _10345_ (.Y(_04447_),
    .A(_04445_),
    .B(_04446_));
 sg13g2_nand3_1 _10346_ (.B(\ChiselTop.wild.cpu.pcReg[4] ),
    .C(_03470_),
    .A(\ChiselTop.wild.cpu.pcReg[5] ),
    .Y(_04448_));
 sg13g2_xor2_1 _10347_ (.B(_03472_),
    .A(net860),
    .X(_04449_));
 sg13g2_o21ai_1 _10348_ (.B1(_04447_),
    .Y(_00776_),
    .A1(net2179),
    .A2(_04449_));
 sg13g2_o21ai_1 _10349_ (.B1(net2176),
    .Y(_04450_),
    .A1(net2543),
    .A2(_01718_));
 sg13g2_a21o_1 _10350_ (.A2(_01707_),
    .A1(net2543),
    .B1(_04450_),
    .X(_04451_));
 sg13g2_nor2_2 _10351_ (.A(_00952_),
    .B(_04448_),
    .Y(_04452_));
 sg13g2_xnor2_1 _10352_ (.Y(_04453_),
    .A(_00952_),
    .B(_04448_));
 sg13g2_o21ai_1 _10353_ (.B1(_04451_),
    .Y(_00777_),
    .A1(net2180),
    .A2(_04453_));
 sg13g2_and2_1 _10354_ (.A(net2539),
    .B(_01639_),
    .X(_04454_));
 sg13g2_o21ai_1 _10355_ (.B1(net2175),
    .Y(_04455_),
    .A1(net2539),
    .A2(_01650_));
 sg13g2_a21oi_1 _10356_ (.A1(net866),
    .A2(_04452_),
    .Y(_04456_),
    .B1(net2180));
 sg13g2_o21ai_1 _10357_ (.B1(_04456_),
    .Y(_04457_),
    .A1(net866),
    .A2(_04452_));
 sg13g2_o21ai_1 _10358_ (.B1(_04457_),
    .Y(_00778_),
    .A1(_04454_),
    .A2(_04455_));
 sg13g2_o21ai_1 _10359_ (.B1(net2175),
    .Y(_04458_),
    .A1(net2539),
    .A2(_02324_));
 sg13g2_a21o_1 _10360_ (.A2(_02322_),
    .A1(net2539),
    .B1(_04458_),
    .X(_04459_));
 sg13g2_a21oi_1 _10361_ (.A1(net866),
    .A2(_04452_),
    .Y(_04460_),
    .B1(net849));
 sg13g2_nand3_1 _10362_ (.B(net849),
    .C(_04452_),
    .A(net1415),
    .Y(_04461_));
 sg13g2_nand2_1 _10363_ (.Y(_04462_),
    .A(net2167),
    .B(_04461_));
 sg13g2_o21ai_1 _10364_ (.B1(_04459_),
    .Y(_00779_),
    .A1(_04460_),
    .A2(_04462_));
 sg13g2_o21ai_1 _10365_ (.B1(net2175),
    .Y(_04463_),
    .A1(net2537),
    .A2(_02371_));
 sg13g2_a21o_1 _10366_ (.A2(_02368_),
    .A1(net2537),
    .B1(_04463_),
    .X(_04464_));
 sg13g2_nor2_2 _10367_ (.A(_00953_),
    .B(_04461_),
    .Y(_04465_));
 sg13g2_xnor2_1 _10368_ (.Y(_04466_),
    .A(_00953_),
    .B(_04461_));
 sg13g2_o21ai_1 _10369_ (.B1(_04464_),
    .Y(_00780_),
    .A1(net2180),
    .A2(_04466_));
 sg13g2_and2_1 _10370_ (.A(net2536),
    .B(_02280_),
    .X(_04467_));
 sg13g2_o21ai_1 _10371_ (.B1(net2175),
    .Y(_04468_),
    .A1(net2537),
    .A2(_02286_));
 sg13g2_a21oi_1 _10372_ (.A1(net863),
    .A2(_04465_),
    .Y(_04469_),
    .B1(net2180));
 sg13g2_o21ai_1 _10373_ (.B1(_04469_),
    .Y(_04470_),
    .A1(net863),
    .A2(_04465_));
 sg13g2_o21ai_1 _10374_ (.B1(_04470_),
    .Y(_00781_),
    .A1(_04467_),
    .A2(_04468_));
 sg13g2_o21ai_1 _10375_ (.B1(net2175),
    .Y(_04471_),
    .A1(net2537),
    .A2(_02419_));
 sg13g2_a21o_1 _10376_ (.A2(_02413_),
    .A1(net2536),
    .B1(_04471_),
    .X(_04472_));
 sg13g2_a21oi_1 _10377_ (.A1(net863),
    .A2(_04465_),
    .Y(_04473_),
    .B1(net838));
 sg13g2_nand3_1 _10378_ (.B(net838),
    .C(_04465_),
    .A(net1516),
    .Y(_04474_));
 sg13g2_nand2_1 _10379_ (.Y(_04475_),
    .A(net2167),
    .B(_04474_));
 sg13g2_o21ai_1 _10380_ (.B1(_04472_),
    .Y(_00782_),
    .A1(_04473_),
    .A2(_04475_));
 sg13g2_o21ai_1 _10381_ (.B1(net2175),
    .Y(_04476_),
    .A1(net2538),
    .A2(_02611_));
 sg13g2_a21oi_1 _10382_ (.A1(net2536),
    .A2(_02609_),
    .Y(_04477_),
    .B1(_04476_));
 sg13g2_nor2_2 _10383_ (.A(_00954_),
    .B(_04474_),
    .Y(_04478_));
 sg13g2_xnor2_1 _10384_ (.Y(_04479_),
    .A(net852),
    .B(_04474_));
 sg13g2_a21o_1 _10385_ (.A2(_04479_),
    .A1(net2167),
    .B1(_04477_),
    .X(_00783_));
 sg13g2_and2_1 _10386_ (.A(net2536),
    .B(_02560_),
    .X(_04480_));
 sg13g2_o21ai_1 _10387_ (.B1(net2175),
    .Y(_04481_),
    .A1(net2537),
    .A2(_02566_));
 sg13g2_a21oi_1 _10388_ (.A1(net865),
    .A2(_04478_),
    .Y(_04482_),
    .B1(net2180));
 sg13g2_o21ai_1 _10389_ (.B1(_04482_),
    .Y(_04483_),
    .A1(net865),
    .A2(_04478_));
 sg13g2_o21ai_1 _10390_ (.B1(_04483_),
    .Y(_00784_),
    .A1(_04480_),
    .A2(_04481_));
 sg13g2_a221oi_1 _10391_ (.B2(net2184),
    .C1(net2540),
    .B1(_02472_),
    .A1(_02467_),
    .Y(_04484_),
    .A2(_02469_));
 sg13g2_a21o_1 _10392_ (.A2(_02468_),
    .A1(net2539),
    .B1(net2189),
    .X(_04485_));
 sg13g2_a21o_1 _10393_ (.A2(_04478_),
    .A1(net865),
    .B1(net836),
    .X(_04486_));
 sg13g2_nand3_1 _10394_ (.B(net836),
    .C(_04478_),
    .A(net865),
    .Y(_04487_));
 sg13g2_nand3_1 _10395_ (.B(_04486_),
    .C(_04487_),
    .A(net2167),
    .Y(_04488_));
 sg13g2_o21ai_1 _10396_ (.B1(_04488_),
    .Y(_00785_),
    .A1(_04484_),
    .A2(_04485_));
 sg13g2_a221oi_1 _10397_ (.B2(_02518_),
    .C1(net2540),
    .B1(_02515_),
    .A1(net2184),
    .Y(_04489_),
    .A2(_02493_));
 sg13g2_a21oi_1 _10398_ (.A1(net2540),
    .A2(_02517_),
    .Y(_04490_),
    .B1(_04489_));
 sg13g2_nand2_1 _10399_ (.Y(_04491_),
    .A(net2175),
    .B(_04490_));
 sg13g2_nor2_1 _10400_ (.A(_00955_),
    .B(_04487_),
    .Y(_04492_));
 sg13g2_xnor2_1 _10401_ (.Y(_04493_),
    .A(_00955_),
    .B(_04487_));
 sg13g2_o21ai_1 _10402_ (.B1(_04491_),
    .Y(_00786_),
    .A1(net2180),
    .A2(_04493_));
 sg13g2_xnor2_1 _10403_ (.Y(_04494_),
    .A(net858),
    .B(_04492_));
 sg13g2_a21oi_1 _10404_ (.A1(net2542),
    .A2(_01546_),
    .Y(_04495_),
    .B1(net2189));
 sg13g2_o21ai_1 _10405_ (.B1(_04495_),
    .Y(_04496_),
    .A1(net2542),
    .A2(_01551_));
 sg13g2_o21ai_1 _10406_ (.B1(_04496_),
    .Y(_00787_),
    .A1(net2180),
    .A2(_04494_));
 sg13g2_a21oi_1 _10407_ (.A1(net858),
    .A2(_04492_),
    .Y(_04497_),
    .B1(net851));
 sg13g2_nand3_1 _10408_ (.B(net851),
    .C(_04492_),
    .A(net858),
    .Y(_04498_));
 sg13g2_nand2_1 _10409_ (.Y(_04499_),
    .A(net2167),
    .B(_04498_));
 sg13g2_a21oi_1 _10410_ (.A1(net2541),
    .A2(_03191_),
    .Y(_04500_),
    .B1(net2189));
 sg13g2_o21ai_1 _10411_ (.B1(_04500_),
    .Y(_04501_),
    .A1(net2541),
    .A2(_03193_));
 sg13g2_o21ai_1 _10412_ (.B1(_04501_),
    .Y(_00788_),
    .A1(_04497_),
    .A2(_04499_));
 sg13g2_nor2_1 _10413_ (.A(_00956_),
    .B(_04498_),
    .Y(_04502_));
 sg13g2_xnor2_1 _10414_ (.Y(_04503_),
    .A(_00956_),
    .B(_04498_));
 sg13g2_o21ai_1 _10415_ (.B1(net2176),
    .Y(_04504_),
    .A1(net2541),
    .A2(_03268_));
 sg13g2_a21o_1 _10416_ (.A2(_03265_),
    .A1(net2542),
    .B1(_04504_),
    .X(_04505_));
 sg13g2_o21ai_1 _10417_ (.B1(_04505_),
    .Y(_00789_),
    .A1(net2181),
    .A2(_04503_));
 sg13g2_and2_1 _10418_ (.A(net841),
    .B(_04502_),
    .X(_04506_));
 sg13g2_nor2_1 _10419_ (.A(net2181),
    .B(_04506_),
    .Y(_04507_));
 sg13g2_o21ai_1 _10420_ (.B1(_04507_),
    .Y(_04508_),
    .A1(net841),
    .A2(_04502_));
 sg13g2_nand2_1 _10421_ (.Y(_04509_),
    .A(net2542),
    .B(_03230_));
 sg13g2_a21oi_1 _10422_ (.A1(net2615),
    .A2(_03232_),
    .Y(_04510_),
    .B1(net2189));
 sg13g2_nand2_1 _10423_ (.Y(_04511_),
    .A(_04509_),
    .B(_04510_));
 sg13g2_nand2_1 _10424_ (.Y(_00790_),
    .A(_04508_),
    .B(_04511_));
 sg13g2_a21oi_1 _10425_ (.A1(net2614),
    .A2(_03155_),
    .Y(_04512_),
    .B1(net2189));
 sg13g2_o21ai_1 _10426_ (.B1(_04512_),
    .Y(_04513_),
    .A1(net2614),
    .A2(_03150_));
 sg13g2_xnor2_1 _10427_ (.Y(_04514_),
    .A(net857),
    .B(_04506_));
 sg13g2_o21ai_1 _10428_ (.B1(_04513_),
    .Y(_00791_),
    .A1(net2181),
    .A2(_04514_));
 sg13g2_and2_1 _10429_ (.A(net2543),
    .B(_03112_),
    .X(_04515_));
 sg13g2_a21oi_1 _10430_ (.A1(net2614),
    .A2(_03116_),
    .Y(_04516_),
    .B1(_04515_));
 sg13g2_a21oi_1 _10431_ (.A1(net857),
    .A2(_04506_),
    .Y(_04517_),
    .B1(net837));
 sg13g2_and3_1 _10432_ (.X(_04518_),
    .A(net857),
    .B(net837),
    .C(_04506_));
 sg13g2_nor3_1 _10433_ (.A(net2181),
    .B(_04517_),
    .C(_04518_),
    .Y(_04519_));
 sg13g2_a21o_1 _10434_ (.A2(_04516_),
    .A1(net2176),
    .B1(_04519_),
    .X(_00792_));
 sg13g2_a21oi_1 _10435_ (.A1(net2543),
    .A2(_03066_),
    .Y(_04520_),
    .B1(net2189));
 sg13g2_o21ai_1 _10436_ (.B1(_04520_),
    .Y(_04521_),
    .A1(net2544),
    .A2(_03070_));
 sg13g2_and2_1 _10437_ (.A(net846),
    .B(_04518_),
    .X(_04522_));
 sg13g2_o21ai_1 _10438_ (.B1(net2167),
    .Y(_04523_),
    .A1(net846),
    .A2(_04518_));
 sg13g2_o21ai_1 _10439_ (.B1(_04521_),
    .Y(_00793_),
    .A1(_04522_),
    .A2(_04523_));
 sg13g2_nand2_1 _10440_ (.Y(_04524_),
    .A(net2545),
    .B(_02995_));
 sg13g2_a21oi_1 _10441_ (.A1(net2614),
    .A2(_02997_),
    .Y(_04525_),
    .B1(net2189));
 sg13g2_nand2_1 _10442_ (.Y(_04526_),
    .A(_04524_),
    .B(_04525_));
 sg13g2_and2_1 _10443_ (.A(net845),
    .B(_04522_),
    .X(_04527_));
 sg13g2_o21ai_1 _10444_ (.B1(net2167),
    .Y(_04528_),
    .A1(net845),
    .A2(_04522_));
 sg13g2_o21ai_1 _10445_ (.B1(_04526_),
    .Y(_00794_),
    .A1(_04527_),
    .A2(_04528_));
 sg13g2_and2_1 _10446_ (.A(net2545),
    .B(_03035_),
    .X(_04529_));
 sg13g2_o21ai_1 _10447_ (.B1(net2176),
    .Y(_04530_),
    .A1(net2545),
    .A2(_03037_));
 sg13g2_and2_1 _10448_ (.A(net842),
    .B(_04527_),
    .X(_04531_));
 sg13g2_nor2_1 _10449_ (.A(net2180),
    .B(_04531_),
    .Y(_04532_));
 sg13g2_o21ai_1 _10450_ (.B1(_04532_),
    .Y(_04533_),
    .A1(net842),
    .A2(_04527_));
 sg13g2_o21ai_1 _10451_ (.B1(_04533_),
    .Y(_00795_),
    .A1(_04529_),
    .A2(_04530_));
 sg13g2_and2_1 _10452_ (.A(net2545),
    .B(_02946_),
    .X(_04534_));
 sg13g2_o21ai_1 _10453_ (.B1(net2176),
    .Y(_04535_),
    .A1(net2545),
    .A2(_02949_));
 sg13g2_and2_1 _10454_ (.A(net850),
    .B(_04531_),
    .X(_04536_));
 sg13g2_nor2_1 _10455_ (.A(net2182),
    .B(_04536_),
    .Y(_04537_));
 sg13g2_o21ai_1 _10456_ (.B1(_04537_),
    .Y(_04538_),
    .A1(net850),
    .A2(_04531_));
 sg13g2_o21ai_1 _10457_ (.B1(_04538_),
    .Y(_00796_),
    .A1(_04534_),
    .A2(_04535_));
 sg13g2_nand2_1 _10458_ (.Y(_04539_),
    .A(net2546),
    .B(_02898_));
 sg13g2_o21ai_1 _10459_ (.B1(_04539_),
    .Y(_04540_),
    .A1(net2546),
    .A2(_02900_));
 sg13g2_and2_1 _10460_ (.A(net848),
    .B(_04536_),
    .X(_04541_));
 sg13g2_nor2_1 _10461_ (.A(net2182),
    .B(_04541_),
    .Y(_04542_));
 sg13g2_o21ai_1 _10462_ (.B1(_04542_),
    .Y(_04543_),
    .A1(net848),
    .A2(_04536_));
 sg13g2_o21ai_1 _10463_ (.B1(_04543_),
    .Y(_00797_),
    .A1(net2190),
    .A2(_04540_));
 sg13g2_nand2_1 _10464_ (.Y(_04544_),
    .A(net2546),
    .B(_02852_));
 sg13g2_a21oi_1 _10465_ (.A1(net2618),
    .A2(_02860_),
    .Y(_04545_),
    .B1(net2190));
 sg13g2_nand2_1 _10466_ (.Y(_04546_),
    .A(_04544_),
    .B(_04545_));
 sg13g2_and2_1 _10467_ (.A(net839),
    .B(_04541_),
    .X(_04547_));
 sg13g2_o21ai_1 _10468_ (.B1(net2168),
    .Y(_04548_),
    .A1(net839),
    .A2(_04541_));
 sg13g2_o21ai_1 _10469_ (.B1(_04546_),
    .Y(_00798_),
    .A1(_04547_),
    .A2(_04548_));
 sg13g2_nand2_1 _10470_ (.Y(_04549_),
    .A(net2546),
    .B(_03357_));
 sg13g2_o21ai_1 _10471_ (.B1(_04549_),
    .Y(_04550_),
    .A1(net2546),
    .A2(_03363_));
 sg13g2_and2_1 _10472_ (.A(net1476),
    .B(_04547_),
    .X(_04551_));
 sg13g2_nor2_1 _10473_ (.A(net2182),
    .B(_04551_),
    .Y(_04552_));
 sg13g2_o21ai_1 _10474_ (.B1(_04552_),
    .Y(_04553_),
    .A1(net843),
    .A2(_04547_));
 sg13g2_o21ai_1 _10475_ (.B1(_04553_),
    .Y(_00799_),
    .A1(net2190),
    .A2(_04550_));
 sg13g2_nand2_1 _10476_ (.Y(_04554_),
    .A(net2548),
    .B(_03319_));
 sg13g2_a21oi_1 _10477_ (.A1(net2618),
    .A2(_03323_),
    .Y(_04555_),
    .B1(net2190));
 sg13g2_o21ai_1 _10478_ (.B1(net2167),
    .Y(_04556_),
    .A1(net855),
    .A2(_04551_));
 sg13g2_a21oi_1 _10479_ (.A1(net855),
    .A2(_04551_),
    .Y(_04557_),
    .B1(_04556_));
 sg13g2_a21o_1 _10480_ (.A2(_04555_),
    .A1(_04554_),
    .B1(_04557_),
    .X(_00800_));
 sg13g2_a21o_1 _10481_ (.A2(_02802_),
    .A1(net2619),
    .B1(net2190),
    .X(_04558_));
 sg13g2_a21oi_1 _10482_ (.A1(net2548),
    .A2(_02797_),
    .Y(_04559_),
    .B1(_04558_));
 sg13g2_nand3_1 _10483_ (.B(net847),
    .C(_04551_),
    .A(net855),
    .Y(_04560_));
 sg13g2_a21oi_1 _10484_ (.A1(net855),
    .A2(_04551_),
    .Y(_04561_),
    .B1(net847));
 sg13g2_nor2_1 _10485_ (.A(net2182),
    .B(_04561_),
    .Y(_04562_));
 sg13g2_a21o_1 _10486_ (.A2(_04562_),
    .A1(_04560_),
    .B1(_04559_),
    .X(_00801_));
 sg13g2_xor2_1 _10487_ (.B(_04560_),
    .A(net840),
    .X(_04563_));
 sg13g2_nand2_1 _10488_ (.Y(_04564_),
    .A(net2548),
    .B(_03409_));
 sg13g2_a21oi_1 _10489_ (.A1(net2619),
    .A2(_03413_),
    .Y(_04565_),
    .B1(net2189));
 sg13g2_nand2_1 _10490_ (.Y(_04566_),
    .A(_04564_),
    .B(_04565_));
 sg13g2_o21ai_1 _10491_ (.B1(_04566_),
    .Y(_00802_),
    .A1(net2182),
    .A2(_04563_));
 sg13g2_and2_1 _10492_ (.A(net2732),
    .B(net897),
    .X(_00835_));
 sg13g2_nor2_1 _10493_ (.A(net1202),
    .B(\ChiselTop.wild.tx.tx.bitsReg[1] ),
    .Y(_04567_));
 sg13g2_nor4_1 _10494_ (.A(net924),
    .B(\ChiselTop.wild.tx.tx.bitsReg[2] ),
    .C(\ChiselTop.wild.tx.tx.bitsReg[1] ),
    .D(\ChiselTop.wild.tx.tx.bitsReg[0] ),
    .Y(_04568_));
 sg13g2_nor2b_1 _10495_ (.A(_03501_),
    .B_N(_04568_),
    .Y(_04569_));
 sg13g2_nand2b_2 _10496_ (.Y(_04570_),
    .B(net1544),
    .A_N(_04569_));
 sg13g2_nor2_1 _10497_ (.A(\ChiselTop.wild.tx.buf_.io_out_valid ),
    .B(_03574_),
    .Y(_04571_));
 sg13g2_nand2_1 _10498_ (.Y(_04572_),
    .A(\ChiselTop.wild.cpu.io_dmem_rdAddress[2] ),
    .B(_04571_));
 sg13g2_or4_1 _10499_ (.A(\ChiselTop.wild.cpu.io_dmem_rdAddress[16] ),
    .B(\ChiselTop.wild.cpu.io_dmem_rdAddress[3] ),
    .C(_04135_),
    .D(_04572_),
    .X(_04573_));
 sg13g2_o21ai_1 _10500_ (.B1(_04570_),
    .Y(_04574_),
    .A1(_03576_),
    .A2(_04573_));
 sg13g2_and2_1 _10501_ (.A(net2734),
    .B(_04574_),
    .X(_00836_));
 sg13g2_nor2b_1 _10502_ (.A(\ChiselTop.wild.tx.buf_.io_out_valid ),
    .B_N(_04568_),
    .Y(_04575_));
 sg13g2_nor3_2 _10503_ (.A(net1448),
    .B(_03501_),
    .C(_04575_),
    .Y(_04576_));
 sg13g2_a21oi_1 _10504_ (.A1(net1448),
    .A2(_03501_),
    .Y(_04577_),
    .B1(_04576_));
 sg13g2_nor2_1 _10505_ (.A(net2726),
    .B(net1449),
    .Y(_00837_));
 sg13g2_nand2b_1 _10506_ (.Y(_04578_),
    .B(_04576_),
    .A_N(net1427));
 sg13g2_o21ai_1 _10507_ (.B1(net1427),
    .Y(_04579_),
    .A1(\ChiselTop.wild.tx.tx.bitsReg[0] ),
    .A2(_03501_));
 sg13g2_a21oi_1 _10508_ (.A1(_04578_),
    .A2(net1428),
    .Y(_00838_),
    .B1(net2726));
 sg13g2_nand2_1 _10509_ (.Y(_04580_),
    .A(_04567_),
    .B(_04576_));
 sg13g2_a22oi_1 _10510_ (.Y(_04581_),
    .B1(_04578_),
    .B2(net1202),
    .A2(_04576_),
    .A1(_04567_));
 sg13g2_a21oi_1 _10511_ (.A1(\ChiselTop.wild.tx.buf_.io_out_valid ),
    .A2(_04569_),
    .Y(_04582_),
    .B1(net2726));
 sg13g2_nor2b_1 _10512_ (.A(net1203),
    .B_N(_04582_),
    .Y(_00839_));
 sg13g2_a22oi_1 _10513_ (.Y(_04583_),
    .B1(_04580_),
    .B2(net924),
    .A2(_04569_),
    .A1(\ChiselTop.wild.tx.buf_.io_out_valid ));
 sg13g2_nor2_1 _10514_ (.A(net2726),
    .B(net925),
    .Y(_00840_));
 sg13g2_and4_1 _10515_ (.A(net854),
    .B(net2192),
    .C(net2448),
    .D(_01811_),
    .X(_04584_));
 sg13g2_nor3_2 _10516_ (.A(net1501),
    .B(\ChiselTop.wild.rx.cntReg[1] ),
    .C(\ChiselTop.wild.rx.cntReg[0] ),
    .Y(_04585_));
 sg13g2_nor2b_1 _10517_ (.A(\ChiselTop.wild.rx.cntReg[3] ),
    .B_N(_04585_),
    .Y(_04586_));
 sg13g2_nand2b_2 _10518_ (.Y(_04587_),
    .B(_04586_),
    .A_N(net1225));
 sg13g2_nor3_2 _10519_ (.A(net1526),
    .B(net1514),
    .C(_04587_),
    .Y(_04588_));
 sg13g2_nand2b_2 _10520_ (.Y(_04589_),
    .B(_04588_),
    .A_N(net1159));
 sg13g2_nor2_1 _10521_ (.A(net1406),
    .B(_04589_),
    .Y(_04590_));
 sg13g2_nor3_2 _10522_ (.A(net1489),
    .B(net1406),
    .C(_04589_),
    .Y(_04591_));
 sg13g2_nand2b_2 _10523_ (.Y(_04592_),
    .B(_04591_),
    .A_N(net1175));
 sg13g2_nor3_2 _10524_ (.A(net1505),
    .B(net1466),
    .C(_04592_),
    .Y(_04593_));
 sg13g2_nand2b_2 _10525_ (.Y(_04594_),
    .B(_04593_),
    .A_N(net1057));
 sg13g2_nor3_1 _10526_ (.A(net1368),
    .B(\ChiselTop.wild.rx.cntReg[14] ),
    .C(_04594_),
    .Y(_04595_));
 sg13g2_nor2b_2 _10527_ (.A(net1411),
    .B_N(_04595_),
    .Y(_04596_));
 sg13g2_nand2b_2 _10528_ (.Y(_04597_),
    .B(_04596_),
    .A_N(net1307));
 sg13g2_nor3_2 _10529_ (.A(net1480),
    .B(\ChiselTop.wild.rx.cntReg[18] ),
    .C(_04597_),
    .Y(_04598_));
 sg13g2_or3_1 _10530_ (.A(\ChiselTop.wild.rx.cntReg[19] ),
    .B(\ChiselTop.wild.rx.cntReg[18] ),
    .C(_04597_),
    .X(_04599_));
 sg13g2_nor4_1 _10531_ (.A(net1287),
    .B(net1358),
    .C(\ChiselTop.wild.rx.bitsReg[1] ),
    .D(_00902_),
    .Y(_04600_));
 sg13g2_a21oi_1 _10532_ (.A1(net2166),
    .A2(net1359),
    .Y(_04601_),
    .B1(net854));
 sg13g2_nor3_1 _10533_ (.A(net2727),
    .B(_04584_),
    .C(_04601_),
    .Y(_00841_));
 sg13g2_nor2_1 _10534_ (.A(\ChiselTop.wild.rx.bitsReg[1] ),
    .B(net1512),
    .Y(_04602_));
 sg13g2_nor4_2 _10535_ (.A(net1287),
    .B(\ChiselTop.wild.rx.bitsReg[2] ),
    .C(\ChiselTop.wild.rx.bitsReg[1] ),
    .Y(_04603_),
    .D(\ChiselTop.wild.rx.bitsReg[0] ));
 sg13g2_nand2b_1 _10536_ (.Y(_04604_),
    .B(net2166),
    .A_N(_04603_));
 sg13g2_nor2_1 _10537_ (.A(net1441),
    .B(net2159),
    .Y(_04605_));
 sg13g2_nand2_1 _10538_ (.Y(_04606_),
    .A(net2744),
    .B(_04599_));
 sg13g2_inv_1 _10539_ (.Y(_04607_),
    .A(net2155));
 sg13g2_a22oi_1 _10540_ (.Y(_04608_),
    .B1(_04607_),
    .B2(net1441),
    .A2(_04605_),
    .A1(net2741));
 sg13g2_inv_1 _10541_ (.Y(_00842_),
    .A(_04608_));
 sg13g2_o21ai_1 _10542_ (.B1(net2741),
    .Y(_04609_),
    .A1(net1388),
    .A2(_04605_));
 sg13g2_a21oi_1 _10543_ (.A1(net1388),
    .A2(_04605_),
    .Y(_00843_),
    .B1(_04609_));
 sg13g2_nand2b_1 _10544_ (.Y(_04610_),
    .B(\ChiselTop.wild.rx.falling_REG ),
    .A_N(\ChiselTop.wild.rx._shiftReg_T_1[7] ));
 sg13g2_nor2_1 _10545_ (.A(_04599_),
    .B(_04610_),
    .Y(_04611_));
 sg13g2_o21ai_1 _10546_ (.B1(net1358),
    .Y(_04612_),
    .A1(_04599_),
    .A2(_04610_));
 sg13g2_xnor2_1 _10547_ (.Y(_04613_),
    .A(net1358),
    .B(net1513));
 sg13g2_a221oi_1 _10548_ (.B2(net2166),
    .C1(net2726),
    .B1(_04613_),
    .A1(net2159),
    .Y(_00844_),
    .A2(_04612_));
 sg13g2_nand3b_1 _10549_ (.B(net2166),
    .C(_04602_),
    .Y(_04614_),
    .A_N(\ChiselTop.wild.rx.bitsReg[2] ));
 sg13g2_a22oi_1 _10550_ (.Y(_04615_),
    .B1(_04614_),
    .B2(net1287),
    .A2(_04611_),
    .A1(_04603_));
 sg13g2_nor2_1 _10551_ (.A(net2726),
    .B(net1288),
    .Y(_00845_));
 sg13g2_o21ai_1 _10552_ (.B1(net2733),
    .Y(_04616_),
    .A1(\ChiselTop.wild.rx._shiftReg_T_1[0] ),
    .A2(net2157));
 sg13g2_a21oi_1 _10553_ (.A1(_00901_),
    .A2(net2157),
    .Y(_00846_),
    .B1(_04616_));
 sg13g2_o21ai_1 _10554_ (.B1(net2733),
    .Y(_04617_),
    .A1(net1276),
    .A2(net2157));
 sg13g2_a21oi_1 _10555_ (.A1(_00900_),
    .A2(net2157),
    .Y(_00847_),
    .B1(_04617_));
 sg13g2_o21ai_1 _10556_ (.B1(net2740),
    .Y(_04618_),
    .A1(\ChiselTop.wild.rx._shiftReg_T_1[2] ),
    .A2(net2157));
 sg13g2_a21oi_1 _10557_ (.A1(_00899_),
    .A2(net2157),
    .Y(_00848_),
    .B1(_04618_));
 sg13g2_o21ai_1 _10558_ (.B1(net2740),
    .Y(_04619_),
    .A1(\ChiselTop.wild.rx._shiftReg_T_1[3] ),
    .A2(net2158));
 sg13g2_a21oi_1 _10559_ (.A1(_00898_),
    .A2(net2159),
    .Y(_00849_),
    .B1(_04619_));
 sg13g2_o21ai_1 _10560_ (.B1(net2740),
    .Y(_04620_),
    .A1(net1387),
    .A2(net2157));
 sg13g2_a21oi_1 _10561_ (.A1(_00897_),
    .A2(net2157),
    .Y(_00850_),
    .B1(_04620_));
 sg13g2_o21ai_1 _10562_ (.B1(net2740),
    .Y(_04621_),
    .A1(net1185),
    .A2(net2158));
 sg13g2_a21oi_1 _10563_ (.A1(_00896_),
    .A2(net2158),
    .Y(_00851_),
    .B1(_04621_));
 sg13g2_o21ai_1 _10564_ (.B1(net2740),
    .Y(_04622_),
    .A1(\ChiselTop.wild.rx._shiftReg_T_1[6] ),
    .A2(net2158));
 sg13g2_a21oi_1 _10565_ (.A1(_00895_),
    .A2(net2158),
    .Y(_00852_),
    .B1(_04622_));
 sg13g2_o21ai_1 _10566_ (.B1(net2740),
    .Y(_04623_),
    .A1(net864),
    .A2(net2158));
 sg13g2_a21oi_1 _10567_ (.A1(_00894_),
    .A2(net2158),
    .Y(_00853_),
    .B1(_04623_));
 sg13g2_and2_1 _10568_ (.A(net2729),
    .B(net2),
    .X(_00854_));
 sg13g2_nand2_1 _10569_ (.Y(_04624_),
    .A(\ChiselTop.wild.cpu.decOut_opcode[5] ),
    .B(_01806_));
 sg13g2_o21ai_1 _10570_ (.B1(net2522),
    .Y(_04625_),
    .A1(net2550),
    .A2(_04624_));
 sg13g2_o21ai_1 _10571_ (.B1(net2731),
    .Y(_04626_),
    .A1(_01813_),
    .A2(_04625_));
 sg13g2_inv_1 _10572_ (.Y(_00855_),
    .A(_04626_));
 sg13g2_and2_2 _10573_ (.A(net2741),
    .B(net2159),
    .X(_04627_));
 sg13g2_o21ai_1 _10574_ (.B1(_04627_),
    .Y(_00856_),
    .A1(_00957_),
    .A2(_04598_));
 sg13g2_xor2_1 _10575_ (.B(net1507),
    .A(\ChiselTop.wild.rx.cntReg[1] ),
    .X(_04628_));
 sg13g2_o21ai_1 _10576_ (.B1(_04627_),
    .Y(_00857_),
    .A1(_04598_),
    .A2(net1508));
 sg13g2_nand3_1 _10577_ (.B(_04603_),
    .C(_04610_),
    .A(net2166),
    .Y(_04629_));
 sg13g2_inv_1 _10578_ (.Y(_04630_),
    .A(_04629_));
 sg13g2_nand2_1 _10579_ (.Y(_04631_),
    .A(_04627_),
    .B(_04629_));
 sg13g2_o21ai_1 _10580_ (.B1(net1501),
    .Y(_04632_),
    .A1(\ChiselTop.wild.rx.cntReg[1] ),
    .A2(\ChiselTop.wild.rx.cntReg[0] ));
 sg13g2_nor2b_1 _10581_ (.A(net1502),
    .B_N(_04632_),
    .Y(_04633_));
 sg13g2_nor2_1 _10582_ (.A(_04631_),
    .B(net1503),
    .Y(_00858_));
 sg13g2_xnor2_1 _10583_ (.Y(_04634_),
    .A(net1374),
    .B(_04585_));
 sg13g2_nor2_1 _10584_ (.A(net2155),
    .B(net1375),
    .Y(_00859_));
 sg13g2_nand2b_1 _10585_ (.Y(_04635_),
    .B(net1225),
    .A_N(_04586_));
 sg13g2_a21oi_1 _10586_ (.A1(_04587_),
    .A2(net1226),
    .Y(_00860_),
    .B1(_04631_));
 sg13g2_xor2_1 _10587_ (.B(_04587_),
    .A(net1514),
    .X(_04636_));
 sg13g2_o21ai_1 _10588_ (.B1(_04627_),
    .Y(_00861_),
    .A1(net2166),
    .A2(net1515));
 sg13g2_o21ai_1 _10589_ (.B1(net1526),
    .Y(_04637_),
    .A1(\ChiselTop.wild.rx.cntReg[5] ),
    .A2(_04587_));
 sg13g2_nor2b_1 _10590_ (.A(_04588_),
    .B_N(_04637_),
    .Y(_04638_));
 sg13g2_o21ai_1 _10591_ (.B1(_04627_),
    .Y(_00862_),
    .A1(net2166),
    .A2(net1527));
 sg13g2_nand2b_1 _10592_ (.Y(_04639_),
    .B(net1159),
    .A_N(_04588_));
 sg13g2_a21oi_1 _10593_ (.A1(_04589_),
    .A2(net1160),
    .Y(_00863_),
    .B1(net2155));
 sg13g2_o21ai_1 _10594_ (.B1(net1406),
    .Y(_04640_),
    .A1(_04589_),
    .A2(_04630_));
 sg13g2_a21oi_1 _10595_ (.A1(_04590_),
    .A2(_04629_),
    .Y(_04641_),
    .B1(net2726));
 sg13g2_nand2_1 _10596_ (.Y(_00864_),
    .A(net1407),
    .B(_04641_));
 sg13g2_xnor2_1 _10597_ (.Y(_04642_),
    .A(net1489),
    .B(_04590_));
 sg13g2_o21ai_1 _10598_ (.B1(_04627_),
    .Y(_00865_),
    .A1(net2166),
    .A2(_04642_));
 sg13g2_nand2b_1 _10599_ (.Y(_04643_),
    .B(net1175),
    .A_N(_04591_));
 sg13g2_a21oi_1 _10600_ (.A1(_04592_),
    .A2(net1176),
    .Y(_00866_),
    .B1(_04631_));
 sg13g2_xor2_1 _10601_ (.B(_04592_),
    .A(net1466),
    .X(_04644_));
 sg13g2_nor2_1 _10602_ (.A(net2156),
    .B(net1467),
    .Y(_00867_));
 sg13g2_o21ai_1 _10603_ (.B1(net1505),
    .Y(_04645_),
    .A1(net1466),
    .A2(_04592_));
 sg13g2_nor2b_1 _10604_ (.A(_04593_),
    .B_N(_04645_),
    .Y(_04646_));
 sg13g2_nor2_1 _10605_ (.A(net2156),
    .B(_04646_),
    .Y(_00868_));
 sg13g2_nand2b_1 _10606_ (.Y(_04647_),
    .B(net1057),
    .A_N(_04593_));
 sg13g2_a21oi_1 _10607_ (.A1(_04594_),
    .A2(net1058),
    .Y(_00869_),
    .B1(net2156));
 sg13g2_nor2_1 _10608_ (.A(_00958_),
    .B(_04594_),
    .Y(_04648_));
 sg13g2_xnor2_1 _10609_ (.Y(_04649_),
    .A(net939),
    .B(_04594_));
 sg13g2_nor2_1 _10610_ (.A(net2156),
    .B(net940),
    .Y(_00870_));
 sg13g2_xnor2_1 _10611_ (.Y(_04650_),
    .A(net1368),
    .B(_04648_));
 sg13g2_nor2_1 _10612_ (.A(net2155),
    .B(net1369),
    .Y(_00871_));
 sg13g2_xnor2_1 _10613_ (.Y(_04651_),
    .A(net1411),
    .B(_04595_));
 sg13g2_nor2_1 _10614_ (.A(net2155),
    .B(net1412),
    .Y(_00872_));
 sg13g2_nand2b_1 _10615_ (.Y(_04652_),
    .B(net1307),
    .A_N(_04596_));
 sg13g2_a21oi_1 _10616_ (.A1(_04597_),
    .A2(net1308),
    .Y(_00873_),
    .B1(net2155));
 sg13g2_nand3b_1 _10617_ (.B(net1022),
    .C(_04596_),
    .Y(_04653_),
    .A_N(net1307));
 sg13g2_xnor2_1 _10618_ (.Y(_04654_),
    .A(net1022),
    .B(_04597_));
 sg13g2_nor2_1 _10619_ (.A(net2155),
    .B(net1023),
    .Y(_00874_));
 sg13g2_xor2_1 _10620_ (.B(_04653_),
    .A(net1480),
    .X(_04655_));
 sg13g2_nor2_1 _10621_ (.A(net2155),
    .B(_04655_),
    .Y(_00875_));
 sg13g2_nand3b_1 _10622_ (.B(net2553),
    .C(_03463_),
    .Y(_04656_),
    .A_N(net2552));
 sg13g2_and2_1 _10623_ (.A(_03474_),
    .B(_04656_),
    .X(_04657_));
 sg13g2_a21oi_1 _10624_ (.A1(_03469_),
    .A2(_04657_),
    .Y(_00880_),
    .B1(net2178));
 sg13g2_nor2_1 _10625_ (.A(_00195_),
    .B(_00880_),
    .Y(_00876_));
 sg13g2_nor2b_1 _10626_ (.A(_03473_),
    .B_N(_03569_),
    .Y(_04658_));
 sg13g2_a21oi_1 _10627_ (.A1(_04657_),
    .A2(_04658_),
    .Y(_00877_),
    .B1(net2178));
 sg13g2_nor3_1 _10628_ (.A(\ChiselTop.wild.cpu.io_imem_data[22] ),
    .B(_03486_),
    .C(net2177),
    .Y(_00878_));
 sg13g2_nor2_1 _10629_ (.A(net2177),
    .B(_04657_),
    .Y(_00879_));
 sg13g2_nor2b_1 _10630_ (.A(net2177),
    .B_N(\ChiselTop.wild.cpu.io_imem_data[15] ),
    .Y(_00881_));
 sg13g2_and2_1 _10631_ (.A(\ChiselTop.wild.cpu.io_imem_data[16] ),
    .B(net2169),
    .X(_00882_));
 sg13g2_nor2b_1 _10632_ (.A(net2177),
    .B_N(\ChiselTop.wild.cpu.io_imem_data[20] ),
    .Y(_00884_));
 sg13g2_nor2_1 _10633_ (.A(_03485_),
    .B(net2177),
    .Y(_00886_));
 sg13g2_nor2b_1 _10634_ (.A(net2177),
    .B_N(\ChiselTop.wild.cpu.io_imem_data[21] ),
    .Y(_00885_));
 sg13g2_a21oi_1 _10635_ (.A1(_03468_),
    .A2(_03478_),
    .Y(_00887_),
    .B1(net2178));
 sg13g2_nor2b_1 _10636_ (.A(net2177),
    .B_N(_03487_),
    .Y(_00888_));
 sg13g2_nor2b_1 _10637_ (.A(_03479_),
    .B_N(_00888_),
    .Y(_00889_));
 sg13g2_o21ai_1 _10638_ (.B1(net2176),
    .Y(_04659_),
    .A1(net2616),
    .A2(_02152_));
 sg13g2_a21oi_1 _10639_ (.A1(net2620),
    .A2(_02165_),
    .Y(_04660_),
    .B1(_04659_));
 sg13g2_a21o_1 _10640_ (.A2(net2168),
    .A1(net829),
    .B1(_04660_),
    .X(_00890_));
 sg13g2_o21ai_1 _10641_ (.B1(net2176),
    .Y(_04661_),
    .A1(net2616),
    .A2(_01969_));
 sg13g2_a21oi_1 _10642_ (.A1(net2616),
    .A2(_01982_),
    .Y(_04662_),
    .B1(_04661_));
 sg13g2_a21o_1 _10643_ (.A2(net2168),
    .A1(net833),
    .B1(_04662_),
    .X(_00891_));
 sg13g2_o21ai_1 _10644_ (.B1(net2729),
    .Y(_04663_),
    .A1(\ChiselTop.ledReg ),
    .A2(_04239_));
 sg13g2_a21oi_1 _10645_ (.A1(_00893_),
    .A2(_04239_),
    .Y(_00892_),
    .B1(_04663_));
 sg13g2_nor2_1 _10646_ (.A(net1454),
    .B(_03528_),
    .Y(_00193_));
 sg13g2_buf_1 _10647_ (.A(net910),
    .X(_00803_));
 sg13g2_buf_1 _10648_ (.A(net932),
    .X(_00804_));
 sg13g2_buf_1 _10649_ (.A(net934),
    .X(_00805_));
 sg13g2_buf_1 _10650_ (.A(net908),
    .X(_00806_));
 sg13g2_buf_1 _10651_ (.A(net909),
    .X(_00807_));
 sg13g2_buf_1 _10652_ (.A(net923),
    .X(_00808_));
 sg13g2_buf_1 _10653_ (.A(net922),
    .X(_00809_));
 sg13g2_buf_1 _10654_ (.A(net911),
    .X(_00810_));
 sg13g2_buf_1 _10655_ (.A(net906),
    .X(_00811_));
 sg13g2_buf_1 _10656_ (.A(net919),
    .X(_00812_));
 sg13g2_buf_1 _10657_ (.A(net917),
    .X(_00813_));
 sg13g2_buf_1 _10658_ (.A(net928),
    .X(_00814_));
 sg13g2_buf_1 _10659_ (.A(net929),
    .X(_00815_));
 sg13g2_buf_1 _10660_ (.A(net907),
    .X(_00816_));
 sg13g2_buf_1 _10661_ (.A(net933),
    .X(_00817_));
 sg13g2_buf_1 _10662_ (.A(net916),
    .X(_00818_));
 sg13g2_buf_1 _10663_ (.A(net920),
    .X(_00819_));
 sg13g2_buf_1 _10664_ (.A(net941),
    .X(_00820_));
 sg13g2_buf_1 _10665_ (.A(net935),
    .X(_00821_));
 sg13g2_buf_1 _10666_ (.A(net914),
    .X(_00822_));
 sg13g2_buf_1 _10667_ (.A(net912),
    .X(_00823_));
 sg13g2_buf_1 _10668_ (.A(net913),
    .X(_00824_));
 sg13g2_buf_1 _10669_ (.A(net921),
    .X(_00825_));
 sg13g2_buf_1 _10670_ (.A(net927),
    .X(_00826_));
 sg13g2_buf_1 _10671_ (.A(net938),
    .X(_00827_));
 sg13g2_buf_1 _10672_ (.A(net905),
    .X(_00828_));
 sg13g2_buf_1 _10673_ (.A(net936),
    .X(_00829_));
 sg13g2_buf_1 _10674_ (.A(net915),
    .X(_00830_));
 sg13g2_buf_1 _10675_ (.A(net942),
    .X(_00831_));
 sg13g2_buf_1 _10676_ (.A(net926),
    .X(_00832_));
 sg13g2_buf_1 _10677_ (.A(net918),
    .X(_00833_));
 sg13g2_buf_1 _10678_ (.A(net904),
    .X(_00834_));
 sg13g2_nor2_1 _10679_ (.A(_03465_),
    .B(net2177),
    .Y(_00883_));
 sg13g2_dfrbp_1 _10680_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net70),
    .D(_00143_),
    .Q_N(_05269_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[2] ));
 sg13g2_dfrbp_1 _10681_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net65),
    .D(_00144_),
    .Q_N(_05268_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[3] ));
 sg13g2_dfrbp_1 _10682_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net64),
    .D(_00145_),
    .Q_N(_05267_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[4] ));
 sg13g2_dfrbp_1 _10683_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net63),
    .D(net1080),
    .Q_N(_05266_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[7] ));
 sg13g2_dfrbp_1 _10684_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net62),
    .D(net1108),
    .Q_N(_05265_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[10] ));
 sg13g2_dfrbp_1 _10685_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net61),
    .D(_00148_),
    .Q_N(_05264_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[11] ));
 sg13g2_dfrbp_1 _10686_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net60),
    .D(_00149_),
    .Q_N(_05263_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[12] ));
 sg13g2_dfrbp_1 _10687_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net59),
    .D(net1140),
    .Q_N(_05262_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[13] ));
 sg13g2_dfrbp_1 _10688_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net58),
    .D(_00151_),
    .Q_N(_05261_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[14] ));
 sg13g2_dfrbp_1 _10689_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net57),
    .D(_00152_),
    .Q_N(_05260_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[15] ));
 sg13g2_dfrbp_1 _10690_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net56),
    .D(net1044),
    .Q_N(_05259_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[16] ));
 sg13g2_dfrbp_1 _10691_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net55),
    .D(_00154_),
    .Q_N(_05258_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[17] ));
 sg13g2_dfrbp_1 _10692_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net54),
    .D(_00155_),
    .Q_N(_05257_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[18] ));
 sg13g2_dfrbp_1 _10693_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net53),
    .D(net931),
    .Q_N(_05256_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[19] ));
 sg13g2_dfrbp_1 _10694_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net52),
    .D(_00157_),
    .Q_N(_00123_),
    .Q(\ChiselTop.wild.cpu.decExReg_csrVal[1] ));
 sg13g2_dfrbp_1 _10695_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net51),
    .D(_00158_),
    .Q_N(_05255_),
    .Q(\ChiselTop.wild.cpu.decExReg_csrVal[2] ));
 sg13g2_dfrbp_1 _10696_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net50),
    .D(_00159_),
    .Q_N(_05254_),
    .Q(\ChiselTop.wild.cpu.regs[1][0] ));
 sg13g2_dfrbp_1 _10697_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net49),
    .D(_00160_),
    .Q_N(_05253_),
    .Q(\ChiselTop.wild.cpu.regs[1][1] ));
 sg13g2_dfrbp_1 _10698_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net48),
    .D(_00161_),
    .Q_N(_05252_),
    .Q(\ChiselTop.wild.cpu.regs[1][2] ));
 sg13g2_dfrbp_1 _10699_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net47),
    .D(_00162_),
    .Q_N(_05251_),
    .Q(\ChiselTop.wild.cpu.regs[1][3] ));
 sg13g2_dfrbp_1 _10700_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net46),
    .D(_00163_),
    .Q_N(_05250_),
    .Q(\ChiselTop.wild.cpu.regs[1][4] ));
 sg13g2_dfrbp_1 _10701_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net45),
    .D(_00164_),
    .Q_N(_05249_),
    .Q(\ChiselTop.wild.cpu.regs[1][5] ));
 sg13g2_dfrbp_1 _10702_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net44),
    .D(_00165_),
    .Q_N(_05248_),
    .Q(\ChiselTop.wild.cpu.regs[1][6] ));
 sg13g2_dfrbp_1 _10703_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net43),
    .D(_00166_),
    .Q_N(_05247_),
    .Q(\ChiselTop.wild.cpu.regs[1][7] ));
 sg13g2_dfrbp_1 _10704_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net42),
    .D(_00167_),
    .Q_N(_05246_),
    .Q(\ChiselTop.wild.cpu.regs[1][8] ));
 sg13g2_dfrbp_1 _10705_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net41),
    .D(_00168_),
    .Q_N(_05245_),
    .Q(\ChiselTop.wild.cpu.regs[1][9] ));
 sg13g2_dfrbp_1 _10706_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net40),
    .D(_00169_),
    .Q_N(_05244_),
    .Q(\ChiselTop.wild.cpu.regs[1][10] ));
 sg13g2_dfrbp_1 _10707_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net39),
    .D(_00170_),
    .Q_N(_05243_),
    .Q(\ChiselTop.wild.cpu.regs[1][11] ));
 sg13g2_dfrbp_1 _10708_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net38),
    .D(_00171_),
    .Q_N(_05242_),
    .Q(\ChiselTop.wild.cpu.regs[1][12] ));
 sg13g2_dfrbp_1 _10709_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net37),
    .D(_00172_),
    .Q_N(_05241_),
    .Q(\ChiselTop.wild.cpu.regs[1][13] ));
 sg13g2_dfrbp_1 _10710_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net36),
    .D(_00173_),
    .Q_N(_05240_),
    .Q(\ChiselTop.wild.cpu.regs[1][14] ));
 sg13g2_dfrbp_1 _10711_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net35),
    .D(_00174_),
    .Q_N(_05239_),
    .Q(\ChiselTop.wild.cpu.regs[1][15] ));
 sg13g2_dfrbp_1 _10712_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net34),
    .D(_00175_),
    .Q_N(_05238_),
    .Q(\ChiselTop.wild.cpu.regs[1][16] ));
 sg13g2_dfrbp_1 _10713_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net33),
    .D(_00176_),
    .Q_N(_05237_),
    .Q(\ChiselTop.wild.cpu.regs[1][17] ));
 sg13g2_dfrbp_1 _10714_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net32),
    .D(_00177_),
    .Q_N(_05236_),
    .Q(\ChiselTop.wild.cpu.regs[1][18] ));
 sg13g2_dfrbp_1 _10715_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net31),
    .D(_00178_),
    .Q_N(_05235_),
    .Q(\ChiselTop.wild.cpu.regs[1][19] ));
 sg13g2_dfrbp_1 _10716_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net30),
    .D(_00179_),
    .Q_N(_05234_),
    .Q(\ChiselTop.wild.cpu.regs[1][20] ));
 sg13g2_dfrbp_1 _10717_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net29),
    .D(_00180_),
    .Q_N(_05233_),
    .Q(\ChiselTop.wild.cpu.regs[1][21] ));
 sg13g2_dfrbp_1 _10718_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net28),
    .D(_00181_),
    .Q_N(_05232_),
    .Q(\ChiselTop.wild.cpu.regs[1][22] ));
 sg13g2_dfrbp_1 _10719_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net27),
    .D(_00182_),
    .Q_N(_05231_),
    .Q(\ChiselTop.wild.cpu.regs[1][23] ));
 sg13g2_dfrbp_1 _10720_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net26),
    .D(_00183_),
    .Q_N(_05230_),
    .Q(\ChiselTop.wild.cpu.regs[1][24] ));
 sg13g2_dfrbp_1 _10721_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net25),
    .D(_00184_),
    .Q_N(_05229_),
    .Q(\ChiselTop.wild.cpu.regs[1][25] ));
 sg13g2_dfrbp_1 _10722_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net24),
    .D(_00185_),
    .Q_N(_05228_),
    .Q(\ChiselTop.wild.cpu.regs[1][26] ));
 sg13g2_dfrbp_1 _10723_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net23),
    .D(_00186_),
    .Q_N(_05227_),
    .Q(\ChiselTop.wild.cpu.regs[1][27] ));
 sg13g2_dfrbp_1 _10724_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net22),
    .D(_00187_),
    .Q_N(_05226_),
    .Q(\ChiselTop.wild.cpu.regs[1][28] ));
 sg13g2_dfrbp_1 _10725_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net21),
    .D(_00188_),
    .Q_N(_05225_),
    .Q(\ChiselTop.wild.cpu.regs[1][29] ));
 sg13g2_dfrbp_1 _10726_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net20),
    .D(_00189_),
    .Q_N(_05224_),
    .Q(\ChiselTop.wild.cpu.regs[1][30] ));
 sg13g2_dfrbp_1 _10727_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net19),
    .D(_00190_),
    .Q_N(_05223_),
    .Q(\ChiselTop.wild.cpu.regs[1][31] ));
 sg13g2_dfrbp_1 _10728_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net71),
    .D(\ChiselTop.wild.cpu.io_imem_data[15] ),
    .Q_N(_05270_),
    .Q(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[0] ));
 sg13g2_dfrbp_1 _10729_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net433),
    .D(\ChiselTop.wild.cpu.io_imem_data[16] ),
    .Q_N(_05271_),
    .Q(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[1] ));
 sg13g2_dfrbp_1 _10730_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net825),
    .D(\ChiselTop.wild.cpu.io_imem_data[13] ),
    .Q_N(_00001_),
    .Q(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[2] ));
 sg13g2_dfrbp_1 _10731_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net824),
    .D(_00191_),
    .Q_N(_05222_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[1] ));
 sg13g2_dfrbp_1 _10732_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net823),
    .D(_00192_),
    .Q_N(_00066_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[2] ));
 sg13g2_dfrbp_1 _10733_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net822),
    .D(net1455),
    .Q_N(_05221_),
    .Q(\ChiselTop.wild.cpu.decExReg_csrVal[3] ));
 sg13g2_dfrbp_1 _10734_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net821),
    .D(_00194_),
    .Q_N(_05220_),
    .Q(\ChiselTop.wild.cpu._GEN_176[5] ));
 sg13g2_dfrbp_1 _10735_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net820),
    .D(_00195_),
    .Q_N(_00113_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[13] ));
 sg13g2_dfrbp_1 _10736_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net819),
    .D(net1536),
    .Q_N(_05219_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[1] ));
 sg13g2_dfrbp_1 _10737_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net818),
    .D(_00197_),
    .Q_N(_05218_),
    .Q(\ChiselTop.wild.cpu.decOut_opcode[5] ));
 sg13g2_dfrbp_1 _10738_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net816),
    .D(_00198_),
    .Q_N(_05217_),
    .Q(\ChiselTop.wild.dmem.MEM_2[0][0] ));
 sg13g2_dfrbp_1 _10739_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net815),
    .D(_00199_),
    .Q_N(_05216_),
    .Q(\ChiselTop.wild.dmem.MEM_2[0][1] ));
 sg13g2_dfrbp_1 _10740_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net814),
    .D(_00200_),
    .Q_N(_05215_),
    .Q(\ChiselTop.wild.dmem.MEM_2[0][2] ));
 sg13g2_dfrbp_1 _10741_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net813),
    .D(_00201_),
    .Q_N(_05214_),
    .Q(\ChiselTop.wild.dmem.MEM_2[0][3] ));
 sg13g2_dfrbp_1 _10742_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net812),
    .D(_00202_),
    .Q_N(_05213_),
    .Q(\ChiselTop.wild.dmem.MEM_2[0][4] ));
 sg13g2_dfrbp_1 _10743_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net811),
    .D(_00203_),
    .Q_N(_05212_),
    .Q(\ChiselTop.wild.dmem.MEM_2[0][5] ));
 sg13g2_dfrbp_1 _10744_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net810),
    .D(_00204_),
    .Q_N(_05211_),
    .Q(\ChiselTop.wild.dmem.MEM_2[0][6] ));
 sg13g2_dfrbp_1 _10745_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net809),
    .D(_00205_),
    .Q_N(_05210_),
    .Q(\ChiselTop.wild.dmem.MEM_2[0][7] ));
 sg13g2_dfrbp_1 _10746_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net808),
    .D(_00206_),
    .Q_N(_05209_),
    .Q(\ChiselTop.wild.dmem.MEM_1[0][0] ));
 sg13g2_dfrbp_1 _10747_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net807),
    .D(_00207_),
    .Q_N(_05208_),
    .Q(\ChiselTop.wild.dmem.MEM_1[0][1] ));
 sg13g2_dfrbp_1 _10748_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net806),
    .D(_00208_),
    .Q_N(_05207_),
    .Q(\ChiselTop.wild.dmem.MEM_1[0][2] ));
 sg13g2_dfrbp_1 _10749_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net805),
    .D(_00209_),
    .Q_N(_05206_),
    .Q(\ChiselTop.wild.dmem.MEM_1[0][3] ));
 sg13g2_dfrbp_1 _10750_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net804),
    .D(_00210_),
    .Q_N(_05205_),
    .Q(\ChiselTop.wild.dmem.MEM_1[0][4] ));
 sg13g2_dfrbp_1 _10751_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net803),
    .D(_00211_),
    .Q_N(_05204_),
    .Q(\ChiselTop.wild.dmem.MEM_1[0][5] ));
 sg13g2_dfrbp_1 _10752_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net802),
    .D(_00212_),
    .Q_N(_05203_),
    .Q(\ChiselTop.wild.dmem.MEM_1[0][6] ));
 sg13g2_dfrbp_1 _10753_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net801),
    .D(_00213_),
    .Q_N(_05202_),
    .Q(\ChiselTop.wild.dmem.MEM_1[0][7] ));
 sg13g2_dfrbp_1 _10754_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net800),
    .D(_00214_),
    .Q_N(_05201_),
    .Q(\ChiselTop.wild.dmem.MEM[0][0] ));
 sg13g2_dfrbp_1 _10755_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net799),
    .D(_00215_),
    .Q_N(_05200_),
    .Q(\ChiselTop.wild.dmem.MEM[0][1] ));
 sg13g2_dfrbp_1 _10756_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net798),
    .D(_00216_),
    .Q_N(_05199_),
    .Q(\ChiselTop.wild.dmem.MEM[0][2] ));
 sg13g2_dfrbp_1 _10757_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net797),
    .D(_00217_),
    .Q_N(_05198_),
    .Q(\ChiselTop.wild.dmem.MEM[0][3] ));
 sg13g2_dfrbp_1 _10758_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net796),
    .D(_00218_),
    .Q_N(_05197_),
    .Q(\ChiselTop.wild.dmem.MEM[0][4] ));
 sg13g2_dfrbp_1 _10759_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net795),
    .D(_00219_),
    .Q_N(_05196_),
    .Q(\ChiselTop.wild.dmem.MEM[0][5] ));
 sg13g2_dfrbp_1 _10760_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net794),
    .D(_00220_),
    .Q_N(_05195_),
    .Q(\ChiselTop.wild.dmem.MEM[0][6] ));
 sg13g2_dfrbp_1 _10761_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net793),
    .D(_00221_),
    .Q_N(_05194_),
    .Q(\ChiselTop.wild.dmem.MEM[0][7] ));
 sg13g2_dfrbp_1 _10762_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net792),
    .D(_00222_),
    .Q_N(_05193_),
    .Q(\ChiselTop.wild.cpu.regs[3][0] ));
 sg13g2_dfrbp_1 _10763_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net791),
    .D(_00223_),
    .Q_N(_05192_),
    .Q(\ChiselTop.wild.cpu.regs[3][1] ));
 sg13g2_dfrbp_1 _10764_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net790),
    .D(_00224_),
    .Q_N(_05191_),
    .Q(\ChiselTop.wild.cpu.regs[3][2] ));
 sg13g2_dfrbp_1 _10765_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net789),
    .D(_00225_),
    .Q_N(_05190_),
    .Q(\ChiselTop.wild.cpu.regs[3][3] ));
 sg13g2_dfrbp_1 _10766_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net788),
    .D(_00226_),
    .Q_N(_05189_),
    .Q(\ChiselTop.wild.cpu.regs[3][4] ));
 sg13g2_dfrbp_1 _10767_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net787),
    .D(_00227_),
    .Q_N(_05188_),
    .Q(\ChiselTop.wild.cpu.regs[3][5] ));
 sg13g2_dfrbp_1 _10768_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net786),
    .D(_00228_),
    .Q_N(_05187_),
    .Q(\ChiselTop.wild.cpu.regs[3][6] ));
 sg13g2_dfrbp_1 _10769_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net785),
    .D(_00229_),
    .Q_N(_05186_),
    .Q(\ChiselTop.wild.cpu.regs[3][7] ));
 sg13g2_dfrbp_1 _10770_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net784),
    .D(_00230_),
    .Q_N(_05185_),
    .Q(\ChiselTop.wild.cpu.regs[3][8] ));
 sg13g2_dfrbp_1 _10771_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net783),
    .D(_00231_),
    .Q_N(_05184_),
    .Q(\ChiselTop.wild.cpu.regs[3][9] ));
 sg13g2_dfrbp_1 _10772_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net782),
    .D(_00232_),
    .Q_N(_05183_),
    .Q(\ChiselTop.wild.cpu.regs[3][10] ));
 sg13g2_dfrbp_1 _10773_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net781),
    .D(_00233_),
    .Q_N(_05182_),
    .Q(\ChiselTop.wild.cpu.regs[3][11] ));
 sg13g2_dfrbp_1 _10774_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net780),
    .D(_00234_),
    .Q_N(_05181_),
    .Q(\ChiselTop.wild.cpu.regs[3][12] ));
 sg13g2_dfrbp_1 _10775_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net779),
    .D(_00235_),
    .Q_N(_05180_),
    .Q(\ChiselTop.wild.cpu.regs[3][13] ));
 sg13g2_dfrbp_1 _10776_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net778),
    .D(_00236_),
    .Q_N(_05179_),
    .Q(\ChiselTop.wild.cpu.regs[3][14] ));
 sg13g2_dfrbp_1 _10777_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net777),
    .D(_00237_),
    .Q_N(_05178_),
    .Q(\ChiselTop.wild.cpu.regs[3][15] ));
 sg13g2_dfrbp_1 _10778_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net776),
    .D(_00238_),
    .Q_N(_05177_),
    .Q(\ChiselTop.wild.cpu.regs[3][16] ));
 sg13g2_dfrbp_1 _10779_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net775),
    .D(_00239_),
    .Q_N(_05176_),
    .Q(\ChiselTop.wild.cpu.regs[3][17] ));
 sg13g2_dfrbp_1 _10780_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net774),
    .D(_00240_),
    .Q_N(_05175_),
    .Q(\ChiselTop.wild.cpu.regs[3][18] ));
 sg13g2_dfrbp_1 _10781_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net773),
    .D(_00241_),
    .Q_N(_05174_),
    .Q(\ChiselTop.wild.cpu.regs[3][19] ));
 sg13g2_dfrbp_1 _10782_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net772),
    .D(_00242_),
    .Q_N(_05173_),
    .Q(\ChiselTop.wild.cpu.regs[3][20] ));
 sg13g2_dfrbp_1 _10783_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net771),
    .D(_00243_),
    .Q_N(_05172_),
    .Q(\ChiselTop.wild.cpu.regs[3][21] ));
 sg13g2_dfrbp_1 _10784_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net770),
    .D(_00244_),
    .Q_N(_05171_),
    .Q(\ChiselTop.wild.cpu.regs[3][22] ));
 sg13g2_dfrbp_1 _10785_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net769),
    .D(_00245_),
    .Q_N(_05170_),
    .Q(\ChiselTop.wild.cpu.regs[3][23] ));
 sg13g2_dfrbp_1 _10786_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net768),
    .D(_00246_),
    .Q_N(_05169_),
    .Q(\ChiselTop.wild.cpu.regs[3][24] ));
 sg13g2_dfrbp_1 _10787_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net767),
    .D(_00247_),
    .Q_N(_05168_),
    .Q(\ChiselTop.wild.cpu.regs[3][25] ));
 sg13g2_dfrbp_1 _10788_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net766),
    .D(_00248_),
    .Q_N(_05167_),
    .Q(\ChiselTop.wild.cpu.regs[3][26] ));
 sg13g2_dfrbp_1 _10789_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net765),
    .D(_00249_),
    .Q_N(_05166_),
    .Q(\ChiselTop.wild.cpu.regs[3][27] ));
 sg13g2_dfrbp_1 _10790_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net764),
    .D(_00250_),
    .Q_N(_05165_),
    .Q(\ChiselTop.wild.cpu.regs[3][28] ));
 sg13g2_dfrbp_1 _10791_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net763),
    .D(_00251_),
    .Q_N(_05164_),
    .Q(\ChiselTop.wild.cpu.regs[3][29] ));
 sg13g2_dfrbp_1 _10792_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net762),
    .D(_00252_),
    .Q_N(_05163_),
    .Q(\ChiselTop.wild.cpu.regs[3][30] ));
 sg13g2_dfrbp_1 _10793_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net761),
    .D(_00253_),
    .Q_N(_05162_),
    .Q(\ChiselTop.wild.cpu.regs[3][31] ));
 sg13g2_dfrbp_1 _10794_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net760),
    .D(_00254_),
    .Q_N(_05161_),
    .Q(\ChiselTop.wild.cpu.regs[31][0] ));
 sg13g2_dfrbp_1 _10795_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net759),
    .D(_00255_),
    .Q_N(_05160_),
    .Q(\ChiselTop.wild.cpu.regs[31][1] ));
 sg13g2_dfrbp_1 _10796_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net758),
    .D(_00256_),
    .Q_N(_05159_),
    .Q(\ChiselTop.wild.cpu.regs[31][2] ));
 sg13g2_dfrbp_1 _10797_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net757),
    .D(_00257_),
    .Q_N(_05158_),
    .Q(\ChiselTop.wild.cpu.regs[31][3] ));
 sg13g2_dfrbp_1 _10798_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net756),
    .D(_00258_),
    .Q_N(_05157_),
    .Q(\ChiselTop.wild.cpu.regs[31][4] ));
 sg13g2_dfrbp_1 _10799_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net755),
    .D(_00259_),
    .Q_N(_05156_),
    .Q(\ChiselTop.wild.cpu.regs[31][5] ));
 sg13g2_dfrbp_1 _10800_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net754),
    .D(_00260_),
    .Q_N(_05155_),
    .Q(\ChiselTop.wild.cpu.regs[31][6] ));
 sg13g2_dfrbp_1 _10801_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net753),
    .D(_00261_),
    .Q_N(_05154_),
    .Q(\ChiselTop.wild.cpu.regs[31][7] ));
 sg13g2_dfrbp_1 _10802_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net752),
    .D(_00262_),
    .Q_N(_05153_),
    .Q(\ChiselTop.wild.cpu.regs[31][8] ));
 sg13g2_dfrbp_1 _10803_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net751),
    .D(_00263_),
    .Q_N(_05152_),
    .Q(\ChiselTop.wild.cpu.regs[31][9] ));
 sg13g2_dfrbp_1 _10804_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net750),
    .D(_00264_),
    .Q_N(_05151_),
    .Q(\ChiselTop.wild.cpu.regs[31][10] ));
 sg13g2_dfrbp_1 _10805_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net749),
    .D(_00265_),
    .Q_N(_05150_),
    .Q(\ChiselTop.wild.cpu.regs[31][11] ));
 sg13g2_dfrbp_1 _10806_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net748),
    .D(_00266_),
    .Q_N(_05149_),
    .Q(\ChiselTop.wild.cpu.regs[31][12] ));
 sg13g2_dfrbp_1 _10807_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net747),
    .D(_00267_),
    .Q_N(_05148_),
    .Q(\ChiselTop.wild.cpu.regs[31][13] ));
 sg13g2_dfrbp_1 _10808_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net746),
    .D(_00268_),
    .Q_N(_05147_),
    .Q(\ChiselTop.wild.cpu.regs[31][14] ));
 sg13g2_dfrbp_1 _10809_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net745),
    .D(_00269_),
    .Q_N(_05146_),
    .Q(\ChiselTop.wild.cpu.regs[31][15] ));
 sg13g2_dfrbp_1 _10810_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net744),
    .D(_00270_),
    .Q_N(_05145_),
    .Q(\ChiselTop.wild.cpu.regs[31][16] ));
 sg13g2_dfrbp_1 _10811_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net743),
    .D(_00271_),
    .Q_N(_05144_),
    .Q(\ChiselTop.wild.cpu.regs[31][17] ));
 sg13g2_dfrbp_1 _10812_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net742),
    .D(_00272_),
    .Q_N(_05143_),
    .Q(\ChiselTop.wild.cpu.regs[31][18] ));
 sg13g2_dfrbp_1 _10813_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net741),
    .D(_00273_),
    .Q_N(_05142_),
    .Q(\ChiselTop.wild.cpu.regs[31][19] ));
 sg13g2_dfrbp_1 _10814_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net740),
    .D(_00274_),
    .Q_N(_05141_),
    .Q(\ChiselTop.wild.cpu.regs[31][20] ));
 sg13g2_dfrbp_1 _10815_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net739),
    .D(_00275_),
    .Q_N(_05140_),
    .Q(\ChiselTop.wild.cpu.regs[31][21] ));
 sg13g2_dfrbp_1 _10816_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net738),
    .D(_00276_),
    .Q_N(_05139_),
    .Q(\ChiselTop.wild.cpu.regs[31][22] ));
 sg13g2_dfrbp_1 _10817_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net737),
    .D(_00277_),
    .Q_N(_05138_),
    .Q(\ChiselTop.wild.cpu.regs[31][23] ));
 sg13g2_dfrbp_1 _10818_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net736),
    .D(_00278_),
    .Q_N(_05137_),
    .Q(\ChiselTop.wild.cpu.regs[31][24] ));
 sg13g2_dfrbp_1 _10819_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net735),
    .D(_00279_),
    .Q_N(_05136_),
    .Q(\ChiselTop.wild.cpu.regs[31][25] ));
 sg13g2_dfrbp_1 _10820_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net734),
    .D(_00280_),
    .Q_N(_05135_),
    .Q(\ChiselTop.wild.cpu.regs[31][26] ));
 sg13g2_dfrbp_1 _10821_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net733),
    .D(_00281_),
    .Q_N(_05134_),
    .Q(\ChiselTop.wild.cpu.regs[31][27] ));
 sg13g2_dfrbp_1 _10822_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net732),
    .D(_00282_),
    .Q_N(_05133_),
    .Q(\ChiselTop.wild.cpu.regs[31][28] ));
 sg13g2_dfrbp_1 _10823_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net731),
    .D(_00283_),
    .Q_N(_05132_),
    .Q(\ChiselTop.wild.cpu.regs[31][29] ));
 sg13g2_dfrbp_1 _10824_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net730),
    .D(_00284_),
    .Q_N(_05131_),
    .Q(\ChiselTop.wild.cpu.regs[31][30] ));
 sg13g2_dfrbp_1 _10825_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net729),
    .D(_00285_),
    .Q_N(_05130_),
    .Q(\ChiselTop.wild.cpu.regs[31][31] ));
 sg13g2_dfrbp_1 _10826_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net728),
    .D(_00286_),
    .Q_N(_05129_),
    .Q(\ChiselTop.wild.cpu.regs[29][0] ));
 sg13g2_dfrbp_1 _10827_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net727),
    .D(_00287_),
    .Q_N(_05128_),
    .Q(\ChiselTop.wild.cpu.regs[29][1] ));
 sg13g2_dfrbp_1 _10828_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net726),
    .D(_00288_),
    .Q_N(_05127_),
    .Q(\ChiselTop.wild.cpu.regs[29][2] ));
 sg13g2_dfrbp_1 _10829_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net725),
    .D(_00289_),
    .Q_N(_05126_),
    .Q(\ChiselTop.wild.cpu.regs[29][3] ));
 sg13g2_dfrbp_1 _10830_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net724),
    .D(_00290_),
    .Q_N(_05125_),
    .Q(\ChiselTop.wild.cpu.regs[29][4] ));
 sg13g2_dfrbp_1 _10831_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net723),
    .D(_00291_),
    .Q_N(_05124_),
    .Q(\ChiselTop.wild.cpu.regs[29][5] ));
 sg13g2_dfrbp_1 _10832_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net722),
    .D(_00292_),
    .Q_N(_05123_),
    .Q(\ChiselTop.wild.cpu.regs[29][6] ));
 sg13g2_dfrbp_1 _10833_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net721),
    .D(_00293_),
    .Q_N(_05122_),
    .Q(\ChiselTop.wild.cpu.regs[29][7] ));
 sg13g2_dfrbp_1 _10834_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net720),
    .D(_00294_),
    .Q_N(_05121_),
    .Q(\ChiselTop.wild.cpu.regs[29][8] ));
 sg13g2_dfrbp_1 _10835_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net719),
    .D(_00295_),
    .Q_N(_05120_),
    .Q(\ChiselTop.wild.cpu.regs[29][9] ));
 sg13g2_dfrbp_1 _10836_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net718),
    .D(_00296_),
    .Q_N(_05119_),
    .Q(\ChiselTop.wild.cpu.regs[29][10] ));
 sg13g2_dfrbp_1 _10837_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net717),
    .D(_00297_),
    .Q_N(_05118_),
    .Q(\ChiselTop.wild.cpu.regs[29][11] ));
 sg13g2_dfrbp_1 _10838_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net716),
    .D(_00298_),
    .Q_N(_05117_),
    .Q(\ChiselTop.wild.cpu.regs[29][12] ));
 sg13g2_dfrbp_1 _10839_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net715),
    .D(_00299_),
    .Q_N(_05116_),
    .Q(\ChiselTop.wild.cpu.regs[29][13] ));
 sg13g2_dfrbp_1 _10840_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net714),
    .D(_00300_),
    .Q_N(_05115_),
    .Q(\ChiselTop.wild.cpu.regs[29][14] ));
 sg13g2_dfrbp_1 _10841_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net713),
    .D(_00301_),
    .Q_N(_05114_),
    .Q(\ChiselTop.wild.cpu.regs[29][15] ));
 sg13g2_dfrbp_1 _10842_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net712),
    .D(_00302_),
    .Q_N(_05113_),
    .Q(\ChiselTop.wild.cpu.regs[29][16] ));
 sg13g2_dfrbp_1 _10843_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net711),
    .D(_00303_),
    .Q_N(_05112_),
    .Q(\ChiselTop.wild.cpu.regs[29][17] ));
 sg13g2_dfrbp_1 _10844_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net710),
    .D(_00304_),
    .Q_N(_05111_),
    .Q(\ChiselTop.wild.cpu.regs[29][18] ));
 sg13g2_dfrbp_1 _10845_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net709),
    .D(_00305_),
    .Q_N(_05110_),
    .Q(\ChiselTop.wild.cpu.regs[29][19] ));
 sg13g2_dfrbp_1 _10846_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net708),
    .D(_00306_),
    .Q_N(_05109_),
    .Q(\ChiselTop.wild.cpu.regs[29][20] ));
 sg13g2_dfrbp_1 _10847_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net707),
    .D(_00307_),
    .Q_N(_05108_),
    .Q(\ChiselTop.wild.cpu.regs[29][21] ));
 sg13g2_dfrbp_1 _10848_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net706),
    .D(_00308_),
    .Q_N(_05107_),
    .Q(\ChiselTop.wild.cpu.regs[29][22] ));
 sg13g2_dfrbp_1 _10849_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net705),
    .D(_00309_),
    .Q_N(_05106_),
    .Q(\ChiselTop.wild.cpu.regs[29][23] ));
 sg13g2_dfrbp_1 _10850_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net704),
    .D(_00310_),
    .Q_N(_05105_),
    .Q(\ChiselTop.wild.cpu.regs[29][24] ));
 sg13g2_dfrbp_1 _10851_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net703),
    .D(_00311_),
    .Q_N(_05104_),
    .Q(\ChiselTop.wild.cpu.regs[29][25] ));
 sg13g2_dfrbp_1 _10852_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net702),
    .D(_00312_),
    .Q_N(_05103_),
    .Q(\ChiselTop.wild.cpu.regs[29][26] ));
 sg13g2_dfrbp_1 _10853_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net701),
    .D(_00313_),
    .Q_N(_05102_),
    .Q(\ChiselTop.wild.cpu.regs[29][27] ));
 sg13g2_dfrbp_1 _10854_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net700),
    .D(_00314_),
    .Q_N(_05101_),
    .Q(\ChiselTop.wild.cpu.regs[29][28] ));
 sg13g2_dfrbp_1 _10855_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net699),
    .D(_00315_),
    .Q_N(_05100_),
    .Q(\ChiselTop.wild.cpu.regs[29][29] ));
 sg13g2_dfrbp_1 _10856_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net698),
    .D(_00316_),
    .Q_N(_05099_),
    .Q(\ChiselTop.wild.cpu.regs[29][30] ));
 sg13g2_dfrbp_1 _10857_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net697),
    .D(_00317_),
    .Q_N(_05098_),
    .Q(\ChiselTop.wild.cpu.regs[29][31] ));
 sg13g2_dfrbp_1 _10858_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net696),
    .D(_00318_),
    .Q_N(_05097_),
    .Q(\ChiselTop.wild.cpu.regs[30][0] ));
 sg13g2_dfrbp_1 _10859_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net695),
    .D(_00319_),
    .Q_N(_05096_),
    .Q(\ChiselTop.wild.cpu.regs[30][1] ));
 sg13g2_dfrbp_1 _10860_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net694),
    .D(_00320_),
    .Q_N(_05095_),
    .Q(\ChiselTop.wild.cpu.regs[30][2] ));
 sg13g2_dfrbp_1 _10861_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net693),
    .D(_00321_),
    .Q_N(_05094_),
    .Q(\ChiselTop.wild.cpu.regs[30][3] ));
 sg13g2_dfrbp_1 _10862_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net692),
    .D(_00322_),
    .Q_N(_05093_),
    .Q(\ChiselTop.wild.cpu.regs[30][4] ));
 sg13g2_dfrbp_1 _10863_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net691),
    .D(_00323_),
    .Q_N(_05092_),
    .Q(\ChiselTop.wild.cpu.regs[30][5] ));
 sg13g2_dfrbp_1 _10864_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net690),
    .D(_00324_),
    .Q_N(_05091_),
    .Q(\ChiselTop.wild.cpu.regs[30][6] ));
 sg13g2_dfrbp_1 _10865_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net689),
    .D(_00325_),
    .Q_N(_05090_),
    .Q(\ChiselTop.wild.cpu.regs[30][7] ));
 sg13g2_dfrbp_1 _10866_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net688),
    .D(_00326_),
    .Q_N(_05089_),
    .Q(\ChiselTop.wild.cpu.regs[30][8] ));
 sg13g2_dfrbp_1 _10867_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net687),
    .D(_00327_),
    .Q_N(_05088_),
    .Q(\ChiselTop.wild.cpu.regs[30][9] ));
 sg13g2_dfrbp_1 _10868_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net686),
    .D(_00328_),
    .Q_N(_05087_),
    .Q(\ChiselTop.wild.cpu.regs[30][10] ));
 sg13g2_dfrbp_1 _10869_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net685),
    .D(_00329_),
    .Q_N(_05086_),
    .Q(\ChiselTop.wild.cpu.regs[30][11] ));
 sg13g2_dfrbp_1 _10870_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net684),
    .D(_00330_),
    .Q_N(_05085_),
    .Q(\ChiselTop.wild.cpu.regs[30][12] ));
 sg13g2_dfrbp_1 _10871_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net683),
    .D(_00331_),
    .Q_N(_05084_),
    .Q(\ChiselTop.wild.cpu.regs[30][13] ));
 sg13g2_dfrbp_1 _10872_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net682),
    .D(_00332_),
    .Q_N(_05083_),
    .Q(\ChiselTop.wild.cpu.regs[30][14] ));
 sg13g2_dfrbp_1 _10873_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net681),
    .D(_00333_),
    .Q_N(_05082_),
    .Q(\ChiselTop.wild.cpu.regs[30][15] ));
 sg13g2_dfrbp_1 _10874_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net680),
    .D(_00334_),
    .Q_N(_05081_),
    .Q(\ChiselTop.wild.cpu.regs[30][16] ));
 sg13g2_dfrbp_1 _10875_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net679),
    .D(_00335_),
    .Q_N(_05080_),
    .Q(\ChiselTop.wild.cpu.regs[30][17] ));
 sg13g2_dfrbp_1 _10876_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net678),
    .D(_00336_),
    .Q_N(_05079_),
    .Q(\ChiselTop.wild.cpu.regs[30][18] ));
 sg13g2_dfrbp_1 _10877_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net677),
    .D(_00337_),
    .Q_N(_05078_),
    .Q(\ChiselTop.wild.cpu.regs[30][19] ));
 sg13g2_dfrbp_1 _10878_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net676),
    .D(_00338_),
    .Q_N(_05077_),
    .Q(\ChiselTop.wild.cpu.regs[30][20] ));
 sg13g2_dfrbp_1 _10879_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net675),
    .D(_00339_),
    .Q_N(_05076_),
    .Q(\ChiselTop.wild.cpu.regs[30][21] ));
 sg13g2_dfrbp_1 _10880_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net674),
    .D(_00340_),
    .Q_N(_05075_),
    .Q(\ChiselTop.wild.cpu.regs[30][22] ));
 sg13g2_dfrbp_1 _10881_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net673),
    .D(_00341_),
    .Q_N(_05074_),
    .Q(\ChiselTop.wild.cpu.regs[30][23] ));
 sg13g2_dfrbp_1 _10882_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net672),
    .D(_00342_),
    .Q_N(_05073_),
    .Q(\ChiselTop.wild.cpu.regs[30][24] ));
 sg13g2_dfrbp_1 _10883_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net671),
    .D(_00343_),
    .Q_N(_05072_),
    .Q(\ChiselTop.wild.cpu.regs[30][25] ));
 sg13g2_dfrbp_1 _10884_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net670),
    .D(_00344_),
    .Q_N(_05071_),
    .Q(\ChiselTop.wild.cpu.regs[30][26] ));
 sg13g2_dfrbp_1 _10885_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net669),
    .D(_00345_),
    .Q_N(_05070_),
    .Q(\ChiselTop.wild.cpu.regs[30][27] ));
 sg13g2_dfrbp_1 _10886_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net668),
    .D(_00346_),
    .Q_N(_05069_),
    .Q(\ChiselTop.wild.cpu.regs[30][28] ));
 sg13g2_dfrbp_1 _10887_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net667),
    .D(_00347_),
    .Q_N(_05068_),
    .Q(\ChiselTop.wild.cpu.regs[30][29] ));
 sg13g2_dfrbp_1 _10888_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net666),
    .D(_00348_),
    .Q_N(_05067_),
    .Q(\ChiselTop.wild.cpu.regs[30][30] ));
 sg13g2_dfrbp_1 _10889_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net665),
    .D(_00349_),
    .Q_N(_05066_),
    .Q(\ChiselTop.wild.cpu.regs[30][31] ));
 sg13g2_dfrbp_1 _10890_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net664),
    .D(_00350_),
    .Q_N(_05065_),
    .Q(\ChiselTop.wild.cpu.regs[4][0] ));
 sg13g2_dfrbp_1 _10891_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net663),
    .D(_00351_),
    .Q_N(_05064_),
    .Q(\ChiselTop.wild.cpu.regs[4][1] ));
 sg13g2_dfrbp_1 _10892_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net662),
    .D(_00352_),
    .Q_N(_05063_),
    .Q(\ChiselTop.wild.cpu.regs[4][2] ));
 sg13g2_dfrbp_1 _10893_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net661),
    .D(_00353_),
    .Q_N(_05062_),
    .Q(\ChiselTop.wild.cpu.regs[4][3] ));
 sg13g2_dfrbp_1 _10894_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net660),
    .D(_00354_),
    .Q_N(_05061_),
    .Q(\ChiselTop.wild.cpu.regs[4][4] ));
 sg13g2_dfrbp_1 _10895_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net659),
    .D(_00355_),
    .Q_N(_05060_),
    .Q(\ChiselTop.wild.cpu.regs[4][5] ));
 sg13g2_dfrbp_1 _10896_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net658),
    .D(_00356_),
    .Q_N(_05059_),
    .Q(\ChiselTop.wild.cpu.regs[4][6] ));
 sg13g2_dfrbp_1 _10897_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net657),
    .D(_00357_),
    .Q_N(_05058_),
    .Q(\ChiselTop.wild.cpu.regs[4][7] ));
 sg13g2_dfrbp_1 _10898_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net656),
    .D(_00358_),
    .Q_N(_05057_),
    .Q(\ChiselTop.wild.cpu.regs[4][8] ));
 sg13g2_dfrbp_1 _10899_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net655),
    .D(_00359_),
    .Q_N(_05056_),
    .Q(\ChiselTop.wild.cpu.regs[4][9] ));
 sg13g2_dfrbp_1 _10900_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net654),
    .D(_00360_),
    .Q_N(_05055_),
    .Q(\ChiselTop.wild.cpu.regs[4][10] ));
 sg13g2_dfrbp_1 _10901_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net653),
    .D(_00361_),
    .Q_N(_05054_),
    .Q(\ChiselTop.wild.cpu.regs[4][11] ));
 sg13g2_dfrbp_1 _10902_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net652),
    .D(_00362_),
    .Q_N(_05053_),
    .Q(\ChiselTop.wild.cpu.regs[4][12] ));
 sg13g2_dfrbp_1 _10903_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net651),
    .D(_00363_),
    .Q_N(_05052_),
    .Q(\ChiselTop.wild.cpu.regs[4][13] ));
 sg13g2_dfrbp_1 _10904_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net650),
    .D(_00364_),
    .Q_N(_05051_),
    .Q(\ChiselTop.wild.cpu.regs[4][14] ));
 sg13g2_dfrbp_1 _10905_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net649),
    .D(_00365_),
    .Q_N(_05050_),
    .Q(\ChiselTop.wild.cpu.regs[4][15] ));
 sg13g2_dfrbp_1 _10906_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net648),
    .D(_00366_),
    .Q_N(_05049_),
    .Q(\ChiselTop.wild.cpu.regs[4][16] ));
 sg13g2_dfrbp_1 _10907_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net647),
    .D(_00367_),
    .Q_N(_05048_),
    .Q(\ChiselTop.wild.cpu.regs[4][17] ));
 sg13g2_dfrbp_1 _10908_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net646),
    .D(_00368_),
    .Q_N(_05047_),
    .Q(\ChiselTop.wild.cpu.regs[4][18] ));
 sg13g2_dfrbp_1 _10909_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net645),
    .D(_00369_),
    .Q_N(_05046_),
    .Q(\ChiselTop.wild.cpu.regs[4][19] ));
 sg13g2_dfrbp_1 _10910_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net644),
    .D(_00370_),
    .Q_N(_05045_),
    .Q(\ChiselTop.wild.cpu.regs[4][20] ));
 sg13g2_dfrbp_1 _10911_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net643),
    .D(_00371_),
    .Q_N(_05044_),
    .Q(\ChiselTop.wild.cpu.regs[4][21] ));
 sg13g2_dfrbp_1 _10912_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net642),
    .D(_00372_),
    .Q_N(_05043_),
    .Q(\ChiselTop.wild.cpu.regs[4][22] ));
 sg13g2_dfrbp_1 _10913_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net641),
    .D(_00373_),
    .Q_N(_05042_),
    .Q(\ChiselTop.wild.cpu.regs[4][23] ));
 sg13g2_dfrbp_1 _10914_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net640),
    .D(_00374_),
    .Q_N(_05041_),
    .Q(\ChiselTop.wild.cpu.regs[4][24] ));
 sg13g2_dfrbp_1 _10915_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net639),
    .D(_00375_),
    .Q_N(_05040_),
    .Q(\ChiselTop.wild.cpu.regs[4][25] ));
 sg13g2_dfrbp_1 _10916_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net638),
    .D(_00376_),
    .Q_N(_05039_),
    .Q(\ChiselTop.wild.cpu.regs[4][26] ));
 sg13g2_dfrbp_1 _10917_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net637),
    .D(_00377_),
    .Q_N(_05038_),
    .Q(\ChiselTop.wild.cpu.regs[4][27] ));
 sg13g2_dfrbp_1 _10918_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net636),
    .D(_00378_),
    .Q_N(_05037_),
    .Q(\ChiselTop.wild.cpu.regs[4][28] ));
 sg13g2_dfrbp_1 _10919_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net635),
    .D(_00379_),
    .Q_N(_05036_),
    .Q(\ChiselTop.wild.cpu.regs[4][29] ));
 sg13g2_dfrbp_1 _10920_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net631),
    .D(_00380_),
    .Q_N(_05035_),
    .Q(\ChiselTop.wild.cpu.regs[4][30] ));
 sg13g2_dfrbp_1 _10921_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net630),
    .D(_00381_),
    .Q_N(_05034_),
    .Q(\ChiselTop.wild.cpu.regs[4][31] ));
 sg13g2_dfrbp_1 _10922_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net629),
    .D(_00382_),
    .Q_N(_05033_),
    .Q(\ChiselTop.wild.cpu.regs[2][0] ));
 sg13g2_dfrbp_1 _10923_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net628),
    .D(_00383_),
    .Q_N(_05032_),
    .Q(\ChiselTop.wild.cpu.regs[2][1] ));
 sg13g2_dfrbp_1 _10924_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net627),
    .D(_00384_),
    .Q_N(_05031_),
    .Q(\ChiselTop.wild.cpu.regs[2][2] ));
 sg13g2_dfrbp_1 _10925_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net626),
    .D(_00385_),
    .Q_N(_05030_),
    .Q(\ChiselTop.wild.cpu.regs[2][3] ));
 sg13g2_dfrbp_1 _10926_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net625),
    .D(_00386_),
    .Q_N(_05029_),
    .Q(\ChiselTop.wild.cpu.regs[2][4] ));
 sg13g2_dfrbp_1 _10927_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net624),
    .D(_00387_),
    .Q_N(_05028_),
    .Q(\ChiselTop.wild.cpu.regs[2][5] ));
 sg13g2_dfrbp_1 _10928_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net623),
    .D(_00388_),
    .Q_N(_05027_),
    .Q(\ChiselTop.wild.cpu.regs[2][6] ));
 sg13g2_dfrbp_1 _10929_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net622),
    .D(_00389_),
    .Q_N(_05026_),
    .Q(\ChiselTop.wild.cpu.regs[2][7] ));
 sg13g2_dfrbp_1 _10930_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net621),
    .D(_00390_),
    .Q_N(_05025_),
    .Q(\ChiselTop.wild.cpu.regs[2][8] ));
 sg13g2_dfrbp_1 _10931_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net620),
    .D(_00391_),
    .Q_N(_05024_),
    .Q(\ChiselTop.wild.cpu.regs[2][9] ));
 sg13g2_dfrbp_1 _10932_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net619),
    .D(_00392_),
    .Q_N(_05023_),
    .Q(\ChiselTop.wild.cpu.regs[2][10] ));
 sg13g2_dfrbp_1 _10933_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net618),
    .D(_00393_),
    .Q_N(_05022_),
    .Q(\ChiselTop.wild.cpu.regs[2][11] ));
 sg13g2_dfrbp_1 _10934_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net617),
    .D(_00394_),
    .Q_N(_05021_),
    .Q(\ChiselTop.wild.cpu.regs[2][12] ));
 sg13g2_dfrbp_1 _10935_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net616),
    .D(_00395_),
    .Q_N(_05020_),
    .Q(\ChiselTop.wild.cpu.regs[2][13] ));
 sg13g2_dfrbp_1 _10936_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net615),
    .D(_00396_),
    .Q_N(_05019_),
    .Q(\ChiselTop.wild.cpu.regs[2][14] ));
 sg13g2_dfrbp_1 _10937_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net614),
    .D(_00397_),
    .Q_N(_05018_),
    .Q(\ChiselTop.wild.cpu.regs[2][15] ));
 sg13g2_dfrbp_1 _10938_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net613),
    .D(_00398_),
    .Q_N(_05017_),
    .Q(\ChiselTop.wild.cpu.regs[2][16] ));
 sg13g2_dfrbp_1 _10939_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net612),
    .D(_00399_),
    .Q_N(_05016_),
    .Q(\ChiselTop.wild.cpu.regs[2][17] ));
 sg13g2_dfrbp_1 _10940_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net611),
    .D(_00400_),
    .Q_N(_05015_),
    .Q(\ChiselTop.wild.cpu.regs[2][18] ));
 sg13g2_dfrbp_1 _10941_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net610),
    .D(_00401_),
    .Q_N(_05014_),
    .Q(\ChiselTop.wild.cpu.regs[2][19] ));
 sg13g2_dfrbp_1 _10942_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net609),
    .D(_00402_),
    .Q_N(_05013_),
    .Q(\ChiselTop.wild.cpu.regs[2][20] ));
 sg13g2_dfrbp_1 _10943_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net608),
    .D(_00403_),
    .Q_N(_05012_),
    .Q(\ChiselTop.wild.cpu.regs[2][21] ));
 sg13g2_dfrbp_1 _10944_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net607),
    .D(_00404_),
    .Q_N(_05011_),
    .Q(\ChiselTop.wild.cpu.regs[2][22] ));
 sg13g2_dfrbp_1 _10945_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net606),
    .D(_00405_),
    .Q_N(_05010_),
    .Q(\ChiselTop.wild.cpu.regs[2][23] ));
 sg13g2_dfrbp_1 _10946_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net605),
    .D(_00406_),
    .Q_N(_05009_),
    .Q(\ChiselTop.wild.cpu.regs[2][24] ));
 sg13g2_dfrbp_1 _10947_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net604),
    .D(_00407_),
    .Q_N(_05008_),
    .Q(\ChiselTop.wild.cpu.regs[2][25] ));
 sg13g2_dfrbp_1 _10948_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net603),
    .D(_00408_),
    .Q_N(_05007_),
    .Q(\ChiselTop.wild.cpu.regs[2][26] ));
 sg13g2_dfrbp_1 _10949_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net602),
    .D(_00409_),
    .Q_N(_05006_),
    .Q(\ChiselTop.wild.cpu.regs[2][27] ));
 sg13g2_dfrbp_1 _10950_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net601),
    .D(_00410_),
    .Q_N(_05005_),
    .Q(\ChiselTop.wild.cpu.regs[2][28] ));
 sg13g2_dfrbp_1 _10951_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net600),
    .D(_00411_),
    .Q_N(_05004_),
    .Q(\ChiselTop.wild.cpu.regs[2][29] ));
 sg13g2_dfrbp_1 _10952_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net599),
    .D(_00412_),
    .Q_N(_05003_),
    .Q(\ChiselTop.wild.cpu.regs[2][30] ));
 sg13g2_dfrbp_1 _10953_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net598),
    .D(_00413_),
    .Q_N(_05002_),
    .Q(\ChiselTop.wild.cpu.regs[2][31] ));
 sg13g2_dfrbp_1 _10954_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net597),
    .D(_00414_),
    .Q_N(_05001_),
    .Q(\ChiselTop.wild.cpu.regs[28][0] ));
 sg13g2_dfrbp_1 _10955_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net596),
    .D(_00415_),
    .Q_N(_05000_),
    .Q(\ChiselTop.wild.cpu.regs[28][1] ));
 sg13g2_dfrbp_1 _10956_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net595),
    .D(_00416_),
    .Q_N(_04999_),
    .Q(\ChiselTop.wild.cpu.regs[28][2] ));
 sg13g2_dfrbp_1 _10957_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net594),
    .D(_00417_),
    .Q_N(_04998_),
    .Q(\ChiselTop.wild.cpu.regs[28][3] ));
 sg13g2_dfrbp_1 _10958_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net593),
    .D(_00418_),
    .Q_N(_04997_),
    .Q(\ChiselTop.wild.cpu.regs[28][4] ));
 sg13g2_dfrbp_1 _10959_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net592),
    .D(_00419_),
    .Q_N(_04996_),
    .Q(\ChiselTop.wild.cpu.regs[28][5] ));
 sg13g2_dfrbp_1 _10960_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net591),
    .D(_00420_),
    .Q_N(_04995_),
    .Q(\ChiselTop.wild.cpu.regs[28][6] ));
 sg13g2_dfrbp_1 _10961_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net590),
    .D(_00421_),
    .Q_N(_04994_),
    .Q(\ChiselTop.wild.cpu.regs[28][7] ));
 sg13g2_dfrbp_1 _10962_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net589),
    .D(_00422_),
    .Q_N(_04993_),
    .Q(\ChiselTop.wild.cpu.regs[28][8] ));
 sg13g2_dfrbp_1 _10963_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net588),
    .D(_00423_),
    .Q_N(_04992_),
    .Q(\ChiselTop.wild.cpu.regs[28][9] ));
 sg13g2_dfrbp_1 _10964_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net587),
    .D(_00424_),
    .Q_N(_04991_),
    .Q(\ChiselTop.wild.cpu.regs[28][10] ));
 sg13g2_dfrbp_1 _10965_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net586),
    .D(_00425_),
    .Q_N(_04990_),
    .Q(\ChiselTop.wild.cpu.regs[28][11] ));
 sg13g2_dfrbp_1 _10966_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net585),
    .D(_00426_),
    .Q_N(_04989_),
    .Q(\ChiselTop.wild.cpu.regs[28][12] ));
 sg13g2_dfrbp_1 _10967_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net584),
    .D(_00427_),
    .Q_N(_04988_),
    .Q(\ChiselTop.wild.cpu.regs[28][13] ));
 sg13g2_dfrbp_1 _10968_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net583),
    .D(_00428_),
    .Q_N(_04987_),
    .Q(\ChiselTop.wild.cpu.regs[28][14] ));
 sg13g2_dfrbp_1 _10969_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net582),
    .D(_00429_),
    .Q_N(_04986_),
    .Q(\ChiselTop.wild.cpu.regs[28][15] ));
 sg13g2_dfrbp_1 _10970_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net581),
    .D(_00430_),
    .Q_N(_04985_),
    .Q(\ChiselTop.wild.cpu.regs[28][16] ));
 sg13g2_dfrbp_1 _10971_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net580),
    .D(_00431_),
    .Q_N(_04984_),
    .Q(\ChiselTop.wild.cpu.regs[28][17] ));
 sg13g2_dfrbp_1 _10972_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net579),
    .D(_00432_),
    .Q_N(_04983_),
    .Q(\ChiselTop.wild.cpu.regs[28][18] ));
 sg13g2_dfrbp_1 _10973_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net578),
    .D(_00433_),
    .Q_N(_04982_),
    .Q(\ChiselTop.wild.cpu.regs[28][19] ));
 sg13g2_dfrbp_1 _10974_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net577),
    .D(_00434_),
    .Q_N(_04981_),
    .Q(\ChiselTop.wild.cpu.regs[28][20] ));
 sg13g2_dfrbp_1 _10975_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net576),
    .D(_00435_),
    .Q_N(_04980_),
    .Q(\ChiselTop.wild.cpu.regs[28][21] ));
 sg13g2_dfrbp_1 _10976_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net575),
    .D(_00436_),
    .Q_N(_04979_),
    .Q(\ChiselTop.wild.cpu.regs[28][22] ));
 sg13g2_dfrbp_1 _10977_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net574),
    .D(_00437_),
    .Q_N(_04978_),
    .Q(\ChiselTop.wild.cpu.regs[28][23] ));
 sg13g2_dfrbp_1 _10978_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net573),
    .D(_00438_),
    .Q_N(_04977_),
    .Q(\ChiselTop.wild.cpu.regs[28][24] ));
 sg13g2_dfrbp_1 _10979_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net572),
    .D(_00439_),
    .Q_N(_04976_),
    .Q(\ChiselTop.wild.cpu.regs[28][25] ));
 sg13g2_dfrbp_1 _10980_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net571),
    .D(_00440_),
    .Q_N(_04975_),
    .Q(\ChiselTop.wild.cpu.regs[28][26] ));
 sg13g2_dfrbp_1 _10981_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net570),
    .D(_00441_),
    .Q_N(_04974_),
    .Q(\ChiselTop.wild.cpu.regs[28][27] ));
 sg13g2_dfrbp_1 _10982_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net569),
    .D(_00442_),
    .Q_N(_04973_),
    .Q(\ChiselTop.wild.cpu.regs[28][28] ));
 sg13g2_dfrbp_1 _10983_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net568),
    .D(_00443_),
    .Q_N(_04972_),
    .Q(\ChiselTop.wild.cpu.regs[28][29] ));
 sg13g2_dfrbp_1 _10984_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net567),
    .D(_00444_),
    .Q_N(_04971_),
    .Q(\ChiselTop.wild.cpu.regs[28][30] ));
 sg13g2_dfrbp_1 _10985_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net566),
    .D(_00445_),
    .Q_N(_04970_),
    .Q(\ChiselTop.wild.cpu.regs[28][31] ));
 sg13g2_dfrbp_1 _10986_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net565),
    .D(_00446_),
    .Q_N(_04969_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[0] ));
 sg13g2_dfrbp_1 _10987_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net564),
    .D(_00447_),
    .Q_N(_04968_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[1] ));
 sg13g2_dfrbp_1 _10988_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net563),
    .D(_00448_),
    .Q_N(_04967_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[5] ));
 sg13g2_dfrbp_1 _10989_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net562),
    .D(_00449_),
    .Q_N(_04966_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[6] ));
 sg13g2_dfrbp_1 _10990_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net561),
    .D(_00450_),
    .Q_N(_04965_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[8] ));
 sg13g2_dfrbp_1 _10991_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net560),
    .D(_00451_),
    .Q_N(_04964_),
    .Q(\ChiselTop.wild.tx.tx.cntReg[9] ));
 sg13g2_dfrbp_1 _10992_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net559),
    .D(_00452_),
    .Q_N(_04963_),
    .Q(\ChiselTop.wild.ledReg[0] ));
 sg13g2_dfrbp_1 _10993_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net557),
    .D(_00453_),
    .Q_N(_04962_),
    .Q(\ChiselTop.wild.ledReg[1] ));
 sg13g2_dfrbp_1 _10994_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net555),
    .D(_00454_),
    .Q_N(_04961_),
    .Q(\ChiselTop.wild.ledReg[2] ));
 sg13g2_dfrbp_1 _10995_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net434),
    .D(_00455_),
    .Q_N(_05272_),
    .Q(\ChiselTop.wild.ledReg[3] ));
 sg13g2_dfrbp_1 _10996_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net435),
    .D(net826),
    .Q_N(_05273_),
    .Q(\ChiselTop.wild.uartStatusReg[0] ));
 sg13g2_dfrbp_1 _10997_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net436),
    .D(net854),
    .Q_N(_05274_),
    .Q(\ChiselTop.wild.uartStatusReg[1] ));
 sg13g2_dfrbp_1 _10998_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net437),
    .D(\ChiselTop.wild.cpu.decEx_memLow[0] ),
    .Q_N(_05275_),
    .Q(\ChiselTop.wild.memAddressReg[0] ));
 sg13g2_dfrbp_1 _10999_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net438),
    .D(\ChiselTop.wild.cpu.decEx_memLow[1] ),
    .Q_N(_05276_),
    .Q(\ChiselTop.wild.memAddressReg[1] ));
 sg13g2_dfrbp_1 _11000_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net439),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[2] ),
    .Q_N(_05277_),
    .Q(\ChiselTop.wild.memAddressReg[2] ));
 sg13g2_dfrbp_1 _11001_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net440),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[3] ),
    .Q_N(_05278_),
    .Q(\ChiselTop.wild.memAddressReg[3] ));
 sg13g2_dfrbp_1 _11002_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net441),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[16] ),
    .Q_N(_05279_),
    .Q(\ChiselTop.wild.memAddressReg[16] ));
 sg13g2_dfrbp_1 _11003_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net442),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[17] ),
    .Q_N(_05280_),
    .Q(\ChiselTop.wild.memAddressReg[17] ));
 sg13g2_dfrbp_1 _11004_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net443),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[18] ),
    .Q_N(_05281_),
    .Q(\ChiselTop.wild.memAddressReg[18] ));
 sg13g2_dfrbp_1 _11005_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net444),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[19] ),
    .Q_N(_05282_),
    .Q(\ChiselTop.wild.memAddressReg[19] ));
 sg13g2_dfrbp_1 _11006_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net445),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[28] ),
    .Q_N(_05283_),
    .Q(\ChiselTop.wild.memAddressReg[28] ));
 sg13g2_dfrbp_1 _11007_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net446),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[29] ),
    .Q_N(_05284_),
    .Q(\ChiselTop.wild.memAddressReg[29] ));
 sg13g2_dfrbp_1 _11008_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net447),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[30] ),
    .Q_N(_05285_),
    .Q(\ChiselTop.wild.memAddressReg[30] ));
 sg13g2_dfrbp_1 _11009_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net448),
    .D(\ChiselTop.wild.cpu.io_dmem_rdAddress[31] ),
    .Q_N(_05286_),
    .Q(\ChiselTop.wild.memAddressReg[31] ));
 sg13g2_dfrbp_1 _11010_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net449),
    .D(net834),
    .Q_N(_05287_),
    .Q(\ChiselTop.dec.counter[0] ));
 sg13g2_dfrbp_1 _11011_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net450),
    .D(net830),
    .Q_N(_05288_),
    .Q(\ChiselTop.dec.counter[1] ));
 sg13g2_dfrbp_1 _11012_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net457),
    .D(net831),
    .Q_N(_05289_),
    .Q(\ChiselTop.dec.counter[2] ));
 sg13g2_dfrbp_1 _11013_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net553),
    .D(net827),
    .Q_N(_04960_),
    .Q(\ChiselTop.dec.counter[3] ));
 sg13g2_dfrbp_1 _11014_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net551),
    .D(_00456_),
    .Q_N(_04959_),
    .Q(\ChiselTop.wild.cpu.decExReg_rd[0] ));
 sg13g2_dfrbp_1 _11015_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net550),
    .D(_00457_),
    .Q_N(_04958_),
    .Q(\ChiselTop.wild.cpu.decExReg_rd[1] ));
 sg13g2_dfrbp_1 _11016_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net549),
    .D(_00458_),
    .Q_N(_00142_),
    .Q(\ChiselTop.wild.cpu.decExReg_rd[2] ));
 sg13g2_dfrbp_1 _11017_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net548),
    .D(_00459_),
    .Q_N(_04957_),
    .Q(\ChiselTop.wild.cpu.decExReg_rd[3] ));
 sg13g2_dfrbp_1 _11018_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net547),
    .D(_00460_),
    .Q_N(_04956_),
    .Q(\ChiselTop.wild.cpu.decOut_opcode[2] ));
 sg13g2_dfrbp_1 _11019_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net458),
    .D(_00461_),
    .Q_N(_05290_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_isImm ));
 sg13g2_dfrbp_1 _11020_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net459),
    .D(net829),
    .Q_N(_05291_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[0] ));
 sg13g2_dfrbp_1 _11021_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net460),
    .D(net833),
    .Q_N(_05292_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[1] ));
 sg13g2_dfrbp_1 _11022_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net461),
    .D(net1260),
    .Q_N(_05293_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[2] ));
 sg13g2_dfrbp_1 _11023_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net462),
    .D(net1038),
    .Q_N(_05294_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[3] ));
 sg13g2_dfrbp_1 _11024_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net463),
    .D(net856),
    .Q_N(_05295_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[4] ));
 sg13g2_dfrbp_1 _11025_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net464),
    .D(net860),
    .Q_N(_05296_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[5] ));
 sg13g2_dfrbp_1 _11026_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net465),
    .D(net832),
    .Q_N(_05297_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[6] ));
 sg13g2_dfrbp_1 _11027_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net466),
    .D(net866),
    .Q_N(_05298_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[7] ));
 sg13g2_dfrbp_1 _11028_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net467),
    .D(net849),
    .Q_N(_05299_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[8] ));
 sg13g2_dfrbp_1 _11029_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net468),
    .D(net844),
    .Q_N(_05300_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[9] ));
 sg13g2_dfrbp_1 _11030_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net469),
    .D(net863),
    .Q_N(_05301_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[10] ));
 sg13g2_dfrbp_1 _11031_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net470),
    .D(net838),
    .Q_N(_05302_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[11] ));
 sg13g2_dfrbp_1 _11032_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net471),
    .D(net852),
    .Q_N(_05303_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[12] ));
 sg13g2_dfrbp_1 _11033_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net472),
    .D(net865),
    .Q_N(_05304_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[13] ));
 sg13g2_dfrbp_1 _11034_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net473),
    .D(net836),
    .Q_N(_05305_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[14] ));
 sg13g2_dfrbp_1 _11035_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net474),
    .D(net835),
    .Q_N(_05306_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[15] ));
 sg13g2_dfrbp_1 _11036_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net475),
    .D(net858),
    .Q_N(_05307_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[16] ));
 sg13g2_dfrbp_1 _11037_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net476),
    .D(net851),
    .Q_N(_05308_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[17] ));
 sg13g2_dfrbp_1 _11038_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net477),
    .D(net828),
    .Q_N(_05309_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[18] ));
 sg13g2_dfrbp_1 _11039_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net478),
    .D(net841),
    .Q_N(_05310_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[19] ));
 sg13g2_dfrbp_1 _11040_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net479),
    .D(net857),
    .Q_N(_05311_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[20] ));
 sg13g2_dfrbp_1 _11041_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net480),
    .D(net837),
    .Q_N(_05312_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[21] ));
 sg13g2_dfrbp_1 _11042_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net481),
    .D(net846),
    .Q_N(_05313_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[22] ));
 sg13g2_dfrbp_1 _11043_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net482),
    .D(net845),
    .Q_N(_05314_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[23] ));
 sg13g2_dfrbp_1 _11044_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net483),
    .D(net842),
    .Q_N(_05315_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[24] ));
 sg13g2_dfrbp_1 _11045_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net484),
    .D(net850),
    .Q_N(_05316_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[25] ));
 sg13g2_dfrbp_1 _11046_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net485),
    .D(net848),
    .Q_N(_05317_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[26] ));
 sg13g2_dfrbp_1 _11047_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net486),
    .D(net839),
    .Q_N(_05318_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[27] ));
 sg13g2_dfrbp_1 _11048_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net487),
    .D(net843),
    .Q_N(_05319_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[28] ));
 sg13g2_dfrbp_1 _11049_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net488),
    .D(net855),
    .Q_N(_05320_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[29] ));
 sg13g2_dfrbp_1 _11050_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net632),
    .D(net847),
    .Q_N(_05321_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[30] ));
 sg13g2_dfrbp_1 _11051_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net546),
    .D(net840),
    .Q_N(_04955_),
    .Q(\ChiselTop.wild.cpu.pcRegReg[31] ));
 sg13g2_dfrbp_1 _11052_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net545),
    .D(_00462_),
    .Q_N(_04954_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[0] ));
 sg13g2_dfrbp_1 _11053_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net544),
    .D(net1498),
    .Q_N(_04953_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_isLui ));
 sg13g2_dfrbp_1 _11054_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net543),
    .D(_00464_),
    .Q_N(_00062_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[0] ));
 sg13g2_dfrbp_1 _11055_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net542),
    .D(_00465_),
    .Q_N(_00058_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[1] ));
 sg13g2_dfrbp_1 _11056_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net541),
    .D(_00466_),
    .Q_N(_00054_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[2] ));
 sg13g2_dfrbp_1 _11057_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net540),
    .D(_00467_),
    .Q_N(_00050_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[3] ));
 sg13g2_dfrbp_1 _11058_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net539),
    .D(_00468_),
    .Q_N(_00118_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[4] ));
 sg13g2_dfrbp_1 _11059_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net538),
    .D(_00469_),
    .Q_N(_00044_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[5] ));
 sg13g2_dfrbp_1 _11060_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net537),
    .D(_00470_),
    .Q_N(_00037_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[6] ));
 sg13g2_dfrbp_1 _11061_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net536),
    .D(_00471_),
    .Q_N(_00027_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[10] ));
 sg13g2_dfrbp_1 _11062_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net535),
    .D(_00472_),
    .Q_N(_00023_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[11] ));
 sg13g2_dfrbp_1 _11063_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net534),
    .D(_00473_),
    .Q_N(_00019_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[12] ));
 sg13g2_dfrbp_1 _11064_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net533),
    .D(_00474_),
    .Q_N(_00015_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[13] ));
 sg13g2_dfrbp_1 _11065_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net532),
    .D(_00475_),
    .Q_N(_00007_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[15] ));
 sg13g2_dfrbp_1 _11066_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net531),
    .D(_00476_),
    .Q_N(_00004_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[16] ));
 sg13g2_dfrbp_1 _11067_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net530),
    .D(_00477_),
    .Q_N(_00133_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[17] ));
 sg13g2_dfrbp_1 _11068_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net529),
    .D(_00478_),
    .Q_N(_00011_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[14] ));
 sg13g2_dfrbp_1 _11069_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net528),
    .D(_00479_),
    .Q_N(_00132_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[20] ));
 sg13g2_dfrbp_1 _11070_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net527),
    .D(_00480_),
    .Q_N(_00131_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[21] ));
 sg13g2_dfrbp_1 _11071_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net526),
    .D(_00481_),
    .Q_N(_00130_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[22] ));
 sg13g2_dfrbp_1 _11072_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net525),
    .D(_00482_),
    .Q_N(_00129_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[25] ));
 sg13g2_dfrbp_1 _11073_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net524),
    .D(_00483_),
    .Q_N(_00128_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[26] ));
 sg13g2_dfrbp_1 _11074_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net523),
    .D(_00484_),
    .Q_N(_00127_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[28] ));
 sg13g2_dfrbp_1 _11075_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net522),
    .D(_00485_),
    .Q_N(_00126_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_imm[31] ));
 sg13g2_dfrbp_1 _11076_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net521),
    .D(_00486_),
    .Q_N(_00124_),
    .Q(\ChiselTop.wild.cpu._wbData_T_1[0] ));
 sg13g2_dfrbp_1 _11077_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net520),
    .D(_00487_),
    .Q_N(_04952_),
    .Q(\ChiselTop.wild.cpu._wbData_T_1[1] ));
 sg13g2_dfrbp_1 _11078_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net519),
    .D(_00488_),
    .Q_N(_00121_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[2] ));
 sg13g2_dfrbp_1 _11079_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net518),
    .D(_00489_),
    .Q_N(_04951_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[3] ));
 sg13g2_dfrbp_1 _11080_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net517),
    .D(_00490_),
    .Q_N(_04950_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[4] ));
 sg13g2_dfrbp_1 _11081_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net516),
    .D(_00491_),
    .Q_N(_04949_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[5] ));
 sg13g2_dfrbp_1 _11082_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net515),
    .D(_00492_),
    .Q_N(_00117_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[6] ));
 sg13g2_dfrbp_1 _11083_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net514),
    .D(_00493_),
    .Q_N(_04948_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[7] ));
 sg13g2_dfrbp_1 _11084_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net513),
    .D(_00494_),
    .Q_N(_00116_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[8] ));
 sg13g2_dfrbp_1 _11085_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net512),
    .D(_00495_),
    .Q_N(_04947_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[9] ));
 sg13g2_dfrbp_1 _11086_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net511),
    .D(_00496_),
    .Q_N(_04946_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[10] ));
 sg13g2_dfrbp_1 _11087_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net510),
    .D(_00497_),
    .Q_N(_04945_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[11] ));
 sg13g2_dfrbp_1 _11088_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net509),
    .D(_00498_),
    .Q_N(_04944_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[12] ));
 sg13g2_dfrbp_1 _11089_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net508),
    .D(_00499_),
    .Q_N(_04943_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[13] ));
 sg13g2_dfrbp_1 _11090_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net507),
    .D(_00500_),
    .Q_N(_04942_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[14] ));
 sg13g2_dfrbp_1 _11091_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net506),
    .D(_00501_),
    .Q_N(_04941_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[15] ));
 sg13g2_dfrbp_1 _11092_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net505),
    .D(_00502_),
    .Q_N(_04940_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[16] ));
 sg13g2_dfrbp_1 _11093_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net504),
    .D(_00503_),
    .Q_N(_04939_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[17] ));
 sg13g2_dfrbp_1 _11094_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net503),
    .D(_00504_),
    .Q_N(_04938_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[18] ));
 sg13g2_dfrbp_1 _11095_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net502),
    .D(_00505_),
    .Q_N(_04937_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[19] ));
 sg13g2_dfrbp_1 _11096_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net501),
    .D(_00506_),
    .Q_N(_04936_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[20] ));
 sg13g2_dfrbp_1 _11097_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net500),
    .D(_00507_),
    .Q_N(_04935_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[21] ));
 sg13g2_dfrbp_1 _11098_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net499),
    .D(_00508_),
    .Q_N(_04934_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[22] ));
 sg13g2_dfrbp_1 _11099_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net498),
    .D(_00509_),
    .Q_N(_04933_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[23] ));
 sg13g2_dfrbp_1 _11100_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net497),
    .D(_00510_),
    .Q_N(_04932_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[24] ));
 sg13g2_dfrbp_1 _11101_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net496),
    .D(_00511_),
    .Q_N(_04931_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[25] ));
 sg13g2_dfrbp_1 _11102_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net495),
    .D(_00512_),
    .Q_N(_04930_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[26] ));
 sg13g2_dfrbp_1 _11103_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net494),
    .D(_00513_),
    .Q_N(_04929_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[27] ));
 sg13g2_dfrbp_1 _11104_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net493),
    .D(_00514_),
    .Q_N(_00135_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[28] ));
 sg13g2_dfrbp_1 _11105_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net492),
    .D(_00515_),
    .Q_N(_04928_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[29] ));
 sg13g2_dfrbp_1 _11106_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net491),
    .D(_00516_),
    .Q_N(_04927_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[30] ));
 sg13g2_dfrbp_1 _11107_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net490),
    .D(_00517_),
    .Q_N(_04926_),
    .Q(\ChiselTop.wild.cpu.decExReg_pc[31] ));
 sg13g2_dfrbp_1 _11108_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net489),
    .D(net1500),
    .Q_N(_04925_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_isAuiPc ));
 sg13g2_dfrbp_1 _11109_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net456),
    .D(_00519_),
    .Q_N(_00125_),
    .Q(\ChiselTop.wild.cpu.decExReg_csrVal[0] ));
 sg13g2_dfrbp_1 _11110_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net455),
    .D(_00520_),
    .Q_N(_00003_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_isCssrw ));
 sg13g2_dfrbp_1 _11111_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net454),
    .D(_00521_),
    .Q_N(_04924_),
    .Q(\ChiselTop.wild.cpu.decExReg_memLow[0] ));
 sg13g2_dfrbp_1 _11112_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net453),
    .D(_00522_),
    .Q_N(_04923_),
    .Q(\ChiselTop.wild.cpu.decExReg_memLow[1] ));
 sg13g2_dfrbp_1 _11113_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net452),
    .D(_00523_),
    .Q_N(_04922_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_isLoad ));
 sg13g2_dfrbp_1 _11114_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net451),
    .D(net2169),
    .Q_N(_04921_),
    .Q(\ChiselTop.wild.cpu.decExReg_valid ));
 sg13g2_dfrbp_1 _11115_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net432),
    .D(net1473),
    .Q_N(_00002_),
    .Q(\ChiselTop.wild.cpu._T_12 ));
 sg13g2_dfrbp_1 _11116_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net431),
    .D(_00526_),
    .Q_N(_04920_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1[0] ));
 sg13g2_dfrbp_1 _11117_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net430),
    .D(_00527_),
    .Q_N(_04919_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1[1] ));
 sg13g2_dfrbp_1 _11118_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net429),
    .D(_00528_),
    .Q_N(_04918_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1[2] ));
 sg13g2_dfrbp_1 _11119_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net428),
    .D(_00529_),
    .Q_N(_04917_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_isBranch ));
 sg13g2_dfrbp_1 _11120_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net427),
    .D(_00530_),
    .Q_N(_00063_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[0] ));
 sg13g2_dfrbp_1 _11121_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net426),
    .D(_00531_),
    .Q_N(_00059_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[1] ));
 sg13g2_dfrbp_1 _11122_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net425),
    .D(_00532_),
    .Q_N(_00055_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[2] ));
 sg13g2_dfrbp_1 _11123_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net424),
    .D(_00533_),
    .Q_N(_00051_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[3] ));
 sg13g2_dfrbp_1 _11124_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net423),
    .D(_00534_),
    .Q_N(_04916_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[4] ));
 sg13g2_dfrbp_1 _11125_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net422),
    .D(_00535_),
    .Q_N(_00045_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[5] ));
 sg13g2_dfrbp_1 _11126_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net421),
    .D(_00536_),
    .Q_N(_00041_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[6] ));
 sg13g2_dfrbp_1 _11127_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net420),
    .D(_00537_),
    .Q_N(_00038_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[7] ));
 sg13g2_dfrbp_1 _11128_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net419),
    .D(_00538_),
    .Q_N(_00034_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[8] ));
 sg13g2_dfrbp_1 _11129_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net418),
    .D(_00539_),
    .Q_N(_00031_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[9] ));
 sg13g2_dfrbp_1 _11130_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net417),
    .D(_00540_),
    .Q_N(_00028_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[10] ));
 sg13g2_dfrbp_1 _11131_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net416),
    .D(_00541_),
    .Q_N(_00024_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[11] ));
 sg13g2_dfrbp_1 _11132_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net415),
    .D(_00542_),
    .Q_N(_00020_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[12] ));
 sg13g2_dfrbp_1 _11133_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net414),
    .D(_00543_),
    .Q_N(_00016_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[13] ));
 sg13g2_dfrbp_1 _11134_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net413),
    .D(_00544_),
    .Q_N(_00012_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[14] ));
 sg13g2_dfrbp_1 _11135_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net412),
    .D(_00545_),
    .Q_N(_00008_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[15] ));
 sg13g2_dfrbp_1 _11136_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net411),
    .D(_00546_),
    .Q_N(_04915_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[16] ));
 sg13g2_dfrbp_1 _11137_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net410),
    .D(_00547_),
    .Q_N(_00109_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[17] ));
 sg13g2_dfrbp_1 _11138_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net409),
    .D(_00548_),
    .Q_N(_00108_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[18] ));
 sg13g2_dfrbp_1 _11139_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net408),
    .D(_00549_),
    .Q_N(_00107_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[19] ));
 sg13g2_dfrbp_1 _11140_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net407),
    .D(_00550_),
    .Q_N(_00106_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[20] ));
 sg13g2_dfrbp_1 _11141_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net406),
    .D(_00551_),
    .Q_N(_00105_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[21] ));
 sg13g2_dfrbp_1 _11142_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net405),
    .D(_00552_),
    .Q_N(_00104_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[22] ));
 sg13g2_dfrbp_1 _11143_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net404),
    .D(_00553_),
    .Q_N(_00103_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[23] ));
 sg13g2_dfrbp_1 _11144_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net403),
    .D(_00554_),
    .Q_N(_00102_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[24] ));
 sg13g2_dfrbp_1 _11145_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net402),
    .D(_00555_),
    .Q_N(_00101_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[25] ));
 sg13g2_dfrbp_1 _11146_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net401),
    .D(_00556_),
    .Q_N(_00100_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[26] ));
 sg13g2_dfrbp_1 _11147_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net400),
    .D(_00557_),
    .Q_N(_00099_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[27] ));
 sg13g2_dfrbp_1 _11148_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net399),
    .D(_00558_),
    .Q_N(_00098_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[28] ));
 sg13g2_dfrbp_1 _11149_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net398),
    .D(_00559_),
    .Q_N(_00097_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[29] ));
 sg13g2_dfrbp_1 _11150_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net397),
    .D(_00560_),
    .Q_N(_00095_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[30] ));
 sg13g2_dfrbp_1 _11151_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net396),
    .D(_00561_),
    .Q_N(_00093_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2Val[31] ));
 sg13g2_dfrbp_1 _11152_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net395),
    .D(_00562_),
    .Q_N(_04914_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2[0] ));
 sg13g2_dfrbp_1 _11153_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net394),
    .D(_00563_),
    .Q_N(_04913_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2[1] ));
 sg13g2_dfrbp_1 _11154_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net393),
    .D(_00564_),
    .Q_N(_04912_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs2[2] ));
 sg13g2_dfrbp_1 _11155_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net392),
    .D(_00565_),
    .Q_N(_00065_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[0] ));
 sg13g2_dfrbp_1 _11156_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net391),
    .D(_00566_),
    .Q_N(_00061_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[1] ));
 sg13g2_dfrbp_1 _11157_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net390),
    .D(_00567_),
    .Q_N(_00057_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[2] ));
 sg13g2_dfrbp_1 _11158_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net389),
    .D(_00568_),
    .Q_N(_00053_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[3] ));
 sg13g2_dfrbp_1 _11159_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net388),
    .D(_00569_),
    .Q_N(_00049_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[4] ));
 sg13g2_dfrbp_1 _11160_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net387),
    .D(_00570_),
    .Q_N(_00047_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[5] ));
 sg13g2_dfrbp_1 _11161_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net386),
    .D(_00571_),
    .Q_N(_00043_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[6] ));
 sg13g2_dfrbp_1 _11162_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net385),
    .D(_00572_),
    .Q_N(_00040_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[7] ));
 sg13g2_dfrbp_1 _11163_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net384),
    .D(_00573_),
    .Q_N(_00036_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[8] ));
 sg13g2_dfrbp_1 _11164_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net383),
    .D(_00574_),
    .Q_N(_00033_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[9] ));
 sg13g2_dfrbp_1 _11165_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net382),
    .D(_00575_),
    .Q_N(_00030_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[10] ));
 sg13g2_dfrbp_1 _11166_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net381),
    .D(_00576_),
    .Q_N(_00026_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[11] ));
 sg13g2_dfrbp_1 _11167_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net380),
    .D(_00577_),
    .Q_N(_00022_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[12] ));
 sg13g2_dfrbp_1 _11168_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net379),
    .D(_00578_),
    .Q_N(_00018_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[13] ));
 sg13g2_dfrbp_1 _11169_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net378),
    .D(_00579_),
    .Q_N(_00014_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[14] ));
 sg13g2_dfrbp_1 _11170_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net377),
    .D(_00580_),
    .Q_N(_00010_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[15] ));
 sg13g2_dfrbp_1 _11171_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net376),
    .D(_00581_),
    .Q_N(_00006_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[16] ));
 sg13g2_dfrbp_1 _11172_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net375),
    .D(_00582_),
    .Q_N(_00068_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[17] ));
 sg13g2_dfrbp_1 _11173_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net374),
    .D(_00583_),
    .Q_N(_00070_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[18] ));
 sg13g2_dfrbp_1 _11174_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net373),
    .D(_00584_),
    .Q_N(_00072_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[19] ));
 sg13g2_dfrbp_1 _11175_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net372),
    .D(_00585_),
    .Q_N(_00074_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[20] ));
 sg13g2_dfrbp_1 _11176_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net371),
    .D(_00586_),
    .Q_N(_00076_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[21] ));
 sg13g2_dfrbp_1 _11177_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net370),
    .D(_00587_),
    .Q_N(_00078_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[22] ));
 sg13g2_dfrbp_1 _11178_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net369),
    .D(_00588_),
    .Q_N(_00080_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[23] ));
 sg13g2_dfrbp_1 _11179_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net368),
    .D(_00589_),
    .Q_N(_00082_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[24] ));
 sg13g2_dfrbp_1 _11180_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net367),
    .D(_00590_),
    .Q_N(_00084_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[25] ));
 sg13g2_dfrbp_1 _11181_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net366),
    .D(_00591_),
    .Q_N(_00086_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[26] ));
 sg13g2_dfrbp_1 _11182_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net365),
    .D(_00592_),
    .Q_N(_00088_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[27] ));
 sg13g2_dfrbp_1 _11183_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net364),
    .D(_00593_),
    .Q_N(_00090_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[28] ));
 sg13g2_dfrbp_1 _11184_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net363),
    .D(_00594_),
    .Q_N(_00092_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[29] ));
 sg13g2_dfrbp_1 _11185_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net362),
    .D(_00595_),
    .Q_N(_04911_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[30] ));
 sg13g2_dfrbp_1 _11186_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net361),
    .D(_00596_),
    .Q_N(_04910_),
    .Q(\ChiselTop.wild.cpu.decExReg_rs1Val[31] ));
 sg13g2_dfrbp_1 _11187_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net360),
    .D(_00597_),
    .Q_N(_04909_),
    .Q(\ChiselTop.wild.cpu.decExReg_func3[0] ));
 sg13g2_dfrbp_1 _11188_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net359),
    .D(_00598_),
    .Q_N(_04908_),
    .Q(\ChiselTop.wild.cpu.decExReg_func3[1] ));
 sg13g2_dfrbp_1 _11189_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net358),
    .D(_00599_),
    .Q_N(_00064_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[0] ));
 sg13g2_dfrbp_1 _11190_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net357),
    .D(_00600_),
    .Q_N(_00060_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[1] ));
 sg13g2_dfrbp_1 _11191_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net356),
    .D(_00601_),
    .Q_N(_00056_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[2] ));
 sg13g2_dfrbp_1 _11192_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net355),
    .D(_00602_),
    .Q_N(_00052_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[3] ));
 sg13g2_dfrbp_1 _11193_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net354),
    .D(_00603_),
    .Q_N(_00048_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[4] ));
 sg13g2_dfrbp_1 _11194_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net353),
    .D(_00604_),
    .Q_N(_00046_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[5] ));
 sg13g2_dfrbp_1 _11195_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net352),
    .D(_00605_),
    .Q_N(_00042_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[6] ));
 sg13g2_dfrbp_1 _11196_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net351),
    .D(_00606_),
    .Q_N(_00039_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[7] ));
 sg13g2_dfrbp_1 _11197_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net350),
    .D(_00607_),
    .Q_N(_00035_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[8] ));
 sg13g2_dfrbp_1 _11198_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net349),
    .D(_00608_),
    .Q_N(_00032_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[9] ));
 sg13g2_dfrbp_1 _11199_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net348),
    .D(_00609_),
    .Q_N(_00029_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[10] ));
 sg13g2_dfrbp_1 _11200_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net347),
    .D(_00610_),
    .Q_N(_00025_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[11] ));
 sg13g2_dfrbp_1 _11201_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net346),
    .D(_00611_),
    .Q_N(_00021_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[12] ));
 sg13g2_dfrbp_1 _11202_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net345),
    .D(_00612_),
    .Q_N(_00017_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[13] ));
 sg13g2_dfrbp_1 _11203_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net344),
    .D(_00613_),
    .Q_N(_00013_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[14] ));
 sg13g2_dfrbp_1 _11204_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net343),
    .D(_00614_),
    .Q_N(_00009_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[15] ));
 sg13g2_dfrbp_1 _11205_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net342),
    .D(_00615_),
    .Q_N(_00005_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[16] ));
 sg13g2_dfrbp_1 _11206_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net341),
    .D(_00616_),
    .Q_N(_00067_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[17] ));
 sg13g2_dfrbp_1 _11207_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net340),
    .D(_00617_),
    .Q_N(_00069_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[18] ));
 sg13g2_dfrbp_1 _11208_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net339),
    .D(_00618_),
    .Q_N(_00071_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[19] ));
 sg13g2_dfrbp_1 _11209_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net338),
    .D(_00619_),
    .Q_N(_00073_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[20] ));
 sg13g2_dfrbp_1 _11210_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net337),
    .D(_00620_),
    .Q_N(_00075_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[21] ));
 sg13g2_dfrbp_1 _11211_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net336),
    .D(_00621_),
    .Q_N(_00077_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[22] ));
 sg13g2_dfrbp_1 _11212_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net335),
    .D(_00622_),
    .Q_N(_00079_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[23] ));
 sg13g2_dfrbp_1 _11213_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net334),
    .D(_00623_),
    .Q_N(_00081_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[24] ));
 sg13g2_dfrbp_1 _11214_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net333),
    .D(_00624_),
    .Q_N(_00083_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[25] ));
 sg13g2_dfrbp_1 _11215_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net332),
    .D(_00625_),
    .Q_N(_00085_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[26] ));
 sg13g2_dfrbp_1 _11216_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net331),
    .D(_00626_),
    .Q_N(_00087_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[27] ));
 sg13g2_dfrbp_1 _11217_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net330),
    .D(_00627_),
    .Q_N(_00089_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[28] ));
 sg13g2_dfrbp_1 _11218_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net329),
    .D(_00628_),
    .Q_N(_00091_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[29] ));
 sg13g2_dfrbp_1 _11219_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net328),
    .D(_00629_),
    .Q_N(_00096_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[30] ));
 sg13g2_dfrbp_1 _11220_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net327),
    .D(_00630_),
    .Q_N(_00094_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbData[31] ));
 sg13g2_dfrbp_1 _11221_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net326),
    .D(_00631_),
    .Q_N(_04907_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbDest[0] ));
 sg13g2_dfrbp_1 _11222_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net325),
    .D(_00632_),
    .Q_N(_04906_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbDest[1] ));
 sg13g2_dfrbp_1 _11223_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net324),
    .D(_00633_),
    .Q_N(_04905_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbDest[2] ));
 sg13g2_dfrbp_1 _11224_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net323),
    .D(_00634_),
    .Q_N(_04904_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbDest[3] ));
 sg13g2_dfrbp_1 _11225_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net322),
    .D(_00635_),
    .Q_N(_04903_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_wbDest[4] ));
 sg13g2_dfrbp_1 _11226_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net321),
    .D(_00636_),
    .Q_N(_04902_),
    .Q(\ChiselTop.wild.cpu.exFwdReg_valid ));
 sg13g2_dfrbp_1 _11227_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net320),
    .D(_00637_),
    .Q_N(\ChiselTop._cntReg_T_1[0] ),
    .Q(\ChiselTop.cntReg[0] ));
 sg13g2_dfrbp_1 _11228_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net319),
    .D(net1462),
    .Q_N(_04901_),
    .Q(\ChiselTop.cntReg[1] ));
 sg13g2_dfrbp_1 _11229_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net318),
    .D(net1402),
    .Q_N(_04900_),
    .Q(\ChiselTop.cntReg[2] ));
 sg13g2_dfrbp_1 _11230_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net317),
    .D(_00640_),
    .Q_N(_04899_),
    .Q(\ChiselTop.cntReg[3] ));
 sg13g2_dfrbp_1 _11231_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net316),
    .D(_00641_),
    .Q_N(_04898_),
    .Q(\ChiselTop.cntReg[4] ));
 sg13g2_dfrbp_1 _11232_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net315),
    .D(_00642_),
    .Q_N(_04897_),
    .Q(\ChiselTop.cntReg[5] ));
 sg13g2_dfrbp_1 _11233_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net314),
    .D(net1164),
    .Q_N(_04896_),
    .Q(\ChiselTop.cntReg[6] ));
 sg13g2_dfrbp_1 _11234_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net313),
    .D(_00644_),
    .Q_N(_04895_),
    .Q(\ChiselTop.cntReg[7] ));
 sg13g2_dfrbp_1 _11235_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net312),
    .D(_00645_),
    .Q_N(_04894_),
    .Q(\ChiselTop.cntReg[8] ));
 sg13g2_dfrbp_1 _11236_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net311),
    .D(_00646_),
    .Q_N(_04893_),
    .Q(\ChiselTop.cntReg[9] ));
 sg13g2_dfrbp_1 _11237_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net310),
    .D(_00647_),
    .Q_N(_04892_),
    .Q(\ChiselTop.cntReg[10] ));
 sg13g2_dfrbp_1 _11238_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net309),
    .D(_00648_),
    .Q_N(_04891_),
    .Q(\ChiselTop.cntReg[11] ));
 sg13g2_dfrbp_1 _11239_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net308),
    .D(_00649_),
    .Q_N(_04890_),
    .Q(\ChiselTop.cntReg[12] ));
 sg13g2_dfrbp_1 _11240_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net307),
    .D(_00650_),
    .Q_N(_04889_),
    .Q(\ChiselTop.cntReg[13] ));
 sg13g2_dfrbp_1 _11241_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net306),
    .D(_00651_),
    .Q_N(_04888_),
    .Q(\ChiselTop.cntReg[14] ));
 sg13g2_dfrbp_1 _11242_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net305),
    .D(_00652_),
    .Q_N(_04887_),
    .Q(\ChiselTop.cntReg[15] ));
 sg13g2_dfrbp_1 _11243_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net304),
    .D(_00653_),
    .Q_N(_04886_),
    .Q(\ChiselTop.cntReg[16] ));
 sg13g2_dfrbp_1 _11244_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net303),
    .D(_00654_),
    .Q_N(_04885_),
    .Q(\ChiselTop.cntReg[17] ));
 sg13g2_dfrbp_1 _11245_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net302),
    .D(_00655_),
    .Q_N(_04884_),
    .Q(\ChiselTop.cntReg[18] ));
 sg13g2_dfrbp_1 _11246_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net301),
    .D(_00656_),
    .Q_N(_04883_),
    .Q(\ChiselTop.cntReg[19] ));
 sg13g2_dfrbp_1 _11247_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net300),
    .D(_00657_),
    .Q_N(_04882_),
    .Q(\ChiselTop.cntReg[20] ));
 sg13g2_dfrbp_1 _11248_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net299),
    .D(net1418),
    .Q_N(_04881_),
    .Q(\ChiselTop.cntReg[21] ));
 sg13g2_dfrbp_1 _11249_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net298),
    .D(_00659_),
    .Q_N(_04880_),
    .Q(\ChiselTop.cntReg[22] ));
 sg13g2_dfrbp_1 _11250_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net297),
    .D(_00660_),
    .Q_N(_04879_),
    .Q(\ChiselTop.cntReg[23] ));
 sg13g2_dfrbp_1 _11251_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net296),
    .D(net1099),
    .Q_N(_04878_),
    .Q(\ChiselTop.cntReg[24] ));
 sg13g2_dfrbp_1 _11252_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net295),
    .D(_00662_),
    .Q_N(_04877_),
    .Q(\ChiselTop.cntReg[25] ));
 sg13g2_dfrbp_1 _11253_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net294),
    .D(_00663_),
    .Q_N(_04876_),
    .Q(\ChiselTop.cntReg[26] ));
 sg13g2_dfrbp_1 _11254_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net293),
    .D(net1156),
    .Q_N(_04875_),
    .Q(\ChiselTop.cntReg[27] ));
 sg13g2_dfrbp_1 _11255_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net292),
    .D(_00665_),
    .Q_N(_04874_),
    .Q(\ChiselTop.cntReg[28] ));
 sg13g2_dfrbp_1 _11256_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net291),
    .D(_00666_),
    .Q_N(_04873_),
    .Q(\ChiselTop.cntReg[29] ));
 sg13g2_dfrbp_1 _11257_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net290),
    .D(net1305),
    .Q_N(_04872_),
    .Q(\ChiselTop.cntReg[30] ));
 sg13g2_dfrbp_1 _11258_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net633),
    .D(_00668_),
    .Q_N(_05322_),
    .Q(\ChiselTop.cntReg[31] ));
 sg13g2_dfrbp_1 _11259_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net634),
    .D(\ChiselTop.wild.cpu.io_imem_data[20] ),
    .Q_N(_05323_),
    .Q(\ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[0] ));
 sg13g2_dfrbp_1 _11260_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net817),
    .D(\ChiselTop.wild.cpu.io_imem_data[21] ),
    .Q_N(_05324_),
    .Q(\ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[1] ));
 sg13g2_dfrbp_1 _11261_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net289),
    .D(\ChiselTop.wild.cpu.io_imem_data[22] ),
    .Q_N(_00138_),
    .Q(\ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[2] ));
 sg13g2_dfrbp_1 _11262_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net288),
    .D(_00669_),
    .Q_N(_04871_),
    .Q(\ChiselTop.wild.cpu.regs[7][0] ));
 sg13g2_dfrbp_1 _11263_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net287),
    .D(_00670_),
    .Q_N(_04870_),
    .Q(\ChiselTop.wild.cpu.regs[7][1] ));
 sg13g2_dfrbp_1 _11264_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net286),
    .D(_00671_),
    .Q_N(_04869_),
    .Q(\ChiselTop.wild.cpu.regs[7][2] ));
 sg13g2_dfrbp_1 _11265_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net285),
    .D(_00672_),
    .Q_N(_04868_),
    .Q(\ChiselTop.wild.cpu.regs[7][3] ));
 sg13g2_dfrbp_1 _11266_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net284),
    .D(_00673_),
    .Q_N(_04867_),
    .Q(\ChiselTop.wild.cpu.regs[7][4] ));
 sg13g2_dfrbp_1 _11267_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net283),
    .D(_00674_),
    .Q_N(_04866_),
    .Q(\ChiselTop.wild.cpu.regs[7][5] ));
 sg13g2_dfrbp_1 _11268_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net282),
    .D(_00675_),
    .Q_N(_04865_),
    .Q(\ChiselTop.wild.cpu.regs[7][6] ));
 sg13g2_dfrbp_1 _11269_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net281),
    .D(_00676_),
    .Q_N(_04864_),
    .Q(\ChiselTop.wild.cpu.regs[7][7] ));
 sg13g2_dfrbp_1 _11270_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net280),
    .D(_00677_),
    .Q_N(_04863_),
    .Q(\ChiselTop.wild.cpu.regs[7][8] ));
 sg13g2_dfrbp_1 _11271_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net279),
    .D(_00678_),
    .Q_N(_04862_),
    .Q(\ChiselTop.wild.cpu.regs[7][9] ));
 sg13g2_dfrbp_1 _11272_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net278),
    .D(_00679_),
    .Q_N(_04861_),
    .Q(\ChiselTop.wild.cpu.regs[7][10] ));
 sg13g2_dfrbp_1 _11273_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net277),
    .D(_00680_),
    .Q_N(_04860_),
    .Q(\ChiselTop.wild.cpu.regs[7][11] ));
 sg13g2_dfrbp_1 _11274_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net276),
    .D(_00681_),
    .Q_N(_04859_),
    .Q(\ChiselTop.wild.cpu.regs[7][12] ));
 sg13g2_dfrbp_1 _11275_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net275),
    .D(_00682_),
    .Q_N(_04858_),
    .Q(\ChiselTop.wild.cpu.regs[7][13] ));
 sg13g2_dfrbp_1 _11276_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net274),
    .D(_00683_),
    .Q_N(_04857_),
    .Q(\ChiselTop.wild.cpu.regs[7][14] ));
 sg13g2_dfrbp_1 _11277_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net273),
    .D(_00684_),
    .Q_N(_04856_),
    .Q(\ChiselTop.wild.cpu.regs[7][15] ));
 sg13g2_dfrbp_1 _11278_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net272),
    .D(_00685_),
    .Q_N(_04855_),
    .Q(\ChiselTop.wild.cpu.regs[7][16] ));
 sg13g2_dfrbp_1 _11279_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net271),
    .D(_00686_),
    .Q_N(_04854_),
    .Q(\ChiselTop.wild.cpu.regs[7][17] ));
 sg13g2_dfrbp_1 _11280_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net270),
    .D(_00687_),
    .Q_N(_04853_),
    .Q(\ChiselTop.wild.cpu.regs[7][18] ));
 sg13g2_dfrbp_1 _11281_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net269),
    .D(_00688_),
    .Q_N(_04852_),
    .Q(\ChiselTop.wild.cpu.regs[7][19] ));
 sg13g2_dfrbp_1 _11282_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net268),
    .D(_00689_),
    .Q_N(_04851_),
    .Q(\ChiselTop.wild.cpu.regs[7][20] ));
 sg13g2_dfrbp_1 _11283_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net267),
    .D(_00690_),
    .Q_N(_04850_),
    .Q(\ChiselTop.wild.cpu.regs[7][21] ));
 sg13g2_dfrbp_1 _11284_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net266),
    .D(_00691_),
    .Q_N(_04849_),
    .Q(\ChiselTop.wild.cpu.regs[7][22] ));
 sg13g2_dfrbp_1 _11285_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net265),
    .D(_00692_),
    .Q_N(_04848_),
    .Q(\ChiselTop.wild.cpu.regs[7][23] ));
 sg13g2_dfrbp_1 _11286_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net264),
    .D(_00693_),
    .Q_N(_04847_),
    .Q(\ChiselTop.wild.cpu.regs[7][24] ));
 sg13g2_dfrbp_1 _11287_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net263),
    .D(_00694_),
    .Q_N(_04846_),
    .Q(\ChiselTop.wild.cpu.regs[7][25] ));
 sg13g2_dfrbp_1 _11288_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net262),
    .D(_00695_),
    .Q_N(_04845_),
    .Q(\ChiselTop.wild.cpu.regs[7][26] ));
 sg13g2_dfrbp_1 _11289_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net261),
    .D(_00696_),
    .Q_N(_04844_),
    .Q(\ChiselTop.wild.cpu.regs[7][27] ));
 sg13g2_dfrbp_1 _11290_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net260),
    .D(_00697_),
    .Q_N(_04843_),
    .Q(\ChiselTop.wild.cpu.regs[7][28] ));
 sg13g2_dfrbp_1 _11291_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net259),
    .D(_00698_),
    .Q_N(_04842_),
    .Q(\ChiselTop.wild.cpu.regs[7][29] ));
 sg13g2_dfrbp_1 _11292_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net258),
    .D(_00699_),
    .Q_N(_04841_),
    .Q(\ChiselTop.wild.cpu.regs[7][30] ));
 sg13g2_dfrbp_1 _11293_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net257),
    .D(_00700_),
    .Q_N(_04840_),
    .Q(\ChiselTop.wild.cpu.regs[7][31] ));
 sg13g2_dfrbp_1 _11294_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net256),
    .D(_00701_),
    .Q_N(_04839_),
    .Q(\ChiselTop.wild.dmem.MEM_3[0][0] ));
 sg13g2_dfrbp_1 _11295_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net255),
    .D(_00702_),
    .Q_N(_04838_),
    .Q(\ChiselTop.wild.dmem.MEM_3[0][1] ));
 sg13g2_dfrbp_1 _11296_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net254),
    .D(_00703_),
    .Q_N(_04837_),
    .Q(\ChiselTop.wild.dmem.MEM_3[0][2] ));
 sg13g2_dfrbp_1 _11297_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net253),
    .D(_00704_),
    .Q_N(_04836_),
    .Q(\ChiselTop.wild.dmem.MEM_3[0][3] ));
 sg13g2_dfrbp_1 _11298_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net252),
    .D(_00705_),
    .Q_N(_04835_),
    .Q(\ChiselTop.wild.dmem.MEM_3[0][4] ));
 sg13g2_dfrbp_1 _11299_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net251),
    .D(_00706_),
    .Q_N(_04834_),
    .Q(\ChiselTop.wild.dmem.MEM_3[0][5] ));
 sg13g2_dfrbp_1 _11300_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net250),
    .D(_00707_),
    .Q_N(_04833_),
    .Q(\ChiselTop.wild.dmem.MEM_3[0][6] ));
 sg13g2_dfrbp_1 _11301_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net249),
    .D(_00708_),
    .Q_N(_04832_),
    .Q(\ChiselTop.wild.dmem.MEM_3[0][7] ));
 sg13g2_dfrbp_1 _11302_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net248),
    .D(_00709_),
    .Q_N(_04831_),
    .Q(\ChiselTop.wild.cpu.regs[6][0] ));
 sg13g2_dfrbp_1 _11303_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net247),
    .D(_00710_),
    .Q_N(_04830_),
    .Q(\ChiselTop.wild.cpu.regs[6][1] ));
 sg13g2_dfrbp_1 _11304_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net246),
    .D(_00711_),
    .Q_N(_04829_),
    .Q(\ChiselTop.wild.cpu.regs[6][2] ));
 sg13g2_dfrbp_1 _11305_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net245),
    .D(_00712_),
    .Q_N(_04828_),
    .Q(\ChiselTop.wild.cpu.regs[6][3] ));
 sg13g2_dfrbp_1 _11306_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net244),
    .D(_00713_),
    .Q_N(_04827_),
    .Q(\ChiselTop.wild.cpu.regs[6][4] ));
 sg13g2_dfrbp_1 _11307_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net243),
    .D(_00714_),
    .Q_N(_04826_),
    .Q(\ChiselTop.wild.cpu.regs[6][5] ));
 sg13g2_dfrbp_1 _11308_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net242),
    .D(_00715_),
    .Q_N(_04825_),
    .Q(\ChiselTop.wild.cpu.regs[6][6] ));
 sg13g2_dfrbp_1 _11309_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net241),
    .D(_00716_),
    .Q_N(_04824_),
    .Q(\ChiselTop.wild.cpu.regs[6][7] ));
 sg13g2_dfrbp_1 _11310_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net240),
    .D(_00717_),
    .Q_N(_04823_),
    .Q(\ChiselTop.wild.cpu.regs[6][8] ));
 sg13g2_dfrbp_1 _11311_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net239),
    .D(_00718_),
    .Q_N(_04822_),
    .Q(\ChiselTop.wild.cpu.regs[6][9] ));
 sg13g2_dfrbp_1 _11312_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net238),
    .D(_00719_),
    .Q_N(_04821_),
    .Q(\ChiselTop.wild.cpu.regs[6][10] ));
 sg13g2_dfrbp_1 _11313_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net237),
    .D(_00720_),
    .Q_N(_04820_),
    .Q(\ChiselTop.wild.cpu.regs[6][11] ));
 sg13g2_dfrbp_1 _11314_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net236),
    .D(_00721_),
    .Q_N(_04819_),
    .Q(\ChiselTop.wild.cpu.regs[6][12] ));
 sg13g2_dfrbp_1 _11315_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net235),
    .D(_00722_),
    .Q_N(_04818_),
    .Q(\ChiselTop.wild.cpu.regs[6][13] ));
 sg13g2_dfrbp_1 _11316_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net234),
    .D(_00723_),
    .Q_N(_04817_),
    .Q(\ChiselTop.wild.cpu.regs[6][14] ));
 sg13g2_dfrbp_1 _11317_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net233),
    .D(_00724_),
    .Q_N(_04816_),
    .Q(\ChiselTop.wild.cpu.regs[6][15] ));
 sg13g2_dfrbp_1 _11318_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net232),
    .D(_00725_),
    .Q_N(_04815_),
    .Q(\ChiselTop.wild.cpu.regs[6][16] ));
 sg13g2_dfrbp_1 _11319_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net231),
    .D(_00726_),
    .Q_N(_04814_),
    .Q(\ChiselTop.wild.cpu.regs[6][17] ));
 sg13g2_dfrbp_1 _11320_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net230),
    .D(_00727_),
    .Q_N(_04813_),
    .Q(\ChiselTop.wild.cpu.regs[6][18] ));
 sg13g2_dfrbp_1 _11321_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net229),
    .D(_00728_),
    .Q_N(_04812_),
    .Q(\ChiselTop.wild.cpu.regs[6][19] ));
 sg13g2_dfrbp_1 _11322_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net228),
    .D(_00729_),
    .Q_N(_04811_),
    .Q(\ChiselTop.wild.cpu.regs[6][20] ));
 sg13g2_dfrbp_1 _11323_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net227),
    .D(_00730_),
    .Q_N(_04810_),
    .Q(\ChiselTop.wild.cpu.regs[6][21] ));
 sg13g2_dfrbp_1 _11324_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net226),
    .D(_00731_),
    .Q_N(_04809_),
    .Q(\ChiselTop.wild.cpu.regs[6][22] ));
 sg13g2_dfrbp_1 _11325_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net225),
    .D(_00732_),
    .Q_N(_04808_),
    .Q(\ChiselTop.wild.cpu.regs[6][23] ));
 sg13g2_dfrbp_1 _11326_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net224),
    .D(_00733_),
    .Q_N(_04807_),
    .Q(\ChiselTop.wild.cpu.regs[6][24] ));
 sg13g2_dfrbp_1 _11327_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net223),
    .D(_00734_),
    .Q_N(_04806_),
    .Q(\ChiselTop.wild.cpu.regs[6][25] ));
 sg13g2_dfrbp_1 _11328_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net222),
    .D(_00735_),
    .Q_N(_04805_),
    .Q(\ChiselTop.wild.cpu.regs[6][26] ));
 sg13g2_dfrbp_1 _11329_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net221),
    .D(_00736_),
    .Q_N(_04804_),
    .Q(\ChiselTop.wild.cpu.regs[6][27] ));
 sg13g2_dfrbp_1 _11330_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net220),
    .D(_00737_),
    .Q_N(_04803_),
    .Q(\ChiselTop.wild.cpu.regs[6][28] ));
 sg13g2_dfrbp_1 _11331_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net219),
    .D(_00738_),
    .Q_N(_04802_),
    .Q(\ChiselTop.wild.cpu.regs[6][29] ));
 sg13g2_dfrbp_1 _11332_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net218),
    .D(_00739_),
    .Q_N(_04801_),
    .Q(\ChiselTop.wild.cpu.regs[6][30] ));
 sg13g2_dfrbp_1 _11333_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net217),
    .D(_00740_),
    .Q_N(_04800_),
    .Q(\ChiselTop.wild.cpu.regs[6][31] ));
 sg13g2_dfrbp_1 _11334_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net216),
    .D(_00741_),
    .Q_N(_04799_),
    .Q(\ChiselTop.wild.cpu.regs[5][0] ));
 sg13g2_dfrbp_1 _11335_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net215),
    .D(_00742_),
    .Q_N(_04798_),
    .Q(\ChiselTop.wild.cpu.regs[5][1] ));
 sg13g2_dfrbp_1 _11336_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net214),
    .D(_00743_),
    .Q_N(_04797_),
    .Q(\ChiselTop.wild.cpu.regs[5][2] ));
 sg13g2_dfrbp_1 _11337_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net213),
    .D(_00744_),
    .Q_N(_04796_),
    .Q(\ChiselTop.wild.cpu.regs[5][3] ));
 sg13g2_dfrbp_1 _11338_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net212),
    .D(_00745_),
    .Q_N(_04795_),
    .Q(\ChiselTop.wild.cpu.regs[5][4] ));
 sg13g2_dfrbp_1 _11339_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net211),
    .D(_00746_),
    .Q_N(_04794_),
    .Q(\ChiselTop.wild.cpu.regs[5][5] ));
 sg13g2_dfrbp_1 _11340_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net210),
    .D(_00747_),
    .Q_N(_04793_),
    .Q(\ChiselTop.wild.cpu.regs[5][6] ));
 sg13g2_dfrbp_1 _11341_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net209),
    .D(_00748_),
    .Q_N(_04792_),
    .Q(\ChiselTop.wild.cpu.regs[5][7] ));
 sg13g2_dfrbp_1 _11342_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net208),
    .D(_00749_),
    .Q_N(_04791_),
    .Q(\ChiselTop.wild.cpu.regs[5][8] ));
 sg13g2_dfrbp_1 _11343_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net207),
    .D(_00750_),
    .Q_N(_04790_),
    .Q(\ChiselTop.wild.cpu.regs[5][9] ));
 sg13g2_dfrbp_1 _11344_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net206),
    .D(_00751_),
    .Q_N(_04789_),
    .Q(\ChiselTop.wild.cpu.regs[5][10] ));
 sg13g2_dfrbp_1 _11345_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net205),
    .D(_00752_),
    .Q_N(_04788_),
    .Q(\ChiselTop.wild.cpu.regs[5][11] ));
 sg13g2_dfrbp_1 _11346_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net204),
    .D(_00753_),
    .Q_N(_04787_),
    .Q(\ChiselTop.wild.cpu.regs[5][12] ));
 sg13g2_dfrbp_1 _11347_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net203),
    .D(_00754_),
    .Q_N(_04786_),
    .Q(\ChiselTop.wild.cpu.regs[5][13] ));
 sg13g2_dfrbp_1 _11348_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net202),
    .D(_00755_),
    .Q_N(_04785_),
    .Q(\ChiselTop.wild.cpu.regs[5][14] ));
 sg13g2_dfrbp_1 _11349_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net201),
    .D(_00756_),
    .Q_N(_04784_),
    .Q(\ChiselTop.wild.cpu.regs[5][15] ));
 sg13g2_dfrbp_1 _11350_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net200),
    .D(_00757_),
    .Q_N(_04783_),
    .Q(\ChiselTop.wild.cpu.regs[5][16] ));
 sg13g2_dfrbp_1 _11351_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net199),
    .D(_00758_),
    .Q_N(_04782_),
    .Q(\ChiselTop.wild.cpu.regs[5][17] ));
 sg13g2_dfrbp_1 _11352_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net198),
    .D(_00759_),
    .Q_N(_04781_),
    .Q(\ChiselTop.wild.cpu.regs[5][18] ));
 sg13g2_dfrbp_1 _11353_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net197),
    .D(_00760_),
    .Q_N(_04780_),
    .Q(\ChiselTop.wild.cpu.regs[5][19] ));
 sg13g2_dfrbp_1 _11354_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net196),
    .D(_00761_),
    .Q_N(_04779_),
    .Q(\ChiselTop.wild.cpu.regs[5][20] ));
 sg13g2_dfrbp_1 _11355_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net195),
    .D(_00762_),
    .Q_N(_04778_),
    .Q(\ChiselTop.wild.cpu.regs[5][21] ));
 sg13g2_dfrbp_1 _11356_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net194),
    .D(_00763_),
    .Q_N(_04777_),
    .Q(\ChiselTop.wild.cpu.regs[5][22] ));
 sg13g2_dfrbp_1 _11357_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net193),
    .D(_00764_),
    .Q_N(_04776_),
    .Q(\ChiselTop.wild.cpu.regs[5][23] ));
 sg13g2_dfrbp_1 _11358_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net192),
    .D(_00765_),
    .Q_N(_04775_),
    .Q(\ChiselTop.wild.cpu.regs[5][24] ));
 sg13g2_dfrbp_1 _11359_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net191),
    .D(_00766_),
    .Q_N(_04774_),
    .Q(\ChiselTop.wild.cpu.regs[5][25] ));
 sg13g2_dfrbp_1 _11360_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net190),
    .D(_00767_),
    .Q_N(_04773_),
    .Q(\ChiselTop.wild.cpu.regs[5][26] ));
 sg13g2_dfrbp_1 _11361_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net189),
    .D(_00768_),
    .Q_N(_04772_),
    .Q(\ChiselTop.wild.cpu.regs[5][27] ));
 sg13g2_dfrbp_1 _11362_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net188),
    .D(_00769_),
    .Q_N(_04771_),
    .Q(\ChiselTop.wild.cpu.regs[5][28] ));
 sg13g2_dfrbp_1 _11363_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net187),
    .D(_00770_),
    .Q_N(_04770_),
    .Q(\ChiselTop.wild.cpu.regs[5][29] ));
 sg13g2_dfrbp_1 _11364_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net186),
    .D(_00771_),
    .Q_N(_04769_),
    .Q(\ChiselTop.wild.cpu.regs[5][30] ));
 sg13g2_dfrbp_1 _11365_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net185),
    .D(_00772_),
    .Q_N(_04768_),
    .Q(\ChiselTop.wild.cpu.regs[5][31] ));
 sg13g2_dfrbp_1 _11366_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net184),
    .D(_00773_),
    .Q_N(_00137_),
    .Q(\ChiselTop.wild.cpu.pcReg[2] ));
 sg13g2_dfrbp_1 _11367_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net183),
    .D(_00774_),
    .Q_N(_04767_),
    .Q(\ChiselTop.wild.cpu.pcReg[3] ));
 sg13g2_dfrbp_1 _11368_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net182),
    .D(_00775_),
    .Q_N(_04766_),
    .Q(\ChiselTop.wild.cpu.pcReg[4] ));
 sg13g2_dfrbp_1 _11369_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net181),
    .D(_00776_),
    .Q_N(_04765_),
    .Q(\ChiselTop.wild.cpu.pcReg[5] ));
 sg13g2_dfrbp_1 _11370_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net180),
    .D(_00777_),
    .Q_N(_04764_),
    .Q(\ChiselTop.wild.cpu.pcReg[6] ));
 sg13g2_dfrbp_1 _11371_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net179),
    .D(_00778_),
    .Q_N(_04763_),
    .Q(\ChiselTop.wild.cpu.pcReg[7] ));
 sg13g2_dfrbp_1 _11372_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net178),
    .D(_00779_),
    .Q_N(_04762_),
    .Q(\ChiselTop.wild.cpu.pcReg[8] ));
 sg13g2_dfrbp_1 _11373_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net177),
    .D(_00780_),
    .Q_N(_04761_),
    .Q(\ChiselTop.wild.cpu.pcReg[9] ));
 sg13g2_dfrbp_1 _11374_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net176),
    .D(_00781_),
    .Q_N(_04760_),
    .Q(\ChiselTop.wild.cpu.pcReg[10] ));
 sg13g2_dfrbp_1 _11375_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net175),
    .D(net1398),
    .Q_N(_04759_),
    .Q(\ChiselTop.wild.cpu.pcReg[11] ));
 sg13g2_dfrbp_1 _11376_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net174),
    .D(_00783_),
    .Q_N(_04758_),
    .Q(\ChiselTop.wild.cpu.pcReg[12] ));
 sg13g2_dfrbp_1 _11377_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net173),
    .D(_00784_),
    .Q_N(_04757_),
    .Q(\ChiselTop.wild.cpu.pcReg[13] ));
 sg13g2_dfrbp_1 _11378_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net172),
    .D(_00785_),
    .Q_N(_04756_),
    .Q(\ChiselTop.wild.cpu.pcReg[14] ));
 sg13g2_dfrbp_1 _11379_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net171),
    .D(_00786_),
    .Q_N(_04755_),
    .Q(\ChiselTop.wild.cpu.pcReg[15] ));
 sg13g2_dfrbp_1 _11380_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net170),
    .D(_00787_),
    .Q_N(_04754_),
    .Q(\ChiselTop.wild.cpu.pcReg[16] ));
 sg13g2_dfrbp_1 _11381_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net169),
    .D(_00788_),
    .Q_N(_04753_),
    .Q(\ChiselTop.wild.cpu.pcReg[17] ));
 sg13g2_dfrbp_1 _11382_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net168),
    .D(_00789_),
    .Q_N(_04752_),
    .Q(\ChiselTop.wild.cpu.pcReg[18] ));
 sg13g2_dfrbp_1 _11383_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net167),
    .D(_00790_),
    .Q_N(_04751_),
    .Q(\ChiselTop.wild.cpu.pcReg[19] ));
 sg13g2_dfrbp_1 _11384_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net166),
    .D(_00791_),
    .Q_N(_04750_),
    .Q(\ChiselTop.wild.cpu.pcReg[20] ));
 sg13g2_dfrbp_1 _11385_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net165),
    .D(_00792_),
    .Q_N(_04749_),
    .Q(\ChiselTop.wild.cpu.pcReg[21] ));
 sg13g2_dfrbp_1 _11386_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net164),
    .D(_00793_),
    .Q_N(_04748_),
    .Q(\ChiselTop.wild.cpu.pcReg[22] ));
 sg13g2_dfrbp_1 _11387_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net163),
    .D(_00794_),
    .Q_N(_04747_),
    .Q(\ChiselTop.wild.cpu.pcReg[23] ));
 sg13g2_dfrbp_1 _11388_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net162),
    .D(_00795_),
    .Q_N(_04746_),
    .Q(\ChiselTop.wild.cpu.pcReg[24] ));
 sg13g2_dfrbp_1 _11389_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net161),
    .D(_00796_),
    .Q_N(_04745_),
    .Q(\ChiselTop.wild.cpu.pcReg[25] ));
 sg13g2_dfrbp_1 _11390_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net160),
    .D(_00797_),
    .Q_N(_04744_),
    .Q(\ChiselTop.wild.cpu.pcReg[26] ));
 sg13g2_dfrbp_1 _11391_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net159),
    .D(_00798_),
    .Q_N(_04743_),
    .Q(\ChiselTop.wild.cpu.pcReg[27] ));
 sg13g2_dfrbp_1 _11392_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net158),
    .D(net1477),
    .Q_N(_04742_),
    .Q(\ChiselTop.wild.cpu.pcReg[28] ));
 sg13g2_dfrbp_1 _11393_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net157),
    .D(_00800_),
    .Q_N(_04741_),
    .Q(\ChiselTop.wild.cpu.pcReg[29] ));
 sg13g2_dfrbp_1 _11394_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net156),
    .D(_00801_),
    .Q_N(_04740_),
    .Q(\ChiselTop.wild.cpu.pcReg[30] ));
 sg13g2_dfrbp_1 _11395_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net155),
    .D(_00802_),
    .Q_N(_04739_),
    .Q(\ChiselTop.wild.cpu.pcReg[31] ));
 sg13g2_dfrbp_1 _11396_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net154),
    .D(_00803_),
    .Q_N(_04738_),
    .Q(\ChiselTop.wild.cpu.regs[0][0] ));
 sg13g2_dfrbp_1 _11397_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net153),
    .D(_00804_),
    .Q_N(_04737_),
    .Q(\ChiselTop.wild.cpu.regs[0][1] ));
 sg13g2_dfrbp_1 _11398_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net152),
    .D(_00805_),
    .Q_N(_04736_),
    .Q(\ChiselTop.wild.cpu.regs[0][2] ));
 sg13g2_dfrbp_1 _11399_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net151),
    .D(_00806_),
    .Q_N(_04735_),
    .Q(\ChiselTop.wild.cpu.regs[0][3] ));
 sg13g2_dfrbp_1 _11400_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net150),
    .D(_00807_),
    .Q_N(_04734_),
    .Q(\ChiselTop.wild.cpu.regs[0][4] ));
 sg13g2_dfrbp_1 _11401_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net149),
    .D(_00808_),
    .Q_N(_04733_),
    .Q(\ChiselTop.wild.cpu.regs[0][5] ));
 sg13g2_dfrbp_1 _11402_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net148),
    .D(_00809_),
    .Q_N(_04732_),
    .Q(\ChiselTop.wild.cpu.regs[0][6] ));
 sg13g2_dfrbp_1 _11403_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net147),
    .D(_00810_),
    .Q_N(_04731_),
    .Q(\ChiselTop.wild.cpu.regs[0][7] ));
 sg13g2_dfrbp_1 _11404_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(_00811_),
    .Q_N(_04730_),
    .Q(\ChiselTop.wild.cpu.regs[0][8] ));
 sg13g2_dfrbp_1 _11405_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net145),
    .D(_00812_),
    .Q_N(_04729_),
    .Q(\ChiselTop.wild.cpu.regs[0][9] ));
 sg13g2_dfrbp_1 _11406_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net144),
    .D(_00813_),
    .Q_N(_04728_),
    .Q(\ChiselTop.wild.cpu.regs[0][10] ));
 sg13g2_dfrbp_1 _11407_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net143),
    .D(_00814_),
    .Q_N(_04727_),
    .Q(\ChiselTop.wild.cpu.regs[0][11] ));
 sg13g2_dfrbp_1 _11408_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net142),
    .D(_00815_),
    .Q_N(_04726_),
    .Q(\ChiselTop.wild.cpu.regs[0][12] ));
 sg13g2_dfrbp_1 _11409_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net141),
    .D(_00816_),
    .Q_N(_04725_),
    .Q(\ChiselTop.wild.cpu.regs[0][13] ));
 sg13g2_dfrbp_1 _11410_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net140),
    .D(_00817_),
    .Q_N(_04724_),
    .Q(\ChiselTop.wild.cpu.regs[0][14] ));
 sg13g2_dfrbp_1 _11411_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net139),
    .D(_00818_),
    .Q_N(_04723_),
    .Q(\ChiselTop.wild.cpu.regs[0][15] ));
 sg13g2_dfrbp_1 _11412_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net138),
    .D(_00819_),
    .Q_N(_04722_),
    .Q(\ChiselTop.wild.cpu.regs[0][16] ));
 sg13g2_dfrbp_1 _11413_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net137),
    .D(_00820_),
    .Q_N(_04721_),
    .Q(\ChiselTop.wild.cpu.regs[0][17] ));
 sg13g2_dfrbp_1 _11414_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net136),
    .D(_00821_),
    .Q_N(_04720_),
    .Q(\ChiselTop.wild.cpu.regs[0][18] ));
 sg13g2_dfrbp_1 _11415_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net135),
    .D(_00822_),
    .Q_N(_04719_),
    .Q(\ChiselTop.wild.cpu.regs[0][19] ));
 sg13g2_dfrbp_1 _11416_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net134),
    .D(_00823_),
    .Q_N(_04718_),
    .Q(\ChiselTop.wild.cpu.regs[0][20] ));
 sg13g2_dfrbp_1 _11417_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net133),
    .D(_00824_),
    .Q_N(_04717_),
    .Q(\ChiselTop.wild.cpu.regs[0][21] ));
 sg13g2_dfrbp_1 _11418_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net132),
    .D(_00825_),
    .Q_N(_04716_),
    .Q(\ChiselTop.wild.cpu.regs[0][22] ));
 sg13g2_dfrbp_1 _11419_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net131),
    .D(_00826_),
    .Q_N(_04715_),
    .Q(\ChiselTop.wild.cpu.regs[0][23] ));
 sg13g2_dfrbp_1 _11420_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net130),
    .D(_00827_),
    .Q_N(_04714_),
    .Q(\ChiselTop.wild.cpu.regs[0][24] ));
 sg13g2_dfrbp_1 _11421_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net129),
    .D(_00828_),
    .Q_N(_04713_),
    .Q(\ChiselTop.wild.cpu.regs[0][25] ));
 sg13g2_dfrbp_1 _11422_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net128),
    .D(_00829_),
    .Q_N(_04712_),
    .Q(\ChiselTop.wild.cpu.regs[0][26] ));
 sg13g2_dfrbp_1 _11423_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net127),
    .D(_00830_),
    .Q_N(_04711_),
    .Q(\ChiselTop.wild.cpu.regs[0][27] ));
 sg13g2_dfrbp_1 _11424_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net126),
    .D(_00831_),
    .Q_N(_04710_),
    .Q(\ChiselTop.wild.cpu.regs[0][28] ));
 sg13g2_dfrbp_1 _11425_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net125),
    .D(_00832_),
    .Q_N(_04709_),
    .Q(\ChiselTop.wild.cpu.regs[0][29] ));
 sg13g2_dfrbp_1 _11426_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net124),
    .D(_00833_),
    .Q_N(_04708_),
    .Q(\ChiselTop.wild.cpu.regs[0][30] ));
 sg13g2_dfrbp_1 _11427_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net123),
    .D(_00834_),
    .Q_N(_04707_),
    .Q(\ChiselTop.wild.cpu.regs[0][31] ));
 sg13g2_dfrbp_1 _11428_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net122),
    .D(_00835_),
    .Q_N(_04706_),
    .Q(\ChiselTop.wild.rx._shiftReg_T_1[7] ));
 sg13g2_dfrbp_1 _11429_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net121),
    .D(_00836_),
    .Q_N(\ChiselTop.wild.tx.buf_.io_in_ready ),
    .Q(\ChiselTop.wild.tx.buf_.io_out_valid ));
 sg13g2_dfrbp_1 _11430_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net120),
    .D(_00837_),
    .Q_N(_04705_),
    .Q(\ChiselTop.wild.tx.tx.bitsReg[0] ));
 sg13g2_dfrbp_1 _11431_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net118),
    .D(net1429),
    .Q_N(_04704_),
    .Q(\ChiselTop.wild.tx.tx.bitsReg[1] ));
 sg13g2_dfrbp_1 _11432_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net116),
    .D(net1204),
    .Q_N(_04703_),
    .Q(\ChiselTop.wild.tx.tx.bitsReg[2] ));
 sg13g2_dfrbp_1 _11433_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net114),
    .D(_00840_),
    .Q_N(_04702_),
    .Q(\ChiselTop.wild.tx.tx.bitsReg[3] ));
 sg13g2_dfrbp_1 _11434_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net112),
    .D(_00841_),
    .Q_N(_04701_),
    .Q(\ChiselTop.wild.rx.io_channel_valid ));
 sg13g2_dfrbp_1 _11435_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net110),
    .D(_00842_),
    .Q_N(_04700_),
    .Q(\ChiselTop.wild.rx.bitsReg[0] ));
 sg13g2_dfrbp_1 _11436_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net108),
    .D(net1389),
    .Q_N(_04699_),
    .Q(\ChiselTop.wild.rx.bitsReg[1] ));
 sg13g2_dfrbp_1 _11437_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net106),
    .D(_00844_),
    .Q_N(_04698_),
    .Q(\ChiselTop.wild.rx.bitsReg[2] ));
 sg13g2_dfrbp_1 _11438_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net104),
    .D(_00845_),
    .Q_N(_04697_),
    .Q(\ChiselTop.wild.rx.bitsReg[3] ));
 sg13g2_dfrbp_1 _11439_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net102),
    .D(net1065),
    .Q_N(_04696_),
    .Q(\ChiselTop.wild.rx.io_channel_bits[0] ));
 sg13g2_dfrbp_1 _11440_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net100),
    .D(_00847_),
    .Q_N(_04695_),
    .Q(\ChiselTop.wild.rx._shiftReg_T_1[0] ));
 sg13g2_dfrbp_1 _11441_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net98),
    .D(net1277),
    .Q_N(_04694_),
    .Q(\ChiselTop.wild.rx._shiftReg_T_1[1] ));
 sg13g2_dfrbp_1 _11442_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net96),
    .D(net1384),
    .Q_N(_04693_),
    .Q(\ChiselTop.wild.rx._shiftReg_T_1[2] ));
 sg13g2_dfrbp_1 _11443_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net94),
    .D(_00850_),
    .Q_N(_04692_),
    .Q(\ChiselTop.wild.rx._shiftReg_T_1[3] ));
 sg13g2_dfrbp_1 _11444_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net92),
    .D(_00851_),
    .Q_N(_04691_),
    .Q(\ChiselTop.wild.rx._shiftReg_T_1[4] ));
 sg13g2_dfrbp_1 _11445_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net90),
    .D(net1186),
    .Q_N(_04690_),
    .Q(\ChiselTop.wild.rx._shiftReg_T_1[5] ));
 sg13g2_dfrbp_1 _11446_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net81),
    .D(_00853_),
    .Q_N(_05325_),
    .Q(\ChiselTop.wild.rx._shiftReg_T_1[6] ));
 sg13g2_dfrbp_1 _11447_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net88),
    .D(net864),
    .Q_N(_04689_),
    .Q(\ChiselTop.wild.rx.falling_REG ));
 sg13g2_dfrbp_1 _11448_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net86),
    .D(_00854_),
    .Q_N(_04688_),
    .Q(\ChiselTop.wild.rx.rxReg_REG ));
 sg13g2_dfrbp_1 _11449_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net85),
    .D(_00855_),
    .Q_N(_04687_),
    .Q(\ChiselTop.wild.cpu.decExReg_decOut_rfWrite ));
 sg13g2_dfrbp_1 _11450_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net84),
    .D(net870),
    .Q_N(_00139_),
    .Q(\ChiselTop.wild.rx.cntReg[0] ));
 sg13g2_dfrbp_1 _11451_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net82),
    .D(net1509),
    .Q_N(_04686_),
    .Q(\ChiselTop.wild.rx.cntReg[1] ));
 sg13g2_dfrbp_1 _11452_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net80),
    .D(_00858_),
    .Q_N(_04685_),
    .Q(\ChiselTop.wild.rx.cntReg[2] ));
 sg13g2_dfrbp_1 _11453_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net78),
    .D(_00859_),
    .Q_N(_04684_),
    .Q(\ChiselTop.wild.rx.cntReg[3] ));
 sg13g2_dfrbp_1 _11454_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net76),
    .D(net1227),
    .Q_N(_04683_),
    .Q(\ChiselTop.wild.rx.cntReg[4] ));
 sg13g2_dfrbp_1 _11455_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net74),
    .D(_00861_),
    .Q_N(_04682_),
    .Q(\ChiselTop.wild.rx.cntReg[5] ));
 sg13g2_dfrbp_1 _11456_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net72),
    .D(_00862_),
    .Q_N(_04681_),
    .Q(\ChiselTop.wild.rx.cntReg[6] ));
 sg13g2_dfrbp_1 _11457_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net68),
    .D(net1161),
    .Q_N(_04680_),
    .Q(\ChiselTop.wild.rx.cntReg[7] ));
 sg13g2_dfrbp_1 _11458_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net66),
    .D(net1408),
    .Q_N(_04679_),
    .Q(\ChiselTop.wild.rx.cntReg[8] ));
 sg13g2_dfrbp_1 _11459_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net556),
    .D(_00865_),
    .Q_N(_04678_),
    .Q(\ChiselTop.wild.rx.cntReg[9] ));
 sg13g2_dfrbp_1 _11460_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net552),
    .D(net1177),
    .Q_N(_04677_),
    .Q(\ChiselTop.wild.rx.cntReg[10] ));
 sg13g2_dfrbp_1 _11461_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net117),
    .D(_00867_),
    .Q_N(_04676_),
    .Q(\ChiselTop.wild.rx.cntReg[11] ));
 sg13g2_dfrbp_1 _11462_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net113),
    .D(_00868_),
    .Q_N(_04675_),
    .Q(\ChiselTop.wild.rx.cntReg[12] ));
 sg13g2_dfrbp_1 _11463_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net109),
    .D(net1059),
    .Q_N(_04674_),
    .Q(\ChiselTop.wild.rx.cntReg[13] ));
 sg13g2_dfrbp_1 _11464_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net105),
    .D(_00870_),
    .Q_N(_00140_),
    .Q(\ChiselTop.wild.rx.cntReg[14] ));
 sg13g2_dfrbp_1 _11465_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net101),
    .D(_00871_),
    .Q_N(_04673_),
    .Q(\ChiselTop.wild.rx.cntReg[15] ));
 sg13g2_dfrbp_1 _11466_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net97),
    .D(_00872_),
    .Q_N(_04672_),
    .Q(\ChiselTop.wild.rx.cntReg[16] ));
 sg13g2_dfrbp_1 _11467_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net93),
    .D(net1309),
    .Q_N(_04671_),
    .Q(\ChiselTop.wild.rx.cntReg[17] ));
 sg13g2_dfrbp_1 _11468_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net89),
    .D(_00874_),
    .Q_N(_00141_),
    .Q(\ChiselTop.wild.rx.cntReg[18] ));
 sg13g2_dfrbp_1 _11469_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net83),
    .D(_00875_),
    .Q_N(_04670_),
    .Q(\ChiselTop.wild.rx.cntReg[19] ));
 sg13g2_dfrbp_1 _11470_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net79),
    .D(_00876_),
    .Q_N(_04669_),
    .Q(\ChiselTop.wild.cpu.decOut_opcode[4] ));
 sg13g2_dfrbp_1 _11471_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net77),
    .D(_00877_),
    .Q_N(_04668_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[0] ));
 sg13g2_dfrbp_1 _11472_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net75),
    .D(_00878_),
    .Q_N(_00122_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[2] ));
 sg13g2_dfrbp_1 _11473_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net73),
    .D(_00879_),
    .Q_N(_00120_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[3] ));
 sg13g2_dfrbp_1 _11474_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net69),
    .D(_00880_),
    .Q_N(_00114_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[4] ));
 sg13g2_dfrbp_1 _11475_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net67),
    .D(_00881_),
    .Q_N(_00112_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[15] ));
 sg13g2_dfrbp_1 _11476_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net558),
    .D(_00882_),
    .Q_N(_00111_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[16] ));
 sg13g2_dfrbp_1 _11477_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net554),
    .D(_00883_),
    .Q_N(_00136_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[17] ));
 sg13g2_dfrbp_1 _11478_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net119),
    .D(_00884_),
    .Q_N(_00115_),
    .Q(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_1[0] ));
 sg13g2_dfrbp_1 _11479_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net115),
    .D(_00885_),
    .Q_N(_04667_),
    .Q(\ChiselTop.wild.cpu._GEN_176[1] ));
 sg13g2_dfrbp_1 _11480_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net111),
    .D(_00886_),
    .Q_N(_00119_),
    .Q(\ChiselTop.wild.cpu._GEN_176[2] ));
 sg13g2_dfrbp_1 _11481_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net107),
    .D(_00887_),
    .Q_N(_04666_),
    .Q(\ChiselTop.wild.cpu._GEN_176[6] ));
 sg13g2_dfrbp_1 _11482_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net103),
    .D(_00888_),
    .Q_N(_00134_),
    .Q(\ChiselTop.wild.cpu._GEN_176[10] ));
 sg13g2_dfrbp_1 _11483_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net99),
    .D(_00889_),
    .Q_N(_00110_),
    .Q(\ChiselTop.wild.cpu._GEN_176[20] ));
 sg13g2_dfrbp_1 _11484_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net95),
    .D(_00890_),
    .Q_N(_04665_),
    .Q(\ChiselTop.wild.cpu._pcNext_T_1[0] ));
 sg13g2_dfrbp_1 _11485_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net87),
    .D(_00891_),
    .Q_N(_04664_),
    .Q(\ChiselTop.wild.cpu._pcNext_T_1[1] ));
 sg13g2_dfrbp_1 _11486_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net91),
    .D(net862),
    .Q_N(_00000_),
    .Q(\ChiselTop.ledReg ));
 sg13g2_tiehi _10726__20 (.L_HI(net20));
 sg13g2_tiehi _10725__21 (.L_HI(net21));
 sg13g2_tiehi _10724__22 (.L_HI(net22));
 sg13g2_tiehi _10723__23 (.L_HI(net23));
 sg13g2_tiehi _10722__24 (.L_HI(net24));
 sg13g2_tiehi _10721__25 (.L_HI(net25));
 sg13g2_tiehi _10720__26 (.L_HI(net26));
 sg13g2_tiehi _10719__27 (.L_HI(net27));
 sg13g2_tiehi _10718__28 (.L_HI(net28));
 sg13g2_tiehi _10717__29 (.L_HI(net29));
 sg13g2_tiehi _10716__30 (.L_HI(net30));
 sg13g2_tiehi _10715__31 (.L_HI(net31));
 sg13g2_tiehi _10714__32 (.L_HI(net32));
 sg13g2_tiehi _10713__33 (.L_HI(net33));
 sg13g2_tiehi _10712__34 (.L_HI(net34));
 sg13g2_tiehi _10711__35 (.L_HI(net35));
 sg13g2_tiehi _10710__36 (.L_HI(net36));
 sg13g2_tiehi _10709__37 (.L_HI(net37));
 sg13g2_tiehi _10708__38 (.L_HI(net38));
 sg13g2_tiehi _10707__39 (.L_HI(net39));
 sg13g2_tiehi _10706__40 (.L_HI(net40));
 sg13g2_tiehi _10705__41 (.L_HI(net41));
 sg13g2_tiehi _10704__42 (.L_HI(net42));
 sg13g2_tiehi _10703__43 (.L_HI(net43));
 sg13g2_tiehi _10702__44 (.L_HI(net44));
 sg13g2_tiehi _10701__45 (.L_HI(net45));
 sg13g2_tiehi _10700__46 (.L_HI(net46));
 sg13g2_tiehi _10699__47 (.L_HI(net47));
 sg13g2_tiehi _10698__48 (.L_HI(net48));
 sg13g2_tiehi _10697__49 (.L_HI(net49));
 sg13g2_tiehi _10696__50 (.L_HI(net50));
 sg13g2_tiehi _10695__51 (.L_HI(net51));
 sg13g2_tiehi _10694__52 (.L_HI(net52));
 sg13g2_tiehi _10693__53 (.L_HI(net53));
 sg13g2_tiehi _10692__54 (.L_HI(net54));
 sg13g2_tiehi _10691__55 (.L_HI(net55));
 sg13g2_tiehi _10690__56 (.L_HI(net56));
 sg13g2_tiehi _10689__57 (.L_HI(net57));
 sg13g2_tiehi _10688__58 (.L_HI(net58));
 sg13g2_tiehi _10687__59 (.L_HI(net59));
 sg13g2_tiehi _10686__60 (.L_HI(net60));
 sg13g2_tiehi _10685__61 (.L_HI(net61));
 sg13g2_tiehi _10684__62 (.L_HI(net62));
 sg13g2_tiehi _10683__63 (.L_HI(net63));
 sg13g2_tiehi _10682__64 (.L_HI(net64));
 sg13g2_tiehi _10681__65 (.L_HI(net65));
 sg13g2_tiehi _11458__66 (.L_HI(net66));
 sg13g2_tiehi _11475__67 (.L_HI(net67));
 sg13g2_tiehi _11457__68 (.L_HI(net68));
 sg13g2_tiehi _11474__69 (.L_HI(net69));
 sg13g2_tiehi _10680__70 (.L_HI(net70));
 sg13g2_tiehi _10728__71 (.L_HI(net71));
 sg13g2_tiehi _11456__72 (.L_HI(net72));
 sg13g2_tiehi _11473__73 (.L_HI(net73));
 sg13g2_tiehi _11455__74 (.L_HI(net74));
 sg13g2_tiehi _11472__75 (.L_HI(net75));
 sg13g2_tiehi _11454__76 (.L_HI(net76));
 sg13g2_tiehi _11471__77 (.L_HI(net77));
 sg13g2_tiehi _11453__78 (.L_HI(net78));
 sg13g2_tiehi _11470__79 (.L_HI(net79));
 sg13g2_tiehi _11452__80 (.L_HI(net80));
 sg13g2_tiehi _11446__81 (.L_HI(net81));
 sg13g2_tiehi _11451__82 (.L_HI(net82));
 sg13g2_tiehi _11469__83 (.L_HI(net83));
 sg13g2_tiehi _11450__84 (.L_HI(net84));
 sg13g2_tiehi _11449__85 (.L_HI(net85));
 sg13g2_tiehi _11448__86 (.L_HI(net86));
 sg13g2_tiehi _11485__87 (.L_HI(net87));
 sg13g2_tiehi _11447__88 (.L_HI(net88));
 sg13g2_tiehi _11468__89 (.L_HI(net89));
 sg13g2_tiehi _11445__90 (.L_HI(net90));
 sg13g2_tiehi _11486__91 (.L_HI(net91));
 sg13g2_tiehi _11444__92 (.L_HI(net92));
 sg13g2_tiehi _11467__93 (.L_HI(net93));
 sg13g2_tiehi _11443__94 (.L_HI(net94));
 sg13g2_tiehi _11484__95 (.L_HI(net95));
 sg13g2_tiehi _11442__96 (.L_HI(net96));
 sg13g2_tiehi _11466__97 (.L_HI(net97));
 sg13g2_tiehi _11441__98 (.L_HI(net98));
 sg13g2_tiehi _11483__99 (.L_HI(net99));
 sg13g2_tiehi _11440__100 (.L_HI(net100));
 sg13g2_tiehi _11465__101 (.L_HI(net101));
 sg13g2_tiehi _11439__102 (.L_HI(net102));
 sg13g2_tiehi _11482__103 (.L_HI(net103));
 sg13g2_tiehi _11438__104 (.L_HI(net104));
 sg13g2_tiehi _11464__105 (.L_HI(net105));
 sg13g2_tiehi _11437__106 (.L_HI(net106));
 sg13g2_tiehi _11481__107 (.L_HI(net107));
 sg13g2_tiehi _11436__108 (.L_HI(net108));
 sg13g2_tiehi _11463__109 (.L_HI(net109));
 sg13g2_tiehi _11435__110 (.L_HI(net110));
 sg13g2_tiehi _11480__111 (.L_HI(net111));
 sg13g2_tiehi _11434__112 (.L_HI(net112));
 sg13g2_tiehi _11462__113 (.L_HI(net113));
 sg13g2_tiehi _11433__114 (.L_HI(net114));
 sg13g2_tiehi _11479__115 (.L_HI(net115));
 sg13g2_tiehi _11432__116 (.L_HI(net116));
 sg13g2_tiehi _11461__117 (.L_HI(net117));
 sg13g2_tiehi _11431__118 (.L_HI(net118));
 sg13g2_tiehi _11478__119 (.L_HI(net119));
 sg13g2_tiehi _11430__120 (.L_HI(net120));
 sg13g2_tiehi _11429__121 (.L_HI(net121));
 sg13g2_tiehi _11428__122 (.L_HI(net122));
 sg13g2_tiehi _11427__123 (.L_HI(net123));
 sg13g2_tiehi _11426__124 (.L_HI(net124));
 sg13g2_tiehi _11425__125 (.L_HI(net125));
 sg13g2_tiehi _11424__126 (.L_HI(net126));
 sg13g2_tiehi _11423__127 (.L_HI(net127));
 sg13g2_tiehi _11422__128 (.L_HI(net128));
 sg13g2_tiehi _11421__129 (.L_HI(net129));
 sg13g2_tiehi _11420__130 (.L_HI(net130));
 sg13g2_tiehi _11419__131 (.L_HI(net131));
 sg13g2_tiehi _11418__132 (.L_HI(net132));
 sg13g2_tiehi _11417__133 (.L_HI(net133));
 sg13g2_tiehi _11416__134 (.L_HI(net134));
 sg13g2_tiehi _11415__135 (.L_HI(net135));
 sg13g2_tiehi _11414__136 (.L_HI(net136));
 sg13g2_tiehi _11413__137 (.L_HI(net137));
 sg13g2_tiehi _11412__138 (.L_HI(net138));
 sg13g2_tiehi _11411__139 (.L_HI(net139));
 sg13g2_tiehi _11410__140 (.L_HI(net140));
 sg13g2_tiehi _11409__141 (.L_HI(net141));
 sg13g2_tiehi _11408__142 (.L_HI(net142));
 sg13g2_tiehi _11407__143 (.L_HI(net143));
 sg13g2_tiehi _11406__144 (.L_HI(net144));
 sg13g2_tiehi _11405__145 (.L_HI(net145));
 sg13g2_tiehi _11404__146 (.L_HI(net146));
 sg13g2_tiehi _11403__147 (.L_HI(net147));
 sg13g2_tiehi _11402__148 (.L_HI(net148));
 sg13g2_tiehi _11401__149 (.L_HI(net149));
 sg13g2_tiehi _11400__150 (.L_HI(net150));
 sg13g2_tiehi _11399__151 (.L_HI(net151));
 sg13g2_tiehi _11398__152 (.L_HI(net152));
 sg13g2_tiehi _11397__153 (.L_HI(net153));
 sg13g2_tiehi _11396__154 (.L_HI(net154));
 sg13g2_tiehi _11395__155 (.L_HI(net155));
 sg13g2_tiehi _11394__156 (.L_HI(net156));
 sg13g2_tiehi _11393__157 (.L_HI(net157));
 sg13g2_tiehi _11392__158 (.L_HI(net158));
 sg13g2_tiehi _11391__159 (.L_HI(net159));
 sg13g2_tiehi _11390__160 (.L_HI(net160));
 sg13g2_tiehi _11389__161 (.L_HI(net161));
 sg13g2_tiehi _11388__162 (.L_HI(net162));
 sg13g2_tiehi _11387__163 (.L_HI(net163));
 sg13g2_tiehi _11386__164 (.L_HI(net164));
 sg13g2_tiehi _11385__165 (.L_HI(net165));
 sg13g2_tiehi _11384__166 (.L_HI(net166));
 sg13g2_tiehi _11383__167 (.L_HI(net167));
 sg13g2_tiehi _11382__168 (.L_HI(net168));
 sg13g2_tiehi _11381__169 (.L_HI(net169));
 sg13g2_tiehi _11380__170 (.L_HI(net170));
 sg13g2_tiehi _11379__171 (.L_HI(net171));
 sg13g2_tiehi _11378__172 (.L_HI(net172));
 sg13g2_tiehi _11377__173 (.L_HI(net173));
 sg13g2_tiehi _11376__174 (.L_HI(net174));
 sg13g2_tiehi _11375__175 (.L_HI(net175));
 sg13g2_tiehi _11374__176 (.L_HI(net176));
 sg13g2_tiehi _11373__177 (.L_HI(net177));
 sg13g2_tiehi _11372__178 (.L_HI(net178));
 sg13g2_tiehi _11371__179 (.L_HI(net179));
 sg13g2_tiehi _11370__180 (.L_HI(net180));
 sg13g2_tiehi _11369__181 (.L_HI(net181));
 sg13g2_tiehi _11368__182 (.L_HI(net182));
 sg13g2_tiehi _11367__183 (.L_HI(net183));
 sg13g2_tiehi _11366__184 (.L_HI(net184));
 sg13g2_tiehi _11365__185 (.L_HI(net185));
 sg13g2_tiehi _11364__186 (.L_HI(net186));
 sg13g2_tiehi _11363__187 (.L_HI(net187));
 sg13g2_tiehi _11362__188 (.L_HI(net188));
 sg13g2_tiehi _11361__189 (.L_HI(net189));
 sg13g2_tiehi _11360__190 (.L_HI(net190));
 sg13g2_tiehi _11359__191 (.L_HI(net191));
 sg13g2_tiehi _11358__192 (.L_HI(net192));
 sg13g2_tiehi _11357__193 (.L_HI(net193));
 sg13g2_tiehi _11356__194 (.L_HI(net194));
 sg13g2_tiehi _11355__195 (.L_HI(net195));
 sg13g2_tiehi _11354__196 (.L_HI(net196));
 sg13g2_tiehi _11353__197 (.L_HI(net197));
 sg13g2_tiehi _11352__198 (.L_HI(net198));
 sg13g2_tiehi _11351__199 (.L_HI(net199));
 sg13g2_tiehi _11350__200 (.L_HI(net200));
 sg13g2_tiehi _11349__201 (.L_HI(net201));
 sg13g2_tiehi _11348__202 (.L_HI(net202));
 sg13g2_tiehi _11347__203 (.L_HI(net203));
 sg13g2_tiehi _11346__204 (.L_HI(net204));
 sg13g2_tiehi _11345__205 (.L_HI(net205));
 sg13g2_tiehi _11344__206 (.L_HI(net206));
 sg13g2_tiehi _11343__207 (.L_HI(net207));
 sg13g2_tiehi _11342__208 (.L_HI(net208));
 sg13g2_tiehi _11341__209 (.L_HI(net209));
 sg13g2_tiehi _11340__210 (.L_HI(net210));
 sg13g2_tiehi _11339__211 (.L_HI(net211));
 sg13g2_tiehi _11338__212 (.L_HI(net212));
 sg13g2_tiehi _11337__213 (.L_HI(net213));
 sg13g2_tiehi _11336__214 (.L_HI(net214));
 sg13g2_tiehi _11335__215 (.L_HI(net215));
 sg13g2_tiehi _11334__216 (.L_HI(net216));
 sg13g2_tiehi _11333__217 (.L_HI(net217));
 sg13g2_tiehi _11332__218 (.L_HI(net218));
 sg13g2_tiehi _11331__219 (.L_HI(net219));
 sg13g2_tiehi _11330__220 (.L_HI(net220));
 sg13g2_tiehi _11329__221 (.L_HI(net221));
 sg13g2_tiehi _11328__222 (.L_HI(net222));
 sg13g2_tiehi _11327__223 (.L_HI(net223));
 sg13g2_tiehi _11326__224 (.L_HI(net224));
 sg13g2_tiehi _11325__225 (.L_HI(net225));
 sg13g2_tiehi _11324__226 (.L_HI(net226));
 sg13g2_tiehi _11323__227 (.L_HI(net227));
 sg13g2_tiehi _11322__228 (.L_HI(net228));
 sg13g2_tiehi _11321__229 (.L_HI(net229));
 sg13g2_tiehi _11320__230 (.L_HI(net230));
 sg13g2_tiehi _11319__231 (.L_HI(net231));
 sg13g2_tiehi _11318__232 (.L_HI(net232));
 sg13g2_tiehi _11317__233 (.L_HI(net233));
 sg13g2_tiehi _11316__234 (.L_HI(net234));
 sg13g2_tiehi _11315__235 (.L_HI(net235));
 sg13g2_tiehi _11314__236 (.L_HI(net236));
 sg13g2_tiehi _11313__237 (.L_HI(net237));
 sg13g2_tiehi _11312__238 (.L_HI(net238));
 sg13g2_tiehi _11311__239 (.L_HI(net239));
 sg13g2_tiehi _11310__240 (.L_HI(net240));
 sg13g2_tiehi _11309__241 (.L_HI(net241));
 sg13g2_tiehi _11308__242 (.L_HI(net242));
 sg13g2_tiehi _11307__243 (.L_HI(net243));
 sg13g2_tiehi _11306__244 (.L_HI(net244));
 sg13g2_tiehi _11305__245 (.L_HI(net245));
 sg13g2_tiehi _11304__246 (.L_HI(net246));
 sg13g2_tiehi _11303__247 (.L_HI(net247));
 sg13g2_tiehi _11302__248 (.L_HI(net248));
 sg13g2_tiehi _11301__249 (.L_HI(net249));
 sg13g2_tiehi _11300__250 (.L_HI(net250));
 sg13g2_tiehi _11299__251 (.L_HI(net251));
 sg13g2_tiehi _11298__252 (.L_HI(net252));
 sg13g2_tiehi _11297__253 (.L_HI(net253));
 sg13g2_tiehi _11296__254 (.L_HI(net254));
 sg13g2_tiehi _11295__255 (.L_HI(net255));
 sg13g2_tiehi _11294__256 (.L_HI(net256));
 sg13g2_tiehi _11293__257 (.L_HI(net257));
 sg13g2_tiehi _11292__258 (.L_HI(net258));
 sg13g2_tiehi _11291__259 (.L_HI(net259));
 sg13g2_tiehi _11290__260 (.L_HI(net260));
 sg13g2_tiehi _11289__261 (.L_HI(net261));
 sg13g2_tiehi _11288__262 (.L_HI(net262));
 sg13g2_tiehi _11287__263 (.L_HI(net263));
 sg13g2_tiehi _11286__264 (.L_HI(net264));
 sg13g2_tiehi _11285__265 (.L_HI(net265));
 sg13g2_tiehi _11284__266 (.L_HI(net266));
 sg13g2_tiehi _11283__267 (.L_HI(net267));
 sg13g2_tiehi _11282__268 (.L_HI(net268));
 sg13g2_tiehi _11281__269 (.L_HI(net269));
 sg13g2_tiehi _11280__270 (.L_HI(net270));
 sg13g2_tiehi _11279__271 (.L_HI(net271));
 sg13g2_tiehi _11278__272 (.L_HI(net272));
 sg13g2_tiehi _11277__273 (.L_HI(net273));
 sg13g2_tiehi _11276__274 (.L_HI(net274));
 sg13g2_tiehi _11275__275 (.L_HI(net275));
 sg13g2_tiehi _11274__276 (.L_HI(net276));
 sg13g2_tiehi _11273__277 (.L_HI(net277));
 sg13g2_tiehi _11272__278 (.L_HI(net278));
 sg13g2_tiehi _11271__279 (.L_HI(net279));
 sg13g2_tiehi _11270__280 (.L_HI(net280));
 sg13g2_tiehi _11269__281 (.L_HI(net281));
 sg13g2_tiehi _11268__282 (.L_HI(net282));
 sg13g2_tiehi _11267__283 (.L_HI(net283));
 sg13g2_tiehi _11266__284 (.L_HI(net284));
 sg13g2_tiehi _11265__285 (.L_HI(net285));
 sg13g2_tiehi _11264__286 (.L_HI(net286));
 sg13g2_tiehi _11263__287 (.L_HI(net287));
 sg13g2_tiehi _11262__288 (.L_HI(net288));
 sg13g2_tiehi _11261__289 (.L_HI(net289));
 sg13g2_tiehi _11257__290 (.L_HI(net290));
 sg13g2_tiehi _11256__291 (.L_HI(net291));
 sg13g2_tiehi _11255__292 (.L_HI(net292));
 sg13g2_tiehi _11254__293 (.L_HI(net293));
 sg13g2_tiehi _11253__294 (.L_HI(net294));
 sg13g2_tiehi _11252__295 (.L_HI(net295));
 sg13g2_tiehi _11251__296 (.L_HI(net296));
 sg13g2_tiehi _11250__297 (.L_HI(net297));
 sg13g2_tiehi _11249__298 (.L_HI(net298));
 sg13g2_tiehi _11248__299 (.L_HI(net299));
 sg13g2_tiehi _11247__300 (.L_HI(net300));
 sg13g2_tiehi _11246__301 (.L_HI(net301));
 sg13g2_tiehi _11245__302 (.L_HI(net302));
 sg13g2_tiehi _11244__303 (.L_HI(net303));
 sg13g2_tiehi _11243__304 (.L_HI(net304));
 sg13g2_tiehi _11242__305 (.L_HI(net305));
 sg13g2_tiehi _11241__306 (.L_HI(net306));
 sg13g2_tiehi _11240__307 (.L_HI(net307));
 sg13g2_tiehi _11239__308 (.L_HI(net308));
 sg13g2_tiehi _11238__309 (.L_HI(net309));
 sg13g2_tiehi _11237__310 (.L_HI(net310));
 sg13g2_tiehi _11236__311 (.L_HI(net311));
 sg13g2_tiehi _11235__312 (.L_HI(net312));
 sg13g2_tiehi _11234__313 (.L_HI(net313));
 sg13g2_tiehi _11233__314 (.L_HI(net314));
 sg13g2_tiehi _11232__315 (.L_HI(net315));
 sg13g2_tiehi _11231__316 (.L_HI(net316));
 sg13g2_tiehi _11230__317 (.L_HI(net317));
 sg13g2_tiehi _11229__318 (.L_HI(net318));
 sg13g2_tiehi _11228__319 (.L_HI(net319));
 sg13g2_tiehi _11227__320 (.L_HI(net320));
 sg13g2_tiehi _11226__321 (.L_HI(net321));
 sg13g2_tiehi _11225__322 (.L_HI(net322));
 sg13g2_tiehi _11224__323 (.L_HI(net323));
 sg13g2_tiehi _11223__324 (.L_HI(net324));
 sg13g2_tiehi _11222__325 (.L_HI(net325));
 sg13g2_tiehi _11221__326 (.L_HI(net326));
 sg13g2_tiehi _11220__327 (.L_HI(net327));
 sg13g2_tiehi _11219__328 (.L_HI(net328));
 sg13g2_tiehi _11218__329 (.L_HI(net329));
 sg13g2_tiehi _11217__330 (.L_HI(net330));
 sg13g2_tiehi _11216__331 (.L_HI(net331));
 sg13g2_tiehi _11215__332 (.L_HI(net332));
 sg13g2_tiehi _11214__333 (.L_HI(net333));
 sg13g2_tiehi _11213__334 (.L_HI(net334));
 sg13g2_tiehi _11212__335 (.L_HI(net335));
 sg13g2_tiehi _11211__336 (.L_HI(net336));
 sg13g2_tiehi _11210__337 (.L_HI(net337));
 sg13g2_tiehi _11209__338 (.L_HI(net338));
 sg13g2_tiehi _11208__339 (.L_HI(net339));
 sg13g2_tiehi _11207__340 (.L_HI(net340));
 sg13g2_tiehi _11206__341 (.L_HI(net341));
 sg13g2_tiehi _11205__342 (.L_HI(net342));
 sg13g2_tiehi _11204__343 (.L_HI(net343));
 sg13g2_tiehi _11203__344 (.L_HI(net344));
 sg13g2_tiehi _11202__345 (.L_HI(net345));
 sg13g2_tiehi _11201__346 (.L_HI(net346));
 sg13g2_tiehi _11200__347 (.L_HI(net347));
 sg13g2_tiehi _11199__348 (.L_HI(net348));
 sg13g2_tiehi _11198__349 (.L_HI(net349));
 sg13g2_tiehi _11197__350 (.L_HI(net350));
 sg13g2_tiehi _11196__351 (.L_HI(net351));
 sg13g2_tiehi _11195__352 (.L_HI(net352));
 sg13g2_tiehi _11194__353 (.L_HI(net353));
 sg13g2_tiehi _11193__354 (.L_HI(net354));
 sg13g2_tiehi _11192__355 (.L_HI(net355));
 sg13g2_tiehi _11191__356 (.L_HI(net356));
 sg13g2_tiehi _11190__357 (.L_HI(net357));
 sg13g2_tiehi _11189__358 (.L_HI(net358));
 sg13g2_tiehi _11188__359 (.L_HI(net359));
 sg13g2_tiehi _11187__360 (.L_HI(net360));
 sg13g2_tiehi _11186__361 (.L_HI(net361));
 sg13g2_tiehi _11185__362 (.L_HI(net362));
 sg13g2_tiehi _11184__363 (.L_HI(net363));
 sg13g2_tiehi _11183__364 (.L_HI(net364));
 sg13g2_tiehi _11182__365 (.L_HI(net365));
 sg13g2_tiehi _11181__366 (.L_HI(net366));
 sg13g2_tiehi _11180__367 (.L_HI(net367));
 sg13g2_tiehi _11179__368 (.L_HI(net368));
 sg13g2_tiehi _11178__369 (.L_HI(net369));
 sg13g2_tiehi _11177__370 (.L_HI(net370));
 sg13g2_tiehi _11176__371 (.L_HI(net371));
 sg13g2_tiehi _11175__372 (.L_HI(net372));
 sg13g2_tiehi _11174__373 (.L_HI(net373));
 sg13g2_tiehi _11173__374 (.L_HI(net374));
 sg13g2_tiehi _11172__375 (.L_HI(net375));
 sg13g2_tiehi _11171__376 (.L_HI(net376));
 sg13g2_tiehi _11170__377 (.L_HI(net377));
 sg13g2_tiehi _11169__378 (.L_HI(net378));
 sg13g2_tiehi _11168__379 (.L_HI(net379));
 sg13g2_tiehi _11167__380 (.L_HI(net380));
 sg13g2_tiehi _11166__381 (.L_HI(net381));
 sg13g2_tiehi _11165__382 (.L_HI(net382));
 sg13g2_tiehi _11164__383 (.L_HI(net383));
 sg13g2_tiehi _11163__384 (.L_HI(net384));
 sg13g2_tiehi _11162__385 (.L_HI(net385));
 sg13g2_tiehi _11161__386 (.L_HI(net386));
 sg13g2_tiehi _11160__387 (.L_HI(net387));
 sg13g2_tiehi _11159__388 (.L_HI(net388));
 sg13g2_tiehi _11158__389 (.L_HI(net389));
 sg13g2_tiehi _11157__390 (.L_HI(net390));
 sg13g2_tiehi _11156__391 (.L_HI(net391));
 sg13g2_tiehi _11155__392 (.L_HI(net392));
 sg13g2_tiehi _11154__393 (.L_HI(net393));
 sg13g2_tiehi _11153__394 (.L_HI(net394));
 sg13g2_tiehi _11152__395 (.L_HI(net395));
 sg13g2_tiehi _11151__396 (.L_HI(net396));
 sg13g2_tiehi _11150__397 (.L_HI(net397));
 sg13g2_tiehi _11149__398 (.L_HI(net398));
 sg13g2_tiehi _11148__399 (.L_HI(net399));
 sg13g2_tiehi _11147__400 (.L_HI(net400));
 sg13g2_tiehi _11146__401 (.L_HI(net401));
 sg13g2_tiehi _11145__402 (.L_HI(net402));
 sg13g2_tiehi _11144__403 (.L_HI(net403));
 sg13g2_tiehi _11143__404 (.L_HI(net404));
 sg13g2_tiehi _11142__405 (.L_HI(net405));
 sg13g2_tiehi _11141__406 (.L_HI(net406));
 sg13g2_tiehi _11140__407 (.L_HI(net407));
 sg13g2_tiehi _11139__408 (.L_HI(net408));
 sg13g2_tiehi _11138__409 (.L_HI(net409));
 sg13g2_tiehi _11137__410 (.L_HI(net410));
 sg13g2_tiehi _11136__411 (.L_HI(net411));
 sg13g2_tiehi _11135__412 (.L_HI(net412));
 sg13g2_tiehi _11134__413 (.L_HI(net413));
 sg13g2_tiehi _11133__414 (.L_HI(net414));
 sg13g2_tiehi _11132__415 (.L_HI(net415));
 sg13g2_tiehi _11131__416 (.L_HI(net416));
 sg13g2_tiehi _11130__417 (.L_HI(net417));
 sg13g2_tiehi _11129__418 (.L_HI(net418));
 sg13g2_tiehi _11128__419 (.L_HI(net419));
 sg13g2_tiehi _11127__420 (.L_HI(net420));
 sg13g2_tiehi _11126__421 (.L_HI(net421));
 sg13g2_tiehi _11125__422 (.L_HI(net422));
 sg13g2_tiehi _11124__423 (.L_HI(net423));
 sg13g2_tiehi _11123__424 (.L_HI(net424));
 sg13g2_tiehi _11122__425 (.L_HI(net425));
 sg13g2_tiehi _11121__426 (.L_HI(net426));
 sg13g2_tiehi _11120__427 (.L_HI(net427));
 sg13g2_tiehi _11119__428 (.L_HI(net428));
 sg13g2_tiehi _11118__429 (.L_HI(net429));
 sg13g2_tiehi _11117__430 (.L_HI(net430));
 sg13g2_tiehi _11116__431 (.L_HI(net431));
 sg13g2_tiehi _11115__432 (.L_HI(net432));
 sg13g2_tiehi _10729__433 (.L_HI(net433));
 sg13g2_tiehi _10995__434 (.L_HI(net434));
 sg13g2_tiehi _10996__435 (.L_HI(net435));
 sg13g2_tiehi _10997__436 (.L_HI(net436));
 sg13g2_tiehi _10998__437 (.L_HI(net437));
 sg13g2_tiehi _10999__438 (.L_HI(net438));
 sg13g2_tiehi _11000__439 (.L_HI(net439));
 sg13g2_tiehi _11001__440 (.L_HI(net440));
 sg13g2_tiehi _11002__441 (.L_HI(net441));
 sg13g2_tiehi _11003__442 (.L_HI(net442));
 sg13g2_tiehi _11004__443 (.L_HI(net443));
 sg13g2_tiehi _11005__444 (.L_HI(net444));
 sg13g2_tiehi _11006__445 (.L_HI(net445));
 sg13g2_tiehi _11007__446 (.L_HI(net446));
 sg13g2_tiehi _11008__447 (.L_HI(net447));
 sg13g2_tiehi _11009__448 (.L_HI(net448));
 sg13g2_tiehi _11010__449 (.L_HI(net449));
 sg13g2_tiehi _11011__450 (.L_HI(net450));
 sg13g2_tiehi _11114__451 (.L_HI(net451));
 sg13g2_tiehi _11113__452 (.L_HI(net452));
 sg13g2_tiehi _11112__453 (.L_HI(net453));
 sg13g2_tiehi _11111__454 (.L_HI(net454));
 sg13g2_tiehi _11110__455 (.L_HI(net455));
 sg13g2_tiehi _11109__456 (.L_HI(net456));
 sg13g2_tiehi _11012__457 (.L_HI(net457));
 sg13g2_tiehi _11019__458 (.L_HI(net458));
 sg13g2_tiehi _11020__459 (.L_HI(net459));
 sg13g2_tiehi _11021__460 (.L_HI(net460));
 sg13g2_tiehi _11022__461 (.L_HI(net461));
 sg13g2_tiehi _11023__462 (.L_HI(net462));
 sg13g2_tiehi _11024__463 (.L_HI(net463));
 sg13g2_tiehi _11025__464 (.L_HI(net464));
 sg13g2_tiehi _11026__465 (.L_HI(net465));
 sg13g2_tiehi _11027__466 (.L_HI(net466));
 sg13g2_tiehi _11028__467 (.L_HI(net467));
 sg13g2_tiehi _11029__468 (.L_HI(net468));
 sg13g2_tiehi _11030__469 (.L_HI(net469));
 sg13g2_tiehi _11031__470 (.L_HI(net470));
 sg13g2_tiehi _11032__471 (.L_HI(net471));
 sg13g2_tiehi _11033__472 (.L_HI(net472));
 sg13g2_tiehi _11034__473 (.L_HI(net473));
 sg13g2_tiehi _11035__474 (.L_HI(net474));
 sg13g2_tiehi _11036__475 (.L_HI(net475));
 sg13g2_tiehi _11037__476 (.L_HI(net476));
 sg13g2_tiehi _11038__477 (.L_HI(net477));
 sg13g2_tiehi _11039__478 (.L_HI(net478));
 sg13g2_tiehi _11040__479 (.L_HI(net479));
 sg13g2_tiehi _11041__480 (.L_HI(net480));
 sg13g2_tiehi _11042__481 (.L_HI(net481));
 sg13g2_tiehi _11043__482 (.L_HI(net482));
 sg13g2_tiehi _11044__483 (.L_HI(net483));
 sg13g2_tiehi _11045__484 (.L_HI(net484));
 sg13g2_tiehi _11046__485 (.L_HI(net485));
 sg13g2_tiehi _11047__486 (.L_HI(net486));
 sg13g2_tiehi _11048__487 (.L_HI(net487));
 sg13g2_tiehi _11049__488 (.L_HI(net488));
 sg13g2_tiehi _11108__489 (.L_HI(net489));
 sg13g2_tiehi _11107__490 (.L_HI(net490));
 sg13g2_tiehi _11106__491 (.L_HI(net491));
 sg13g2_tiehi _11105__492 (.L_HI(net492));
 sg13g2_tiehi _11104__493 (.L_HI(net493));
 sg13g2_tiehi _11103__494 (.L_HI(net494));
 sg13g2_tiehi _11102__495 (.L_HI(net495));
 sg13g2_tiehi _11101__496 (.L_HI(net496));
 sg13g2_tiehi _11100__497 (.L_HI(net497));
 sg13g2_tiehi _11099__498 (.L_HI(net498));
 sg13g2_tiehi _11098__499 (.L_HI(net499));
 sg13g2_tiehi _11097__500 (.L_HI(net500));
 sg13g2_tiehi _11096__501 (.L_HI(net501));
 sg13g2_tiehi _11095__502 (.L_HI(net502));
 sg13g2_tiehi _11094__503 (.L_HI(net503));
 sg13g2_tiehi _11093__504 (.L_HI(net504));
 sg13g2_tiehi _11092__505 (.L_HI(net505));
 sg13g2_tiehi _11091__506 (.L_HI(net506));
 sg13g2_tiehi _11090__507 (.L_HI(net507));
 sg13g2_tiehi _11089__508 (.L_HI(net508));
 sg13g2_tiehi _11088__509 (.L_HI(net509));
 sg13g2_tiehi _11087__510 (.L_HI(net510));
 sg13g2_tiehi _11086__511 (.L_HI(net511));
 sg13g2_tiehi _11085__512 (.L_HI(net512));
 sg13g2_tiehi _11084__513 (.L_HI(net513));
 sg13g2_tiehi _11083__514 (.L_HI(net514));
 sg13g2_tiehi _11082__515 (.L_HI(net515));
 sg13g2_tiehi _11081__516 (.L_HI(net516));
 sg13g2_tiehi _11080__517 (.L_HI(net517));
 sg13g2_tiehi _11079__518 (.L_HI(net518));
 sg13g2_tiehi _11078__519 (.L_HI(net519));
 sg13g2_tiehi _11077__520 (.L_HI(net520));
 sg13g2_tiehi _11076__521 (.L_HI(net521));
 sg13g2_tiehi _11075__522 (.L_HI(net522));
 sg13g2_tiehi _11074__523 (.L_HI(net523));
 sg13g2_tiehi _11073__524 (.L_HI(net524));
 sg13g2_tiehi _11072__525 (.L_HI(net525));
 sg13g2_tiehi _11071__526 (.L_HI(net526));
 sg13g2_tiehi _11070__527 (.L_HI(net527));
 sg13g2_tiehi _11069__528 (.L_HI(net528));
 sg13g2_tiehi _11068__529 (.L_HI(net529));
 sg13g2_tiehi _11067__530 (.L_HI(net530));
 sg13g2_tiehi _11066__531 (.L_HI(net531));
 sg13g2_tiehi _11065__532 (.L_HI(net532));
 sg13g2_tiehi _11064__533 (.L_HI(net533));
 sg13g2_tiehi _11063__534 (.L_HI(net534));
 sg13g2_tiehi _11062__535 (.L_HI(net535));
 sg13g2_tiehi _11061__536 (.L_HI(net536));
 sg13g2_tiehi _11060__537 (.L_HI(net537));
 sg13g2_tiehi _11059__538 (.L_HI(net538));
 sg13g2_tiehi _11058__539 (.L_HI(net539));
 sg13g2_tiehi _11057__540 (.L_HI(net540));
 sg13g2_tiehi _11056__541 (.L_HI(net541));
 sg13g2_tiehi _11055__542 (.L_HI(net542));
 sg13g2_tiehi _11054__543 (.L_HI(net543));
 sg13g2_tiehi _11053__544 (.L_HI(net544));
 sg13g2_tiehi _11052__545 (.L_HI(net545));
 sg13g2_tiehi _11051__546 (.L_HI(net546));
 sg13g2_tiehi _11018__547 (.L_HI(net547));
 sg13g2_tiehi _11017__548 (.L_HI(net548));
 sg13g2_tiehi _11016__549 (.L_HI(net549));
 sg13g2_tiehi _11015__550 (.L_HI(net550));
 sg13g2_tiehi _11014__551 (.L_HI(net551));
 sg13g2_tiehi _11460__552 (.L_HI(net552));
 sg13g2_tiehi _11013__553 (.L_HI(net553));
 sg13g2_tiehi _11477__554 (.L_HI(net554));
 sg13g2_tiehi _10994__555 (.L_HI(net555));
 sg13g2_tiehi _11459__556 (.L_HI(net556));
 sg13g2_tiehi _10993__557 (.L_HI(net557));
 sg13g2_tiehi _11476__558 (.L_HI(net558));
 sg13g2_tiehi _10992__559 (.L_HI(net559));
 sg13g2_tiehi _10991__560 (.L_HI(net560));
 sg13g2_tiehi _10990__561 (.L_HI(net561));
 sg13g2_tiehi _10989__562 (.L_HI(net562));
 sg13g2_tiehi _10988__563 (.L_HI(net563));
 sg13g2_tiehi _10987__564 (.L_HI(net564));
 sg13g2_tiehi _10986__565 (.L_HI(net565));
 sg13g2_tiehi _10985__566 (.L_HI(net566));
 sg13g2_tiehi _10984__567 (.L_HI(net567));
 sg13g2_tiehi _10983__568 (.L_HI(net568));
 sg13g2_tiehi _10982__569 (.L_HI(net569));
 sg13g2_tiehi _10981__570 (.L_HI(net570));
 sg13g2_tiehi _10980__571 (.L_HI(net571));
 sg13g2_tiehi _10979__572 (.L_HI(net572));
 sg13g2_tiehi _10978__573 (.L_HI(net573));
 sg13g2_tiehi _10977__574 (.L_HI(net574));
 sg13g2_tiehi _10976__575 (.L_HI(net575));
 sg13g2_tiehi _10975__576 (.L_HI(net576));
 sg13g2_tiehi _10974__577 (.L_HI(net577));
 sg13g2_tiehi _10973__578 (.L_HI(net578));
 sg13g2_tiehi _10972__579 (.L_HI(net579));
 sg13g2_tiehi _10971__580 (.L_HI(net580));
 sg13g2_tiehi _10970__581 (.L_HI(net581));
 sg13g2_tiehi _10969__582 (.L_HI(net582));
 sg13g2_tiehi _10968__583 (.L_HI(net583));
 sg13g2_tiehi _10967__584 (.L_HI(net584));
 sg13g2_tiehi _10966__585 (.L_HI(net585));
 sg13g2_tiehi _10965__586 (.L_HI(net586));
 sg13g2_tiehi _10964__587 (.L_HI(net587));
 sg13g2_tiehi _10963__588 (.L_HI(net588));
 sg13g2_tiehi _10962__589 (.L_HI(net589));
 sg13g2_tiehi _10961__590 (.L_HI(net590));
 sg13g2_tiehi _10960__591 (.L_HI(net591));
 sg13g2_tiehi _10959__592 (.L_HI(net592));
 sg13g2_tiehi _10958__593 (.L_HI(net593));
 sg13g2_tiehi _10957__594 (.L_HI(net594));
 sg13g2_tiehi _10956__595 (.L_HI(net595));
 sg13g2_tiehi _10955__596 (.L_HI(net596));
 sg13g2_tiehi _10954__597 (.L_HI(net597));
 sg13g2_tiehi _10953__598 (.L_HI(net598));
 sg13g2_tiehi _10952__599 (.L_HI(net599));
 sg13g2_tiehi _10951__600 (.L_HI(net600));
 sg13g2_tiehi _10950__601 (.L_HI(net601));
 sg13g2_tiehi _10949__602 (.L_HI(net602));
 sg13g2_tiehi _10948__603 (.L_HI(net603));
 sg13g2_tiehi _10947__604 (.L_HI(net604));
 sg13g2_tiehi _10946__605 (.L_HI(net605));
 sg13g2_tiehi _10945__606 (.L_HI(net606));
 sg13g2_tiehi _10944__607 (.L_HI(net607));
 sg13g2_tiehi _10943__608 (.L_HI(net608));
 sg13g2_tiehi _10942__609 (.L_HI(net609));
 sg13g2_tiehi _10941__610 (.L_HI(net610));
 sg13g2_tiehi _10940__611 (.L_HI(net611));
 sg13g2_tiehi _10939__612 (.L_HI(net612));
 sg13g2_tiehi _10938__613 (.L_HI(net613));
 sg13g2_tiehi _10937__614 (.L_HI(net614));
 sg13g2_tiehi _10936__615 (.L_HI(net615));
 sg13g2_tiehi _10935__616 (.L_HI(net616));
 sg13g2_tiehi _10934__617 (.L_HI(net617));
 sg13g2_tiehi _10933__618 (.L_HI(net618));
 sg13g2_tiehi _10932__619 (.L_HI(net619));
 sg13g2_tiehi _10931__620 (.L_HI(net620));
 sg13g2_tiehi _10930__621 (.L_HI(net621));
 sg13g2_tiehi _10929__622 (.L_HI(net622));
 sg13g2_tiehi _10928__623 (.L_HI(net623));
 sg13g2_tiehi _10927__624 (.L_HI(net624));
 sg13g2_tiehi _10926__625 (.L_HI(net625));
 sg13g2_tiehi _10925__626 (.L_HI(net626));
 sg13g2_tiehi _10924__627 (.L_HI(net627));
 sg13g2_tiehi _10923__628 (.L_HI(net628));
 sg13g2_tiehi _10922__629 (.L_HI(net629));
 sg13g2_tiehi _10921__630 (.L_HI(net630));
 sg13g2_tiehi _10920__631 (.L_HI(net631));
 sg13g2_tiehi _11050__632 (.L_HI(net632));
 sg13g2_tiehi _11258__633 (.L_HI(net633));
 sg13g2_tiehi _11259__634 (.L_HI(net634));
 sg13g2_tiehi _10919__635 (.L_HI(net635));
 sg13g2_tiehi _10918__636 (.L_HI(net636));
 sg13g2_tiehi _10917__637 (.L_HI(net637));
 sg13g2_tiehi _10916__638 (.L_HI(net638));
 sg13g2_tiehi _10915__639 (.L_HI(net639));
 sg13g2_tiehi _10914__640 (.L_HI(net640));
 sg13g2_tiehi _10913__641 (.L_HI(net641));
 sg13g2_tiehi _10912__642 (.L_HI(net642));
 sg13g2_tiehi _10911__643 (.L_HI(net643));
 sg13g2_tiehi _10910__644 (.L_HI(net644));
 sg13g2_tiehi _10909__645 (.L_HI(net645));
 sg13g2_tiehi _10908__646 (.L_HI(net646));
 sg13g2_tiehi _10907__647 (.L_HI(net647));
 sg13g2_tiehi _10906__648 (.L_HI(net648));
 sg13g2_tiehi _10905__649 (.L_HI(net649));
 sg13g2_tiehi _10904__650 (.L_HI(net650));
 sg13g2_tiehi _10903__651 (.L_HI(net651));
 sg13g2_tiehi _10902__652 (.L_HI(net652));
 sg13g2_tiehi _10901__653 (.L_HI(net653));
 sg13g2_tiehi _10900__654 (.L_HI(net654));
 sg13g2_tiehi _10899__655 (.L_HI(net655));
 sg13g2_tiehi _10898__656 (.L_HI(net656));
 sg13g2_tiehi _10897__657 (.L_HI(net657));
 sg13g2_tiehi _10896__658 (.L_HI(net658));
 sg13g2_tiehi _10895__659 (.L_HI(net659));
 sg13g2_tiehi _10894__660 (.L_HI(net660));
 sg13g2_tiehi _10893__661 (.L_HI(net661));
 sg13g2_tiehi _10892__662 (.L_HI(net662));
 sg13g2_tiehi _10891__663 (.L_HI(net663));
 sg13g2_tiehi _10890__664 (.L_HI(net664));
 sg13g2_tiehi _10889__665 (.L_HI(net665));
 sg13g2_tiehi _10888__666 (.L_HI(net666));
 sg13g2_tiehi _10887__667 (.L_HI(net667));
 sg13g2_tiehi _10886__668 (.L_HI(net668));
 sg13g2_tiehi _10885__669 (.L_HI(net669));
 sg13g2_tiehi _10884__670 (.L_HI(net670));
 sg13g2_tiehi _10883__671 (.L_HI(net671));
 sg13g2_tiehi _10882__672 (.L_HI(net672));
 sg13g2_tiehi _10881__673 (.L_HI(net673));
 sg13g2_tiehi _10880__674 (.L_HI(net674));
 sg13g2_tiehi _10879__675 (.L_HI(net675));
 sg13g2_tiehi _10878__676 (.L_HI(net676));
 sg13g2_tiehi _10877__677 (.L_HI(net677));
 sg13g2_tiehi _10876__678 (.L_HI(net678));
 sg13g2_tiehi _10875__679 (.L_HI(net679));
 sg13g2_tiehi _10874__680 (.L_HI(net680));
 sg13g2_tiehi _10873__681 (.L_HI(net681));
 sg13g2_tiehi _10872__682 (.L_HI(net682));
 sg13g2_tiehi _10871__683 (.L_HI(net683));
 sg13g2_tiehi _10870__684 (.L_HI(net684));
 sg13g2_tiehi _10869__685 (.L_HI(net685));
 sg13g2_tiehi _10868__686 (.L_HI(net686));
 sg13g2_tiehi _10867__687 (.L_HI(net687));
 sg13g2_tiehi _10866__688 (.L_HI(net688));
 sg13g2_tiehi _10865__689 (.L_HI(net689));
 sg13g2_tiehi _10864__690 (.L_HI(net690));
 sg13g2_tiehi _10863__691 (.L_HI(net691));
 sg13g2_tiehi _10862__692 (.L_HI(net692));
 sg13g2_tiehi _10861__693 (.L_HI(net693));
 sg13g2_tiehi _10860__694 (.L_HI(net694));
 sg13g2_tiehi _10859__695 (.L_HI(net695));
 sg13g2_tiehi _10858__696 (.L_HI(net696));
 sg13g2_tiehi _10857__697 (.L_HI(net697));
 sg13g2_tiehi _10856__698 (.L_HI(net698));
 sg13g2_tiehi _10855__699 (.L_HI(net699));
 sg13g2_tiehi _10854__700 (.L_HI(net700));
 sg13g2_tiehi _10853__701 (.L_HI(net701));
 sg13g2_tiehi _10852__702 (.L_HI(net702));
 sg13g2_tiehi _10851__703 (.L_HI(net703));
 sg13g2_tiehi _10850__704 (.L_HI(net704));
 sg13g2_tiehi _10849__705 (.L_HI(net705));
 sg13g2_tiehi _10848__706 (.L_HI(net706));
 sg13g2_tiehi _10847__707 (.L_HI(net707));
 sg13g2_tiehi _10846__708 (.L_HI(net708));
 sg13g2_tiehi _10845__709 (.L_HI(net709));
 sg13g2_tiehi _10844__710 (.L_HI(net710));
 sg13g2_tiehi _10843__711 (.L_HI(net711));
 sg13g2_tiehi _10842__712 (.L_HI(net712));
 sg13g2_tiehi _10841__713 (.L_HI(net713));
 sg13g2_tiehi _10840__714 (.L_HI(net714));
 sg13g2_tiehi _10839__715 (.L_HI(net715));
 sg13g2_tiehi _10838__716 (.L_HI(net716));
 sg13g2_tiehi _10837__717 (.L_HI(net717));
 sg13g2_tiehi _10836__718 (.L_HI(net718));
 sg13g2_tiehi _10835__719 (.L_HI(net719));
 sg13g2_tiehi _10834__720 (.L_HI(net720));
 sg13g2_tiehi _10833__721 (.L_HI(net721));
 sg13g2_tiehi _10832__722 (.L_HI(net722));
 sg13g2_tiehi _10831__723 (.L_HI(net723));
 sg13g2_tiehi _10830__724 (.L_HI(net724));
 sg13g2_tiehi _10829__725 (.L_HI(net725));
 sg13g2_tiehi _10828__726 (.L_HI(net726));
 sg13g2_tiehi _10827__727 (.L_HI(net727));
 sg13g2_tiehi _10826__728 (.L_HI(net728));
 sg13g2_tiehi _10825__729 (.L_HI(net729));
 sg13g2_tiehi _10824__730 (.L_HI(net730));
 sg13g2_tiehi _10823__731 (.L_HI(net731));
 sg13g2_tiehi _10822__732 (.L_HI(net732));
 sg13g2_tiehi _10821__733 (.L_HI(net733));
 sg13g2_tiehi _10820__734 (.L_HI(net734));
 sg13g2_tiehi _10819__735 (.L_HI(net735));
 sg13g2_tiehi _10818__736 (.L_HI(net736));
 sg13g2_tiehi _10817__737 (.L_HI(net737));
 sg13g2_tiehi _10816__738 (.L_HI(net738));
 sg13g2_tiehi _10815__739 (.L_HI(net739));
 sg13g2_tiehi _10814__740 (.L_HI(net740));
 sg13g2_tiehi _10813__741 (.L_HI(net741));
 sg13g2_tiehi _10812__742 (.L_HI(net742));
 sg13g2_tiehi _10811__743 (.L_HI(net743));
 sg13g2_tiehi _10810__744 (.L_HI(net744));
 sg13g2_tiehi _10809__745 (.L_HI(net745));
 sg13g2_tiehi _10808__746 (.L_HI(net746));
 sg13g2_tiehi _10807__747 (.L_HI(net747));
 sg13g2_tiehi _10806__748 (.L_HI(net748));
 sg13g2_tiehi _10805__749 (.L_HI(net749));
 sg13g2_tiehi _10804__750 (.L_HI(net750));
 sg13g2_tiehi _10803__751 (.L_HI(net751));
 sg13g2_tiehi _10802__752 (.L_HI(net752));
 sg13g2_tiehi _10801__753 (.L_HI(net753));
 sg13g2_tiehi _10800__754 (.L_HI(net754));
 sg13g2_tiehi _10799__755 (.L_HI(net755));
 sg13g2_tiehi _10798__756 (.L_HI(net756));
 sg13g2_tiehi _10797__757 (.L_HI(net757));
 sg13g2_tiehi _10796__758 (.L_HI(net758));
 sg13g2_tiehi _10795__759 (.L_HI(net759));
 sg13g2_tiehi _10794__760 (.L_HI(net760));
 sg13g2_tiehi _10793__761 (.L_HI(net761));
 sg13g2_tiehi _10792__762 (.L_HI(net762));
 sg13g2_tiehi _10791__763 (.L_HI(net763));
 sg13g2_tiehi _10790__764 (.L_HI(net764));
 sg13g2_tiehi _10789__765 (.L_HI(net765));
 sg13g2_tiehi _10788__766 (.L_HI(net766));
 sg13g2_tiehi _10787__767 (.L_HI(net767));
 sg13g2_tiehi _10786__768 (.L_HI(net768));
 sg13g2_tiehi _10785__769 (.L_HI(net769));
 sg13g2_tiehi _10784__770 (.L_HI(net770));
 sg13g2_tiehi _10783__771 (.L_HI(net771));
 sg13g2_tiehi _10782__772 (.L_HI(net772));
 sg13g2_tiehi _10781__773 (.L_HI(net773));
 sg13g2_tiehi _10780__774 (.L_HI(net774));
 sg13g2_tiehi _10779__775 (.L_HI(net775));
 sg13g2_tiehi _10778__776 (.L_HI(net776));
 sg13g2_tiehi _10777__777 (.L_HI(net777));
 sg13g2_tiehi _10776__778 (.L_HI(net778));
 sg13g2_tiehi _10775__779 (.L_HI(net779));
 sg13g2_tiehi _10774__780 (.L_HI(net780));
 sg13g2_tiehi _10773__781 (.L_HI(net781));
 sg13g2_tiehi _10772__782 (.L_HI(net782));
 sg13g2_tiehi _10771__783 (.L_HI(net783));
 sg13g2_tiehi _10770__784 (.L_HI(net784));
 sg13g2_tiehi _10769__785 (.L_HI(net785));
 sg13g2_tiehi _10768__786 (.L_HI(net786));
 sg13g2_tiehi _10767__787 (.L_HI(net787));
 sg13g2_tiehi _10766__788 (.L_HI(net788));
 sg13g2_tiehi _10765__789 (.L_HI(net789));
 sg13g2_tiehi _10764__790 (.L_HI(net790));
 sg13g2_tiehi _10763__791 (.L_HI(net791));
 sg13g2_tiehi _10762__792 (.L_HI(net792));
 sg13g2_tiehi _10761__793 (.L_HI(net793));
 sg13g2_tiehi _10760__794 (.L_HI(net794));
 sg13g2_tiehi _10759__795 (.L_HI(net795));
 sg13g2_tiehi _10758__796 (.L_HI(net796));
 sg13g2_tiehi _10757__797 (.L_HI(net797));
 sg13g2_tiehi _10756__798 (.L_HI(net798));
 sg13g2_tiehi _10755__799 (.L_HI(net799));
 sg13g2_tiehi _10754__800 (.L_HI(net800));
 sg13g2_tiehi _10753__801 (.L_HI(net801));
 sg13g2_tiehi _10752__802 (.L_HI(net802));
 sg13g2_tiehi _10751__803 (.L_HI(net803));
 sg13g2_tiehi _10750__804 (.L_HI(net804));
 sg13g2_tiehi _10749__805 (.L_HI(net805));
 sg13g2_tiehi _10748__806 (.L_HI(net806));
 sg13g2_tiehi _10747__807 (.L_HI(net807));
 sg13g2_tiehi _10746__808 (.L_HI(net808));
 sg13g2_tiehi _10745__809 (.L_HI(net809));
 sg13g2_tiehi _10744__810 (.L_HI(net810));
 sg13g2_tiehi _10743__811 (.L_HI(net811));
 sg13g2_tiehi _10742__812 (.L_HI(net812));
 sg13g2_tiehi _10741__813 (.L_HI(net813));
 sg13g2_tiehi _10740__814 (.L_HI(net814));
 sg13g2_tiehi _10739__815 (.L_HI(net815));
 sg13g2_tiehi _10738__816 (.L_HI(net816));
 sg13g2_tiehi _11260__817 (.L_HI(net817));
 sg13g2_tiehi _10737__818 (.L_HI(net818));
 sg13g2_tiehi _10736__819 (.L_HI(net819));
 sg13g2_tiehi _10735__820 (.L_HI(net820));
 sg13g2_tiehi _10734__821 (.L_HI(net821));
 sg13g2_tiehi _10733__822 (.L_HI(net822));
 sg13g2_tiehi _10732__823 (.L_HI(net823));
 sg13g2_tiehi _10731__824 (.L_HI(net824));
 sg13g2_tiehi _10730__825 (.L_HI(net825));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_schoeberl_wildcat_4 (.L_LO(net4));
 sg13g2_tielo tt_um_schoeberl_wildcat_5 (.L_LO(net5));
 sg13g2_tielo tt_um_schoeberl_wildcat_6 (.L_LO(net6));
 sg13g2_tielo tt_um_schoeberl_wildcat_7 (.L_LO(net7));
 sg13g2_tielo tt_um_schoeberl_wildcat_8 (.L_LO(net8));
 sg13g2_tielo tt_um_schoeberl_wildcat_9 (.L_LO(net9));
 sg13g2_tielo tt_um_schoeberl_wildcat_10 (.L_LO(net10));
 sg13g2_tielo tt_um_schoeberl_wildcat_11 (.L_LO(net11));
 sg13g2_tielo tt_um_schoeberl_wildcat_12 (.L_LO(net12));
 sg13g2_tielo tt_um_schoeberl_wildcat_13 (.L_LO(net13));
 sg13g2_tielo tt_um_schoeberl_wildcat_14 (.L_LO(net14));
 sg13g2_tielo tt_um_schoeberl_wildcat_15 (.L_LO(net15));
 sg13g2_tielo tt_um_schoeberl_wildcat_16 (.L_LO(net16));
 sg13g2_tielo tt_um_schoeberl_wildcat_17 (.L_LO(net17));
 sg13g2_tielo tt_um_schoeberl_wildcat_18 (.L_LO(net18));
 sg13g2_tiehi _10727__19 (.L_HI(net19));
 sg13g2_buf_1 _12310_ (.A(\ChiselTop.led ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout2072 (.X(net2072),
    .A(_03900_));
 sg13g2_buf_2 fanout2073 (.A(net2074),
    .X(net2073));
 sg13g2_buf_4 fanout2074 (.X(net2074),
    .A(_03416_));
 sg13g2_buf_2 fanout2075 (.A(net2076),
    .X(net2075));
 sg13g2_buf_2 fanout2076 (.A(_02803_),
    .X(net2076));
 sg13g2_buf_4 fanout2077 (.X(net2077),
    .A(net2078));
 sg13g2_buf_4 fanout2078 (.X(net2078),
    .A(_03368_));
 sg13g2_buf_2 fanout2079 (.A(net2080),
    .X(net2079));
 sg13g2_buf_4 fanout2080 (.X(net2080),
    .A(_03325_));
 sg13g2_buf_2 fanout2081 (.A(net2082),
    .X(net2081));
 sg13g2_buf_1 fanout2082 (.A(net2083),
    .X(net2082));
 sg13g2_buf_4 fanout2083 (.X(net2083),
    .A(_02950_));
 sg13g2_buf_4 fanout2084 (.X(net2084),
    .A(net2086));
 sg13g2_buf_1 fanout2085 (.A(net2086),
    .X(net2085));
 sg13g2_buf_4 fanout2086 (.X(net2086),
    .A(_02903_));
 sg13g2_buf_2 fanout2087 (.A(net2088),
    .X(net2087));
 sg13g2_buf_1 fanout2088 (.A(net2089),
    .X(net2088));
 sg13g2_buf_4 fanout2089 (.X(net2089),
    .A(_02862_));
 sg13g2_buf_2 fanout2090 (.A(net2091),
    .X(net2090));
 sg13g2_buf_2 fanout2091 (.A(net2092),
    .X(net2091));
 sg13g2_buf_4 fanout2092 (.X(net2092),
    .A(_03000_));
 sg13g2_buf_2 fanout2093 (.A(net2094),
    .X(net2093));
 sg13g2_buf_2 fanout2094 (.A(net2095),
    .X(net2094));
 sg13g2_buf_4 fanout2095 (.X(net2095),
    .A(_03073_));
 sg13g2_buf_4 fanout2096 (.X(net2096),
    .A(net2098));
 sg13g2_buf_1 fanout2097 (.A(net2098),
    .X(net2097));
 sg13g2_buf_2 fanout2098 (.A(_03039_),
    .X(net2098));
 sg13g2_buf_2 fanout2099 (.A(net2100),
    .X(net2099));
 sg13g2_buf_1 fanout2100 (.A(net2101),
    .X(net2100));
 sg13g2_buf_4 fanout2101 (.X(net2101),
    .A(_03156_));
 sg13g2_buf_4 fanout2102 (.X(net2102),
    .A(net2104));
 sg13g2_buf_2 fanout2103 (.A(net2104),
    .X(net2103));
 sg13g2_buf_4 fanout2104 (.X(net2104),
    .A(_03117_));
 sg13g2_buf_2 fanout2105 (.A(net2106),
    .X(net2105));
 sg13g2_buf_1 fanout2106 (.A(net2107),
    .X(net2106));
 sg13g2_buf_4 fanout2107 (.X(net2107),
    .A(_03271_));
 sg13g2_buf_2 fanout2108 (.A(net2109),
    .X(net2108));
 sg13g2_buf_2 fanout2109 (.A(net2110),
    .X(net2109));
 sg13g2_buf_2 fanout2110 (.A(_03235_),
    .X(net2110));
 sg13g2_buf_2 fanout2111 (.A(net2112),
    .X(net2111));
 sg13g2_buf_1 fanout2112 (.A(net2113),
    .X(net2112));
 sg13g2_buf_4 fanout2113 (.X(net2113),
    .A(_01553_));
 sg13g2_buf_2 fanout2114 (.A(net2115),
    .X(net2114));
 sg13g2_buf_1 fanout2115 (.A(net2116),
    .X(net2115));
 sg13g2_buf_4 fanout2116 (.X(net2116),
    .A(_03195_));
 sg13g2_buf_2 fanout2117 (.A(_02520_),
    .X(net2117));
 sg13g2_buf_1 fanout2118 (.A(_02520_),
    .X(net2118));
 sg13g2_buf_4 fanout2119 (.X(net2119),
    .A(net2120));
 sg13g2_buf_2 fanout2120 (.A(_02474_),
    .X(net2120));
 sg13g2_buf_4 fanout2121 (.X(net2121),
    .A(net2122));
 sg13g2_buf_2 fanout2122 (.A(_02568_),
    .X(net2122));
 sg13g2_buf_4 fanout2123 (.X(net2123),
    .A(net2124));
 sg13g2_buf_4 fanout2124 (.X(net2124),
    .A(_02421_));
 sg13g2_buf_4 fanout2125 (.X(net2125),
    .A(net2126));
 sg13g2_buf_4 fanout2126 (.X(net2126),
    .A(_02612_));
 sg13g2_buf_2 fanout2127 (.A(net2128),
    .X(net2127));
 sg13g2_buf_1 fanout2128 (.A(net2129),
    .X(net2128));
 sg13g2_buf_4 fanout2129 (.X(net2129),
    .A(_02372_));
 sg13g2_buf_2 fanout2130 (.A(net2131),
    .X(net2130));
 sg13g2_buf_4 fanout2131 (.X(net2131),
    .A(_02328_));
 sg13g2_buf_2 fanout2132 (.A(net2133),
    .X(net2132));
 sg13g2_buf_2 fanout2133 (.A(_02288_),
    .X(net2133));
 sg13g2_buf_2 fanout2134 (.A(net2135),
    .X(net2134));
 sg13g2_buf_4 fanout2135 (.X(net2135),
    .A(_02236_));
 sg13g2_buf_2 fanout2136 (.A(_02168_),
    .X(net2136));
 sg13g2_buf_1 fanout2137 (.A(_02168_),
    .X(net2137));
 sg13g2_buf_2 fanout2138 (.A(net2140),
    .X(net2138));
 sg13g2_buf_1 fanout2139 (.A(net2140),
    .X(net2139));
 sg13g2_buf_4 fanout2140 (.X(net2140),
    .A(_01927_));
 sg13g2_buf_2 fanout2141 (.A(net2142),
    .X(net2141));
 sg13g2_buf_2 fanout2142 (.A(_01789_),
    .X(net2142));
 sg13g2_buf_4 fanout2143 (.X(net2143),
    .A(_01721_));
 sg13g2_buf_2 fanout2144 (.A(_01721_),
    .X(net2144));
 sg13g2_buf_2 fanout2145 (.A(net2146),
    .X(net2145));
 sg13g2_buf_4 fanout2146 (.X(net2146),
    .A(_01651_));
 sg13g2_buf_4 fanout2147 (.X(net2147),
    .A(net2149));
 sg13g2_buf_1 fanout2148 (.A(net2149),
    .X(net2148));
 sg13g2_buf_2 fanout2149 (.A(_01984_),
    .X(net2149));
 sg13g2_buf_2 fanout2150 (.A(net2151),
    .X(net2150));
 sg13g2_buf_1 fanout2151 (.A(net2152),
    .X(net2151));
 sg13g2_buf_4 fanout2152 (.X(net2152),
    .A(_01864_));
 sg13g2_buf_2 fanout2153 (.A(net2154),
    .X(net2153));
 sg13g2_buf_2 fanout2154 (.A(_03502_),
    .X(net2154));
 sg13g2_buf_2 fanout2155 (.A(_04606_),
    .X(net2155));
 sg13g2_buf_1 fanout2156 (.A(_04606_),
    .X(net2156));
 sg13g2_buf_2 fanout2157 (.A(net2158),
    .X(net2157));
 sg13g2_buf_2 fanout2158 (.A(net2159),
    .X(net2158));
 sg13g2_buf_2 fanout2159 (.A(_04604_),
    .X(net2159));
 sg13g2_buf_2 fanout2160 (.A(net2161),
    .X(net2160));
 sg13g2_buf_1 fanout2161 (.A(net2162),
    .X(net2161));
 sg13g2_buf_2 fanout2162 (.A(net2163),
    .X(net2162));
 sg13g2_buf_2 fanout2163 (.A(net2165),
    .X(net2163));
 sg13g2_buf_2 fanout2164 (.A(net2165),
    .X(net2164));
 sg13g2_buf_2 fanout2165 (.A(_03585_),
    .X(net2165));
 sg13g2_buf_2 fanout2166 (.A(_04598_),
    .X(net2166));
 sg13g2_buf_4 fanout2167 (.X(net2167),
    .A(net2169));
 sg13g2_buf_2 fanout2168 (.A(net2169),
    .X(net2168));
 sg13g2_buf_4 fanout2169 (.X(net2169),
    .A(_00524_));
 sg13g2_buf_2 fanout2170 (.A(net2174),
    .X(net2170));
 sg13g2_buf_1 fanout2171 (.A(net2174),
    .X(net2171));
 sg13g2_buf_2 fanout2172 (.A(net2174),
    .X(net2172));
 sg13g2_buf_1 fanout2173 (.A(net2174),
    .X(net2173));
 sg13g2_buf_2 fanout2174 (.A(_01548_),
    .X(net2174));
 sg13g2_buf_2 fanout2175 (.A(net2176),
    .X(net2175));
 sg13g2_buf_4 fanout2176 (.X(net2176),
    .A(_04436_));
 sg13g2_buf_2 fanout2177 (.A(net2179),
    .X(net2177));
 sg13g2_buf_1 fanout2178 (.A(net2179),
    .X(net2178));
 sg13g2_buf_1 fanout2179 (.A(_03565_),
    .X(net2179));
 sg13g2_buf_4 fanout2180 (.X(net2180),
    .A(net2182));
 sg13g2_buf_1 fanout2181 (.A(net2182),
    .X(net2181));
 sg13g2_buf_4 fanout2182 (.X(net2182),
    .A(_03565_));
 sg13g2_buf_2 fanout2183 (.A(net2184),
    .X(net2183));
 sg13g2_buf_4 fanout2184 (.X(net2184),
    .A(_01215_));
 sg13g2_buf_2 fanout2185 (.A(net2188),
    .X(net2185));
 sg13g2_buf_2 fanout2186 (.A(net2187),
    .X(net2186));
 sg13g2_buf_1 fanout2187 (.A(net2188),
    .X(net2187));
 sg13g2_buf_2 fanout2188 (.A(_01215_),
    .X(net2188));
 sg13g2_buf_4 fanout2189 (.X(net2189),
    .A(_04437_));
 sg13g2_buf_2 fanout2190 (.A(_04437_),
    .X(net2190));
 sg13g2_buf_2 fanout2191 (.A(_01214_),
    .X(net2191));
 sg13g2_buf_2 fanout2192 (.A(_01214_),
    .X(net2192));
 sg13g2_buf_2 fanout2193 (.A(net2194),
    .X(net2193));
 sg13g2_buf_4 fanout2194 (.X(net2194),
    .A(net2202));
 sg13g2_buf_2 fanout2195 (.A(net2196),
    .X(net2195));
 sg13g2_buf_4 fanout2196 (.X(net2196),
    .A(net2202));
 sg13g2_buf_2 fanout2197 (.A(net2201),
    .X(net2197));
 sg13g2_buf_2 fanout2198 (.A(net2201),
    .X(net2198));
 sg13g2_buf_4 fanout2199 (.X(net2199),
    .A(net2200));
 sg13g2_buf_4 fanout2200 (.X(net2200),
    .A(net2201));
 sg13g2_buf_2 fanout2201 (.A(net2202),
    .X(net2201));
 sg13g2_buf_4 fanout2202 (.X(net2202),
    .A(_04403_));
 sg13g2_buf_2 fanout2203 (.A(net2204),
    .X(net2203));
 sg13g2_buf_4 fanout2204 (.X(net2204),
    .A(net2212));
 sg13g2_buf_2 fanout2205 (.A(net2206),
    .X(net2205));
 sg13g2_buf_4 fanout2206 (.X(net2206),
    .A(net2212));
 sg13g2_buf_4 fanout2207 (.X(net2207),
    .A(net2208));
 sg13g2_buf_2 fanout2208 (.A(net2212),
    .X(net2208));
 sg13g2_buf_2 fanout2209 (.A(net2212),
    .X(net2209));
 sg13g2_buf_4 fanout2210 (.X(net2210),
    .A(net2211));
 sg13g2_buf_2 fanout2211 (.A(net2212),
    .X(net2211));
 sg13g2_buf_8 fanout2212 (.A(_04371_),
    .X(net2212));
 sg13g2_buf_2 fanout2213 (.A(net2214),
    .X(net2213));
 sg13g2_buf_4 fanout2214 (.X(net2214),
    .A(net2222));
 sg13g2_buf_2 fanout2215 (.A(net2216),
    .X(net2215));
 sg13g2_buf_4 fanout2216 (.X(net2216),
    .A(net2222));
 sg13g2_buf_2 fanout2217 (.A(net2218),
    .X(net2217));
 sg13g2_buf_2 fanout2218 (.A(net2222),
    .X(net2218));
 sg13g2_buf_2 fanout2219 (.A(net2222),
    .X(net2219));
 sg13g2_buf_4 fanout2220 (.X(net2220),
    .A(net2221));
 sg13g2_buf_2 fanout2221 (.A(net2222),
    .X(net2221));
 sg13g2_buf_8 fanout2222 (.A(_04297_),
    .X(net2222));
 sg13g2_buf_2 fanout2223 (.A(net2225),
    .X(net2223));
 sg13g2_buf_1 fanout2224 (.A(net2225),
    .X(net2224));
 sg13g2_buf_4 fanout2225 (.X(net2225),
    .A(net2233));
 sg13g2_buf_2 fanout2226 (.A(net2227),
    .X(net2226));
 sg13g2_buf_4 fanout2227 (.X(net2227),
    .A(net2233));
 sg13g2_buf_1 fanout2228 (.A(net2233),
    .X(net2228));
 sg13g2_buf_4 fanout2229 (.X(net2229),
    .A(net2232));
 sg13g2_buf_2 fanout2230 (.A(net2232),
    .X(net2230));
 sg13g2_buf_4 fanout2231 (.X(net2231),
    .A(net2232));
 sg13g2_buf_2 fanout2232 (.A(net2233),
    .X(net2232));
 sg13g2_buf_2 fanout2233 (.A(_04097_),
    .X(net2233));
 sg13g2_buf_2 fanout2234 (.A(net2238),
    .X(net2234));
 sg13g2_buf_4 fanout2235 (.X(net2235),
    .A(net2238));
 sg13g2_buf_2 fanout2236 (.A(net2237),
    .X(net2236));
 sg13g2_buf_4 fanout2237 (.X(net2237),
    .A(net2238));
 sg13g2_buf_4 fanout2238 (.X(net2238),
    .A(_04065_));
 sg13g2_buf_2 fanout2239 (.A(net2243),
    .X(net2239));
 sg13g2_buf_4 fanout2240 (.X(net2240),
    .A(net2243));
 sg13g2_buf_4 fanout2241 (.X(net2241),
    .A(net2243));
 sg13g2_buf_1 fanout2242 (.A(net2243),
    .X(net2242));
 sg13g2_buf_2 fanout2243 (.A(_04065_),
    .X(net2243));
 sg13g2_buf_2 fanout2244 (.A(net2254),
    .X(net2244));
 sg13g2_buf_2 fanout2245 (.A(net2254),
    .X(net2245));
 sg13g2_buf_2 fanout2246 (.A(net2247),
    .X(net2246));
 sg13g2_buf_4 fanout2247 (.X(net2247),
    .A(net2254));
 sg13g2_buf_4 fanout2248 (.X(net2248),
    .A(net2253));
 sg13g2_buf_2 fanout2249 (.A(net2253),
    .X(net2249));
 sg13g2_buf_2 fanout2250 (.A(net2253),
    .X(net2250));
 sg13g2_buf_4 fanout2251 (.X(net2251),
    .A(net2253));
 sg13g2_buf_2 fanout2252 (.A(net2253),
    .X(net2252));
 sg13g2_buf_2 fanout2253 (.A(net2254),
    .X(net2253));
 sg13g2_buf_4 fanout2254 (.X(net2254),
    .A(_04033_));
 sg13g2_buf_2 fanout2255 (.A(net2256),
    .X(net2255));
 sg13g2_buf_4 fanout2256 (.X(net2256),
    .A(net2259));
 sg13g2_buf_2 fanout2257 (.A(net2259),
    .X(net2257));
 sg13g2_buf_2 fanout2258 (.A(net2259),
    .X(net2258));
 sg13g2_buf_4 fanout2259 (.X(net2259),
    .A(net2265));
 sg13g2_buf_2 fanout2260 (.A(net2262),
    .X(net2260));
 sg13g2_buf_2 fanout2261 (.A(net2262),
    .X(net2261));
 sg13g2_buf_2 fanout2262 (.A(net2265),
    .X(net2262));
 sg13g2_buf_4 fanout2263 (.X(net2263),
    .A(net2265));
 sg13g2_buf_2 fanout2264 (.A(net2265),
    .X(net2264));
 sg13g2_buf_2 fanout2265 (.A(_04000_),
    .X(net2265));
 sg13g2_buf_2 fanout2266 (.A(net2268),
    .X(net2266));
 sg13g2_buf_1 fanout2267 (.A(net2268),
    .X(net2267));
 sg13g2_buf_4 fanout2268 (.X(net2268),
    .A(net2276));
 sg13g2_buf_2 fanout2269 (.A(net2270),
    .X(net2269));
 sg13g2_buf_4 fanout2270 (.X(net2270),
    .A(net2276));
 sg13g2_buf_1 fanout2271 (.A(net2276),
    .X(net2271));
 sg13g2_buf_2 fanout2272 (.A(net2273),
    .X(net2272));
 sg13g2_buf_4 fanout2273 (.X(net2273),
    .A(net2275));
 sg13g2_buf_2 fanout2274 (.A(net2275),
    .X(net2274));
 sg13g2_buf_4 fanout2275 (.X(net2275),
    .A(net2276));
 sg13g2_buf_2 fanout2276 (.A(_03968_),
    .X(net2276));
 sg13g2_buf_2 fanout2277 (.A(net2278),
    .X(net2277));
 sg13g2_buf_4 fanout2278 (.X(net2278),
    .A(net2282));
 sg13g2_buf_2 fanout2279 (.A(net2281),
    .X(net2279));
 sg13g2_buf_1 fanout2280 (.A(net2281),
    .X(net2280));
 sg13g2_buf_4 fanout2281 (.X(net2281),
    .A(net2282));
 sg13g2_buf_2 fanout2282 (.A(_03936_),
    .X(net2282));
 sg13g2_buf_2 fanout2283 (.A(net2287),
    .X(net2283));
 sg13g2_buf_2 fanout2284 (.A(net2287),
    .X(net2284));
 sg13g2_buf_2 fanout2285 (.A(net2287),
    .X(net2285));
 sg13g2_buf_1 fanout2286 (.A(net2287),
    .X(net2286));
 sg13g2_buf_2 fanout2287 (.A(_03936_),
    .X(net2287));
 sg13g2_buf_2 fanout2288 (.A(net2292),
    .X(net2288));
 sg13g2_buf_2 fanout2289 (.A(net2292),
    .X(net2289));
 sg13g2_buf_2 fanout2290 (.A(net2291),
    .X(net2290));
 sg13g2_buf_4 fanout2291 (.X(net2291),
    .A(net2292));
 sg13g2_buf_4 fanout2292 (.X(net2292),
    .A(_03903_));
 sg13g2_buf_4 fanout2293 (.X(net2293),
    .A(net2294));
 sg13g2_buf_4 fanout2294 (.X(net2294),
    .A(net2296));
 sg13g2_buf_4 fanout2295 (.X(net2295),
    .A(net2296));
 sg13g2_buf_4 fanout2296 (.X(net2296),
    .A(_03903_));
 sg13g2_buf_4 fanout2297 (.X(net2297),
    .A(net2301));
 sg13g2_buf_2 fanout2298 (.A(net2301),
    .X(net2298));
 sg13g2_buf_2 fanout2299 (.A(net2300),
    .X(net2299));
 sg13g2_buf_4 fanout2300 (.X(net2300),
    .A(net2301));
 sg13g2_buf_4 fanout2301 (.X(net2301),
    .A(_03531_));
 sg13g2_buf_4 fanout2302 (.X(net2302),
    .A(net2306));
 sg13g2_buf_4 fanout2303 (.X(net2303),
    .A(net2306));
 sg13g2_buf_4 fanout2304 (.X(net2304),
    .A(net2306));
 sg13g2_buf_1 fanout2305 (.A(net2306),
    .X(net2305));
 sg13g2_buf_2 fanout2306 (.A(_03531_),
    .X(net2306));
 sg13g2_buf_2 fanout2307 (.A(net2308),
    .X(net2307));
 sg13g2_buf_2 fanout2308 (.A(_02722_),
    .X(net2308));
 sg13g2_buf_2 fanout2309 (.A(_02721_),
    .X(net2309));
 sg13g2_buf_2 fanout2310 (.A(_02721_),
    .X(net2310));
 sg13g2_buf_2 fanout2311 (.A(_02023_),
    .X(net2311));
 sg13g2_buf_2 fanout2312 (.A(_02018_),
    .X(net2312));
 sg13g2_buf_2 fanout2313 (.A(_01485_),
    .X(net2313));
 sg13g2_buf_2 fanout2314 (.A(_01479_),
    .X(net2314));
 sg13g2_buf_2 fanout2315 (.A(_01479_),
    .X(net2315));
 sg13g2_buf_2 fanout2316 (.A(net2317),
    .X(net2316));
 sg13g2_buf_2 fanout2317 (.A(_01478_),
    .X(net2317));
 sg13g2_buf_4 fanout2318 (.X(net2318),
    .A(_01456_));
 sg13g2_buf_2 fanout2319 (.A(_01453_),
    .X(net2319));
 sg13g2_buf_1 fanout2320 (.A(_01453_),
    .X(net2320));
 sg13g2_buf_2 fanout2321 (.A(_01277_),
    .X(net2321));
 sg13g2_buf_2 fanout2322 (.A(_01238_),
    .X(net2322));
 sg13g2_buf_2 fanout2323 (.A(net2324),
    .X(net2323));
 sg13g2_buf_2 fanout2324 (.A(net2327),
    .X(net2324));
 sg13g2_buf_2 fanout2325 (.A(net2326),
    .X(net2325));
 sg13g2_buf_2 fanout2326 (.A(net2327),
    .X(net2326));
 sg13g2_buf_1 fanout2327 (.A(_04240_),
    .X(net2327));
 sg13g2_buf_4 fanout2328 (.X(net2328),
    .A(net2331));
 sg13g2_buf_2 fanout2329 (.A(net2331),
    .X(net2329));
 sg13g2_buf_4 fanout2330 (.X(net2330),
    .A(net2331));
 sg13g2_buf_2 fanout2331 (.A(net2332),
    .X(net2331));
 sg13g2_buf_2 fanout2332 (.A(net2341),
    .X(net2332));
 sg13g2_buf_2 fanout2333 (.A(net2334),
    .X(net2333));
 sg13g2_buf_2 fanout2334 (.A(net2337),
    .X(net2334));
 sg13g2_buf_2 fanout2335 (.A(net2337),
    .X(net2335));
 sg13g2_buf_1 fanout2336 (.A(net2337),
    .X(net2336));
 sg13g2_buf_2 fanout2337 (.A(net2341),
    .X(net2337));
 sg13g2_buf_4 fanout2338 (.X(net2338),
    .A(net2341));
 sg13g2_buf_2 fanout2339 (.A(net2340),
    .X(net2339));
 sg13g2_buf_2 fanout2340 (.A(net2341),
    .X(net2340));
 sg13g2_buf_2 fanout2341 (.A(_01355_),
    .X(net2341));
 sg13g2_buf_4 fanout2342 (.X(net2342),
    .A(net2347));
 sg13g2_buf_2 fanout2343 (.A(net2347),
    .X(net2343));
 sg13g2_buf_4 fanout2344 (.X(net2344),
    .A(net2345));
 sg13g2_buf_4 fanout2345 (.X(net2345),
    .A(net2346));
 sg13g2_buf_2 fanout2346 (.A(net2347),
    .X(net2346));
 sg13g2_buf_2 fanout2347 (.A(_01345_),
    .X(net2347));
 sg13g2_buf_2 fanout2348 (.A(net2349),
    .X(net2348));
 sg13g2_buf_4 fanout2349 (.X(net2349),
    .A(_01345_));
 sg13g2_buf_4 fanout2350 (.X(net2350),
    .A(net2352));
 sg13g2_buf_2 fanout2351 (.A(net2352),
    .X(net2351));
 sg13g2_buf_4 fanout2352 (.X(net2352),
    .A(net2355));
 sg13g2_buf_2 fanout2353 (.A(net2354),
    .X(net2353));
 sg13g2_buf_4 fanout2354 (.X(net2354),
    .A(net2355));
 sg13g2_buf_2 fanout2355 (.A(_01344_),
    .X(net2355));
 sg13g2_buf_4 fanout2356 (.X(net2356),
    .A(net2357));
 sg13g2_buf_2 fanout2357 (.A(net2364),
    .X(net2357));
 sg13g2_buf_2 fanout2358 (.A(net2359),
    .X(net2358));
 sg13g2_buf_2 fanout2359 (.A(net2364),
    .X(net2359));
 sg13g2_buf_2 fanout2360 (.A(net2361),
    .X(net2360));
 sg13g2_buf_1 fanout2361 (.A(net2362),
    .X(net2361));
 sg13g2_buf_1 fanout2362 (.A(net2363),
    .X(net2362));
 sg13g2_buf_4 fanout2363 (.X(net2363),
    .A(net2364));
 sg13g2_buf_2 fanout2364 (.A(_01335_),
    .X(net2364));
 sg13g2_buf_4 fanout2365 (.X(net2365),
    .A(net2374));
 sg13g2_buf_1 fanout2366 (.A(net2374),
    .X(net2366));
 sg13g2_buf_4 fanout2367 (.X(net2367),
    .A(net2368));
 sg13g2_buf_2 fanout2368 (.A(net2369),
    .X(net2368));
 sg13g2_buf_2 fanout2369 (.A(net2374),
    .X(net2369));
 sg13g2_buf_2 fanout2370 (.A(net2371),
    .X(net2370));
 sg13g2_buf_2 fanout2371 (.A(net2374),
    .X(net2371));
 sg13g2_buf_2 fanout2372 (.A(net2374),
    .X(net2372));
 sg13g2_buf_2 fanout2373 (.A(net2374),
    .X(net2373));
 sg13g2_buf_4 fanout2374 (.X(net2374),
    .A(_01334_));
 sg13g2_buf_2 fanout2375 (.A(net2377),
    .X(net2375));
 sg13g2_buf_1 fanout2376 (.A(net2377),
    .X(net2376));
 sg13g2_buf_2 fanout2377 (.A(net2384),
    .X(net2377));
 sg13g2_buf_2 fanout2378 (.A(net2379),
    .X(net2378));
 sg13g2_buf_2 fanout2379 (.A(net2380),
    .X(net2379));
 sg13g2_buf_2 fanout2380 (.A(net2384),
    .X(net2380));
 sg13g2_buf_2 fanout2381 (.A(net2383),
    .X(net2381));
 sg13g2_buf_2 fanout2382 (.A(net2383),
    .X(net2382));
 sg13g2_buf_2 fanout2383 (.A(net2384),
    .X(net2383));
 sg13g2_buf_2 fanout2384 (.A(_01329_),
    .X(net2384));
 sg13g2_buf_2 fanout2385 (.A(net2386),
    .X(net2385));
 sg13g2_buf_2 fanout2386 (.A(net2389),
    .X(net2386));
 sg13g2_buf_2 fanout2387 (.A(net2388),
    .X(net2387));
 sg13g2_buf_2 fanout2388 (.A(net2389),
    .X(net2388));
 sg13g2_buf_1 fanout2389 (.A(net2396),
    .X(net2389));
 sg13g2_buf_2 fanout2390 (.A(net2393),
    .X(net2390));
 sg13g2_buf_2 fanout2391 (.A(net2393),
    .X(net2391));
 sg13g2_buf_2 fanout2392 (.A(net2393),
    .X(net2392));
 sg13g2_buf_2 fanout2393 (.A(net2396),
    .X(net2393));
 sg13g2_buf_2 fanout2394 (.A(net2395),
    .X(net2394));
 sg13g2_buf_2 fanout2395 (.A(net2396),
    .X(net2395));
 sg13g2_buf_2 fanout2396 (.A(_01328_),
    .X(net2396));
 sg13g2_buf_2 fanout2397 (.A(net2401),
    .X(net2397));
 sg13g2_buf_2 fanout2398 (.A(net2399),
    .X(net2398));
 sg13g2_buf_2 fanout2399 (.A(net2400),
    .X(net2399));
 sg13g2_buf_2 fanout2400 (.A(net2401),
    .X(net2400));
 sg13g2_buf_2 fanout2401 (.A(_01320_),
    .X(net2401));
 sg13g2_buf_2 fanout2402 (.A(net2403),
    .X(net2402));
 sg13g2_buf_4 fanout2403 (.X(net2403),
    .A(_01319_));
 sg13g2_buf_4 fanout2404 (.X(net2404),
    .A(net2405));
 sg13g2_buf_4 fanout2405 (.X(net2405),
    .A(net2413));
 sg13g2_buf_4 fanout2406 (.X(net2406),
    .A(net2408));
 sg13g2_buf_4 fanout2407 (.X(net2407),
    .A(net2408));
 sg13g2_buf_2 fanout2408 (.A(net2413),
    .X(net2408));
 sg13g2_buf_2 fanout2409 (.A(net2410),
    .X(net2409));
 sg13g2_buf_2 fanout2410 (.A(net2411),
    .X(net2410));
 sg13g2_buf_2 fanout2411 (.A(net2412),
    .X(net2411));
 sg13g2_buf_4 fanout2412 (.X(net2412),
    .A(net2413));
 sg13g2_buf_4 fanout2413 (.X(net2413),
    .A(_03584_));
 sg13g2_buf_4 fanout2414 (.X(net2414),
    .A(_01167_));
 sg13g2_buf_4 fanout2415 (.X(net2415),
    .A(_01160_));
 sg13g2_buf_4 fanout2416 (.X(net2416),
    .A(_01152_));
 sg13g2_buf_4 fanout2417 (.X(net2417),
    .A(_01134_));
 sg13g2_buf_2 fanout2418 (.A(_01134_),
    .X(net2418));
 sg13g2_buf_4 fanout2419 (.X(net2419),
    .A(_01125_));
 sg13g2_buf_4 fanout2420 (.X(net2420),
    .A(_01108_));
 sg13g2_buf_4 fanout2421 (.X(net2421),
    .A(_01105_));
 sg13g2_buf_4 fanout2422 (.X(net2422),
    .A(_01088_));
 sg13g2_buf_2 fanout2423 (.A(_01088_),
    .X(net2423));
 sg13g2_buf_4 fanout2424 (.X(net2424),
    .A(_01085_));
 sg13g2_buf_2 fanout2425 (.A(_01085_),
    .X(net2425));
 sg13g2_buf_4 fanout2426 (.X(net2426),
    .A(_01082_));
 sg13g2_buf_2 fanout2427 (.A(_01071_),
    .X(net2427));
 sg13g2_buf_4 fanout2428 (.X(net2428),
    .A(net2429));
 sg13g2_buf_4 fanout2429 (.X(net2429),
    .A(_01068_));
 sg13g2_buf_4 fanout2430 (.X(net2430),
    .A(_01059_));
 sg13g2_buf_4 fanout2431 (.X(net2431),
    .A(net2432));
 sg13g2_buf_4 fanout2432 (.X(net2432),
    .A(_01055_));
 sg13g2_buf_4 fanout2433 (.X(net2433),
    .A(net2434));
 sg13g2_buf_4 fanout2434 (.X(net2434),
    .A(_01043_));
 sg13g2_buf_4 fanout2435 (.X(net2435),
    .A(_01027_));
 sg13g2_buf_4 fanout2436 (.X(net2436),
    .A(_01023_));
 sg13g2_buf_4 fanout2437 (.X(net2437),
    .A(_01014_));
 sg13g2_buf_4 fanout2438 (.X(net2438),
    .A(net2447));
 sg13g2_buf_2 fanout2439 (.A(net2447),
    .X(net2439));
 sg13g2_buf_2 fanout2440 (.A(net2442),
    .X(net2440));
 sg13g2_buf_2 fanout2441 (.A(net2442),
    .X(net2441));
 sg13g2_buf_2 fanout2442 (.A(net2447),
    .X(net2442));
 sg13g2_buf_2 fanout2443 (.A(net2446),
    .X(net2443));
 sg13g2_buf_2 fanout2444 (.A(net2446),
    .X(net2444));
 sg13g2_buf_4 fanout2445 (.X(net2445),
    .A(net2446));
 sg13g2_buf_2 fanout2446 (.A(net2447),
    .X(net2446));
 sg13g2_buf_2 fanout2447 (.A(_00975_),
    .X(net2447));
 sg13g2_buf_2 fanout2448 (.A(_01226_),
    .X(net2448));
 sg13g2_buf_4 fanout2449 (.X(net2449),
    .A(net2450));
 sg13g2_buf_4 fanout2450 (.X(net2450),
    .A(_01009_));
 sg13g2_buf_2 fanout2451 (.A(_01009_),
    .X(net2451));
 sg13g2_buf_4 fanout2452 (.X(net2452),
    .A(net2453));
 sg13g2_buf_4 fanout2453 (.X(net2453),
    .A(net2458));
 sg13g2_buf_4 fanout2454 (.X(net2454),
    .A(net2458));
 sg13g2_buf_2 fanout2455 (.A(net2458),
    .X(net2455));
 sg13g2_buf_4 fanout2456 (.X(net2456),
    .A(net2457));
 sg13g2_buf_2 fanout2457 (.A(net2458),
    .X(net2457));
 sg13g2_buf_2 fanout2458 (.A(_00996_),
    .X(net2458));
 sg13g2_buf_4 fanout2459 (.X(net2459),
    .A(net2460));
 sg13g2_buf_4 fanout2460 (.X(net2460),
    .A(net2463));
 sg13g2_buf_4 fanout2461 (.X(net2461),
    .A(net2463));
 sg13g2_buf_4 fanout2462 (.X(net2462),
    .A(net2463));
 sg13g2_buf_4 fanout2463 (.X(net2463),
    .A(_03595_));
 sg13g2_buf_2 fanout2464 (.A(_01815_),
    .X(net2464));
 sg13g2_buf_1 fanout2465 (.A(_01815_),
    .X(net2465));
 sg13g2_buf_4 fanout2466 (.X(net2466),
    .A(net2467));
 sg13g2_buf_4 fanout2467 (.X(net2467),
    .A(net2470));
 sg13g2_buf_4 fanout2468 (.X(net2468),
    .A(net2469));
 sg13g2_buf_4 fanout2469 (.X(net2469),
    .A(net2470));
 sg13g2_buf_4 fanout2470 (.X(net2470),
    .A(_01557_));
 sg13g2_buf_2 fanout2471 (.A(net2472),
    .X(net2471));
 sg13g2_buf_2 fanout2472 (.A(net2473),
    .X(net2472));
 sg13g2_buf_4 fanout2473 (.X(net2473),
    .A(_01484_));
 sg13g2_buf_2 fanout2474 (.A(net2477),
    .X(net2474));
 sg13g2_buf_2 fanout2475 (.A(net2477),
    .X(net2475));
 sg13g2_buf_2 fanout2476 (.A(net2477),
    .X(net2476));
 sg13g2_buf_2 fanout2477 (.A(_01483_),
    .X(net2477));
 sg13g2_buf_2 fanout2478 (.A(net2479),
    .X(net2478));
 sg13g2_buf_2 fanout2479 (.A(_01483_),
    .X(net2479));
 sg13g2_buf_4 fanout2480 (.X(net2480),
    .A(_01450_));
 sg13g2_buf_2 fanout2481 (.A(net2482),
    .X(net2481));
 sg13g2_buf_2 fanout2482 (.A(net2483),
    .X(net2482));
 sg13g2_buf_2 fanout2483 (.A(_01447_),
    .X(net2483));
 sg13g2_buf_2 fanout2484 (.A(net2486),
    .X(net2484));
 sg13g2_buf_2 fanout2485 (.A(net2486),
    .X(net2485));
 sg13g2_buf_2 fanout2486 (.A(_01446_),
    .X(net2486));
 sg13g2_buf_2 fanout2487 (.A(net2488),
    .X(net2487));
 sg13g2_buf_2 fanout2488 (.A(net2489),
    .X(net2488));
 sg13g2_buf_4 fanout2489 (.X(net2489),
    .A(_01426_));
 sg13g2_buf_4 fanout2490 (.X(net2490),
    .A(net2491));
 sg13g2_buf_2 fanout2491 (.A(_01425_),
    .X(net2491));
 sg13g2_buf_2 fanout2492 (.A(net2494),
    .X(net2492));
 sg13g2_buf_1 fanout2493 (.A(net2494),
    .X(net2493));
 sg13g2_buf_2 fanout2494 (.A(_01425_),
    .X(net2494));
 sg13g2_buf_4 fanout2495 (.X(net2495),
    .A(net2496));
 sg13g2_buf_4 fanout2496 (.X(net2496),
    .A(_01388_));
 sg13g2_buf_2 fanout2497 (.A(net2498),
    .X(net2497));
 sg13g2_buf_2 fanout2498 (.A(net2499),
    .X(net2498));
 sg13g2_buf_2 fanout2499 (.A(_01387_),
    .X(net2499));
 sg13g2_buf_2 fanout2500 (.A(net2504),
    .X(net2500));
 sg13g2_buf_2 fanout2501 (.A(net2503),
    .X(net2501));
 sg13g2_buf_2 fanout2502 (.A(net2503),
    .X(net2502));
 sg13g2_buf_2 fanout2503 (.A(net2504),
    .X(net2503));
 sg13g2_buf_2 fanout2504 (.A(net2505),
    .X(net2504));
 sg13g2_buf_2 fanout2505 (.A(_01219_),
    .X(net2505));
 sg13g2_buf_2 fanout2506 (.A(net2507),
    .X(net2506));
 sg13g2_buf_1 fanout2507 (.A(_01219_),
    .X(net2507));
 sg13g2_buf_4 fanout2508 (.X(net2508),
    .A(_01008_));
 sg13g2_buf_2 fanout2509 (.A(net2512),
    .X(net2509));
 sg13g2_buf_2 fanout2510 (.A(net2512),
    .X(net2510));
 sg13g2_buf_2 fanout2511 (.A(net2512),
    .X(net2511));
 sg13g2_buf_2 fanout2512 (.A(_01007_),
    .X(net2512));
 sg13g2_buf_4 fanout2513 (.X(net2513),
    .A(_01005_));
 sg13g2_buf_2 fanout2514 (.A(net2517),
    .X(net2514));
 sg13g2_buf_2 fanout2515 (.A(net2517),
    .X(net2515));
 sg13g2_buf_2 fanout2516 (.A(net2517),
    .X(net2516));
 sg13g2_buf_2 fanout2517 (.A(_01004_),
    .X(net2517));
 sg13g2_buf_2 fanout2518 (.A(_00994_),
    .X(net2518));
 sg13g2_buf_2 fanout2519 (.A(_00994_),
    .X(net2519));
 sg13g2_buf_2 fanout2520 (.A(_00989_),
    .X(net2520));
 sg13g2_buf_2 fanout2521 (.A(_00989_),
    .X(net2521));
 sg13g2_buf_2 fanout2522 (.A(net2523),
    .X(net2522));
 sg13g2_buf_4 fanout2523 (.X(net2523),
    .A(_00962_));
 sg13g2_buf_2 fanout2524 (.A(_03563_),
    .X(net2524));
 sg13g2_buf_2 fanout2525 (.A(net2526),
    .X(net2525));
 sg13g2_buf_1 fanout2526 (.A(_01175_),
    .X(net2526));
 sg13g2_buf_2 fanout2527 (.A(net2528),
    .X(net2527));
 sg13g2_buf_2 fanout2528 (.A(_00928_),
    .X(net2528));
 sg13g2_buf_4 fanout2529 (.X(net2529),
    .A(_00925_));
 sg13g2_buf_2 fanout2530 (.A(net2531),
    .X(net2530));
 sg13g2_buf_4 fanout2531 (.X(net2531),
    .A(_00923_));
 sg13g2_buf_2 fanout2532 (.A(net2535),
    .X(net2532));
 sg13g2_buf_4 fanout2533 (.X(net2533),
    .A(net2535));
 sg13g2_buf_4 fanout2534 (.X(net2534),
    .A(net2535));
 sg13g2_buf_2 fanout2535 (.A(_00908_),
    .X(net2535));
 sg13g2_buf_2 fanout2536 (.A(net2537),
    .X(net2536));
 sg13g2_buf_2 fanout2537 (.A(net2538),
    .X(net2537));
 sg13g2_buf_1 fanout2538 (.A(net2539),
    .X(net2538));
 sg13g2_buf_2 fanout2539 (.A(net2540),
    .X(net2539));
 sg13g2_buf_2 fanout2540 (.A(net2549),
    .X(net2540));
 sg13g2_buf_2 fanout2541 (.A(net2542),
    .X(net2541));
 sg13g2_buf_2 fanout2542 (.A(net2544),
    .X(net2542));
 sg13g2_buf_2 fanout2543 (.A(net2544),
    .X(net2543));
 sg13g2_buf_1 fanout2544 (.A(net2549),
    .X(net2544));
 sg13g2_buf_2 fanout2545 (.A(net2549),
    .X(net2545));
 sg13g2_buf_2 fanout2546 (.A(net2549),
    .X(net2546));
 sg13g2_buf_2 fanout2547 (.A(net2548),
    .X(net2547));
 sg13g2_buf_2 fanout2548 (.A(net2549),
    .X(net2548));
 sg13g2_buf_2 fanout2549 (.A(_00907_),
    .X(net2549));
 sg13g2_buf_4 fanout2550 (.X(net2550),
    .A(net1522));
 sg13g2_buf_2 fanout2551 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[4] ),
    .X(net2551));
 sg13g2_buf_2 fanout2552 (.A(net860),
    .X(net2552));
 sg13g2_buf_2 fanout2553 (.A(net856),
    .X(net2553));
 sg13g2_buf_4 fanout2554 (.X(net2554),
    .A(net2555));
 sg13g2_buf_4 fanout2555 (.X(net2555),
    .A(net2559));
 sg13g2_buf_2 fanout2556 (.A(net2558),
    .X(net2556));
 sg13g2_buf_1 fanout2557 (.A(net2558),
    .X(net2557));
 sg13g2_buf_4 fanout2558 (.X(net2558),
    .A(net2559));
 sg13g2_buf_4 fanout2559 (.X(net2559),
    .A(\ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[2] ));
 sg13g2_buf_4 fanout2560 (.X(net2560),
    .A(net2564));
 sg13g2_buf_4 fanout2561 (.X(net2561),
    .A(net2564));
 sg13g2_buf_4 fanout2562 (.X(net2562),
    .A(net2564));
 sg13g2_buf_2 fanout2563 (.A(net2564),
    .X(net2563));
 sg13g2_buf_2 fanout2564 (.A(\ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[2] ),
    .X(net2564));
 sg13g2_buf_4 fanout2565 (.X(net2565),
    .A(net2569));
 sg13g2_buf_2 fanout2566 (.A(net2569),
    .X(net2566));
 sg13g2_buf_4 fanout2567 (.X(net2567),
    .A(net2569));
 sg13g2_buf_2 fanout2568 (.A(net2569),
    .X(net2568));
 sg13g2_buf_2 fanout2569 (.A(net2582),
    .X(net2569));
 sg13g2_buf_4 fanout2570 (.X(net2570),
    .A(net2571));
 sg13g2_buf_4 fanout2571 (.X(net2571),
    .A(net2573));
 sg13g2_buf_4 fanout2572 (.X(net2572),
    .A(net2573));
 sg13g2_buf_2 fanout2573 (.A(net2582),
    .X(net2573));
 sg13g2_buf_4 fanout2574 (.X(net2574),
    .A(net2578));
 sg13g2_buf_2 fanout2575 (.A(net2578),
    .X(net2575));
 sg13g2_buf_4 fanout2576 (.X(net2576),
    .A(net2578));
 sg13g2_buf_2 fanout2577 (.A(net2578),
    .X(net2577));
 sg13g2_buf_2 fanout2578 (.A(net2582),
    .X(net2578));
 sg13g2_buf_4 fanout2579 (.X(net2579),
    .A(net2581));
 sg13g2_buf_2 fanout2580 (.A(net2581),
    .X(net2580));
 sg13g2_buf_4 fanout2581 (.X(net2581),
    .A(net2582));
 sg13g2_buf_4 fanout2582 (.X(net2582),
    .A(\ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[1] ));
 sg13g2_buf_4 fanout2583 (.X(net2583),
    .A(net2590));
 sg13g2_buf_2 fanout2584 (.A(net2585),
    .X(net2584));
 sg13g2_buf_2 fanout2585 (.A(net2590),
    .X(net2585));
 sg13g2_buf_2 fanout2586 (.A(net2589),
    .X(net2586));
 sg13g2_buf_2 fanout2587 (.A(net2589),
    .X(net2587));
 sg13g2_buf_4 fanout2588 (.X(net2588),
    .A(net2589));
 sg13g2_buf_4 fanout2589 (.X(net2589),
    .A(net2590));
 sg13g2_buf_2 fanout2590 (.A(net2610),
    .X(net2590));
 sg13g2_buf_2 fanout2591 (.A(net2592),
    .X(net2591));
 sg13g2_buf_2 fanout2592 (.A(net2597),
    .X(net2592));
 sg13g2_buf_2 fanout2593 (.A(net2594),
    .X(net2593));
 sg13g2_buf_4 fanout2594 (.X(net2594),
    .A(net2597));
 sg13g2_buf_4 fanout2595 (.X(net2595),
    .A(net2596));
 sg13g2_buf_2 fanout2596 (.A(net2597),
    .X(net2596));
 sg13g2_buf_2 fanout2597 (.A(net2610),
    .X(net2597));
 sg13g2_buf_2 fanout2598 (.A(net2601),
    .X(net2598));
 sg13g2_buf_2 fanout2599 (.A(net2601),
    .X(net2599));
 sg13g2_buf_4 fanout2600 (.X(net2600),
    .A(net2601));
 sg13g2_buf_1 fanout2601 (.A(net2610),
    .X(net2601));
 sg13g2_buf_2 fanout2602 (.A(net2604),
    .X(net2602));
 sg13g2_buf_4 fanout2603 (.X(net2603),
    .A(net2604));
 sg13g2_buf_2 fanout2604 (.A(net2610),
    .X(net2604));
 sg13g2_buf_4 fanout2605 (.X(net2605),
    .A(net2609));
 sg13g2_buf_4 fanout2606 (.X(net2606),
    .A(net2608));
 sg13g2_buf_4 fanout2607 (.X(net2607),
    .A(net2608));
 sg13g2_buf_2 fanout2608 (.A(net2609),
    .X(net2608));
 sg13g2_buf_1 fanout2609 (.A(net2610),
    .X(net2609));
 sg13g2_buf_4 fanout2610 (.X(net2610),
    .A(\ChiselTop.wild.cpu.regs_rs2Val_MPORT_addr[0] ));
 sg13g2_buf_2 fanout2611 (.A(\ChiselTop.wild.cpu.decExReg_func3[1] ),
    .X(net2611));
 sg13g2_buf_4 fanout2612 (.X(net2612),
    .A(net1520));
 sg13g2_buf_2 fanout2613 (.A(net2614),
    .X(net2613));
 sg13g2_buf_2 fanout2614 (.A(net2615),
    .X(net2614));
 sg13g2_buf_2 fanout2615 (.A(net1470),
    .X(net2615));
 sg13g2_buf_2 fanout2616 (.A(net2617),
    .X(net2616));
 sg13g2_buf_1 fanout2617 (.A(net2620),
    .X(net2617));
 sg13g2_buf_2 fanout2618 (.A(net2619),
    .X(net2618));
 sg13g2_buf_2 fanout2619 (.A(net2620),
    .X(net2619));
 sg13g2_buf_2 fanout2620 (.A(net1046),
    .X(net2620));
 sg13g2_buf_2 fanout2621 (.A(\ChiselTop.wild.cpu.decExReg_memLow[0] ),
    .X(net2621));
 sg13g2_buf_2 fanout2622 (.A(\ChiselTop.wild.cpu.decExReg_decOut_isCssrw ),
    .X(net2622));
 sg13g2_buf_2 fanout2623 (.A(net2626),
    .X(net2623));
 sg13g2_buf_2 fanout2624 (.A(net2625),
    .X(net2624));
 sg13g2_buf_2 fanout2625 (.A(net2626),
    .X(net2625));
 sg13g2_buf_2 fanout2626 (.A(\ChiselTop.wild.cpu.decExReg_decOut_isAuiPc ),
    .X(net2626));
 sg13g2_buf_2 fanout2627 (.A(net2631),
    .X(net2627));
 sg13g2_buf_2 fanout2628 (.A(net2631),
    .X(net2628));
 sg13g2_buf_2 fanout2629 (.A(net2631),
    .X(net2629));
 sg13g2_buf_2 fanout2630 (.A(net2631),
    .X(net2630));
 sg13g2_buf_1 fanout2631 (.A(\ChiselTop.wild.cpu.decExReg_decOut_isAuiPc ),
    .X(net2631));
 sg13g2_buf_2 fanout2632 (.A(net2634),
    .X(net2632));
 sg13g2_buf_2 fanout2633 (.A(net2634),
    .X(net2633));
 sg13g2_buf_2 fanout2634 (.A(net2637),
    .X(net2634));
 sg13g2_buf_4 fanout2635 (.X(net2635),
    .A(net2637));
 sg13g2_buf_1 fanout2636 (.A(net2637),
    .X(net2636));
 sg13g2_buf_2 fanout2637 (.A(\ChiselTop.wild.cpu.decExReg_decOut_isLui ),
    .X(net2637));
 sg13g2_buf_2 fanout2638 (.A(net2639),
    .X(net2638));
 sg13g2_buf_2 fanout2639 (.A(\ChiselTop.wild.cpu.decExReg_decOut_isLui ),
    .X(net2639));
 sg13g2_buf_4 fanout2640 (.X(net2640),
    .A(\ChiselTop.wild.cpu.decExReg_decOut_aluOp[0] ));
 sg13g2_buf_2 fanout2641 (.A(net2642),
    .X(net2641));
 sg13g2_buf_2 fanout2642 (.A(net2647),
    .X(net2642));
 sg13g2_buf_2 fanout2643 (.A(net2647),
    .X(net2643));
 sg13g2_buf_1 fanout2644 (.A(net2647),
    .X(net2644));
 sg13g2_buf_4 fanout2645 (.X(net2645),
    .A(net2646));
 sg13g2_buf_2 fanout2646 (.A(net2647),
    .X(net2646));
 sg13g2_buf_2 fanout2647 (.A(\ChiselTop.wild.cpu.decExReg_decOut_isImm ),
    .X(net2647));
 sg13g2_buf_4 fanout2648 (.X(net2648),
    .A(net1517));
 sg13g2_buf_4 fanout2649 (.X(net2649),
    .A(net1529));
 sg13g2_buf_2 fanout2650 (.A(\ChiselTop.dec.counter[3] ),
    .X(net2650));
 sg13g2_buf_4 fanout2651 (.X(net2651),
    .A(net2652));
 sg13g2_buf_4 fanout2652 (.X(net2652),
    .A(net2656));
 sg13g2_buf_4 fanout2653 (.X(net2653),
    .A(net2655));
 sg13g2_buf_1 fanout2654 (.A(net2655),
    .X(net2654));
 sg13g2_buf_2 fanout2655 (.A(net2656),
    .X(net2655));
 sg13g2_buf_4 fanout2656 (.X(net2656),
    .A(net1537));
 sg13g2_buf_4 fanout2657 (.X(net2657),
    .A(net2661));
 sg13g2_buf_2 fanout2658 (.A(net2661),
    .X(net2658));
 sg13g2_buf_4 fanout2659 (.X(net2659),
    .A(net2661));
 sg13g2_buf_4 fanout2660 (.X(net2660),
    .A(net2661));
 sg13g2_buf_4 fanout2661 (.X(net2661),
    .A(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[2] ));
 sg13g2_buf_4 fanout2662 (.X(net2662),
    .A(net2665));
 sg13g2_buf_4 fanout2663 (.X(net2663),
    .A(net2664));
 sg13g2_buf_4 fanout2664 (.X(net2664),
    .A(net2665));
 sg13g2_buf_2 fanout2665 (.A(net2669),
    .X(net2665));
 sg13g2_buf_2 fanout2666 (.A(net2667),
    .X(net2666));
 sg13g2_buf_4 fanout2667 (.X(net2667),
    .A(net2668));
 sg13g2_buf_4 fanout2668 (.X(net2668),
    .A(net2669));
 sg13g2_buf_4 fanout2669 (.X(net2669),
    .A(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[1] ));
 sg13g2_buf_4 fanout2670 (.X(net2670),
    .A(net2674));
 sg13g2_buf_2 fanout2671 (.A(net2674),
    .X(net2671));
 sg13g2_buf_4 fanout2672 (.X(net2672),
    .A(net2674));
 sg13g2_buf_4 fanout2673 (.X(net2673),
    .A(net2674));
 sg13g2_buf_2 fanout2674 (.A(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[1] ),
    .X(net2674));
 sg13g2_buf_4 fanout2675 (.X(net2675),
    .A(net2676));
 sg13g2_buf_4 fanout2676 (.X(net2676),
    .A(net2677));
 sg13g2_buf_2 fanout2677 (.A(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[1] ),
    .X(net2677));
 sg13g2_buf_2 fanout2678 (.A(net2679),
    .X(net2678));
 sg13g2_buf_4 fanout2679 (.X(net2679),
    .A(net2691));
 sg13g2_buf_4 fanout2680 (.X(net2680),
    .A(net2681));
 sg13g2_buf_2 fanout2681 (.A(net2682),
    .X(net2681));
 sg13g2_buf_4 fanout2682 (.X(net2682),
    .A(net2691));
 sg13g2_buf_1 fanout2683 (.A(net2691),
    .X(net2683));
 sg13g2_buf_2 fanout2684 (.A(net2688),
    .X(net2684));
 sg13g2_buf_1 fanout2685 (.A(net2688),
    .X(net2685));
 sg13g2_buf_2 fanout2686 (.A(net2688),
    .X(net2686));
 sg13g2_buf_4 fanout2687 (.X(net2687),
    .A(net2688));
 sg13g2_buf_4 fanout2688 (.X(net2688),
    .A(net2690));
 sg13g2_buf_4 fanout2689 (.X(net2689),
    .A(net2690));
 sg13g2_buf_2 fanout2690 (.A(net2691),
    .X(net2690));
 sg13g2_buf_4 fanout2691 (.X(net2691),
    .A(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[0] ));
 sg13g2_buf_4 fanout2692 (.X(net2692),
    .A(net2694));
 sg13g2_buf_1 fanout2693 (.A(net2694),
    .X(net2693));
 sg13g2_buf_4 fanout2694 (.X(net2694),
    .A(net2699));
 sg13g2_buf_4 fanout2695 (.X(net2695),
    .A(net2696));
 sg13g2_buf_2 fanout2696 (.A(net2699),
    .X(net2696));
 sg13g2_buf_4 fanout2697 (.X(net2697),
    .A(net2699));
 sg13g2_buf_1 fanout2698 (.A(net2699),
    .X(net2698));
 sg13g2_buf_4 fanout2699 (.X(net2699),
    .A(net2705));
 sg13g2_buf_4 fanout2700 (.X(net2700),
    .A(net2705));
 sg13g2_buf_2 fanout2701 (.A(net2702),
    .X(net2701));
 sg13g2_buf_4 fanout2702 (.X(net2702),
    .A(net2704));
 sg13g2_buf_4 fanout2703 (.X(net2703),
    .A(net2704));
 sg13g2_buf_1 fanout2704 (.A(net2705),
    .X(net2704));
 sg13g2_buf_2 fanout2705 (.A(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[0] ),
    .X(net2705));
 sg13g2_buf_4 fanout2706 (.X(net2706),
    .A(net2713));
 sg13g2_buf_2 fanout2707 (.A(net2713),
    .X(net2707));
 sg13g2_buf_2 fanout2708 (.A(net2709),
    .X(net2708));
 sg13g2_buf_4 fanout2709 (.X(net2709),
    .A(net2713));
 sg13g2_buf_4 fanout2710 (.X(net2710),
    .A(net2712));
 sg13g2_buf_2 fanout2711 (.A(net2712),
    .X(net2711));
 sg13g2_buf_2 fanout2712 (.A(net2713),
    .X(net2712));
 sg13g2_buf_2 fanout2713 (.A(net2728),
    .X(net2713));
 sg13g2_buf_4 fanout2714 (.X(net2714),
    .A(net2716));
 sg13g2_buf_4 fanout2715 (.X(net2715),
    .A(net2716));
 sg13g2_buf_2 fanout2716 (.A(net2728),
    .X(net2716));
 sg13g2_buf_4 fanout2717 (.X(net2717),
    .A(net2719));
 sg13g2_buf_4 fanout2718 (.X(net2718),
    .A(net2719));
 sg13g2_buf_4 fanout2719 (.X(net2719),
    .A(net2728));
 sg13g2_buf_4 fanout2720 (.X(net2720),
    .A(net2727));
 sg13g2_buf_2 fanout2721 (.A(net2727),
    .X(net2721));
 sg13g2_buf_4 fanout2722 (.X(net2722),
    .A(net2725));
 sg13g2_buf_2 fanout2723 (.A(net2724),
    .X(net2723));
 sg13g2_buf_2 fanout2724 (.A(net2725),
    .X(net2724));
 sg13g2_buf_2 fanout2725 (.A(net2727),
    .X(net2725));
 sg13g2_buf_4 fanout2726 (.X(net2726),
    .A(net2727));
 sg13g2_buf_4 fanout2727 (.X(net2727),
    .A(net2728));
 sg13g2_buf_4 fanout2728 (.X(net2728),
    .A(_00943_));
 sg13g2_buf_4 fanout2729 (.X(net2729),
    .A(net2745));
 sg13g2_buf_2 fanout2730 (.A(net2731),
    .X(net2730));
 sg13g2_buf_2 fanout2731 (.A(net2732),
    .X(net2731));
 sg13g2_buf_2 fanout2732 (.A(net2735),
    .X(net2732));
 sg13g2_buf_2 fanout2733 (.A(net2734),
    .X(net2733));
 sg13g2_buf_2 fanout2734 (.A(net2735),
    .X(net2734));
 sg13g2_buf_4 fanout2735 (.X(net2735),
    .A(net2745));
 sg13g2_buf_2 fanout2736 (.A(net2738),
    .X(net2736));
 sg13g2_buf_2 fanout2737 (.A(net2738),
    .X(net2737));
 sg13g2_buf_2 fanout2738 (.A(net2739),
    .X(net2738));
 sg13g2_buf_2 fanout2739 (.A(net2744),
    .X(net2739));
 sg13g2_buf_2 fanout2740 (.A(net2742),
    .X(net2740));
 sg13g2_buf_1 fanout2741 (.A(net2742),
    .X(net2741));
 sg13g2_buf_2 fanout2742 (.A(net2744),
    .X(net2742));
 sg13g2_buf_4 fanout2743 (.X(net2743),
    .A(net2744));
 sg13g2_buf_2 fanout2744 (.A(net2745),
    .X(net2744));
 sg13g2_buf_2 fanout2745 (.A(rst_n),
    .X(net2745));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_schoeberl_wildcat_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_leaf_97_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_2 clkbuf_leaf_98_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_2 clkbuf_leaf_99_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_2 clkbuf_leaf_100_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_2 clkbuf_leaf_101_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_2 clkbuf_leaf_102_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_2 clkbuf_leaf_103_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_2 clkbuf_leaf_104_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_2 clkbuf_leaf_105_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_2 clkbuf_leaf_106_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_2 clkbuf_leaf_107_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_2 clkbuf_leaf_108_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_2 clkbuf_leaf_109_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_4_8_0_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload10 (.A(clknet_4_12_0_clk));
 sg13g2_buf_1 clkload11 (.A(clknet_4_13_0_clk));
 sg13g2_buf_1 clkload12 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_108_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_109_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_101_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_104_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_90_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_12_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_93_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_82_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_83_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_84_clk));
 sg13g2_inv_8 clkload27 (.A(clknet_leaf_85_clk));
 sg13g2_inv_8 clkload28 (.A(clknet_leaf_73_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_78_clk));
 sg13g2_inv_4 clkload30 (.A(clknet_leaf_44_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_47_clk));
 sg13g2_inv_4 clkload32 (.A(clknet_leaf_39_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_50_clk));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_63_clk));
 sg13g2_inv_2 clkload35 (.A(clknet_leaf_58_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ChiselTop.wild.tx.buf_.io_in_ready ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ChiselTop.wild.ledReg[3] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold3 (.A(\ChiselTop.wild.cpu.pcReg[18] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold4 (.A(\ChiselTop.wild.cpu._pcNext_T_1[0] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ChiselTop.wild.ledReg[1] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold6 (.A(\ChiselTop.wild.ledReg[2] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold7 (.A(\ChiselTop.wild.cpu.pcReg[6] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold8 (.A(\ChiselTop.wild.cpu._pcNext_T_1[1] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold9 (.A(\ChiselTop.wild.ledReg[0] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold10 (.A(\ChiselTop.wild.cpu.pcReg[15] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold11 (.A(\ChiselTop.wild.cpu.pcReg[14] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold12 (.A(\ChiselTop.wild.cpu.pcReg[21] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ChiselTop.wild.cpu.pcReg[11] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold14 (.A(\ChiselTop.wild.cpu.pcReg[27] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold15 (.A(\ChiselTop.wild.cpu.pcReg[31] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ChiselTop.wild.cpu.pcReg[19] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold17 (.A(\ChiselTop.wild.cpu.pcReg[24] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold18 (.A(\ChiselTop.wild.cpu.pcReg[28] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold19 (.A(\ChiselTop.wild.cpu.pcReg[9] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold20 (.A(\ChiselTop.wild.cpu.pcReg[23] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold21 (.A(\ChiselTop.wild.cpu.pcReg[22] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ChiselTop.wild.cpu.pcReg[30] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold23 (.A(\ChiselTop.wild.cpu.pcReg[26] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ChiselTop.wild.cpu.pcReg[8] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold25 (.A(\ChiselTop.wild.cpu.pcReg[25] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ChiselTop.wild.cpu.pcReg[17] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold27 (.A(\ChiselTop.wild.cpu.pcReg[12] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold28 (.A(\ChiselTop._cntReg_T_1[0] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ChiselTop.wild.rx.io_channel_valid ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ChiselTop.wild.cpu.pcReg[29] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold31 (.A(\ChiselTop.wild.cpu.pcReg[4] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold32 (.A(\ChiselTop.wild.cpu.pcReg[20] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold33 (.A(\ChiselTop.wild.cpu.pcReg[16] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold34 (.A(_00137_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold35 (.A(\ChiselTop.wild.cpu.pcReg[5] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold36 (.A(_00000_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold37 (.A(_00892_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold38 (.A(\ChiselTop.wild.cpu.pcReg[10] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold39 (.A(\ChiselTop.wild.rx._shiftReg_T_1[7] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold40 (.A(\ChiselTop.wild.cpu.pcReg[13] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold41 (.A(\ChiselTop.wild.cpu.pcReg[7] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold42 (.A(\ChiselTop.wild.cpu.pcRegReg[10] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold43 (.A(\ChiselTop.wild.cpu.pcRegReg[30] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold44 (.A(_00139_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold45 (.A(_00856_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold46 (.A(\ChiselTop.wild.cpu.pcRegReg[9] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold47 (.A(\ChiselTop.wild.cpu.pcRegReg[17] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold48 (.A(\ChiselTop.wild.cpu.pcRegReg[18] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold49 (.A(\ChiselTop.wild.cpu.pcRegReg[28] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold50 (.A(\ChiselTop.wild.cpu.pcRegReg[7] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold51 (.A(\ChiselTop.wild.cpu.pcRegReg[13] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ChiselTop.wild.cpu.pcRegReg[14] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold53 (.A(\ChiselTop.wild.cpu.pcRegReg[11] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ChiselTop.wild.cpu.pcRegReg[16] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold55 (.A(\ChiselTop.wild.cpu.pcRegReg[20] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold56 (.A(\ChiselTop.wild.cpu.pcRegReg[5] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold57 (.A(\ChiselTop.wild.cpu.pcRegReg[3] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold58 (.A(\ChiselTop.wild.cpu.pcRegReg[23] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold59 (.A(\ChiselTop.wild.cpu.pcRegReg[31] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold60 (.A(\ChiselTop.wild.cpu.pcRegReg[27] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold61 (.A(\ChiselTop.wild.cpu.pcRegReg[22] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ChiselTop.wild.cpu.pcRegReg[1] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold63 (.A(\ChiselTop.wild.cpu.pcRegReg[8] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ChiselTop.wild.cpu.pcRegReg[4] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold65 (.A(\ChiselTop.wild.cpu.pcRegReg[12] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold66 (.A(\ChiselTop.wild.cpu.pcRegReg[25] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold67 (.A(\ChiselTop.wild.cpu.pcRegReg[26] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold68 (.A(\ChiselTop.wild.cpu.pcRegReg[29] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[3] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold70 (.A(\ChiselTop.wild.cpu.pcRegReg[0] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ChiselTop.wild.cpu.pcRegReg[21] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold72 (.A(\ChiselTop.wild.rx.rxReg_REG ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ChiselTop.wild.cpu.pcRegReg[2] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold74 (.A(\ChiselTop.wild.cpu.pcRegReg[19] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold75 (.A(\ChiselTop.wild.cpu.pcRegReg[6] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold76 (.A(\ChiselTop.wild.cpu.pcRegReg[24] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold77 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[2] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold78 (.A(\ChiselTop.wild.cpu.pcRegReg[15] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold79 (.A(\ChiselTop.wild.cpu.regs[0][31] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold80 (.A(\ChiselTop.wild.cpu.regs[0][25] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold81 (.A(\ChiselTop.wild.cpu.regs[0][8] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold82 (.A(\ChiselTop.wild.cpu.regs[0][13] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold83 (.A(\ChiselTop.wild.cpu.regs[0][3] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold84 (.A(\ChiselTop.wild.cpu.regs[0][4] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold85 (.A(\ChiselTop.wild.cpu.regs[0][0] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold86 (.A(\ChiselTop.wild.cpu.regs[0][7] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold87 (.A(\ChiselTop.wild.cpu.regs[0][20] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold88 (.A(\ChiselTop.wild.cpu.regs[0][21] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold89 (.A(\ChiselTop.wild.cpu.regs[0][19] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold90 (.A(\ChiselTop.wild.cpu.regs[0][27] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold91 (.A(\ChiselTop.wild.cpu.regs[0][15] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold92 (.A(\ChiselTop.wild.cpu.regs[0][10] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold93 (.A(\ChiselTop.wild.cpu.regs[0][30] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold94 (.A(\ChiselTop.wild.cpu.regs[0][9] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold95 (.A(\ChiselTop.wild.cpu.regs[0][16] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold96 (.A(\ChiselTop.wild.cpu.regs[0][22] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold97 (.A(\ChiselTop.wild.cpu.regs[0][6] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold98 (.A(\ChiselTop.wild.cpu.regs[0][5] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold99 (.A(\ChiselTop.wild.tx.tx.bitsReg[3] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold100 (.A(_04583_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold101 (.A(\ChiselTop.wild.cpu.regs[0][29] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold102 (.A(\ChiselTop.wild.cpu.regs[0][23] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold103 (.A(\ChiselTop.wild.cpu.regs[0][11] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold104 (.A(\ChiselTop.wild.cpu.regs[0][12] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold105 (.A(\ChiselTop.wild.tx.tx.cntReg[19] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold106 (.A(_00156_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold107 (.A(\ChiselTop.wild.cpu.regs[0][1] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold108 (.A(\ChiselTop.wild.cpu.regs[0][14] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold109 (.A(\ChiselTop.wild.cpu.regs[0][2] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold110 (.A(\ChiselTop.wild.cpu.regs[0][18] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold111 (.A(\ChiselTop.wild.cpu.regs[0][26] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold112 (.A(\ChiselTop.wild.tx.tx.cntReg[0] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold113 (.A(\ChiselTop.wild.cpu.regs[0][24] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold114 (.A(_00140_),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold115 (.A(_04649_),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold116 (.A(\ChiselTop.wild.cpu.regs[0][17] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold117 (.A(\ChiselTop.wild.cpu.regs[0][28] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold118 (.A(\ChiselTop.wild.cpu.regs[29][10] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold119 (.A(\ChiselTop.wild.cpu.regs[28][4] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ChiselTop.wild.cpu.regs[5][10] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold121 (.A(\ChiselTop.wild.cpu.regs[28][31] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold122 (.A(\ChiselTop.wild.cpu.regs[31][25] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold123 (.A(\ChiselTop.wild.cpu.regs[5][22] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold124 (.A(\ChiselTop.wild.cpu.regs[29][24] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold125 (.A(\ChiselTop.wild.cpu.regs[5][24] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold126 (.A(\ChiselTop.wild.cpu.regs[29][14] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold127 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[16] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold128 (.A(\ChiselTop.wild.cpu.regs[7][28] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold129 (.A(\ChiselTop.wild.cpu.regs[31][23] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold130 (.A(\ChiselTop.wild.cpu.regs[28][18] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold131 (.A(\ChiselTop.wild.cpu.regs[31][22] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold132 (.A(\ChiselTop.wild.cpu.regs[29][21] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold133 (.A(\ChiselTop.wild.cpu.regs[6][1] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold134 (.A(\ChiselTop.wild.cpu.regs[29][5] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold135 (.A(\ChiselTop.wild.cpu.regs[28][28] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ChiselTop.wild.cpu.regs[7][29] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold137 (.A(\ChiselTop.wild.cpu.regs[31][4] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold138 (.A(\ChiselTop.wild.cpu.regs[31][0] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold139 (.A(\ChiselTop.wild.cpu.regs[5][17] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold140 (.A(\ChiselTop.wild.cpu.regs[28][23] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold141 (.A(\ChiselTop.wild.cpu.regs[7][20] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold142 (.A(\ChiselTop.wild.cpu.regs[7][4] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold143 (.A(\ChiselTop.wild.cpu.regs[4][0] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold144 (.A(\ChiselTop.wild.cpu.regs[29][0] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold145 (.A(\ChiselTop.wild.cpu.regs[28][0] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold146 (.A(\ChiselTop.wild.cpu.regs[5][30] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold147 (.A(\ChiselTop.wild.cpu.regs[6][3] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold148 (.A(\ChiselTop.wild.cpu.regs[4][3] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold149 (.A(\ChiselTop.wild.cpu.regs[29][7] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold150 (.A(\ChiselTop.wild.cpu.regs[29][1] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold151 (.A(\ChiselTop.wild.cpu.regs[29][12] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold152 (.A(\ChiselTop.wild.cpu.regs[7][25] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold153 (.A(\ChiselTop.wild.cpu.regs[29][27] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold154 (.A(\ChiselTop.wild.cpu.regs[29][31] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold155 (.A(\ChiselTop.wild.cpu.regs[7][14] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold156 (.A(\ChiselTop.wild.cpu.regs[6][30] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold157 (.A(\ChiselTop.wild.cpu.regs[4][2] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold158 (.A(\ChiselTop.wild.cpu.regs[29][2] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold159 (.A(\ChiselTop.wild.cpu.regs[7][0] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold160 (.A(\ChiselTop.wild.cpu.regs[28][10] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold161 (.A(\ChiselTop.wild.cpu.regs[31][24] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold162 (.A(\ChiselTop.wild.cpu.regs[30][9] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold163 (.A(\ChiselTop.wild.cpu.regs[30][16] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold164 (.A(\ChiselTop.wild.cpu.regs[28][1] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold165 (.A(\ChiselTop.wild.cpu.regs[5][0] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold166 (.A(\ChiselTop.wild.cpu.regs[4][4] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold167 (.A(\ChiselTop.wild.cpu.regs[6][24] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold168 (.A(\ChiselTop.wild.dmem.MEM[0][3] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold169 (.A(\ChiselTop.wild.cpu.regs[5][27] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold170 (.A(\ChiselTop.wild.cpu.regs[5][6] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold171 (.A(\ChiselTop.wild.cpu.regs[4][9] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold172 (.A(\ChiselTop.wild.cpu.regs[28][30] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold173 (.A(\ChiselTop.wild.cpu.regs[6][18] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold174 (.A(\ChiselTop.wild.cpu.regs[29][29] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold175 (.A(\ChiselTop.wild.cpu.regs[31][29] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold176 (.A(\ChiselTop.wild.cpu.regs[5][13] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold177 (.A(\ChiselTop.wild.cpu.regs[28][19] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold178 (.A(\ChiselTop.wild.cpu.regs[7][3] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold179 (.A(\ChiselTop.wild.cpu.regs[4][18] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold180 (.A(\ChiselTop.wild.cpu.regs[7][9] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold181 (.A(\ChiselTop.wild.cpu.regs[4][26] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold182 (.A(\ChiselTop.wild.cpu.regs[4][16] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold183 (.A(\ChiselTop.wild.cpu.regs[5][12] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold184 (.A(\ChiselTop.wild.cpu.regs[30][0] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold185 (.A(\ChiselTop.wild.cpu.regs[4][13] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold186 (.A(\ChiselTop.wild.cpu.regs[31][10] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold187 (.A(\ChiselTop.wild.cpu.regs[4][8] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold188 (.A(\ChiselTop.wild.cpu.regs[28][25] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold189 (.A(\ChiselTop.wild.cpu.regs[7][12] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold190 (.A(\ChiselTop.wild.cpu.regs[5][25] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold191 (.A(\ChiselTop.wild.cpu.regs[29][25] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold192 (.A(\ChiselTop.wild.cpu.regs[28][5] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold193 (.A(\ChiselTop.wild.cpu.regs[29][6] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold194 (.A(\ChiselTop.wild.cpu.regs[7][16] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold195 (.A(\ChiselTop.wild.cpu.regs[30][12] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold196 (.A(\ChiselTop.wild.cpu.regs[30][25] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold197 (.A(_00141_),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold198 (.A(_04654_),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold199 (.A(\ChiselTop.wild.cpu.regs[31][31] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold200 (.A(\ChiselTop.wild.cpu.regs[5][4] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold201 (.A(\ChiselTop.wild.cpu.regs[30][14] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold202 (.A(\ChiselTop.wild.cpu.regs[30][2] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold203 (.A(\ChiselTop.wild.cpu.regs[4][23] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold204 (.A(\ChiselTop.wild.cpu.regs[30][6] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold205 (.A(\ChiselTop.wild.cpu.regs[6][14] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold206 (.A(\ChiselTop.wild.cpu.regs[29][20] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold207 (.A(\ChiselTop.wild.cpu.regs[5][29] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold208 (.A(\ChiselTop.wild.cpu.regs[4][21] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold209 (.A(\ChiselTop.wild.cpu.regs[6][29] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold210 (.A(\ChiselTop.wild.cpu.regs[30][10] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold211 (.A(\ChiselTop.wild.cpu.regs[7][19] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold212 (.A(\ChiselTop.wild.cpu.regs[31][9] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold213 (.A(\ChiselTop.wild.cpu.pcReg[3] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold214 (.A(\ChiselTop.wild.cpu.regs[29][9] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold215 (.A(\ChiselTop.wild.cpu.regs[4][17] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold216 (.A(\ChiselTop.wild.cpu.regs[30][3] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold217 (.A(\ChiselTop.wild.tx.tx.cntReg[16] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold218 (.A(_03516_),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold219 (.A(_00153_),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold220 (.A(\ChiselTop.wild.cpu.regs[29][17] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold221 (.A(\ChiselTop.wild.cpu._T_12 ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold222 (.A(\ChiselTop.wild.cpu.regs[6][12] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold223 (.A(\ChiselTop.wild.cpu.regs[4][14] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold224 (.A(\ChiselTop.wild.cpu.regs[31][3] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold225 (.A(\ChiselTop.wild.cpu.regs[7][7] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold226 (.A(\ChiselTop.wild.cpu.regs[28][9] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold227 (.A(\ChiselTop.wild.cpu.regs[4][15] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold228 (.A(\ChiselTop.wild.cpu.regs[29][11] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold229 (.A(\ChiselTop.wild.cpu.regs[5][23] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold230 (.A(\ChiselTop.wild.cpu.regs[28][14] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold231 (.A(\ChiselTop.wild.cpu.regs[29][30] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold232 (.A(\ChiselTop.wild.rx.cntReg[13] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold233 (.A(_04647_),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold234 (.A(_00869_),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold235 (.A(\ChiselTop.wild.cpu.regs[28][27] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold236 (.A(\ChiselTop.wild.cpu.regs[7][2] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold237 (.A(\ChiselTop.wild.cpu.regs[31][30] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold238 (.A(\ChiselTop.wild.cpu.regs[6][19] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold239 (.A(\ChiselTop.wild.rx.io_channel_bits[0] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold240 (.A(_00846_),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold241 (.A(\ChiselTop.wild.cpu.regs[28][7] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold242 (.A(\ChiselTop.wild.cpu.regs[7][8] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold243 (.A(\ChiselTop.wild.cpu.regs[29][3] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold244 (.A(\ChiselTop.wild.cpu.regs[7][13] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold245 (.A(\ChiselTop.wild.cpu.regs[5][1] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold246 (.A(\ChiselTop.wild.cpu.regs[5][16] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold247 (.A(\ChiselTop.wild.cpu.regs[31][19] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold248 (.A(\ChiselTop.wild.cpu.regs[31][1] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold249 (.A(\ChiselTop.wild.cpu.regs[29][4] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold250 (.A(\ChiselTop.wild.cpu.regs[4][19] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold251 (.A(\ChiselTop.wild.cpu.regs[28][22] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold252 (.A(\ChiselTop.wild.cpu.regs[5][5] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold253 (.A(\ChiselTop.wild.tx.tx.cntReg[7] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold254 (.A(_03507_),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold255 (.A(_00146_),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold256 (.A(\ChiselTop.wild.cpu.regs[6][23] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold257 (.A(\ChiselTop.wild.cpu.regs[6][15] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold258 (.A(\ChiselTop.wild.cpu.regs[4][24] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold259 (.A(\ChiselTop.wild.cpu.regs[7][6] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold260 (.A(\ChiselTop.wild.cpu.regs[30][24] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold261 (.A(\ChiselTop.wild.cpu.regs[4][22] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold262 (.A(\ChiselTop.wild.cpu.regs[5][11] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold263 (.A(\ChiselTop.wild.cpu.regs[5][8] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold264 (.A(\ChiselTop.wild.cpu.regs[31][28] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold265 (.A(\ChiselTop.wild.cpu.regs[7][17] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold266 (.A(\ChiselTop.wild.cpu.regs[7][23] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold267 (.A(\ChiselTop.wild.cpu.regs[6][10] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold268 (.A(\ChiselTop.wild.cpu.regs[6][13] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold269 (.A(\ChiselTop.wild.cpu.regs[28][20] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold270 (.A(\ChiselTop.wild.cpu.regs[5][21] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold271 (.A(\ChiselTop.wild.cpu.regs[31][11] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold272 (.A(\ChiselTop.cntReg[24] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold273 (.A(_04284_),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold274 (.A(_00661_),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold275 (.A(\ChiselTop.wild.cpu.regs[5][2] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold276 (.A(\ChiselTop.wild.cpu.regs[31][26] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold277 (.A(\ChiselTop.wild.cpu.regs[31][27] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold278 (.A(\ChiselTop.wild.cpu.regs[31][18] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold279 (.A(\ChiselTop.wild.cpu.regs[6][5] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold280 (.A(\ChiselTop.wild.cpu.regs[6][25] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold281 (.A(\ChiselTop.wild.tx.tx.cntReg[10] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold282 (.A(_03508_),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold283 (.A(_00147_),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold284 (.A(\ChiselTop.wild.cpu.regs[28][13] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold285 (.A(\ChiselTop.wild.cpu.regs[30][13] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold286 (.A(\ChiselTop.wild.cpu.regs[7][18] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold287 (.A(\ChiselTop.wild.dmem.MEM[0][4] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold288 (.A(\ChiselTop.wild.cpu.regs[6][8] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold289 (.A(\ChiselTop.wild.cpu.regs[31][17] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold290 (.A(\ChiselTop.wild.cpu.regs[31][7] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold291 (.A(\ChiselTop.wild.cpu.regs[4][6] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold292 (.A(\ChiselTop.wild.cpu.regs[28][11] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold293 (.A(\ChiselTop.wild.cpu.regs[4][27] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold294 (.A(\ChiselTop.wild.cpu.regs[6][28] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold295 (.A(\ChiselTop.wild.dmem.MEM[0][5] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold296 (.A(\ChiselTop.wild.cpu.regs[5][31] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold297 (.A(\ChiselTop.wild.cpu.regs[31][2] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold298 (.A(\ChiselTop.wild.cpu.regs[30][26] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold299 (.A(\ChiselTop.wild.cpu.regs[7][22] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold300 (.A(_00123_),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold301 (.A(\ChiselTop.wild.cpu.regs[6][2] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold302 (.A(\ChiselTop.wild.cpu.regs[6][4] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold303 (.A(\ChiselTop.wild.cpu.regs[7][26] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold304 (.A(\ChiselTop.wild.cpu.regs[29][19] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold305 (.A(\ChiselTop.wild.cpu.regs[7][27] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold306 (.A(\ChiselTop.wild.cpu.regs[7][11] ),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold307 (.A(\ChiselTop.wild.cpu.regs[30][19] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold308 (.A(\ChiselTop.wild.cpu.regs[28][17] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold309 (.A(\ChiselTop.wild.cpu.regs[4][7] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold310 (.A(\ChiselTop.wild.cpu.regs[28][8] ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold311 (.A(\ChiselTop.wild.cpu.regs[7][1] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold312 (.A(\ChiselTop.wild.cpu.regs[31][6] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold313 (.A(\ChiselTop.wild.tx.tx.cntReg[13] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold314 (.A(_03512_),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold315 (.A(_00150_),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold316 (.A(\ChiselTop.wild.cpu.regs[30][15] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold317 (.A(\ChiselTop.wild.cpu.regs[4][10] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold318 (.A(\ChiselTop.wild.cpu.regs[31][13] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold319 (.A(\ChiselTop.wild.cpu.regs[31][20] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold320 (.A(\ChiselTop.wild.cpu.regs[5][28] ),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold321 (.A(\ChiselTop.wild.cpu.regs[30][27] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold322 (.A(\ChiselTop.wild.cpu.regs[29][8] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold323 (.A(\ChiselTop.wild.cpu.regs[30][7] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold324 (.A(\ChiselTop.wild.dmem.MEM[0][2] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold325 (.A(\ChiselTop.wild.cpu.regs[5][18] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold326 (.A(\ChiselTop.wild.cpu.regs[4][11] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold327 (.A(\ChiselTop.wild.cpu.regs[28][6] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold328 (.A(\ChiselTop.wild.cpu.regs[29][18] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold329 (.A(\ChiselTop.cntReg[27] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold330 (.A(_04289_),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold331 (.A(_00664_),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold332 (.A(\ChiselTop.wild.cpu.regs[30][22] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold333 (.A(\ChiselTop.wild.cpu.regs[30][11] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold334 (.A(\ChiselTop.wild.rx.cntReg[7] ),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold335 (.A(_04639_),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold336 (.A(_00863_),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold337 (.A(\ChiselTop.cntReg[6] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold338 (.A(_04249_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold339 (.A(_00643_),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold340 (.A(\ChiselTop.wild.cpu.regs[5][26] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold341 (.A(\ChiselTop.wild.cpu.regs[29][16] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold342 (.A(\ChiselTop.wild.cpu.regs[28][21] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold343 (.A(\ChiselTop.wild.cpu.regs[31][16] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold344 (.A(\ChiselTop.wild.cpu.regs[5][19] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold345 (.A(\ChiselTop.wild.cpu.regs[6][6] ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold346 (.A(\ChiselTop.wild.cpu.regs[29][23] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold347 (.A(\ChiselTop.wild.cpu.regs[31][15] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold348 (.A(\ChiselTop.wild.cpu.regs[5][9] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold349 (.A(\ChiselTop.wild.cpu.regs[31][12] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold350 (.A(\ChiselTop.wild.rx.cntReg[10] ),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold351 (.A(_04643_),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold352 (.A(_00866_),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold353 (.A(\ChiselTop.wild.cpu.regs[5][20] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold354 (.A(\ChiselTop.wild.cpu.regs[28][12] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold355 (.A(\ChiselTop.wild.cpu.regs[28][2] ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold356 (.A(\ChiselTop.wild.cpu.regs[30][5] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold357 (.A(\ChiselTop.wild.cpu.regs[4][12] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold358 (.A(\ChiselTop.wild.cpu.regs[6][31] ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold359 (.A(\ChiselTop.wild.cpu.regs[4][5] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold360 (.A(\ChiselTop.wild.rx._shiftReg_T_1[5] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold361 (.A(_00852_),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold362 (.A(\ChiselTop.wild.cpu.regs[6][11] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold363 (.A(\ChiselTop.wild.cpu.regs[31][14] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold364 (.A(\ChiselTop.wild.cpu.regs[1][31] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold365 (.A(\ChiselTop.wild.cpu.regs[2][25] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold366 (.A(\ChiselTop.wild.cpu.regs[28][3] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold367 (.A(\ChiselTop.wild.cpu.regs[4][31] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold368 (.A(\ChiselTop.wild.cpu.regs[30][20] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold369 (.A(\ChiselTop.wild.cpu.regs[30][29] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold370 (.A(\ChiselTop.wild.cpu.regs[30][23] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold371 (.A(\ChiselTop.wild.cpu.regs[3][15] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold372 (.A(\ChiselTop.wild.cpu.regs[2][8] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold373 (.A(\ChiselTop.wild.cpu.regs[7][31] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold374 (.A(\ChiselTop.wild.cpu.regs[5][15] ),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold375 (.A(\ChiselTop.wild.cpu.regs[4][28] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold376 (.A(\ChiselTop.wild.cpu.regs[6][21] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold377 (.A(\ChiselTop.wild.tx.tx.bitsReg[2] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold378 (.A(_04581_),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold379 (.A(_00839_),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold380 (.A(\ChiselTop.wild.cpu.regs[6][16] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold381 (.A(\ChiselTop.wild.cpu.regs[30][30] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold382 (.A(\ChiselTop.wild.cpu.regs[1][6] ),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold383 (.A(\ChiselTop.wild.cpu.regs[30][18] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold384 (.A(\ChiselTop.wild.cpu.regs[1][21] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold385 (.A(\ChiselTop.wild.cpu.regs[4][25] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold386 (.A(\ChiselTop.wild.cpu.regs[7][15] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold387 (.A(\ChiselTop.wild.cpu.regs[1][1] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold388 (.A(\ChiselTop.wild.cpu.regs[30][1] ),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold389 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[0] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold390 (.A(\ChiselTop.wild.cpu.regs[1][0] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold391 (.A(\ChiselTop.wild.cpu.regs[29][26] ),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold392 (.A(\ChiselTop.wild.cpu.regs[31][8] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold393 (.A(\ChiselTop.wild.cpu.regs[30][28] ),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold394 (.A(\ChiselTop.wild.cpu.regs[7][21] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold395 (.A(\ChiselTop.wild.rx._shiftReg_T_1[6] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold396 (.A(\ChiselTop.wild.cpu.regs[31][21] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold397 (.A(\ChiselTop.wild.cpu.regs[7][5] ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold398 (.A(\ChiselTop.wild.cpu.regs[1][22] ),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold399 (.A(\ChiselTop.wild.cpu.regs[31][5] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold400 (.A(\ChiselTop.wild.rx.cntReg[4] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold401 (.A(_04635_),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold402 (.A(_00860_),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold403 (.A(\ChiselTop.wild.cpu.regs[30][31] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold404 (.A(\ChiselTop.wild.cpu.regs[2][22] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold405 (.A(\ChiselTop.wild.cpu.regs[6][9] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold406 (.A(\ChiselTop.wild.cpu.regs[7][10] ),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold407 (.A(\ChiselTop.wild.cpu.regs[29][28] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold408 (.A(\ChiselTop.wild.cpu.regs[28][29] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold409 (.A(\ChiselTop.wild.cpu.regs[6][26] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold410 (.A(\ChiselTop.wild.cpu.regs[1][18] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold411 (.A(\ChiselTop.wild.cpu.regs[28][26] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold412 (.A(\ChiselTop.wild.cpu.regs[4][30] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold413 (.A(\ChiselTop.wild.cpu.regs[2][1] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold414 (.A(\ChiselTop.wild.cpu.regs[6][7] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold415 (.A(\ChiselTop.wild.cpu.regs[4][20] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold416 (.A(\ChiselTop.wild.cpu.regs[2][29] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold417 (.A(\ChiselTop.wild.dmem.MEM[0][6] ),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold418 (.A(\ChiselTop.wild.cpu.regs[1][19] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold419 (.A(\ChiselTop.wild.cpu.regs[28][16] ),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold420 (.A(\ChiselTop.wild.cpu.regs[5][3] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold421 (.A(\ChiselTop.wild.cpu.regs[6][17] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold422 (.A(\ChiselTop.wild.cpu.regs[1][12] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold423 (.A(\ChiselTop.wild.cpu.regs[3][26] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold424 (.A(\ChiselTop.wild.dmem.MEM[0][7] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold425 (.A(\ChiselTop.wild.cpu.regs[7][30] ),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold426 (.A(\ChiselTop.wild.cpu.regs[3][19] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold427 (.A(\ChiselTop.wild.cpu.regs[30][8] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold428 (.A(\ChiselTop.wild.cpu.regs[1][7] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold429 (.A(\ChiselTop.wild.cpu.regs[2][28] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold430 (.A(\ChiselTop.wild.cpu.regs[30][17] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold431 (.A(\ChiselTop.wild.cpu.regs[5][7] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold432 (.A(\ChiselTop.wild.cpu.regs[30][4] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold433 (.A(\ChiselTop.wild.cpu.regs[2][20] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold434 (.A(\ChiselTop.wild.cpu.regs[6][0] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold435 (.A(\ChiselTop.wild.cpu.pcReg[2] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold436 (.A(\ChiselTop.wild.cpu.regs[6][27] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold437 (.A(\ChiselTop.wild.cpu.regs[2][18] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold438 (.A(\ChiselTop.wild.cpu.regs[1][14] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold439 (.A(\ChiselTop.wild.cpu.regs[28][24] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold440 (.A(\ChiselTop.wild.cpu.regs[3][27] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold441 (.A(\ChiselTop.wild.cpu.regs[2][31] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold442 (.A(\ChiselTop.wild.cpu.regs[1][25] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold443 (.A(\ChiselTop.wild.cpu.regs[3][30] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold444 (.A(\ChiselTop.wild.cpu.regs[7][24] ),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold445 (.A(\ChiselTop.wild.cpu.regs[3][22] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold446 (.A(\ChiselTop.wild.cpu.regs[2][24] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold447 (.A(\ChiselTop.wild.cpu.regs[2][16] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold448 (.A(\ChiselTop.wild.cpu.regs[1][30] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold449 (.A(\ChiselTop.wild.cpu.regs[1][13] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold450 (.A(\ChiselTop.wild.cpu.regs[3][14] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold451 (.A(\ChiselTop.wild.rx._shiftReg_T_1[1] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold452 (.A(_00848_),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold453 (.A(\ChiselTop.wild.cpu.regs[6][22] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold454 (.A(\ChiselTop.wild.rx._shiftReg_T_1[0] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold455 (.A(\ChiselTop.wild.cpu.regs[2][13] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold456 (.A(\ChiselTop.wild.cpu.regs[3][7] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold457 (.A(\ChiselTop.wild.cpu.regs[3][9] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold458 (.A(\ChiselTop.wild.cpu.regs[30][21] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold459 (.A(\ChiselTop.wild.cpu.regs[6][20] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold460 (.A(\ChiselTop.wild.cpu.regs[3][3] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold461 (.A(\ChiselTop.wild.cpu.regs[2][30] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold462 (.A(\ChiselTop.wild.rx.bitsReg[3] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold463 (.A(_04615_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold464 (.A(\ChiselTop.wild.cpu.regs[2][21] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold465 (.A(\ChiselTop.wild.cpu.regs[1][15] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold466 (.A(\ChiselTop.wild.cpu.regs[3][31] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold467 (.A(\ChiselTop.wild.cpu.regs[29][15] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold468 (.A(\ChiselTop.wild.cpu.regs[2][27] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold469 (.A(\ChiselTop.wild.cpu.regs[3][28] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold470 (.A(\ChiselTop.wild.cpu.regs[3][21] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold471 (.A(\ChiselTop.wild.cpu.regs[3][4] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold472 (.A(\ChiselTop.wild.cpu.regs[28][15] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold473 (.A(\ChiselTop.wild.cpu.regs[2][14] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold474 (.A(\ChiselTop.wild.cpu.regs[2][12] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold475 (.A(\ChiselTop.wild.cpu.regs[2][5] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold476 (.A(\ChiselTop.wild.cpu.regs[3][23] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold477 (.A(\ChiselTop.wild.cpu.regs[4][29] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold478 (.A(\ChiselTop.cntReg[30] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold479 (.A(_04294_),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold480 (.A(_00667_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold481 (.A(\ChiselTop.wild.cpu.regs[2][0] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold482 (.A(\ChiselTop.wild.rx.cntReg[17] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold483 (.A(_04652_),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold484 (.A(_00873_),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold485 (.A(\ChiselTop.wild.cpu.regs[3][13] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold486 (.A(\ChiselTop.wild.cpu.regs[29][13] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold487 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[15] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold488 (.A(\ChiselTop.wild.cpu.regs[2][10] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold489 (.A(\ChiselTop.wild.cpu.regs[2][6] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold490 (.A(\ChiselTop.wild.cpu.regs[3][5] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold491 (.A(\ChiselTop.wild.cpu.regs[3][20] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold492 (.A(\ChiselTop.wild.cpu.regs[4][1] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold493 (.A(\ChiselTop.wild.cpu.regs[1][10] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold494 (.A(\ChiselTop.wild.cpu.regs[1][9] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold495 (.A(\ChiselTop.wild.cpu.regs[2][15] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold496 (.A(\ChiselTop.wild.cpu.regs[3][17] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold497 (.A(\ChiselTop.wild.cpu.regs[1][3] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold498 (.A(\ChiselTop.wild.cpu.regs[3][25] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold499 (.A(\ChiselTop.wild.cpu.regs[1][20] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold500 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[1] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold501 (.A(\ChiselTop.wild.cpu.regs[5][14] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold502 (.A(\ChiselTop.wild.cpu.regs[2][17] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold503 (.A(\ChiselTop.wild.cpu.regs[1][27] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold504 (.A(\ChiselTop.wild.cpu.regs[1][24] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold505 (.A(\ChiselTop.wild.cpu.regs[1][29] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold506 (.A(\ChiselTop.wild.tx.tx.cntReg[5] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold507 (.A(_04130_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold508 (.A(\ChiselTop.wild.cpu.regs[2][23] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold509 (.A(\ChiselTop.wild.cpu.regs[1][11] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold510 (.A(\ChiselTop.wild.cpu.regs[3][6] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold511 (.A(\ChiselTop.wild.cpu.regs[2][2] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold512 (.A(\ChiselTop.wild.dmem.MEM[0][1] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold513 (.A(\ChiselTop.wild.cpu.regs[3][11] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold514 (.A(\ChiselTop.wild.cpu.regs[3][10] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold515 (.A(\ChiselTop.wild.cpu.regs[2][3] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold516 (.A(\ChiselTop.wild.cpu.regs[1][4] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold517 (.A(\ChiselTop.wild.tx.tx.cntReg[3] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold518 (.A(_03505_),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold519 (.A(\ChiselTop.wild.cpu.regs[3][8] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold520 (.A(\ChiselTop.wild.cpu.regs[1][23] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold521 (.A(\ChiselTop.wild.dmem.MEM_2[0][3] ),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold522 (.A(\ChiselTop.wild.cpu.regs[1][5] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold523 (.A(\ChiselTop.cntReg[4] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold524 (.A(_04247_),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold525 (.A(\ChiselTop.wild.cpu.regs[2][7] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold526 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[17] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold527 (.A(\ChiselTop.wild.cpu.regs[2][19] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold528 (.A(\ChiselTop.wild.dmem.MEM[0][0] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold529 (.A(\ChiselTop.wild.cpu.regs[29][22] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold530 (.A(\ChiselTop.wild.tx.tx.cntReg[4] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold531 (.A(_03506_),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold532 (.A(\ChiselTop.wild.cpu.regs[1][8] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold533 (.A(\ChiselTop.wild.rx.bitsReg[2] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold534 (.A(_04600_),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold535 (.A(\ChiselTop.cntReg[11] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold536 (.A(_04259_),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold537 (.A(\ChiselTop.cntReg[12] ),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold538 (.A(\ChiselTop.wild.cpu.regs[1][17] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold539 (.A(\ChiselTop.cntReg[10] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold540 (.A(_04257_),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold541 (.A(\ChiselTop.wild.cpu.regs[2][11] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold542 (.A(\ChiselTop.wild.tx.tx.cntReg[6] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold543 (.A(\ChiselTop.wild.rx.cntReg[15] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold544 (.A(_04650_),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold545 (.A(\ChiselTop.wild.cpu.regs[2][9] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold546 (.A(\ChiselTop.wild.cpu.regs[3][29] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold547 (.A(\ChiselTop.cntReg[18] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold548 (.A(_04273_),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold549 (.A(\ChiselTop.wild.rx.cntReg[3] ),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold550 (.A(_04634_),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold551 (.A(\ChiselTop.wild.cpu.regs[2][26] ),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold552 (.A(\ChiselTop.wild.cpu.regs[3][1] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold553 (.A(\ChiselTop.wild.cpu.regs[2][4] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold554 (.A(\ChiselTop.wild.cpu.regs[1][16] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold555 (.A(\ChiselTop.wild.cpu.regs[3][2] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold556 (.A(\ChiselTop.wild.cpu.regs[1][28] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold557 (.A(\ChiselTop.wild.cpu.regs[3][0] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold558 (.A(\ChiselTop.wild.rx._shiftReg_T_1[2] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold559 (.A(_00849_),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold560 (.A(\ChiselTop.wild.cpu.regs[1][2] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold561 (.A(\ChiselTop.wild.cpu.regs[3][12] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold562 (.A(\ChiselTop.wild.rx._shiftReg_T_1[4] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold563 (.A(\ChiselTop.wild.rx.bitsReg[1] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold564 (.A(_00843_),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold565 (.A(\ChiselTop.cntReg[15] ),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold566 (.A(_04267_),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold567 (.A(\ChiselTop.wild.dmem.MEM_3[0][3] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold568 (.A(\ChiselTop.cntReg[17] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold569 (.A(_04271_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold570 (.A(\ChiselTop.cntReg[19] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold571 (.A(\ChiselTop.wild.cpu.regs[1][26] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold572 (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[11] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold573 (.A(_00782_),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold574 (.A(\ChiselTop.wild.dmem.MEM_2[0][0] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold575 (.A(\ChiselTop.cntReg[2] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold576 (.A(_04243_),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold577 (.A(_00639_),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold578 (.A(\ChiselTop.wild.cpu.regs[3][16] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold579 (.A(\ChiselTop.cntReg[13] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold580 (.A(\ChiselTop.wild.dmem.MEM_2[0][2] ),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold581 (.A(\ChiselTop.wild.rx.cntReg[8] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold582 (.A(_04640_),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold583 (.A(_00864_),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold584 (.A(\ChiselTop.cntReg[22] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold585 (.A(_04281_),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold586 (.A(\ChiselTop.wild.rx.cntReg[16] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold587 (.A(_04651_),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold588 (.A(\ChiselTop.wild.rx._shiftReg_T_1[3] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold589 (.A(\ChiselTop.wild.cpu.regs[3][18] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold590 (.A(\ChiselTop.wild.cpu.pcReg[7] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold591 (.A(\ChiselTop.cntReg[21] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold592 (.A(_04279_),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold593 (.A(_00658_),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold594 (.A(\ChiselTop.cntReg[25] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold595 (.A(_04286_),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold596 (.A(\ChiselTop.cntReg[14] ),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold597 (.A(\ChiselTop.cntReg[16] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold598 (.A(\ChiselTop.wild.dmem.MEM_1[0][0] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold599 (.A(\ChiselTop.wild.dmem.MEM_2[0][1] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold600 (.A(\ChiselTop.cntReg[31] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold601 (.A(_04296_),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold602 (.A(\ChiselTop.wild.tx.tx.bitsReg[1] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold603 (.A(_04579_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold604 (.A(_00838_),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold605 (.A(\ChiselTop.cntReg[20] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold606 (.A(\ChiselTop.wild.cpu.regs[3][24] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold607 (.A(\ChiselTop.wild.dmem.MEM_3[0][0] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold608 (.A(\ChiselTop.cntReg[7] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold609 (.A(_04251_),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold610 (.A(\ChiselTop.cntReg[9] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold611 (.A(_04255_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold612 (.A(\ChiselTop.wild.dmem.MEM_3[0][4] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold613 (.A(\ChiselTop.wild.dmem.MEM_3[0][2] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold614 (.A(\ChiselTop.wild.dmem.MEM_1[0][1] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold615 (.A(\ChiselTop.wild.dmem.MEM_3[0][7] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold616 (.A(\ChiselTop.wild.rx.bitsReg[0] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold617 (.A(\ChiselTop.cntReg[3] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold618 (.A(\ChiselTop.wild.dmem.MEM_3[0][5] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold619 (.A(\ChiselTop.cntReg[8] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold620 (.A(\ChiselTop.wild.dmem.MEM_3[0][1] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold621 (.A(\ChiselTop.wild.dmem.MEM_2[0][4] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold622 (.A(\ChiselTop.cntReg[23] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold623 (.A(\ChiselTop.wild.tx.tx.bitsReg[0] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold624 (.A(_04577_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold625 (.A(\ChiselTop.wild.cpu.decExReg_rd[2] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold626 (.A(\ChiselTop.wild.dmem.MEM_2[0][5] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold627 (.A(\ChiselTop.cntReg[26] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold628 (.A(\ChiselTop.wild.cpu._GEN_176[10] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold629 (.A(_03526_),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold630 (.A(_00193_),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold631 (.A(\ChiselTop.cntReg[28] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold632 (.A(\ChiselTop.cntReg[5] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold633 (.A(\ChiselTop.wild.cpu._GEN_176[2] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold634 (.A(\ChiselTop.wild.dmem.MEM_2[0][7] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold635 (.A(\ChiselTop.cntReg[0] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold636 (.A(_04237_),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold637 (.A(_00638_),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold638 (.A(\ChiselTop.cntReg[29] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold639 (.A(\ChiselTop.wild.tx.tx.cntReg[1] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold640 (.A(\ChiselTop.wild.dmem.MEM_1[0][6] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold641 (.A(\ChiselTop.wild.rx.cntReg[11] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold642 (.A(_04644_),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold643 (.A(\ChiselTop.wild.tx.tx.cntReg[14] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold644 (.A(_03513_),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold645 (.A(\ChiselTop.wild.cpu._T_12 ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold646 (.A(\ChiselTop.wild.dmem.MEM_1[0][3] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold647 (.A(\ChiselTop.wild.cpu.decOut_opcode[2] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold648 (.A(_00525_),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold649 (.A(\ChiselTop.wild.dmem.MEM_2[0][6] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold650 (.A(\ChiselTop.wild.cpu.decExReg_rd[3] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold651 (.A(\ChiselTop.wild.cpu.pcReg[28] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold652 (.A(_00799_),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold653 (.A(_00134_),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold654 (.A(\ChiselTop.wild.tx.tx.cntReg[8] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold655 (.A(\ChiselTop.wild.rx.cntReg[19] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold656 (.A(\ChiselTop.wild.tx.tx.cntReg[17] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold657 (.A(_03517_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold658 (.A(\ChiselTop.wild.dmem.MEM_3[0][6] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold659 (.A(\ChiselTop.wild.tx.tx.cntReg[11] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold660 (.A(_03509_),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold661 (.A(\ChiselTop.wild.tx.tx.cntReg[15] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold662 (.A(_03498_),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold663 (.A(\ChiselTop.wild.cpu.decExReg_valid ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold664 (.A(\ChiselTop.wild.rx.cntReg[9] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold665 (.A(\ChiselTop.wild.dmem.MEM_1[0][4] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold666 (.A(\ChiselTop.wild.dmem.MEM_1[0][7] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold667 (.A(\ChiselTop.wild.dmem.MEM_1[0][2] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold668 (.A(\ChiselTop.wild.dmem.MEM_1[0][5] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold669 (.A(_00004_),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold670 (.A(\ChiselTop.wild.tx.tx.cntReg[2] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold671 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_1[0] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold672 (.A(\ChiselTop.wild.cpu.decOut_opcode[4] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold673 (.A(_00463_),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold674 (.A(\ChiselTop.wild.cpu.decOut_opcode[5] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold675 (.A(_00518_),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold676 (.A(\ChiselTop.wild.rx.cntReg[2] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold677 (.A(_04585_),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold678 (.A(_04633_),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold679 (.A(\ChiselTop.wild.tx.tx.cntReg[9] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold680 (.A(\ChiselTop.wild.rx.cntReg[12] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold681 (.A(\ChiselTop.wild.tx.tx.cntReg[18] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold682 (.A(\ChiselTop.wild.rx.cntReg[0] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold683 (.A(_04628_),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold684 (.A(_00857_),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold685 (.A(\ChiselTop.wild.tx.tx.cntReg[12] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold686 (.A(_03511_),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold687 (.A(\ChiselTop.wild.rx.bitsReg[0] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold688 (.A(_04602_),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold689 (.A(\ChiselTop.wild.rx.cntReg[5] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold690 (.A(_04636_),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold691 (.A(\ChiselTop.wild.cpu.pcReg[10] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold692 (.A(\ChiselTop.wild.cpu.decExReg_rd[1] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold693 (.A(_00119_),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold694 (.A(\ChiselTop.wild.cpu.decExReg_decOut_rfWrite ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold695 (.A(\ChiselTop.wild.cpu.decExReg_func3[0] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold696 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_30[13] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold697 (.A(\ChiselTop.wild.cpu._decOut_decOut_imm_imm_T_15[4] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold698 (.A(\ChiselTop.wild.cpu._GEN_176[1] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold699 (.A(_00124_),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold700 (.A(\ChiselTop.wild.cpu._GEN_176[20] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold701 (.A(\ChiselTop.wild.rx.cntReg[6] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold702 (.A(_04638_),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold703 (.A(\ChiselTop.wild.cpu._GEN_176[5] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold704 (.A(\ChiselTop.wild.cpu.decExReg_rd[0] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold705 (.A(\ChiselTop.wild.cpu.decExReg_decOut_imm[11] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold706 (.A(\ChiselTop.wild.cpu.pcReg[3] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold707 (.A(_03470_),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold708 (.A(_00136_),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold709 (.A(\ChiselTop.wild.cpu.decOut_opcode[2] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold710 (.A(\ChiselTop.wild.cpu.pcReg[2] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold711 (.A(_00196_),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold712 (.A(\ChiselTop.wild.cpu.regs_rs1Val_MPORT_addr[2] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold713 (.A(_00121_),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold714 (.A(_00001_),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold715 (.A(\ChiselTop.wild.cpu.regs[5][8] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold716 (.A(_00112_),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold717 (.A(\ChiselTop.wild.cpu._wbData_T_1[1] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold718 (.A(\ChiselTop.wild.cpu.regs[31][14] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold719 (.A(\ChiselTop.wild.tx.buf_.io_out_valid ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold720 (.A(\ChiselTop.wild.cpu.regs[29][12] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold721 (.A(\ChiselTop.wild.cpu.pcReg[3] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold722 (.A(_00116_),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold723 (.A(_00115_),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold724 (.A(\ChiselTop.wild.cpu.regs[28][9] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold725 (.A(\ChiselTop.wild.cpu.regs[29][10] ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold726 (.A(_03827_),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold727 (.A(\ChiselTop.wild.cpu.regs[4][19] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold728 (.A(\ChiselTop.wild.cpu.regs[4][18] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold729 (.A(\ChiselTop.wild.cpu.regs[28][28] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold730 (.A(_04192_),
    .X(net1555));
 sg13g2_antennanp ANTENNA_1 (.A(_00192_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(rst_n));
 sg13g2_antennanp ANTENNA_4 (.A(rst_n));
 sg13g2_antennanp ANTENNA_5 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_6 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_7 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_8 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_9 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_10 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_11 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_12 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_13 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_14 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_15 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_16 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_17 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_18 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_19 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_20 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_21 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_22 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_23 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_24 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_25 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_26 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_27 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_28 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_29 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_30 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_31 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_32 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_33 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_34 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_35 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_36 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_37 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_38 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_39 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_40 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_41 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_42 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_43 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_44 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_45 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_46 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_47 (.A(clk));
 sg13g2_antennanp ANTENNA_48 (.A(clk));
 sg13g2_antennanp ANTENNA_49 (.A(rst_n));
 sg13g2_antennanp ANTENNA_50 (.A(rst_n));
 sg13g2_antennanp ANTENNA_51 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_52 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_53 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_54 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_55 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_56 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_57 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_58 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_59 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_60 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_61 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_62 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_63 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_64 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_65 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_66 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_67 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_68 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_69 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_70 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_71 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_72 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_73 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_74 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_75 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_76 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_77 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_78 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_79 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_80 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_81 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_82 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_83 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_84 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_85 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_86 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_87 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_88 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_89 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_90 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_91 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_92 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_93 (.A(clk));
 sg13g2_antennanp ANTENNA_94 (.A(clk));
 sg13g2_antennanp ANTENNA_95 (.A(rst_n));
 sg13g2_antennanp ANTENNA_96 (.A(rst_n));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_fill_2 FILLER_0_343 ();
 sg13g2_fill_1 FILLER_0_371 ();
 sg13g2_fill_2 FILLER_0_398 ();
 sg13g2_fill_2 FILLER_0_409 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_1 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_472 ();
 sg13g2_fill_2 FILLER_0_478 ();
 sg13g2_fill_1 FILLER_0_480 ();
 sg13g2_decap_8 FILLER_0_485 ();
 sg13g2_decap_8 FILLER_0_492 ();
 sg13g2_decap_8 FILLER_0_499 ();
 sg13g2_decap_4 FILLER_0_506 ();
 sg13g2_fill_2 FILLER_0_510 ();
 sg13g2_fill_2 FILLER_0_546 ();
 sg13g2_fill_2 FILLER_0_557 ();
 sg13g2_fill_1 FILLER_0_569 ();
 sg13g2_decap_4 FILLER_0_593 ();
 sg13g2_decap_8 FILLER_0_610 ();
 sg13g2_decap_8 FILLER_0_617 ();
 sg13g2_decap_8 FILLER_0_624 ();
 sg13g2_decap_8 FILLER_0_631 ();
 sg13g2_decap_8 FILLER_0_638 ();
 sg13g2_decap_8 FILLER_0_645 ();
 sg13g2_decap_8 FILLER_0_652 ();
 sg13g2_decap_8 FILLER_0_659 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_8 FILLER_0_673 ();
 sg13g2_decap_4 FILLER_0_680 ();
 sg13g2_fill_1 FILLER_0_684 ();
 sg13g2_fill_2 FILLER_0_713 ();
 sg13g2_fill_2 FILLER_0_744 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_4 FILLER_0_763 ();
 sg13g2_fill_1 FILLER_0_767 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_fill_2 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_fill_1 FILLER_0_808 ();
 sg13g2_decap_4 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_827 ();
 sg13g2_fill_2 FILLER_0_834 ();
 sg13g2_fill_1 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_842 ();
 sg13g2_decap_4 FILLER_0_849 ();
 sg13g2_fill_1 FILLER_0_853 ();
 sg13g2_decap_8 FILLER_0_858 ();
 sg13g2_decap_4 FILLER_0_865 ();
 sg13g2_fill_2 FILLER_0_873 ();
 sg13g2_decap_8 FILLER_0_878 ();
 sg13g2_decap_8 FILLER_0_885 ();
 sg13g2_decap_8 FILLER_0_892 ();
 sg13g2_decap_8 FILLER_0_899 ();
 sg13g2_decap_8 FILLER_0_906 ();
 sg13g2_decap_8 FILLER_0_913 ();
 sg13g2_decap_8 FILLER_0_920 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_8 FILLER_0_1025 ();
 sg13g2_decap_8 FILLER_0_1032 ();
 sg13g2_decap_8 FILLER_0_1039 ();
 sg13g2_decap_8 FILLER_0_1046 ();
 sg13g2_decap_8 FILLER_0_1053 ();
 sg13g2_decap_8 FILLER_0_1060 ();
 sg13g2_decap_8 FILLER_0_1067 ();
 sg13g2_decap_8 FILLER_0_1074 ();
 sg13g2_decap_8 FILLER_0_1081 ();
 sg13g2_decap_8 FILLER_0_1088 ();
 sg13g2_decap_8 FILLER_0_1095 ();
 sg13g2_decap_8 FILLER_0_1102 ();
 sg13g2_decap_8 FILLER_0_1109 ();
 sg13g2_decap_8 FILLER_0_1116 ();
 sg13g2_decap_8 FILLER_0_1123 ();
 sg13g2_decap_8 FILLER_0_1130 ();
 sg13g2_decap_8 FILLER_0_1137 ();
 sg13g2_decap_8 FILLER_0_1144 ();
 sg13g2_decap_8 FILLER_0_1151 ();
 sg13g2_decap_8 FILLER_0_1158 ();
 sg13g2_decap_8 FILLER_0_1165 ();
 sg13g2_decap_8 FILLER_0_1172 ();
 sg13g2_decap_8 FILLER_0_1179 ();
 sg13g2_decap_8 FILLER_0_1186 ();
 sg13g2_decap_8 FILLER_0_1193 ();
 sg13g2_decap_8 FILLER_0_1200 ();
 sg13g2_decap_8 FILLER_0_1207 ();
 sg13g2_decap_8 FILLER_0_1214 ();
 sg13g2_decap_8 FILLER_0_1221 ();
 sg13g2_decap_8 FILLER_0_1228 ();
 sg13g2_decap_8 FILLER_0_1235 ();
 sg13g2_decap_8 FILLER_0_1242 ();
 sg13g2_decap_8 FILLER_0_1249 ();
 sg13g2_decap_8 FILLER_0_1256 ();
 sg13g2_decap_8 FILLER_0_1263 ();
 sg13g2_decap_8 FILLER_0_1270 ();
 sg13g2_decap_8 FILLER_0_1277 ();
 sg13g2_decap_8 FILLER_0_1284 ();
 sg13g2_decap_8 FILLER_0_1291 ();
 sg13g2_decap_8 FILLER_0_1298 ();
 sg13g2_decap_8 FILLER_0_1305 ();
 sg13g2_fill_2 FILLER_0_1312 ();
 sg13g2_fill_1 FILLER_0_1314 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_fill_1 FILLER_1_336 ();
 sg13g2_fill_1 FILLER_1_441 ();
 sg13g2_fill_2 FILLER_1_452 ();
 sg13g2_fill_2 FILLER_1_515 ();
 sg13g2_fill_1 FILLER_1_526 ();
 sg13g2_decap_8 FILLER_1_618 ();
 sg13g2_decap_8 FILLER_1_625 ();
 sg13g2_decap_8 FILLER_1_632 ();
 sg13g2_decap_8 FILLER_1_639 ();
 sg13g2_decap_8 FILLER_1_646 ();
 sg13g2_decap_8 FILLER_1_653 ();
 sg13g2_fill_1 FILLER_1_660 ();
 sg13g2_decap_4 FILLER_1_703 ();
 sg13g2_decap_4 FILLER_1_728 ();
 sg13g2_fill_1 FILLER_1_732 ();
 sg13g2_decap_4 FILLER_1_742 ();
 sg13g2_fill_1 FILLER_1_761 ();
 sg13g2_fill_2 FILLER_1_805 ();
 sg13g2_fill_1 FILLER_1_807 ();
 sg13g2_fill_2 FILLER_1_825 ();
 sg13g2_fill_1 FILLER_1_827 ();
 sg13g2_fill_1 FILLER_1_838 ();
 sg13g2_decap_8 FILLER_1_886 ();
 sg13g2_decap_8 FILLER_1_893 ();
 sg13g2_decap_8 FILLER_1_900 ();
 sg13g2_decap_8 FILLER_1_907 ();
 sg13g2_decap_8 FILLER_1_914 ();
 sg13g2_decap_8 FILLER_1_921 ();
 sg13g2_decap_8 FILLER_1_928 ();
 sg13g2_decap_8 FILLER_1_935 ();
 sg13g2_decap_8 FILLER_1_942 ();
 sg13g2_decap_8 FILLER_1_949 ();
 sg13g2_decap_8 FILLER_1_956 ();
 sg13g2_decap_8 FILLER_1_963 ();
 sg13g2_decap_8 FILLER_1_970 ();
 sg13g2_decap_8 FILLER_1_977 ();
 sg13g2_decap_8 FILLER_1_984 ();
 sg13g2_decap_8 FILLER_1_991 ();
 sg13g2_decap_8 FILLER_1_998 ();
 sg13g2_decap_8 FILLER_1_1005 ();
 sg13g2_decap_8 FILLER_1_1012 ();
 sg13g2_decap_8 FILLER_1_1019 ();
 sg13g2_decap_8 FILLER_1_1026 ();
 sg13g2_decap_8 FILLER_1_1033 ();
 sg13g2_decap_8 FILLER_1_1040 ();
 sg13g2_decap_8 FILLER_1_1047 ();
 sg13g2_decap_8 FILLER_1_1054 ();
 sg13g2_decap_8 FILLER_1_1061 ();
 sg13g2_decap_8 FILLER_1_1068 ();
 sg13g2_decap_8 FILLER_1_1075 ();
 sg13g2_decap_8 FILLER_1_1082 ();
 sg13g2_decap_8 FILLER_1_1089 ();
 sg13g2_decap_8 FILLER_1_1096 ();
 sg13g2_decap_8 FILLER_1_1103 ();
 sg13g2_decap_8 FILLER_1_1110 ();
 sg13g2_decap_8 FILLER_1_1117 ();
 sg13g2_decap_8 FILLER_1_1124 ();
 sg13g2_decap_8 FILLER_1_1131 ();
 sg13g2_decap_8 FILLER_1_1138 ();
 sg13g2_decap_8 FILLER_1_1145 ();
 sg13g2_decap_8 FILLER_1_1152 ();
 sg13g2_decap_8 FILLER_1_1159 ();
 sg13g2_decap_8 FILLER_1_1166 ();
 sg13g2_decap_8 FILLER_1_1173 ();
 sg13g2_decap_8 FILLER_1_1180 ();
 sg13g2_decap_8 FILLER_1_1187 ();
 sg13g2_decap_8 FILLER_1_1194 ();
 sg13g2_decap_8 FILLER_1_1201 ();
 sg13g2_decap_8 FILLER_1_1208 ();
 sg13g2_decap_8 FILLER_1_1215 ();
 sg13g2_decap_8 FILLER_1_1222 ();
 sg13g2_decap_8 FILLER_1_1229 ();
 sg13g2_decap_8 FILLER_1_1236 ();
 sg13g2_decap_8 FILLER_1_1243 ();
 sg13g2_decap_8 FILLER_1_1250 ();
 sg13g2_decap_8 FILLER_1_1257 ();
 sg13g2_decap_8 FILLER_1_1264 ();
 sg13g2_decap_8 FILLER_1_1271 ();
 sg13g2_decap_8 FILLER_1_1278 ();
 sg13g2_decap_8 FILLER_1_1285 ();
 sg13g2_decap_8 FILLER_1_1292 ();
 sg13g2_decap_8 FILLER_1_1299 ();
 sg13g2_decap_8 FILLER_1_1306 ();
 sg13g2_fill_2 FILLER_1_1313 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_4 FILLER_2_329 ();
 sg13g2_fill_1 FILLER_2_333 ();
 sg13g2_fill_2 FILLER_2_374 ();
 sg13g2_fill_1 FILLER_2_376 ();
 sg13g2_fill_2 FILLER_2_390 ();
 sg13g2_fill_1 FILLER_2_392 ();
 sg13g2_fill_2 FILLER_2_397 ();
 sg13g2_fill_1 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_478 ();
 sg13g2_fill_2 FILLER_2_493 ();
 sg13g2_fill_1 FILLER_2_500 ();
 sg13g2_fill_1 FILLER_2_515 ();
 sg13g2_fill_1 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_625 ();
 sg13g2_fill_1 FILLER_2_632 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_4 FILLER_2_651 ();
 sg13g2_fill_2 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_678 ();
 sg13g2_decap_8 FILLER_2_685 ();
 sg13g2_fill_1 FILLER_2_692 ();
 sg13g2_fill_2 FILLER_2_703 ();
 sg13g2_fill_1 FILLER_2_705 ();
 sg13g2_decap_8 FILLER_2_726 ();
 sg13g2_decap_4 FILLER_2_738 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_4 FILLER_2_779 ();
 sg13g2_fill_1 FILLER_2_783 ();
 sg13g2_fill_1 FILLER_2_795 ();
 sg13g2_decap_4 FILLER_2_811 ();
 sg13g2_fill_2 FILLER_2_815 ();
 sg13g2_fill_2 FILLER_2_822 ();
 sg13g2_fill_2 FILLER_2_838 ();
 sg13g2_fill_2 FILLER_2_845 ();
 sg13g2_fill_1 FILLER_2_847 ();
 sg13g2_fill_2 FILLER_2_855 ();
 sg13g2_fill_1 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_2_894 ();
 sg13g2_decap_8 FILLER_2_901 ();
 sg13g2_decap_8 FILLER_2_908 ();
 sg13g2_decap_8 FILLER_2_915 ();
 sg13g2_decap_8 FILLER_2_922 ();
 sg13g2_decap_8 FILLER_2_929 ();
 sg13g2_decap_8 FILLER_2_936 ();
 sg13g2_decap_8 FILLER_2_943 ();
 sg13g2_decap_8 FILLER_2_950 ();
 sg13g2_decap_8 FILLER_2_957 ();
 sg13g2_decap_8 FILLER_2_964 ();
 sg13g2_decap_8 FILLER_2_971 ();
 sg13g2_decap_8 FILLER_2_978 ();
 sg13g2_decap_8 FILLER_2_985 ();
 sg13g2_decap_8 FILLER_2_992 ();
 sg13g2_decap_8 FILLER_2_999 ();
 sg13g2_decap_8 FILLER_2_1006 ();
 sg13g2_decap_8 FILLER_2_1013 ();
 sg13g2_decap_8 FILLER_2_1020 ();
 sg13g2_decap_8 FILLER_2_1027 ();
 sg13g2_decap_8 FILLER_2_1034 ();
 sg13g2_decap_8 FILLER_2_1041 ();
 sg13g2_decap_8 FILLER_2_1048 ();
 sg13g2_decap_8 FILLER_2_1055 ();
 sg13g2_decap_8 FILLER_2_1062 ();
 sg13g2_decap_8 FILLER_2_1069 ();
 sg13g2_decap_8 FILLER_2_1076 ();
 sg13g2_decap_8 FILLER_2_1083 ();
 sg13g2_decap_8 FILLER_2_1090 ();
 sg13g2_decap_8 FILLER_2_1097 ();
 sg13g2_decap_8 FILLER_2_1104 ();
 sg13g2_decap_8 FILLER_2_1111 ();
 sg13g2_decap_8 FILLER_2_1118 ();
 sg13g2_decap_8 FILLER_2_1125 ();
 sg13g2_decap_8 FILLER_2_1132 ();
 sg13g2_decap_8 FILLER_2_1139 ();
 sg13g2_decap_8 FILLER_2_1146 ();
 sg13g2_decap_8 FILLER_2_1153 ();
 sg13g2_decap_8 FILLER_2_1160 ();
 sg13g2_decap_8 FILLER_2_1167 ();
 sg13g2_decap_8 FILLER_2_1174 ();
 sg13g2_decap_8 FILLER_2_1181 ();
 sg13g2_decap_8 FILLER_2_1188 ();
 sg13g2_decap_8 FILLER_2_1195 ();
 sg13g2_decap_8 FILLER_2_1202 ();
 sg13g2_decap_8 FILLER_2_1209 ();
 sg13g2_decap_8 FILLER_2_1216 ();
 sg13g2_decap_8 FILLER_2_1223 ();
 sg13g2_decap_8 FILLER_2_1230 ();
 sg13g2_decap_8 FILLER_2_1237 ();
 sg13g2_decap_8 FILLER_2_1244 ();
 sg13g2_decap_8 FILLER_2_1251 ();
 sg13g2_decap_8 FILLER_2_1258 ();
 sg13g2_decap_8 FILLER_2_1265 ();
 sg13g2_decap_8 FILLER_2_1272 ();
 sg13g2_decap_8 FILLER_2_1279 ();
 sg13g2_decap_8 FILLER_2_1286 ();
 sg13g2_decap_8 FILLER_2_1293 ();
 sg13g2_decap_8 FILLER_2_1300 ();
 sg13g2_decap_8 FILLER_2_1307 ();
 sg13g2_fill_1 FILLER_2_1314 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_fill_2 FILLER_3_329 ();
 sg13g2_fill_1 FILLER_3_360 ();
 sg13g2_fill_2 FILLER_3_438 ();
 sg13g2_fill_1 FILLER_3_440 ();
 sg13g2_fill_2 FILLER_3_455 ();
 sg13g2_fill_1 FILLER_3_465 ();
 sg13g2_fill_2 FILLER_3_484 ();
 sg13g2_fill_1 FILLER_3_495 ();
 sg13g2_fill_1 FILLER_3_522 ();
 sg13g2_fill_1 FILLER_3_550 ();
 sg13g2_fill_2 FILLER_3_587 ();
 sg13g2_fill_2 FILLER_3_608 ();
 sg13g2_decap_4 FILLER_3_614 ();
 sg13g2_decap_4 FILLER_3_648 ();
 sg13g2_fill_1 FILLER_3_652 ();
 sg13g2_fill_2 FILLER_3_674 ();
 sg13g2_decap_8 FILLER_3_718 ();
 sg13g2_decap_8 FILLER_3_725 ();
 sg13g2_decap_4 FILLER_3_732 ();
 sg13g2_decap_8 FILLER_3_746 ();
 sg13g2_decap_4 FILLER_3_753 ();
 sg13g2_fill_2 FILLER_3_757 ();
 sg13g2_decap_4 FILLER_3_764 ();
 sg13g2_fill_2 FILLER_3_786 ();
 sg13g2_fill_1 FILLER_3_788 ();
 sg13g2_fill_1 FILLER_3_850 ();
 sg13g2_fill_2 FILLER_3_863 ();
 sg13g2_fill_2 FILLER_3_870 ();
 sg13g2_fill_1 FILLER_3_872 ();
 sg13g2_fill_1 FILLER_3_878 ();
 sg13g2_decap_4 FILLER_3_891 ();
 sg13g2_decap_8 FILLER_3_908 ();
 sg13g2_decap_8 FILLER_3_915 ();
 sg13g2_decap_8 FILLER_3_922 ();
 sg13g2_decap_8 FILLER_3_929 ();
 sg13g2_decap_8 FILLER_3_936 ();
 sg13g2_decap_8 FILLER_3_943 ();
 sg13g2_decap_8 FILLER_3_950 ();
 sg13g2_decap_8 FILLER_3_957 ();
 sg13g2_decap_8 FILLER_3_964 ();
 sg13g2_decap_8 FILLER_3_971 ();
 sg13g2_decap_8 FILLER_3_978 ();
 sg13g2_decap_8 FILLER_3_985 ();
 sg13g2_decap_8 FILLER_3_992 ();
 sg13g2_decap_8 FILLER_3_999 ();
 sg13g2_decap_8 FILLER_3_1006 ();
 sg13g2_decap_8 FILLER_3_1013 ();
 sg13g2_decap_8 FILLER_3_1020 ();
 sg13g2_decap_8 FILLER_3_1027 ();
 sg13g2_decap_8 FILLER_3_1034 ();
 sg13g2_decap_8 FILLER_3_1041 ();
 sg13g2_decap_8 FILLER_3_1048 ();
 sg13g2_decap_8 FILLER_3_1055 ();
 sg13g2_decap_8 FILLER_3_1062 ();
 sg13g2_decap_8 FILLER_3_1069 ();
 sg13g2_decap_8 FILLER_3_1076 ();
 sg13g2_decap_8 FILLER_3_1083 ();
 sg13g2_decap_8 FILLER_3_1090 ();
 sg13g2_decap_8 FILLER_3_1097 ();
 sg13g2_decap_8 FILLER_3_1104 ();
 sg13g2_decap_8 FILLER_3_1111 ();
 sg13g2_decap_8 FILLER_3_1118 ();
 sg13g2_decap_8 FILLER_3_1125 ();
 sg13g2_decap_8 FILLER_3_1132 ();
 sg13g2_decap_8 FILLER_3_1139 ();
 sg13g2_decap_8 FILLER_3_1146 ();
 sg13g2_decap_8 FILLER_3_1153 ();
 sg13g2_decap_8 FILLER_3_1160 ();
 sg13g2_decap_8 FILLER_3_1167 ();
 sg13g2_decap_8 FILLER_3_1174 ();
 sg13g2_decap_8 FILLER_3_1181 ();
 sg13g2_decap_8 FILLER_3_1188 ();
 sg13g2_decap_8 FILLER_3_1195 ();
 sg13g2_decap_8 FILLER_3_1202 ();
 sg13g2_decap_8 FILLER_3_1209 ();
 sg13g2_decap_8 FILLER_3_1216 ();
 sg13g2_decap_8 FILLER_3_1223 ();
 sg13g2_decap_8 FILLER_3_1230 ();
 sg13g2_decap_8 FILLER_3_1237 ();
 sg13g2_decap_8 FILLER_3_1244 ();
 sg13g2_decap_8 FILLER_3_1251 ();
 sg13g2_decap_8 FILLER_3_1258 ();
 sg13g2_decap_8 FILLER_3_1265 ();
 sg13g2_decap_8 FILLER_3_1272 ();
 sg13g2_decap_8 FILLER_3_1279 ();
 sg13g2_decap_8 FILLER_3_1286 ();
 sg13g2_decap_8 FILLER_3_1293 ();
 sg13g2_decap_8 FILLER_3_1300 ();
 sg13g2_decap_8 FILLER_3_1307 ();
 sg13g2_fill_1 FILLER_3_1314 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_fill_2 FILLER_4_266 ();
 sg13g2_fill_1 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_fill_1 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_285 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_fill_1 FILLER_4_299 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_fill_1 FILLER_4_359 ();
 sg13g2_fill_2 FILLER_4_370 ();
 sg13g2_fill_2 FILLER_4_382 ();
 sg13g2_fill_2 FILLER_4_394 ();
 sg13g2_fill_1 FILLER_4_396 ();
 sg13g2_fill_2 FILLER_4_402 ();
 sg13g2_fill_2 FILLER_4_409 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_fill_2 FILLER_4_444 ();
 sg13g2_decap_4 FILLER_4_456 ();
 sg13g2_fill_2 FILLER_4_516 ();
 sg13g2_fill_1 FILLER_4_518 ();
 sg13g2_fill_2 FILLER_4_560 ();
 sg13g2_fill_1 FILLER_4_562 ();
 sg13g2_fill_1 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_694 ();
 sg13g2_decap_8 FILLER_4_701 ();
 sg13g2_decap_8 FILLER_4_708 ();
 sg13g2_fill_2 FILLER_4_715 ();
 sg13g2_fill_1 FILLER_4_717 ();
 sg13g2_fill_1 FILLER_4_738 ();
 sg13g2_fill_2 FILLER_4_775 ();
 sg13g2_fill_1 FILLER_4_777 ();
 sg13g2_fill_2 FILLER_4_817 ();
 sg13g2_fill_1 FILLER_4_819 ();
 sg13g2_fill_1 FILLER_4_828 ();
 sg13g2_fill_1 FILLER_4_846 ();
 sg13g2_fill_2 FILLER_4_862 ();
 sg13g2_decap_4 FILLER_4_879 ();
 sg13g2_fill_2 FILLER_4_883 ();
 sg13g2_fill_2 FILLER_4_894 ();
 sg13g2_decap_8 FILLER_4_906 ();
 sg13g2_decap_8 FILLER_4_913 ();
 sg13g2_decap_8 FILLER_4_920 ();
 sg13g2_decap_8 FILLER_4_927 ();
 sg13g2_decap_8 FILLER_4_934 ();
 sg13g2_decap_8 FILLER_4_941 ();
 sg13g2_decap_8 FILLER_4_948 ();
 sg13g2_decap_8 FILLER_4_955 ();
 sg13g2_decap_8 FILLER_4_962 ();
 sg13g2_decap_8 FILLER_4_969 ();
 sg13g2_decap_8 FILLER_4_976 ();
 sg13g2_decap_8 FILLER_4_983 ();
 sg13g2_decap_8 FILLER_4_990 ();
 sg13g2_decap_8 FILLER_4_997 ();
 sg13g2_decap_8 FILLER_4_1004 ();
 sg13g2_decap_8 FILLER_4_1011 ();
 sg13g2_decap_8 FILLER_4_1018 ();
 sg13g2_decap_8 FILLER_4_1025 ();
 sg13g2_decap_8 FILLER_4_1032 ();
 sg13g2_decap_8 FILLER_4_1039 ();
 sg13g2_decap_8 FILLER_4_1046 ();
 sg13g2_decap_8 FILLER_4_1053 ();
 sg13g2_decap_8 FILLER_4_1060 ();
 sg13g2_decap_8 FILLER_4_1067 ();
 sg13g2_decap_8 FILLER_4_1074 ();
 sg13g2_decap_8 FILLER_4_1081 ();
 sg13g2_decap_8 FILLER_4_1088 ();
 sg13g2_decap_8 FILLER_4_1095 ();
 sg13g2_decap_8 FILLER_4_1102 ();
 sg13g2_decap_8 FILLER_4_1109 ();
 sg13g2_decap_8 FILLER_4_1116 ();
 sg13g2_decap_8 FILLER_4_1123 ();
 sg13g2_decap_8 FILLER_4_1130 ();
 sg13g2_decap_8 FILLER_4_1137 ();
 sg13g2_decap_8 FILLER_4_1144 ();
 sg13g2_decap_8 FILLER_4_1151 ();
 sg13g2_decap_8 FILLER_4_1158 ();
 sg13g2_decap_8 FILLER_4_1165 ();
 sg13g2_decap_8 FILLER_4_1172 ();
 sg13g2_decap_8 FILLER_4_1179 ();
 sg13g2_decap_8 FILLER_4_1186 ();
 sg13g2_decap_8 FILLER_4_1193 ();
 sg13g2_decap_8 FILLER_4_1200 ();
 sg13g2_decap_8 FILLER_4_1207 ();
 sg13g2_decap_8 FILLER_4_1214 ();
 sg13g2_decap_8 FILLER_4_1221 ();
 sg13g2_decap_8 FILLER_4_1228 ();
 sg13g2_decap_8 FILLER_4_1235 ();
 sg13g2_decap_8 FILLER_4_1242 ();
 sg13g2_decap_8 FILLER_4_1249 ();
 sg13g2_decap_8 FILLER_4_1256 ();
 sg13g2_decap_8 FILLER_4_1263 ();
 sg13g2_decap_8 FILLER_4_1270 ();
 sg13g2_decap_8 FILLER_4_1277 ();
 sg13g2_decap_8 FILLER_4_1284 ();
 sg13g2_decap_8 FILLER_4_1291 ();
 sg13g2_decap_8 FILLER_4_1298 ();
 sg13g2_decap_8 FILLER_4_1305 ();
 sg13g2_fill_2 FILLER_4_1312 ();
 sg13g2_fill_1 FILLER_4_1314 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_4 FILLER_5_259 ();
 sg13g2_fill_2 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_fill_1 FILLER_5_335 ();
 sg13g2_fill_2 FILLER_5_377 ();
 sg13g2_fill_2 FILLER_5_405 ();
 sg13g2_fill_2 FILLER_5_412 ();
 sg13g2_fill_1 FILLER_5_414 ();
 sg13g2_fill_1 FILLER_5_446 ();
 sg13g2_fill_1 FILLER_5_477 ();
 sg13g2_fill_2 FILLER_5_491 ();
 sg13g2_fill_1 FILLER_5_502 ();
 sg13g2_fill_2 FILLER_5_520 ();
 sg13g2_fill_1 FILLER_5_527 ();
 sg13g2_fill_1 FILLER_5_553 ();
 sg13g2_fill_1 FILLER_5_629 ();
 sg13g2_decap_4 FILLER_5_664 ();
 sg13g2_fill_1 FILLER_5_668 ();
 sg13g2_decap_4 FILLER_5_690 ();
 sg13g2_fill_1 FILLER_5_715 ();
 sg13g2_fill_2 FILLER_5_737 ();
 sg13g2_fill_1 FILLER_5_739 ();
 sg13g2_fill_2 FILLER_5_763 ();
 sg13g2_fill_1 FILLER_5_765 ();
 sg13g2_decap_4 FILLER_5_780 ();
 sg13g2_decap_8 FILLER_5_792 ();
 sg13g2_fill_1 FILLER_5_799 ();
 sg13g2_decap_4 FILLER_5_805 ();
 sg13g2_fill_1 FILLER_5_809 ();
 sg13g2_fill_2 FILLER_5_815 ();
 sg13g2_fill_1 FILLER_5_817 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_4 FILLER_5_861 ();
 sg13g2_fill_1 FILLER_5_869 ();
 sg13g2_fill_2 FILLER_5_880 ();
 sg13g2_fill_1 FILLER_5_882 ();
 sg13g2_decap_8 FILLER_5_891 ();
 sg13g2_fill_2 FILLER_5_898 ();
 sg13g2_fill_1 FILLER_5_900 ();
 sg13g2_decap_8 FILLER_5_905 ();
 sg13g2_decap_8 FILLER_5_912 ();
 sg13g2_decap_8 FILLER_5_919 ();
 sg13g2_decap_8 FILLER_5_926 ();
 sg13g2_decap_8 FILLER_5_933 ();
 sg13g2_decap_8 FILLER_5_940 ();
 sg13g2_decap_8 FILLER_5_947 ();
 sg13g2_decap_8 FILLER_5_954 ();
 sg13g2_decap_8 FILLER_5_961 ();
 sg13g2_decap_8 FILLER_5_968 ();
 sg13g2_decap_8 FILLER_5_975 ();
 sg13g2_decap_8 FILLER_5_982 ();
 sg13g2_decap_8 FILLER_5_989 ();
 sg13g2_decap_8 FILLER_5_996 ();
 sg13g2_decap_8 FILLER_5_1003 ();
 sg13g2_decap_8 FILLER_5_1010 ();
 sg13g2_decap_8 FILLER_5_1017 ();
 sg13g2_decap_8 FILLER_5_1024 ();
 sg13g2_decap_8 FILLER_5_1031 ();
 sg13g2_decap_8 FILLER_5_1038 ();
 sg13g2_decap_8 FILLER_5_1045 ();
 sg13g2_decap_8 FILLER_5_1052 ();
 sg13g2_decap_8 FILLER_5_1059 ();
 sg13g2_decap_8 FILLER_5_1066 ();
 sg13g2_decap_8 FILLER_5_1073 ();
 sg13g2_decap_8 FILLER_5_1080 ();
 sg13g2_decap_8 FILLER_5_1087 ();
 sg13g2_decap_8 FILLER_5_1094 ();
 sg13g2_decap_8 FILLER_5_1101 ();
 sg13g2_decap_8 FILLER_5_1108 ();
 sg13g2_decap_8 FILLER_5_1115 ();
 sg13g2_decap_8 FILLER_5_1122 ();
 sg13g2_decap_8 FILLER_5_1129 ();
 sg13g2_decap_8 FILLER_5_1136 ();
 sg13g2_decap_8 FILLER_5_1143 ();
 sg13g2_decap_8 FILLER_5_1150 ();
 sg13g2_decap_8 FILLER_5_1157 ();
 sg13g2_decap_8 FILLER_5_1164 ();
 sg13g2_decap_8 FILLER_5_1171 ();
 sg13g2_decap_8 FILLER_5_1178 ();
 sg13g2_decap_8 FILLER_5_1185 ();
 sg13g2_decap_8 FILLER_5_1192 ();
 sg13g2_decap_8 FILLER_5_1199 ();
 sg13g2_decap_8 FILLER_5_1206 ();
 sg13g2_decap_8 FILLER_5_1213 ();
 sg13g2_decap_8 FILLER_5_1220 ();
 sg13g2_decap_8 FILLER_5_1227 ();
 sg13g2_decap_8 FILLER_5_1234 ();
 sg13g2_decap_8 FILLER_5_1241 ();
 sg13g2_decap_8 FILLER_5_1248 ();
 sg13g2_decap_8 FILLER_5_1255 ();
 sg13g2_decap_8 FILLER_5_1262 ();
 sg13g2_decap_8 FILLER_5_1269 ();
 sg13g2_decap_8 FILLER_5_1276 ();
 sg13g2_decap_8 FILLER_5_1283 ();
 sg13g2_decap_8 FILLER_5_1290 ();
 sg13g2_decap_8 FILLER_5_1297 ();
 sg13g2_decap_8 FILLER_5_1304 ();
 sg13g2_decap_4 FILLER_5_1311 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_fill_2 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_237 ();
 sg13g2_fill_1 FILLER_6_244 ();
 sg13g2_fill_2 FILLER_6_253 ();
 sg13g2_fill_1 FILLER_6_281 ();
 sg13g2_fill_2 FILLER_6_313 ();
 sg13g2_fill_1 FILLER_6_315 ();
 sg13g2_fill_2 FILLER_6_342 ();
 sg13g2_fill_1 FILLER_6_344 ();
 sg13g2_fill_2 FILLER_6_349 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_fill_2 FILLER_6_377 ();
 sg13g2_fill_1 FILLER_6_379 ();
 sg13g2_fill_2 FILLER_6_410 ();
 sg13g2_decap_4 FILLER_6_425 ();
 sg13g2_fill_2 FILLER_6_442 ();
 sg13g2_fill_2 FILLER_6_453 ();
 sg13g2_fill_1 FILLER_6_455 ();
 sg13g2_fill_1 FILLER_6_472 ();
 sg13g2_fill_1 FILLER_6_508 ();
 sg13g2_fill_1 FILLER_6_519 ();
 sg13g2_fill_2 FILLER_6_558 ();
 sg13g2_fill_1 FILLER_6_560 ();
 sg13g2_decap_4 FILLER_6_582 ();
 sg13g2_fill_1 FILLER_6_610 ();
 sg13g2_decap_4 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_645 ();
 sg13g2_fill_1 FILLER_6_652 ();
 sg13g2_decap_8 FILLER_6_673 ();
 sg13g2_decap_4 FILLER_6_680 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_fill_1 FILLER_6_704 ();
 sg13g2_fill_2 FILLER_6_732 ();
 sg13g2_decap_4 FILLER_6_744 ();
 sg13g2_decap_4 FILLER_6_752 ();
 sg13g2_fill_2 FILLER_6_756 ();
 sg13g2_fill_2 FILLER_6_785 ();
 sg13g2_fill_2 FILLER_6_795 ();
 sg13g2_fill_1 FILLER_6_797 ();
 sg13g2_fill_2 FILLER_6_808 ();
 sg13g2_decap_8 FILLER_6_815 ();
 sg13g2_fill_2 FILLER_6_822 ();
 sg13g2_fill_2 FILLER_6_828 ();
 sg13g2_decap_4 FILLER_6_850 ();
 sg13g2_fill_1 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_862 ();
 sg13g2_fill_1 FILLER_6_888 ();
 sg13g2_decap_8 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_914 ();
 sg13g2_decap_8 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_6_928 ();
 sg13g2_decap_8 FILLER_6_935 ();
 sg13g2_decap_8 FILLER_6_942 ();
 sg13g2_decap_8 FILLER_6_949 ();
 sg13g2_decap_8 FILLER_6_956 ();
 sg13g2_decap_8 FILLER_6_963 ();
 sg13g2_decap_8 FILLER_6_970 ();
 sg13g2_decap_8 FILLER_6_977 ();
 sg13g2_decap_8 FILLER_6_984 ();
 sg13g2_decap_8 FILLER_6_991 ();
 sg13g2_decap_8 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_8 FILLER_6_1019 ();
 sg13g2_decap_8 FILLER_6_1026 ();
 sg13g2_decap_8 FILLER_6_1033 ();
 sg13g2_decap_8 FILLER_6_1040 ();
 sg13g2_decap_8 FILLER_6_1047 ();
 sg13g2_decap_8 FILLER_6_1054 ();
 sg13g2_decap_8 FILLER_6_1061 ();
 sg13g2_decap_8 FILLER_6_1068 ();
 sg13g2_decap_8 FILLER_6_1075 ();
 sg13g2_decap_8 FILLER_6_1082 ();
 sg13g2_decap_8 FILLER_6_1089 ();
 sg13g2_decap_8 FILLER_6_1096 ();
 sg13g2_decap_8 FILLER_6_1103 ();
 sg13g2_decap_8 FILLER_6_1110 ();
 sg13g2_decap_8 FILLER_6_1117 ();
 sg13g2_decap_8 FILLER_6_1124 ();
 sg13g2_decap_8 FILLER_6_1131 ();
 sg13g2_decap_8 FILLER_6_1138 ();
 sg13g2_decap_8 FILLER_6_1145 ();
 sg13g2_decap_8 FILLER_6_1152 ();
 sg13g2_decap_8 FILLER_6_1159 ();
 sg13g2_decap_8 FILLER_6_1166 ();
 sg13g2_decap_8 FILLER_6_1173 ();
 sg13g2_decap_8 FILLER_6_1180 ();
 sg13g2_decap_8 FILLER_6_1187 ();
 sg13g2_decap_8 FILLER_6_1194 ();
 sg13g2_decap_8 FILLER_6_1201 ();
 sg13g2_decap_8 FILLER_6_1208 ();
 sg13g2_decap_8 FILLER_6_1215 ();
 sg13g2_decap_8 FILLER_6_1222 ();
 sg13g2_decap_8 FILLER_6_1229 ();
 sg13g2_decap_8 FILLER_6_1236 ();
 sg13g2_decap_8 FILLER_6_1243 ();
 sg13g2_decap_8 FILLER_6_1250 ();
 sg13g2_decap_8 FILLER_6_1257 ();
 sg13g2_decap_8 FILLER_6_1264 ();
 sg13g2_decap_8 FILLER_6_1271 ();
 sg13g2_decap_8 FILLER_6_1278 ();
 sg13g2_decap_8 FILLER_6_1285 ();
 sg13g2_decap_8 FILLER_6_1292 ();
 sg13g2_decap_8 FILLER_6_1299 ();
 sg13g2_decap_8 FILLER_6_1306 ();
 sg13g2_fill_2 FILLER_6_1313 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_4 FILLER_7_217 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_fill_1 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_288 ();
 sg13g2_fill_2 FILLER_7_315 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_fill_2 FILLER_7_459 ();
 sg13g2_fill_1 FILLER_7_461 ();
 sg13g2_fill_2 FILLER_7_471 ();
 sg13g2_fill_2 FILLER_7_478 ();
 sg13g2_fill_1 FILLER_7_480 ();
 sg13g2_fill_2 FILLER_7_502 ();
 sg13g2_fill_1 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_540 ();
 sg13g2_fill_1 FILLER_7_547 ();
 sg13g2_fill_2 FILLER_7_552 ();
 sg13g2_decap_4 FILLER_7_582 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_fill_2 FILLER_7_602 ();
 sg13g2_fill_1 FILLER_7_604 ();
 sg13g2_decap_8 FILLER_7_613 ();
 sg13g2_fill_2 FILLER_7_624 ();
 sg13g2_fill_1 FILLER_7_626 ();
 sg13g2_decap_8 FILLER_7_653 ();
 sg13g2_decap_8 FILLER_7_670 ();
 sg13g2_decap_8 FILLER_7_677 ();
 sg13g2_fill_2 FILLER_7_744 ();
 sg13g2_decap_4 FILLER_7_758 ();
 sg13g2_fill_2 FILLER_7_762 ();
 sg13g2_fill_1 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_776 ();
 sg13g2_fill_2 FILLER_7_810 ();
 sg13g2_fill_2 FILLER_7_817 ();
 sg13g2_fill_2 FILLER_7_824 ();
 sg13g2_fill_2 FILLER_7_845 ();
 sg13g2_fill_1 FILLER_7_880 ();
 sg13g2_fill_1 FILLER_7_889 ();
 sg13g2_decap_8 FILLER_7_910 ();
 sg13g2_decap_8 FILLER_7_917 ();
 sg13g2_decap_8 FILLER_7_924 ();
 sg13g2_decap_8 FILLER_7_931 ();
 sg13g2_decap_8 FILLER_7_938 ();
 sg13g2_decap_8 FILLER_7_945 ();
 sg13g2_decap_8 FILLER_7_952 ();
 sg13g2_decap_8 FILLER_7_959 ();
 sg13g2_decap_8 FILLER_7_966 ();
 sg13g2_decap_8 FILLER_7_973 ();
 sg13g2_decap_8 FILLER_7_980 ();
 sg13g2_decap_8 FILLER_7_987 ();
 sg13g2_decap_8 FILLER_7_994 ();
 sg13g2_decap_8 FILLER_7_1001 ();
 sg13g2_decap_8 FILLER_7_1008 ();
 sg13g2_decap_8 FILLER_7_1015 ();
 sg13g2_decap_8 FILLER_7_1022 ();
 sg13g2_decap_8 FILLER_7_1029 ();
 sg13g2_decap_8 FILLER_7_1036 ();
 sg13g2_decap_8 FILLER_7_1043 ();
 sg13g2_decap_8 FILLER_7_1050 ();
 sg13g2_decap_8 FILLER_7_1057 ();
 sg13g2_decap_8 FILLER_7_1064 ();
 sg13g2_decap_8 FILLER_7_1071 ();
 sg13g2_decap_8 FILLER_7_1078 ();
 sg13g2_decap_8 FILLER_7_1085 ();
 sg13g2_decap_8 FILLER_7_1092 ();
 sg13g2_decap_8 FILLER_7_1099 ();
 sg13g2_decap_8 FILLER_7_1106 ();
 sg13g2_decap_8 FILLER_7_1113 ();
 sg13g2_decap_8 FILLER_7_1120 ();
 sg13g2_decap_8 FILLER_7_1127 ();
 sg13g2_decap_8 FILLER_7_1134 ();
 sg13g2_decap_8 FILLER_7_1141 ();
 sg13g2_decap_8 FILLER_7_1148 ();
 sg13g2_decap_8 FILLER_7_1155 ();
 sg13g2_decap_8 FILLER_7_1162 ();
 sg13g2_decap_8 FILLER_7_1169 ();
 sg13g2_decap_8 FILLER_7_1176 ();
 sg13g2_decap_8 FILLER_7_1183 ();
 sg13g2_decap_8 FILLER_7_1190 ();
 sg13g2_decap_8 FILLER_7_1197 ();
 sg13g2_decap_8 FILLER_7_1204 ();
 sg13g2_decap_8 FILLER_7_1211 ();
 sg13g2_decap_8 FILLER_7_1218 ();
 sg13g2_decap_8 FILLER_7_1225 ();
 sg13g2_decap_8 FILLER_7_1232 ();
 sg13g2_decap_8 FILLER_7_1239 ();
 sg13g2_decap_8 FILLER_7_1246 ();
 sg13g2_decap_8 FILLER_7_1253 ();
 sg13g2_decap_8 FILLER_7_1260 ();
 sg13g2_decap_8 FILLER_7_1267 ();
 sg13g2_decap_8 FILLER_7_1274 ();
 sg13g2_decap_8 FILLER_7_1281 ();
 sg13g2_decap_8 FILLER_7_1288 ();
 sg13g2_decap_8 FILLER_7_1295 ();
 sg13g2_decap_8 FILLER_7_1302 ();
 sg13g2_decap_4 FILLER_7_1309 ();
 sg13g2_fill_2 FILLER_7_1313 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_283 ();
 sg13g2_decap_4 FILLER_8_298 ();
 sg13g2_fill_1 FILLER_8_302 ();
 sg13g2_fill_2 FILLER_8_308 ();
 sg13g2_fill_1 FILLER_8_310 ();
 sg13g2_fill_1 FILLER_8_360 ();
 sg13g2_fill_2 FILLER_8_383 ();
 sg13g2_fill_1 FILLER_8_385 ();
 sg13g2_fill_1 FILLER_8_399 ();
 sg13g2_fill_1 FILLER_8_409 ();
 sg13g2_fill_1 FILLER_8_436 ();
 sg13g2_fill_2 FILLER_8_459 ();
 sg13g2_fill_1 FILLER_8_461 ();
 sg13g2_fill_2 FILLER_8_467 ();
 sg13g2_fill_1 FILLER_8_469 ();
 sg13g2_fill_1 FILLER_8_517 ();
 sg13g2_fill_2 FILLER_8_523 ();
 sg13g2_fill_1 FILLER_8_525 ();
 sg13g2_fill_1 FILLER_8_531 ();
 sg13g2_fill_2 FILLER_8_571 ();
 sg13g2_fill_1 FILLER_8_573 ();
 sg13g2_decap_8 FILLER_8_605 ();
 sg13g2_decap_8 FILLER_8_612 ();
 sg13g2_fill_2 FILLER_8_619 ();
 sg13g2_decap_8 FILLER_8_625 ();
 sg13g2_fill_1 FILLER_8_632 ();
 sg13g2_decap_4 FILLER_8_647 ();
 sg13g2_fill_2 FILLER_8_659 ();
 sg13g2_decap_8 FILLER_8_671 ();
 sg13g2_decap_8 FILLER_8_678 ();
 sg13g2_decap_8 FILLER_8_685 ();
 sg13g2_decap_4 FILLER_8_692 ();
 sg13g2_fill_1 FILLER_8_696 ();
 sg13g2_decap_4 FILLER_8_712 ();
 sg13g2_fill_2 FILLER_8_730 ();
 sg13g2_fill_1 FILLER_8_747 ();
 sg13g2_fill_2 FILLER_8_763 ();
 sg13g2_fill_1 FILLER_8_765 ();
 sg13g2_fill_2 FILLER_8_779 ();
 sg13g2_decap_4 FILLER_8_812 ();
 sg13g2_fill_2 FILLER_8_816 ();
 sg13g2_fill_2 FILLER_8_828 ();
 sg13g2_fill_1 FILLER_8_830 ();
 sg13g2_decap_4 FILLER_8_834 ();
 sg13g2_fill_1 FILLER_8_838 ();
 sg13g2_fill_2 FILLER_8_844 ();
 sg13g2_fill_1 FILLER_8_855 ();
 sg13g2_decap_8 FILLER_8_902 ();
 sg13g2_decap_8 FILLER_8_909 ();
 sg13g2_decap_8 FILLER_8_916 ();
 sg13g2_decap_8 FILLER_8_923 ();
 sg13g2_decap_8 FILLER_8_930 ();
 sg13g2_decap_8 FILLER_8_937 ();
 sg13g2_decap_8 FILLER_8_944 ();
 sg13g2_decap_8 FILLER_8_951 ();
 sg13g2_decap_8 FILLER_8_958 ();
 sg13g2_decap_8 FILLER_8_965 ();
 sg13g2_decap_8 FILLER_8_972 ();
 sg13g2_decap_8 FILLER_8_979 ();
 sg13g2_decap_8 FILLER_8_986 ();
 sg13g2_decap_8 FILLER_8_993 ();
 sg13g2_decap_8 FILLER_8_1000 ();
 sg13g2_decap_8 FILLER_8_1007 ();
 sg13g2_decap_8 FILLER_8_1014 ();
 sg13g2_decap_8 FILLER_8_1021 ();
 sg13g2_decap_8 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_8_1035 ();
 sg13g2_decap_8 FILLER_8_1042 ();
 sg13g2_decap_8 FILLER_8_1049 ();
 sg13g2_decap_8 FILLER_8_1056 ();
 sg13g2_decap_8 FILLER_8_1063 ();
 sg13g2_decap_8 FILLER_8_1070 ();
 sg13g2_decap_8 FILLER_8_1077 ();
 sg13g2_decap_8 FILLER_8_1084 ();
 sg13g2_decap_8 FILLER_8_1091 ();
 sg13g2_decap_8 FILLER_8_1098 ();
 sg13g2_decap_8 FILLER_8_1105 ();
 sg13g2_decap_8 FILLER_8_1112 ();
 sg13g2_decap_8 FILLER_8_1119 ();
 sg13g2_decap_8 FILLER_8_1126 ();
 sg13g2_decap_8 FILLER_8_1133 ();
 sg13g2_decap_8 FILLER_8_1140 ();
 sg13g2_decap_8 FILLER_8_1147 ();
 sg13g2_decap_8 FILLER_8_1154 ();
 sg13g2_decap_8 FILLER_8_1161 ();
 sg13g2_decap_8 FILLER_8_1168 ();
 sg13g2_decap_8 FILLER_8_1175 ();
 sg13g2_decap_8 FILLER_8_1182 ();
 sg13g2_decap_8 FILLER_8_1189 ();
 sg13g2_decap_8 FILLER_8_1196 ();
 sg13g2_decap_8 FILLER_8_1203 ();
 sg13g2_decap_8 FILLER_8_1210 ();
 sg13g2_decap_8 FILLER_8_1217 ();
 sg13g2_decap_8 FILLER_8_1224 ();
 sg13g2_decap_8 FILLER_8_1231 ();
 sg13g2_decap_8 FILLER_8_1238 ();
 sg13g2_decap_8 FILLER_8_1245 ();
 sg13g2_decap_8 FILLER_8_1252 ();
 sg13g2_decap_8 FILLER_8_1259 ();
 sg13g2_decap_8 FILLER_8_1266 ();
 sg13g2_decap_8 FILLER_8_1273 ();
 sg13g2_decap_8 FILLER_8_1280 ();
 sg13g2_decap_8 FILLER_8_1287 ();
 sg13g2_decap_8 FILLER_8_1294 ();
 sg13g2_decap_8 FILLER_8_1301 ();
 sg13g2_decap_8 FILLER_8_1308 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_fill_2 FILLER_9_210 ();
 sg13g2_fill_1 FILLER_9_212 ();
 sg13g2_decap_8 FILLER_9_248 ();
 sg13g2_fill_2 FILLER_9_255 ();
 sg13g2_fill_1 FILLER_9_257 ();
 sg13g2_fill_1 FILLER_9_272 ();
 sg13g2_fill_2 FILLER_9_297 ();
 sg13g2_fill_1 FILLER_9_299 ();
 sg13g2_fill_1 FILLER_9_386 ();
 sg13g2_decap_4 FILLER_9_410 ();
 sg13g2_fill_1 FILLER_9_414 ();
 sg13g2_fill_1 FILLER_9_454 ();
 sg13g2_decap_8 FILLER_9_485 ();
 sg13g2_fill_2 FILLER_9_513 ();
 sg13g2_fill_2 FILLER_9_586 ();
 sg13g2_fill_1 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_641 ();
 sg13g2_decap_4 FILLER_9_710 ();
 sg13g2_fill_2 FILLER_9_729 ();
 sg13g2_fill_1 FILLER_9_731 ();
 sg13g2_decap_8 FILLER_9_737 ();
 sg13g2_decap_4 FILLER_9_744 ();
 sg13g2_fill_2 FILLER_9_748 ();
 sg13g2_fill_2 FILLER_9_765 ();
 sg13g2_decap_4 FILLER_9_780 ();
 sg13g2_fill_2 FILLER_9_789 ();
 sg13g2_fill_2 FILLER_9_796 ();
 sg13g2_fill_2 FILLER_9_824 ();
 sg13g2_decap_4 FILLER_9_861 ();
 sg13g2_fill_2 FILLER_9_865 ();
 sg13g2_decap_4 FILLER_9_877 ();
 sg13g2_fill_2 FILLER_9_897 ();
 sg13g2_fill_1 FILLER_9_899 ();
 sg13g2_decap_8 FILLER_9_912 ();
 sg13g2_decap_8 FILLER_9_919 ();
 sg13g2_decap_8 FILLER_9_926 ();
 sg13g2_decap_8 FILLER_9_933 ();
 sg13g2_decap_8 FILLER_9_940 ();
 sg13g2_decap_8 FILLER_9_947 ();
 sg13g2_decap_8 FILLER_9_954 ();
 sg13g2_decap_8 FILLER_9_961 ();
 sg13g2_decap_8 FILLER_9_968 ();
 sg13g2_decap_8 FILLER_9_975 ();
 sg13g2_decap_8 FILLER_9_982 ();
 sg13g2_decap_8 FILLER_9_989 ();
 sg13g2_decap_8 FILLER_9_996 ();
 sg13g2_decap_8 FILLER_9_1003 ();
 sg13g2_decap_8 FILLER_9_1010 ();
 sg13g2_decap_8 FILLER_9_1017 ();
 sg13g2_decap_8 FILLER_9_1024 ();
 sg13g2_decap_8 FILLER_9_1031 ();
 sg13g2_decap_8 FILLER_9_1038 ();
 sg13g2_decap_8 FILLER_9_1045 ();
 sg13g2_decap_8 FILLER_9_1052 ();
 sg13g2_decap_8 FILLER_9_1059 ();
 sg13g2_decap_8 FILLER_9_1066 ();
 sg13g2_decap_8 FILLER_9_1073 ();
 sg13g2_decap_8 FILLER_9_1080 ();
 sg13g2_decap_8 FILLER_9_1087 ();
 sg13g2_decap_8 FILLER_9_1094 ();
 sg13g2_decap_8 FILLER_9_1101 ();
 sg13g2_decap_8 FILLER_9_1108 ();
 sg13g2_decap_8 FILLER_9_1115 ();
 sg13g2_decap_8 FILLER_9_1122 ();
 sg13g2_decap_8 FILLER_9_1129 ();
 sg13g2_decap_8 FILLER_9_1136 ();
 sg13g2_decap_8 FILLER_9_1143 ();
 sg13g2_decap_8 FILLER_9_1150 ();
 sg13g2_decap_8 FILLER_9_1157 ();
 sg13g2_decap_8 FILLER_9_1164 ();
 sg13g2_decap_8 FILLER_9_1171 ();
 sg13g2_decap_8 FILLER_9_1178 ();
 sg13g2_decap_8 FILLER_9_1185 ();
 sg13g2_decap_8 FILLER_9_1192 ();
 sg13g2_decap_8 FILLER_9_1199 ();
 sg13g2_decap_8 FILLER_9_1206 ();
 sg13g2_decap_8 FILLER_9_1213 ();
 sg13g2_decap_8 FILLER_9_1220 ();
 sg13g2_decap_8 FILLER_9_1227 ();
 sg13g2_decap_8 FILLER_9_1234 ();
 sg13g2_decap_8 FILLER_9_1241 ();
 sg13g2_decap_8 FILLER_9_1248 ();
 sg13g2_decap_8 FILLER_9_1255 ();
 sg13g2_decap_8 FILLER_9_1262 ();
 sg13g2_decap_8 FILLER_9_1269 ();
 sg13g2_decap_8 FILLER_9_1276 ();
 sg13g2_decap_8 FILLER_9_1283 ();
 sg13g2_decap_8 FILLER_9_1290 ();
 sg13g2_decap_8 FILLER_9_1297 ();
 sg13g2_decap_8 FILLER_9_1304 ();
 sg13g2_decap_4 FILLER_9_1311 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_fill_2 FILLER_10_217 ();
 sg13g2_fill_2 FILLER_10_251 ();
 sg13g2_fill_1 FILLER_10_253 ();
 sg13g2_decap_4 FILLER_10_280 ();
 sg13g2_fill_1 FILLER_10_293 ();
 sg13g2_fill_1 FILLER_10_334 ();
 sg13g2_fill_1 FILLER_10_354 ();
 sg13g2_fill_2 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_373 ();
 sg13g2_fill_1 FILLER_10_500 ();
 sg13g2_fill_2 FILLER_10_510 ();
 sg13g2_fill_1 FILLER_10_512 ();
 sg13g2_fill_1 FILLER_10_529 ();
 sg13g2_fill_2 FILLER_10_535 ();
 sg13g2_fill_1 FILLER_10_537 ();
 sg13g2_fill_1 FILLER_10_547 ();
 sg13g2_fill_2 FILLER_10_556 ();
 sg13g2_fill_1 FILLER_10_558 ();
 sg13g2_decap_8 FILLER_10_611 ();
 sg13g2_decap_8 FILLER_10_618 ();
 sg13g2_fill_1 FILLER_10_625 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_4 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_649 ();
 sg13g2_decap_8 FILLER_10_666 ();
 sg13g2_fill_2 FILLER_10_673 ();
 sg13g2_decap_8 FILLER_10_685 ();
 sg13g2_decap_8 FILLER_10_692 ();
 sg13g2_fill_2 FILLER_10_699 ();
 sg13g2_fill_1 FILLER_10_701 ();
 sg13g2_fill_2 FILLER_10_711 ();
 sg13g2_fill_1 FILLER_10_713 ();
 sg13g2_fill_1 FILLER_10_735 ();
 sg13g2_fill_1 FILLER_10_741 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_fill_1 FILLER_10_785 ();
 sg13g2_decap_4 FILLER_10_791 ();
 sg13g2_fill_2 FILLER_10_803 ();
 sg13g2_decap_4 FILLER_10_811 ();
 sg13g2_fill_1 FILLER_10_815 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_fill_1 FILLER_10_851 ();
 sg13g2_decap_4 FILLER_10_861 ();
 sg13g2_fill_1 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_871 ();
 sg13g2_fill_1 FILLER_10_878 ();
 sg13g2_decap_4 FILLER_10_888 ();
 sg13g2_fill_2 FILLER_10_892 ();
 sg13g2_decap_8 FILLER_10_914 ();
 sg13g2_decap_8 FILLER_10_921 ();
 sg13g2_decap_8 FILLER_10_928 ();
 sg13g2_decap_8 FILLER_10_935 ();
 sg13g2_decap_8 FILLER_10_942 ();
 sg13g2_decap_8 FILLER_10_949 ();
 sg13g2_decap_8 FILLER_10_956 ();
 sg13g2_decap_8 FILLER_10_963 ();
 sg13g2_decap_8 FILLER_10_970 ();
 sg13g2_decap_8 FILLER_10_977 ();
 sg13g2_decap_8 FILLER_10_984 ();
 sg13g2_decap_8 FILLER_10_991 ();
 sg13g2_decap_8 FILLER_10_998 ();
 sg13g2_decap_8 FILLER_10_1005 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_decap_8 FILLER_10_1026 ();
 sg13g2_decap_8 FILLER_10_1033 ();
 sg13g2_decap_8 FILLER_10_1040 ();
 sg13g2_decap_8 FILLER_10_1047 ();
 sg13g2_decap_8 FILLER_10_1054 ();
 sg13g2_decap_8 FILLER_10_1061 ();
 sg13g2_decap_8 FILLER_10_1068 ();
 sg13g2_decap_8 FILLER_10_1075 ();
 sg13g2_decap_8 FILLER_10_1082 ();
 sg13g2_decap_8 FILLER_10_1089 ();
 sg13g2_decap_8 FILLER_10_1096 ();
 sg13g2_decap_8 FILLER_10_1103 ();
 sg13g2_decap_8 FILLER_10_1110 ();
 sg13g2_decap_8 FILLER_10_1117 ();
 sg13g2_decap_8 FILLER_10_1124 ();
 sg13g2_decap_8 FILLER_10_1131 ();
 sg13g2_decap_8 FILLER_10_1138 ();
 sg13g2_decap_8 FILLER_10_1145 ();
 sg13g2_decap_8 FILLER_10_1152 ();
 sg13g2_decap_8 FILLER_10_1159 ();
 sg13g2_decap_8 FILLER_10_1166 ();
 sg13g2_decap_8 FILLER_10_1173 ();
 sg13g2_decap_8 FILLER_10_1180 ();
 sg13g2_decap_8 FILLER_10_1187 ();
 sg13g2_decap_8 FILLER_10_1194 ();
 sg13g2_decap_8 FILLER_10_1201 ();
 sg13g2_decap_8 FILLER_10_1208 ();
 sg13g2_decap_8 FILLER_10_1215 ();
 sg13g2_decap_8 FILLER_10_1222 ();
 sg13g2_decap_8 FILLER_10_1229 ();
 sg13g2_decap_8 FILLER_10_1236 ();
 sg13g2_decap_8 FILLER_10_1243 ();
 sg13g2_decap_8 FILLER_10_1250 ();
 sg13g2_decap_8 FILLER_10_1257 ();
 sg13g2_decap_8 FILLER_10_1264 ();
 sg13g2_decap_8 FILLER_10_1271 ();
 sg13g2_decap_8 FILLER_10_1278 ();
 sg13g2_decap_8 FILLER_10_1285 ();
 sg13g2_decap_8 FILLER_10_1292 ();
 sg13g2_decap_8 FILLER_10_1299 ();
 sg13g2_decap_8 FILLER_10_1306 ();
 sg13g2_fill_2 FILLER_10_1313 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_4 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_214 ();
 sg13g2_fill_2 FILLER_11_276 ();
 sg13g2_fill_1 FILLER_11_278 ();
 sg13g2_fill_2 FILLER_11_318 ();
 sg13g2_fill_1 FILLER_11_320 ();
 sg13g2_fill_2 FILLER_11_329 ();
 sg13g2_fill_1 FILLER_11_331 ();
 sg13g2_fill_1 FILLER_11_372 ();
 sg13g2_fill_1 FILLER_11_400 ();
 sg13g2_decap_4 FILLER_11_426 ();
 sg13g2_decap_8 FILLER_11_439 ();
 sg13g2_fill_2 FILLER_11_446 ();
 sg13g2_fill_1 FILLER_11_448 ();
 sg13g2_fill_2 FILLER_11_467 ();
 sg13g2_decap_4 FILLER_11_474 ();
 sg13g2_fill_2 FILLER_11_483 ();
 sg13g2_fill_1 FILLER_11_498 ();
 sg13g2_decap_4 FILLER_11_512 ();
 sg13g2_decap_4 FILLER_11_534 ();
 sg13g2_decap_8 FILLER_11_564 ();
 sg13g2_decap_8 FILLER_11_571 ();
 sg13g2_decap_4 FILLER_11_645 ();
 sg13g2_fill_2 FILLER_11_649 ();
 sg13g2_fill_1 FILLER_11_671 ();
 sg13g2_fill_1 FILLER_11_682 ();
 sg13g2_fill_2 FILLER_11_776 ();
 sg13g2_decap_8 FILLER_11_786 ();
 sg13g2_fill_2 FILLER_11_793 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_fill_2 FILLER_11_805 ();
 sg13g2_fill_1 FILLER_11_807 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_fill_1 FILLER_11_879 ();
 sg13g2_fill_1 FILLER_11_891 ();
 sg13g2_fill_2 FILLER_11_897 ();
 sg13g2_decap_8 FILLER_11_909 ();
 sg13g2_decap_8 FILLER_11_916 ();
 sg13g2_decap_4 FILLER_11_923 ();
 sg13g2_fill_2 FILLER_11_927 ();
 sg13g2_fill_1 FILLER_11_937 ();
 sg13g2_decap_4 FILLER_11_968 ();
 sg13g2_decap_8 FILLER_11_977 ();
 sg13g2_fill_1 FILLER_11_984 ();
 sg13g2_decap_8 FILLER_11_993 ();
 sg13g2_decap_8 FILLER_11_1000 ();
 sg13g2_decap_8 FILLER_11_1007 ();
 sg13g2_decap_8 FILLER_11_1014 ();
 sg13g2_decap_8 FILLER_11_1021 ();
 sg13g2_decap_8 FILLER_11_1028 ();
 sg13g2_decap_8 FILLER_11_1035 ();
 sg13g2_decap_8 FILLER_11_1042 ();
 sg13g2_decap_8 FILLER_11_1049 ();
 sg13g2_decap_8 FILLER_11_1056 ();
 sg13g2_decap_8 FILLER_11_1063 ();
 sg13g2_decap_8 FILLER_11_1070 ();
 sg13g2_decap_8 FILLER_11_1077 ();
 sg13g2_decap_8 FILLER_11_1084 ();
 sg13g2_decap_8 FILLER_11_1091 ();
 sg13g2_decap_8 FILLER_11_1098 ();
 sg13g2_decap_8 FILLER_11_1105 ();
 sg13g2_decap_8 FILLER_11_1112 ();
 sg13g2_decap_8 FILLER_11_1119 ();
 sg13g2_decap_8 FILLER_11_1126 ();
 sg13g2_decap_8 FILLER_11_1133 ();
 sg13g2_decap_8 FILLER_11_1140 ();
 sg13g2_decap_8 FILLER_11_1147 ();
 sg13g2_decap_8 FILLER_11_1154 ();
 sg13g2_decap_8 FILLER_11_1161 ();
 sg13g2_decap_8 FILLER_11_1168 ();
 sg13g2_decap_8 FILLER_11_1175 ();
 sg13g2_decap_8 FILLER_11_1182 ();
 sg13g2_decap_8 FILLER_11_1189 ();
 sg13g2_decap_8 FILLER_11_1196 ();
 sg13g2_decap_8 FILLER_11_1203 ();
 sg13g2_decap_8 FILLER_11_1210 ();
 sg13g2_decap_8 FILLER_11_1217 ();
 sg13g2_decap_8 FILLER_11_1224 ();
 sg13g2_decap_8 FILLER_11_1231 ();
 sg13g2_decap_8 FILLER_11_1238 ();
 sg13g2_decap_8 FILLER_11_1245 ();
 sg13g2_decap_8 FILLER_11_1252 ();
 sg13g2_decap_8 FILLER_11_1259 ();
 sg13g2_decap_8 FILLER_11_1266 ();
 sg13g2_decap_8 FILLER_11_1273 ();
 sg13g2_decap_8 FILLER_11_1280 ();
 sg13g2_decap_8 FILLER_11_1287 ();
 sg13g2_decap_8 FILLER_11_1294 ();
 sg13g2_decap_8 FILLER_11_1301 ();
 sg13g2_decap_8 FILLER_11_1308 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_4 FILLER_12_210 ();
 sg13g2_fill_2 FILLER_12_214 ();
 sg13g2_fill_2 FILLER_12_252 ();
 sg13g2_fill_1 FILLER_12_254 ();
 sg13g2_fill_2 FILLER_12_259 ();
 sg13g2_fill_1 FILLER_12_265 ();
 sg13g2_fill_2 FILLER_12_275 ();
 sg13g2_fill_2 FILLER_12_282 ();
 sg13g2_fill_2 FILLER_12_293 ();
 sg13g2_fill_1 FILLER_12_295 ();
 sg13g2_fill_2 FILLER_12_348 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_2 FILLER_12_423 ();
 sg13g2_fill_1 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_449 ();
 sg13g2_fill_1 FILLER_12_484 ();
 sg13g2_fill_2 FILLER_12_511 ();
 sg13g2_fill_1 FILLER_12_513 ();
 sg13g2_decap_8 FILLER_12_540 ();
 sg13g2_decap_4 FILLER_12_547 ();
 sg13g2_fill_1 FILLER_12_551 ();
 sg13g2_decap_8 FILLER_12_569 ();
 sg13g2_fill_2 FILLER_12_576 ();
 sg13g2_fill_1 FILLER_12_582 ();
 sg13g2_fill_2 FILLER_12_587 ();
 sg13g2_decap_4 FILLER_12_615 ();
 sg13g2_fill_1 FILLER_12_619 ();
 sg13g2_decap_8 FILLER_12_624 ();
 sg13g2_decap_8 FILLER_12_631 ();
 sg13g2_decap_4 FILLER_12_638 ();
 sg13g2_decap_4 FILLER_12_655 ();
 sg13g2_fill_2 FILLER_12_680 ();
 sg13g2_decap_8 FILLER_12_692 ();
 sg13g2_fill_2 FILLER_12_699 ();
 sg13g2_fill_2 FILLER_12_709 ();
 sg13g2_decap_8 FILLER_12_720 ();
 sg13g2_decap_8 FILLER_12_727 ();
 sg13g2_decap_8 FILLER_12_734 ();
 sg13g2_fill_2 FILLER_12_745 ();
 sg13g2_fill_1 FILLER_12_747 ();
 sg13g2_fill_2 FILLER_12_753 ();
 sg13g2_fill_1 FILLER_12_771 ();
 sg13g2_fill_1 FILLER_12_781 ();
 sg13g2_fill_2 FILLER_12_793 ();
 sg13g2_fill_2 FILLER_12_863 ();
 sg13g2_decap_8 FILLER_12_874 ();
 sg13g2_fill_1 FILLER_12_881 ();
 sg13g2_decap_8 FILLER_12_913 ();
 sg13g2_decap_8 FILLER_12_920 ();
 sg13g2_decap_8 FILLER_12_927 ();
 sg13g2_decap_8 FILLER_12_934 ();
 sg13g2_decap_4 FILLER_12_941 ();
 sg13g2_fill_2 FILLER_12_953 ();
 sg13g2_decap_8 FILLER_12_1000 ();
 sg13g2_decap_8 FILLER_12_1007 ();
 sg13g2_decap_8 FILLER_12_1014 ();
 sg13g2_decap_8 FILLER_12_1021 ();
 sg13g2_decap_8 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_12_1035 ();
 sg13g2_decap_8 FILLER_12_1042 ();
 sg13g2_decap_8 FILLER_12_1049 ();
 sg13g2_decap_8 FILLER_12_1056 ();
 sg13g2_decap_8 FILLER_12_1063 ();
 sg13g2_decap_8 FILLER_12_1070 ();
 sg13g2_decap_8 FILLER_12_1077 ();
 sg13g2_decap_8 FILLER_12_1084 ();
 sg13g2_decap_8 FILLER_12_1091 ();
 sg13g2_decap_8 FILLER_12_1098 ();
 sg13g2_decap_8 FILLER_12_1105 ();
 sg13g2_decap_8 FILLER_12_1112 ();
 sg13g2_decap_8 FILLER_12_1119 ();
 sg13g2_decap_8 FILLER_12_1126 ();
 sg13g2_decap_8 FILLER_12_1133 ();
 sg13g2_decap_8 FILLER_12_1140 ();
 sg13g2_decap_8 FILLER_12_1147 ();
 sg13g2_decap_8 FILLER_12_1154 ();
 sg13g2_decap_8 FILLER_12_1161 ();
 sg13g2_decap_8 FILLER_12_1168 ();
 sg13g2_decap_8 FILLER_12_1175 ();
 sg13g2_decap_8 FILLER_12_1182 ();
 sg13g2_decap_8 FILLER_12_1189 ();
 sg13g2_decap_8 FILLER_12_1196 ();
 sg13g2_decap_8 FILLER_12_1203 ();
 sg13g2_decap_8 FILLER_12_1210 ();
 sg13g2_decap_8 FILLER_12_1217 ();
 sg13g2_decap_8 FILLER_12_1224 ();
 sg13g2_decap_8 FILLER_12_1231 ();
 sg13g2_decap_8 FILLER_12_1238 ();
 sg13g2_decap_8 FILLER_12_1245 ();
 sg13g2_decap_8 FILLER_12_1252 ();
 sg13g2_decap_8 FILLER_12_1259 ();
 sg13g2_decap_8 FILLER_12_1266 ();
 sg13g2_decap_8 FILLER_12_1273 ();
 sg13g2_decap_8 FILLER_12_1280 ();
 sg13g2_decap_8 FILLER_12_1287 ();
 sg13g2_decap_8 FILLER_12_1294 ();
 sg13g2_decap_8 FILLER_12_1301 ();
 sg13g2_decap_8 FILLER_12_1308 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_4 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_179 ();
 sg13g2_decap_4 FILLER_13_184 ();
 sg13g2_fill_1 FILLER_13_188 ();
 sg13g2_decap_8 FILLER_13_198 ();
 sg13g2_decap_4 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_336 ();
 sg13g2_fill_2 FILLER_13_364 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_fill_2 FILLER_13_376 ();
 sg13g2_fill_2 FILLER_13_392 ();
 sg13g2_fill_1 FILLER_13_403 ();
 sg13g2_fill_1 FILLER_13_461 ();
 sg13g2_decap_8 FILLER_13_479 ();
 sg13g2_decap_4 FILLER_13_486 ();
 sg13g2_fill_2 FILLER_13_490 ();
 sg13g2_fill_1 FILLER_13_504 ();
 sg13g2_fill_2 FILLER_13_599 ();
 sg13g2_fill_1 FILLER_13_601 ();
 sg13g2_fill_1 FILLER_13_606 ();
 sg13g2_fill_2 FILLER_13_633 ();
 sg13g2_fill_2 FILLER_13_646 ();
 sg13g2_decap_4 FILLER_13_664 ();
 sg13g2_fill_2 FILLER_13_700 ();
 sg13g2_fill_1 FILLER_13_702 ();
 sg13g2_fill_2 FILLER_13_723 ();
 sg13g2_fill_1 FILLER_13_733 ();
 sg13g2_fill_2 FILLER_13_743 ();
 sg13g2_fill_1 FILLER_13_745 ();
 sg13g2_fill_2 FILLER_13_751 ();
 sg13g2_fill_1 FILLER_13_753 ();
 sg13g2_decap_4 FILLER_13_762 ();
 sg13g2_fill_1 FILLER_13_766 ();
 sg13g2_fill_2 FILLER_13_772 ();
 sg13g2_decap_4 FILLER_13_790 ();
 sg13g2_fill_1 FILLER_13_794 ();
 sg13g2_decap_8 FILLER_13_816 ();
 sg13g2_decap_8 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_8 FILLER_13_844 ();
 sg13g2_decap_4 FILLER_13_851 ();
 sg13g2_fill_1 FILLER_13_855 ();
 sg13g2_fill_2 FILLER_13_865 ();
 sg13g2_fill_1 FILLER_13_867 ();
 sg13g2_fill_1 FILLER_13_881 ();
 sg13g2_decap_8 FILLER_13_927 ();
 sg13g2_decap_4 FILLER_13_934 ();
 sg13g2_fill_2 FILLER_13_977 ();
 sg13g2_fill_1 FILLER_13_979 ();
 sg13g2_decap_8 FILLER_13_1014 ();
 sg13g2_decap_8 FILLER_13_1021 ();
 sg13g2_decap_8 FILLER_13_1028 ();
 sg13g2_decap_8 FILLER_13_1035 ();
 sg13g2_decap_8 FILLER_13_1042 ();
 sg13g2_decap_8 FILLER_13_1049 ();
 sg13g2_decap_8 FILLER_13_1056 ();
 sg13g2_decap_8 FILLER_13_1063 ();
 sg13g2_decap_8 FILLER_13_1070 ();
 sg13g2_decap_8 FILLER_13_1077 ();
 sg13g2_decap_8 FILLER_13_1084 ();
 sg13g2_decap_8 FILLER_13_1091 ();
 sg13g2_decap_8 FILLER_13_1098 ();
 sg13g2_decap_8 FILLER_13_1105 ();
 sg13g2_decap_8 FILLER_13_1112 ();
 sg13g2_decap_8 FILLER_13_1119 ();
 sg13g2_decap_8 FILLER_13_1126 ();
 sg13g2_decap_8 FILLER_13_1133 ();
 sg13g2_decap_8 FILLER_13_1140 ();
 sg13g2_decap_8 FILLER_13_1147 ();
 sg13g2_decap_8 FILLER_13_1154 ();
 sg13g2_decap_8 FILLER_13_1161 ();
 sg13g2_decap_8 FILLER_13_1168 ();
 sg13g2_decap_8 FILLER_13_1175 ();
 sg13g2_decap_8 FILLER_13_1182 ();
 sg13g2_decap_8 FILLER_13_1189 ();
 sg13g2_decap_8 FILLER_13_1196 ();
 sg13g2_decap_8 FILLER_13_1203 ();
 sg13g2_decap_8 FILLER_13_1210 ();
 sg13g2_decap_8 FILLER_13_1217 ();
 sg13g2_decap_8 FILLER_13_1224 ();
 sg13g2_decap_8 FILLER_13_1231 ();
 sg13g2_decap_8 FILLER_13_1238 ();
 sg13g2_decap_8 FILLER_13_1245 ();
 sg13g2_decap_8 FILLER_13_1252 ();
 sg13g2_decap_8 FILLER_13_1259 ();
 sg13g2_decap_8 FILLER_13_1266 ();
 sg13g2_decap_8 FILLER_13_1273 ();
 sg13g2_decap_8 FILLER_13_1280 ();
 sg13g2_decap_8 FILLER_13_1287 ();
 sg13g2_decap_8 FILLER_13_1294 ();
 sg13g2_decap_8 FILLER_13_1301 ();
 sg13g2_decap_8 FILLER_13_1308 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_170 ();
 sg13g2_fill_2 FILLER_14_237 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_250 ();
 sg13g2_fill_1 FILLER_14_259 ();
 sg13g2_fill_1 FILLER_14_274 ();
 sg13g2_fill_1 FILLER_14_283 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_fill_2 FILLER_14_352 ();
 sg13g2_fill_1 FILLER_14_354 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_fill_2 FILLER_14_392 ();
 sg13g2_fill_2 FILLER_14_452 ();
 sg13g2_fill_2 FILLER_14_459 ();
 sg13g2_fill_1 FILLER_14_461 ();
 sg13g2_fill_1 FILLER_14_488 ();
 sg13g2_fill_2 FILLER_14_530 ();
 sg13g2_fill_2 FILLER_14_553 ();
 sg13g2_fill_1 FILLER_14_555 ();
 sg13g2_fill_2 FILLER_14_565 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_4 FILLER_14_595 ();
 sg13g2_fill_1 FILLER_14_599 ();
 sg13g2_decap_8 FILLER_14_604 ();
 sg13g2_fill_1 FILLER_14_611 ();
 sg13g2_fill_1 FILLER_14_642 ();
 sg13g2_decap_4 FILLER_14_661 ();
 sg13g2_fill_2 FILLER_14_665 ();
 sg13g2_fill_1 FILLER_14_697 ();
 sg13g2_decap_4 FILLER_14_703 ();
 sg13g2_fill_1 FILLER_14_707 ();
 sg13g2_fill_2 FILLER_14_713 ();
 sg13g2_decap_4 FILLER_14_759 ();
 sg13g2_fill_1 FILLER_14_763 ();
 sg13g2_fill_2 FILLER_14_799 ();
 sg13g2_fill_2 FILLER_14_806 ();
 sg13g2_decap_8 FILLER_14_818 ();
 sg13g2_fill_2 FILLER_14_825 ();
 sg13g2_fill_1 FILLER_14_827 ();
 sg13g2_fill_2 FILLER_14_840 ();
 sg13g2_decap_4 FILLER_14_852 ();
 sg13g2_fill_2 FILLER_14_856 ();
 sg13g2_decap_8 FILLER_14_867 ();
 sg13g2_fill_2 FILLER_14_874 ();
 sg13g2_fill_1 FILLER_14_876 ();
 sg13g2_decap_4 FILLER_14_881 ();
 sg13g2_fill_1 FILLER_14_885 ();
 sg13g2_decap_8 FILLER_14_894 ();
 sg13g2_fill_1 FILLER_14_901 ();
 sg13g2_decap_8 FILLER_14_921 ();
 sg13g2_decap_8 FILLER_14_928 ();
 sg13g2_decap_8 FILLER_14_935 ();
 sg13g2_decap_8 FILLER_14_942 ();
 sg13g2_fill_2 FILLER_14_949 ();
 sg13g2_fill_1 FILLER_14_951 ();
 sg13g2_fill_1 FILLER_14_970 ();
 sg13g2_decap_8 FILLER_14_1030 ();
 sg13g2_decap_8 FILLER_14_1037 ();
 sg13g2_decap_8 FILLER_14_1044 ();
 sg13g2_decap_8 FILLER_14_1051 ();
 sg13g2_decap_8 FILLER_14_1058 ();
 sg13g2_decap_8 FILLER_14_1065 ();
 sg13g2_decap_8 FILLER_14_1072 ();
 sg13g2_decap_8 FILLER_14_1079 ();
 sg13g2_decap_8 FILLER_14_1086 ();
 sg13g2_decap_8 FILLER_14_1093 ();
 sg13g2_decap_8 FILLER_14_1100 ();
 sg13g2_decap_8 FILLER_14_1107 ();
 sg13g2_decap_8 FILLER_14_1114 ();
 sg13g2_decap_8 FILLER_14_1121 ();
 sg13g2_decap_8 FILLER_14_1128 ();
 sg13g2_decap_8 FILLER_14_1135 ();
 sg13g2_decap_8 FILLER_14_1142 ();
 sg13g2_decap_8 FILLER_14_1149 ();
 sg13g2_decap_8 FILLER_14_1156 ();
 sg13g2_decap_8 FILLER_14_1163 ();
 sg13g2_decap_8 FILLER_14_1170 ();
 sg13g2_decap_8 FILLER_14_1177 ();
 sg13g2_decap_8 FILLER_14_1184 ();
 sg13g2_decap_8 FILLER_14_1191 ();
 sg13g2_decap_8 FILLER_14_1198 ();
 sg13g2_decap_8 FILLER_14_1205 ();
 sg13g2_decap_8 FILLER_14_1212 ();
 sg13g2_decap_8 FILLER_14_1219 ();
 sg13g2_decap_8 FILLER_14_1226 ();
 sg13g2_decap_8 FILLER_14_1233 ();
 sg13g2_decap_8 FILLER_14_1240 ();
 sg13g2_decap_8 FILLER_14_1247 ();
 sg13g2_decap_8 FILLER_14_1254 ();
 sg13g2_decap_8 FILLER_14_1261 ();
 sg13g2_decap_8 FILLER_14_1268 ();
 sg13g2_decap_8 FILLER_14_1275 ();
 sg13g2_decap_8 FILLER_14_1282 ();
 sg13g2_decap_8 FILLER_14_1289 ();
 sg13g2_decap_8 FILLER_14_1296 ();
 sg13g2_decap_8 FILLER_14_1303 ();
 sg13g2_decap_4 FILLER_14_1310 ();
 sg13g2_fill_1 FILLER_14_1314 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_166 ();
 sg13g2_decap_4 FILLER_15_181 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_333 ();
 sg13g2_decap_4 FILLER_15_340 ();
 sg13g2_fill_1 FILLER_15_344 ();
 sg13g2_decap_4 FILLER_15_354 ();
 sg13g2_fill_2 FILLER_15_358 ();
 sg13g2_fill_1 FILLER_15_386 ();
 sg13g2_fill_2 FILLER_15_396 ();
 sg13g2_fill_1 FILLER_15_398 ();
 sg13g2_fill_1 FILLER_15_418 ();
 sg13g2_fill_2 FILLER_15_468 ();
 sg13g2_fill_1 FILLER_15_470 ();
 sg13g2_fill_2 FILLER_15_480 ();
 sg13g2_decap_4 FILLER_15_496 ();
 sg13g2_fill_2 FILLER_15_528 ();
 sg13g2_fill_1 FILLER_15_530 ();
 sg13g2_fill_2 FILLER_15_557 ();
 sg13g2_fill_1 FILLER_15_559 ();
 sg13g2_fill_2 FILLER_15_608 ();
 sg13g2_decap_8 FILLER_15_614 ();
 sg13g2_decap_4 FILLER_15_621 ();
 sg13g2_fill_2 FILLER_15_625 ();
 sg13g2_decap_8 FILLER_15_631 ();
 sg13g2_fill_1 FILLER_15_638 ();
 sg13g2_decap_8 FILLER_15_647 ();
 sg13g2_fill_2 FILLER_15_659 ();
 sg13g2_fill_1 FILLER_15_661 ();
 sg13g2_decap_4 FILLER_15_676 ();
 sg13g2_fill_2 FILLER_15_680 ();
 sg13g2_fill_2 FILLER_15_702 ();
 sg13g2_decap_4 FILLER_15_719 ();
 sg13g2_fill_2 FILLER_15_723 ();
 sg13g2_decap_8 FILLER_15_730 ();
 sg13g2_fill_2 FILLER_15_737 ();
 sg13g2_fill_1 FILLER_15_739 ();
 sg13g2_fill_1 FILLER_15_744 ();
 sg13g2_fill_1 FILLER_15_758 ();
 sg13g2_decap_8 FILLER_15_764 ();
 sg13g2_decap_4 FILLER_15_779 ();
 sg13g2_fill_1 FILLER_15_783 ();
 sg13g2_fill_1 FILLER_15_789 ();
 sg13g2_fill_2 FILLER_15_804 ();
 sg13g2_fill_1 FILLER_15_806 ();
 sg13g2_fill_2 FILLER_15_874 ();
 sg13g2_fill_2 FILLER_15_889 ();
 sg13g2_fill_1 FILLER_15_891 ();
 sg13g2_fill_1 FILLER_15_901 ();
 sg13g2_fill_2 FILLER_15_907 ();
 sg13g2_decap_8 FILLER_15_924 ();
 sg13g2_decap_8 FILLER_15_931 ();
 sg13g2_decap_8 FILLER_15_938 ();
 sg13g2_fill_2 FILLER_15_945 ();
 sg13g2_fill_1 FILLER_15_947 ();
 sg13g2_fill_1 FILLER_15_1004 ();
 sg13g2_decap_8 FILLER_15_1036 ();
 sg13g2_decap_8 FILLER_15_1043 ();
 sg13g2_decap_8 FILLER_15_1050 ();
 sg13g2_decap_8 FILLER_15_1057 ();
 sg13g2_decap_8 FILLER_15_1064 ();
 sg13g2_decap_8 FILLER_15_1071 ();
 sg13g2_decap_8 FILLER_15_1078 ();
 sg13g2_decap_8 FILLER_15_1085 ();
 sg13g2_decap_8 FILLER_15_1092 ();
 sg13g2_decap_8 FILLER_15_1099 ();
 sg13g2_decap_8 FILLER_15_1106 ();
 sg13g2_decap_8 FILLER_15_1113 ();
 sg13g2_decap_8 FILLER_15_1120 ();
 sg13g2_decap_8 FILLER_15_1127 ();
 sg13g2_decap_8 FILLER_15_1134 ();
 sg13g2_decap_8 FILLER_15_1141 ();
 sg13g2_decap_8 FILLER_15_1148 ();
 sg13g2_decap_8 FILLER_15_1155 ();
 sg13g2_decap_8 FILLER_15_1162 ();
 sg13g2_decap_8 FILLER_15_1169 ();
 sg13g2_decap_8 FILLER_15_1176 ();
 sg13g2_decap_8 FILLER_15_1183 ();
 sg13g2_decap_8 FILLER_15_1190 ();
 sg13g2_decap_8 FILLER_15_1197 ();
 sg13g2_decap_8 FILLER_15_1204 ();
 sg13g2_decap_8 FILLER_15_1211 ();
 sg13g2_decap_8 FILLER_15_1218 ();
 sg13g2_decap_8 FILLER_15_1225 ();
 sg13g2_decap_8 FILLER_15_1232 ();
 sg13g2_decap_8 FILLER_15_1239 ();
 sg13g2_decap_8 FILLER_15_1246 ();
 sg13g2_decap_8 FILLER_15_1253 ();
 sg13g2_decap_8 FILLER_15_1260 ();
 sg13g2_decap_8 FILLER_15_1267 ();
 sg13g2_decap_8 FILLER_15_1274 ();
 sg13g2_decap_8 FILLER_15_1281 ();
 sg13g2_decap_8 FILLER_15_1288 ();
 sg13g2_decap_8 FILLER_15_1295 ();
 sg13g2_decap_8 FILLER_15_1302 ();
 sg13g2_decap_4 FILLER_15_1309 ();
 sg13g2_fill_2 FILLER_15_1313 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_4 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_219 ();
 sg13g2_fill_2 FILLER_16_241 ();
 sg13g2_fill_1 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_fill_2 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_333 ();
 sg13g2_fill_2 FILLER_16_357 ();
 sg13g2_fill_1 FILLER_16_359 ();
 sg13g2_fill_1 FILLER_16_386 ();
 sg13g2_fill_2 FILLER_16_413 ();
 sg13g2_fill_2 FILLER_16_429 ();
 sg13g2_fill_1 FILLER_16_431 ();
 sg13g2_fill_2 FILLER_16_454 ();
 sg13g2_fill_1 FILLER_16_456 ();
 sg13g2_fill_1 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_decap_4 FILLER_16_506 ();
 sg13g2_fill_2 FILLER_16_510 ();
 sg13g2_fill_2 FILLER_16_517 ();
 sg13g2_fill_1 FILLER_16_519 ();
 sg13g2_fill_2 FILLER_16_525 ();
 sg13g2_fill_1 FILLER_16_531 ();
 sg13g2_fill_2 FILLER_16_536 ();
 sg13g2_fill_2 FILLER_16_547 ();
 sg13g2_fill_1 FILLER_16_575 ();
 sg13g2_fill_2 FILLER_16_616 ();
 sg13g2_decap_4 FILLER_16_647 ();
 sg13g2_decap_8 FILLER_16_662 ();
 sg13g2_decap_4 FILLER_16_669 ();
 sg13g2_fill_2 FILLER_16_677 ();
 sg13g2_fill_1 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_697 ();
 sg13g2_fill_2 FILLER_16_709 ();
 sg13g2_fill_1 FILLER_16_722 ();
 sg13g2_fill_1 FILLER_16_733 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_fill_1 FILLER_16_751 ();
 sg13g2_fill_2 FILLER_16_765 ();
 sg13g2_fill_1 FILLER_16_767 ();
 sg13g2_fill_2 FILLER_16_781 ();
 sg13g2_fill_1 FILLER_16_783 ();
 sg13g2_fill_1 FILLER_16_808 ();
 sg13g2_fill_1 FILLER_16_819 ();
 sg13g2_decap_4 FILLER_16_825 ();
 sg13g2_fill_1 FILLER_16_829 ();
 sg13g2_fill_1 FILLER_16_834 ();
 sg13g2_fill_2 FILLER_16_848 ();
 sg13g2_fill_1 FILLER_16_850 ();
 sg13g2_fill_2 FILLER_16_878 ();
 sg13g2_fill_1 FILLER_16_880 ();
 sg13g2_decap_4 FILLER_16_894 ();
 sg13g2_fill_2 FILLER_16_908 ();
 sg13g2_fill_2 FILLER_16_918 ();
 sg13g2_decap_8 FILLER_16_934 ();
 sg13g2_decap_8 FILLER_16_941 ();
 sg13g2_decap_8 FILLER_16_948 ();
 sg13g2_decap_4 FILLER_16_955 ();
 sg13g2_fill_2 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_1046 ();
 sg13g2_decap_8 FILLER_16_1053 ();
 sg13g2_decap_8 FILLER_16_1060 ();
 sg13g2_decap_8 FILLER_16_1067 ();
 sg13g2_decap_8 FILLER_16_1074 ();
 sg13g2_decap_8 FILLER_16_1081 ();
 sg13g2_decap_8 FILLER_16_1088 ();
 sg13g2_decap_8 FILLER_16_1095 ();
 sg13g2_decap_8 FILLER_16_1102 ();
 sg13g2_decap_8 FILLER_16_1109 ();
 sg13g2_decap_8 FILLER_16_1116 ();
 sg13g2_decap_8 FILLER_16_1123 ();
 sg13g2_decap_8 FILLER_16_1130 ();
 sg13g2_decap_8 FILLER_16_1137 ();
 sg13g2_decap_8 FILLER_16_1144 ();
 sg13g2_decap_8 FILLER_16_1151 ();
 sg13g2_decap_8 FILLER_16_1158 ();
 sg13g2_decap_8 FILLER_16_1165 ();
 sg13g2_decap_8 FILLER_16_1172 ();
 sg13g2_decap_8 FILLER_16_1179 ();
 sg13g2_decap_8 FILLER_16_1186 ();
 sg13g2_decap_8 FILLER_16_1193 ();
 sg13g2_decap_8 FILLER_16_1200 ();
 sg13g2_decap_8 FILLER_16_1207 ();
 sg13g2_decap_8 FILLER_16_1214 ();
 sg13g2_decap_8 FILLER_16_1221 ();
 sg13g2_decap_8 FILLER_16_1228 ();
 sg13g2_decap_8 FILLER_16_1235 ();
 sg13g2_decap_8 FILLER_16_1242 ();
 sg13g2_decap_8 FILLER_16_1249 ();
 sg13g2_decap_8 FILLER_16_1256 ();
 sg13g2_decap_8 FILLER_16_1263 ();
 sg13g2_decap_8 FILLER_16_1270 ();
 sg13g2_decap_8 FILLER_16_1277 ();
 sg13g2_decap_8 FILLER_16_1284 ();
 sg13g2_decap_8 FILLER_16_1291 ();
 sg13g2_decap_8 FILLER_16_1298 ();
 sg13g2_decap_8 FILLER_16_1305 ();
 sg13g2_fill_2 FILLER_16_1312 ();
 sg13g2_fill_1 FILLER_16_1314 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_135 ();
 sg13g2_fill_1 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_168 ();
 sg13g2_fill_1 FILLER_17_204 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_fill_2 FILLER_17_239 ();
 sg13g2_fill_1 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_fill_2 FILLER_17_274 ();
 sg13g2_fill_1 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_302 ();
 sg13g2_decap_4 FILLER_17_312 ();
 sg13g2_fill_2 FILLER_17_333 ();
 sg13g2_fill_1 FILLER_17_335 ();
 sg13g2_fill_2 FILLER_17_340 ();
 sg13g2_fill_2 FILLER_17_366 ();
 sg13g2_fill_1 FILLER_17_368 ();
 sg13g2_fill_2 FILLER_17_382 ();
 sg13g2_decap_4 FILLER_17_394 ();
 sg13g2_decap_4 FILLER_17_402 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_413 ();
 sg13g2_fill_1 FILLER_17_475 ();
 sg13g2_decap_8 FILLER_17_531 ();
 sg13g2_decap_4 FILLER_17_538 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_564 ();
 sg13g2_decap_8 FILLER_17_571 ();
 sg13g2_decap_8 FILLER_17_591 ();
 sg13g2_decap_4 FILLER_17_598 ();
 sg13g2_fill_1 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_640 ();
 sg13g2_fill_2 FILLER_17_647 ();
 sg13g2_fill_1 FILLER_17_649 ();
 sg13g2_decap_4 FILLER_17_661 ();
 sg13g2_fill_2 FILLER_17_665 ();
 sg13g2_fill_1 FILLER_17_691 ();
 sg13g2_fill_1 FILLER_17_702 ();
 sg13g2_decap_8 FILLER_17_717 ();
 sg13g2_decap_4 FILLER_17_754 ();
 sg13g2_decap_4 FILLER_17_768 ();
 sg13g2_decap_8 FILLER_17_780 ();
 sg13g2_decap_8 FILLER_17_787 ();
 sg13g2_decap_8 FILLER_17_799 ();
 sg13g2_fill_2 FILLER_17_821 ();
 sg13g2_fill_1 FILLER_17_823 ();
 sg13g2_decap_4 FILLER_17_868 ();
 sg13g2_fill_1 FILLER_17_872 ();
 sg13g2_fill_1 FILLER_17_882 ();
 sg13g2_decap_4 FILLER_17_888 ();
 sg13g2_fill_1 FILLER_17_892 ();
 sg13g2_fill_1 FILLER_17_910 ();
 sg13g2_fill_2 FILLER_17_915 ();
 sg13g2_fill_2 FILLER_17_927 ();
 sg13g2_fill_1 FILLER_17_929 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_fill_2 FILLER_17_945 ();
 sg13g2_fill_2 FILLER_17_990 ();
 sg13g2_fill_2 FILLER_17_1001 ();
 sg13g2_fill_1 FILLER_17_1003 ();
 sg13g2_decap_8 FILLER_17_1043 ();
 sg13g2_decap_8 FILLER_17_1050 ();
 sg13g2_decap_8 FILLER_17_1057 ();
 sg13g2_decap_8 FILLER_17_1064 ();
 sg13g2_decap_8 FILLER_17_1071 ();
 sg13g2_decap_8 FILLER_17_1078 ();
 sg13g2_decap_8 FILLER_17_1085 ();
 sg13g2_decap_8 FILLER_17_1092 ();
 sg13g2_decap_8 FILLER_17_1099 ();
 sg13g2_decap_8 FILLER_17_1106 ();
 sg13g2_decap_8 FILLER_17_1113 ();
 sg13g2_decap_8 FILLER_17_1120 ();
 sg13g2_decap_8 FILLER_17_1127 ();
 sg13g2_decap_8 FILLER_17_1134 ();
 sg13g2_decap_8 FILLER_17_1141 ();
 sg13g2_decap_8 FILLER_17_1148 ();
 sg13g2_decap_8 FILLER_17_1155 ();
 sg13g2_decap_8 FILLER_17_1162 ();
 sg13g2_decap_8 FILLER_17_1169 ();
 sg13g2_decap_8 FILLER_17_1176 ();
 sg13g2_decap_8 FILLER_17_1183 ();
 sg13g2_decap_8 FILLER_17_1190 ();
 sg13g2_decap_8 FILLER_17_1197 ();
 sg13g2_decap_8 FILLER_17_1204 ();
 sg13g2_decap_8 FILLER_17_1211 ();
 sg13g2_decap_8 FILLER_17_1218 ();
 sg13g2_decap_8 FILLER_17_1225 ();
 sg13g2_decap_8 FILLER_17_1232 ();
 sg13g2_decap_8 FILLER_17_1239 ();
 sg13g2_decap_8 FILLER_17_1246 ();
 sg13g2_decap_8 FILLER_17_1253 ();
 sg13g2_decap_8 FILLER_17_1260 ();
 sg13g2_decap_8 FILLER_17_1267 ();
 sg13g2_decap_8 FILLER_17_1274 ();
 sg13g2_decap_8 FILLER_17_1281 ();
 sg13g2_decap_8 FILLER_17_1288 ();
 sg13g2_decap_8 FILLER_17_1295 ();
 sg13g2_decap_8 FILLER_17_1302 ();
 sg13g2_decap_4 FILLER_17_1309 ();
 sg13g2_fill_2 FILLER_17_1313 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_126 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_2 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_fill_2 FILLER_18_219 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_4 FILLER_18_402 ();
 sg13g2_decap_4 FILLER_18_412 ();
 sg13g2_fill_1 FILLER_18_416 ();
 sg13g2_fill_1 FILLER_18_422 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_decap_8 FILLER_18_438 ();
 sg13g2_decap_4 FILLER_18_445 ();
 sg13g2_fill_1 FILLER_18_449 ();
 sg13g2_fill_1 FILLER_18_459 ();
 sg13g2_fill_1 FILLER_18_490 ();
 sg13g2_fill_1 FILLER_18_500 ();
 sg13g2_fill_1 FILLER_18_505 ();
 sg13g2_decap_8 FILLER_18_524 ();
 sg13g2_decap_4 FILLER_18_531 ();
 sg13g2_fill_1 FILLER_18_535 ();
 sg13g2_decap_4 FILLER_18_576 ();
 sg13g2_decap_4 FILLER_18_606 ();
 sg13g2_decap_4 FILLER_18_614 ();
 sg13g2_decap_4 FILLER_18_622 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_fill_1 FILLER_18_651 ();
 sg13g2_decap_4 FILLER_18_657 ();
 sg13g2_fill_1 FILLER_18_661 ();
 sg13g2_fill_1 FILLER_18_670 ();
 sg13g2_fill_2 FILLER_18_675 ();
 sg13g2_fill_1 FILLER_18_677 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_fill_1 FILLER_18_689 ();
 sg13g2_decap_8 FILLER_18_704 ();
 sg13g2_fill_2 FILLER_18_711 ();
 sg13g2_fill_2 FILLER_18_736 ();
 sg13g2_fill_1 FILLER_18_738 ();
 sg13g2_fill_1 FILLER_18_744 ();
 sg13g2_decap_8 FILLER_18_767 ();
 sg13g2_fill_1 FILLER_18_792 ();
 sg13g2_decap_8 FILLER_18_806 ();
 sg13g2_decap_4 FILLER_18_813 ();
 sg13g2_decap_8 FILLER_18_831 ();
 sg13g2_decap_4 FILLER_18_847 ();
 sg13g2_fill_1 FILLER_18_866 ();
 sg13g2_fill_2 FILLER_18_872 ();
 sg13g2_fill_1 FILLER_18_874 ();
 sg13g2_decap_8 FILLER_18_885 ();
 sg13g2_decap_4 FILLER_18_892 ();
 sg13g2_fill_2 FILLER_18_896 ();
 sg13g2_decap_4 FILLER_18_903 ();
 sg13g2_fill_2 FILLER_18_907 ();
 sg13g2_fill_1 FILLER_18_926 ();
 sg13g2_decap_8 FILLER_18_945 ();
 sg13g2_fill_2 FILLER_18_952 ();
 sg13g2_fill_1 FILLER_18_954 ();
 sg13g2_fill_2 FILLER_18_959 ();
 sg13g2_fill_2 FILLER_18_974 ();
 sg13g2_fill_1 FILLER_18_999 ();
 sg13g2_fill_1 FILLER_18_1016 ();
 sg13g2_fill_2 FILLER_18_1026 ();
 sg13g2_decap_8 FILLER_18_1051 ();
 sg13g2_decap_8 FILLER_18_1058 ();
 sg13g2_decap_8 FILLER_18_1065 ();
 sg13g2_decap_8 FILLER_18_1072 ();
 sg13g2_decap_8 FILLER_18_1079 ();
 sg13g2_decap_8 FILLER_18_1086 ();
 sg13g2_decap_8 FILLER_18_1093 ();
 sg13g2_decap_8 FILLER_18_1100 ();
 sg13g2_decap_8 FILLER_18_1107 ();
 sg13g2_decap_8 FILLER_18_1114 ();
 sg13g2_decap_8 FILLER_18_1121 ();
 sg13g2_decap_8 FILLER_18_1128 ();
 sg13g2_decap_8 FILLER_18_1135 ();
 sg13g2_decap_8 FILLER_18_1142 ();
 sg13g2_decap_8 FILLER_18_1149 ();
 sg13g2_decap_8 FILLER_18_1156 ();
 sg13g2_decap_8 FILLER_18_1163 ();
 sg13g2_decap_8 FILLER_18_1170 ();
 sg13g2_decap_8 FILLER_18_1177 ();
 sg13g2_decap_8 FILLER_18_1184 ();
 sg13g2_decap_8 FILLER_18_1191 ();
 sg13g2_decap_8 FILLER_18_1198 ();
 sg13g2_decap_8 FILLER_18_1205 ();
 sg13g2_decap_8 FILLER_18_1212 ();
 sg13g2_decap_8 FILLER_18_1219 ();
 sg13g2_decap_8 FILLER_18_1226 ();
 sg13g2_decap_8 FILLER_18_1233 ();
 sg13g2_decap_8 FILLER_18_1240 ();
 sg13g2_decap_8 FILLER_18_1247 ();
 sg13g2_decap_8 FILLER_18_1254 ();
 sg13g2_decap_8 FILLER_18_1261 ();
 sg13g2_decap_8 FILLER_18_1268 ();
 sg13g2_decap_8 FILLER_18_1275 ();
 sg13g2_decap_8 FILLER_18_1282 ();
 sg13g2_decap_8 FILLER_18_1289 ();
 sg13g2_decap_8 FILLER_18_1296 ();
 sg13g2_decap_8 FILLER_18_1303 ();
 sg13g2_decap_4 FILLER_18_1310 ();
 sg13g2_fill_1 FILLER_18_1314 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_fill_1 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_299 ();
 sg13g2_fill_2 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_308 ();
 sg13g2_fill_1 FILLER_19_337 ();
 sg13g2_fill_1 FILLER_19_348 ();
 sg13g2_fill_2 FILLER_19_357 ();
 sg13g2_fill_1 FILLER_19_359 ();
 sg13g2_fill_2 FILLER_19_364 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_378 ();
 sg13g2_fill_1 FILLER_19_380 ();
 sg13g2_decap_4 FILLER_19_385 ();
 sg13g2_fill_2 FILLER_19_389 ();
 sg13g2_fill_2 FILLER_19_422 ();
 sg13g2_decap_8 FILLER_19_443 ();
 sg13g2_decap_4 FILLER_19_450 ();
 sg13g2_fill_1 FILLER_19_454 ();
 sg13g2_fill_2 FILLER_19_460 ();
 sg13g2_fill_1 FILLER_19_462 ();
 sg13g2_fill_2 FILLER_19_472 ();
 sg13g2_fill_1 FILLER_19_474 ();
 sg13g2_fill_2 FILLER_19_479 ();
 sg13g2_fill_1 FILLER_19_481 ();
 sg13g2_fill_2 FILLER_19_538 ();
 sg13g2_fill_1 FILLER_19_540 ();
 sg13g2_decap_4 FILLER_19_555 ();
 sg13g2_fill_2 FILLER_19_589 ();
 sg13g2_fill_2 FILLER_19_625 ();
 sg13g2_fill_1 FILLER_19_627 ();
 sg13g2_decap_8 FILLER_19_663 ();
 sg13g2_fill_1 FILLER_19_695 ();
 sg13g2_fill_1 FILLER_19_706 ();
 sg13g2_decap_4 FILLER_19_726 ();
 sg13g2_fill_2 FILLER_19_740 ();
 sg13g2_fill_1 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_752 ();
 sg13g2_fill_2 FILLER_19_759 ();
 sg13g2_fill_1 FILLER_19_761 ();
 sg13g2_fill_1 FILLER_19_780 ();
 sg13g2_decap_8 FILLER_19_794 ();
 sg13g2_fill_2 FILLER_19_801 ();
 sg13g2_fill_1 FILLER_19_803 ();
 sg13g2_fill_2 FILLER_19_813 ();
 sg13g2_fill_2 FILLER_19_820 ();
 sg13g2_fill_1 FILLER_19_822 ();
 sg13g2_fill_2 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_845 ();
 sg13g2_decap_4 FILLER_19_852 ();
 sg13g2_decap_4 FILLER_19_863 ();
 sg13g2_decap_4 FILLER_19_886 ();
 sg13g2_fill_2 FILLER_19_890 ();
 sg13g2_fill_1 FILLER_19_915 ();
 sg13g2_fill_2 FILLER_19_928 ();
 sg13g2_fill_2 FILLER_19_950 ();
 sg13g2_fill_1 FILLER_19_952 ();
 sg13g2_decap_8 FILLER_19_1044 ();
 sg13g2_decap_8 FILLER_19_1051 ();
 sg13g2_decap_8 FILLER_19_1058 ();
 sg13g2_decap_8 FILLER_19_1065 ();
 sg13g2_decap_8 FILLER_19_1072 ();
 sg13g2_decap_8 FILLER_19_1079 ();
 sg13g2_decap_8 FILLER_19_1086 ();
 sg13g2_decap_8 FILLER_19_1093 ();
 sg13g2_decap_8 FILLER_19_1100 ();
 sg13g2_decap_8 FILLER_19_1107 ();
 sg13g2_decap_8 FILLER_19_1114 ();
 sg13g2_decap_8 FILLER_19_1121 ();
 sg13g2_decap_8 FILLER_19_1128 ();
 sg13g2_decap_8 FILLER_19_1135 ();
 sg13g2_decap_8 FILLER_19_1142 ();
 sg13g2_decap_8 FILLER_19_1149 ();
 sg13g2_decap_8 FILLER_19_1156 ();
 sg13g2_decap_8 FILLER_19_1163 ();
 sg13g2_decap_8 FILLER_19_1170 ();
 sg13g2_decap_8 FILLER_19_1177 ();
 sg13g2_decap_8 FILLER_19_1184 ();
 sg13g2_decap_8 FILLER_19_1191 ();
 sg13g2_decap_8 FILLER_19_1198 ();
 sg13g2_decap_8 FILLER_19_1205 ();
 sg13g2_decap_8 FILLER_19_1212 ();
 sg13g2_decap_8 FILLER_19_1219 ();
 sg13g2_decap_8 FILLER_19_1226 ();
 sg13g2_decap_8 FILLER_19_1233 ();
 sg13g2_decap_8 FILLER_19_1240 ();
 sg13g2_decap_8 FILLER_19_1247 ();
 sg13g2_decap_8 FILLER_19_1254 ();
 sg13g2_decap_8 FILLER_19_1261 ();
 sg13g2_decap_8 FILLER_19_1268 ();
 sg13g2_decap_8 FILLER_19_1275 ();
 sg13g2_decap_8 FILLER_19_1282 ();
 sg13g2_decap_8 FILLER_19_1289 ();
 sg13g2_decap_8 FILLER_19_1296 ();
 sg13g2_decap_8 FILLER_19_1303 ();
 sg13g2_decap_4 FILLER_19_1310 ();
 sg13g2_fill_1 FILLER_19_1314 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_4 FILLER_20_119 ();
 sg13g2_fill_2 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_142 ();
 sg13g2_fill_1 FILLER_20_149 ();
 sg13g2_fill_2 FILLER_20_154 ();
 sg13g2_fill_1 FILLER_20_156 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_fill_1 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_fill_2 FILLER_20_314 ();
 sg13g2_fill_1 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_340 ();
 sg13g2_fill_1 FILLER_20_342 ();
 sg13g2_fill_1 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_20_396 ();
 sg13g2_fill_1 FILLER_20_398 ();
 sg13g2_fill_2 FILLER_20_403 ();
 sg13g2_fill_1 FILLER_20_405 ();
 sg13g2_fill_2 FILLER_20_410 ();
 sg13g2_fill_1 FILLER_20_412 ();
 sg13g2_fill_1 FILLER_20_476 ();
 sg13g2_fill_2 FILLER_20_485 ();
 sg13g2_fill_1 FILLER_20_497 ();
 sg13g2_decap_4 FILLER_20_532 ();
 sg13g2_fill_2 FILLER_20_536 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_562 ();
 sg13g2_decap_4 FILLER_20_569 ();
 sg13g2_fill_1 FILLER_20_573 ();
 sg13g2_fill_1 FILLER_20_578 ();
 sg13g2_fill_1 FILLER_20_583 ();
 sg13g2_fill_2 FILLER_20_632 ();
 sg13g2_fill_1 FILLER_20_634 ();
 sg13g2_decap_8 FILLER_20_646 ();
 sg13g2_decap_4 FILLER_20_653 ();
 sg13g2_fill_2 FILLER_20_657 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_fill_1 FILLER_20_679 ();
 sg13g2_fill_2 FILLER_20_685 ();
 sg13g2_fill_2 FILLER_20_711 ();
 sg13g2_fill_1 FILLER_20_713 ();
 sg13g2_decap_8 FILLER_20_718 ();
 sg13g2_decap_4 FILLER_20_725 ();
 sg13g2_fill_2 FILLER_20_729 ();
 sg13g2_fill_2 FILLER_20_736 ();
 sg13g2_fill_1 FILLER_20_738 ();
 sg13g2_decap_8 FILLER_20_743 ();
 sg13g2_decap_4 FILLER_20_750 ();
 sg13g2_fill_1 FILLER_20_754 ();
 sg13g2_decap_4 FILLER_20_775 ();
 sg13g2_fill_2 FILLER_20_813 ();
 sg13g2_fill_1 FILLER_20_815 ();
 sg13g2_fill_2 FILLER_20_846 ();
 sg13g2_fill_2 FILLER_20_853 ();
 sg13g2_fill_1 FILLER_20_855 ();
 sg13g2_decap_4 FILLER_20_886 ();
 sg13g2_fill_2 FILLER_20_895 ();
 sg13g2_fill_1 FILLER_20_897 ();
 sg13g2_fill_2 FILLER_20_910 ();
 sg13g2_fill_1 FILLER_20_912 ();
 sg13g2_fill_2 FILLER_20_936 ();
 sg13g2_decap_8 FILLER_20_947 ();
 sg13g2_decap_8 FILLER_20_954 ();
 sg13g2_fill_1 FILLER_20_982 ();
 sg13g2_fill_1 FILLER_20_1000 ();
 sg13g2_decap_8 FILLER_20_1041 ();
 sg13g2_decap_8 FILLER_20_1048 ();
 sg13g2_decap_8 FILLER_20_1055 ();
 sg13g2_decap_8 FILLER_20_1062 ();
 sg13g2_decap_8 FILLER_20_1069 ();
 sg13g2_decap_8 FILLER_20_1076 ();
 sg13g2_decap_8 FILLER_20_1083 ();
 sg13g2_decap_8 FILLER_20_1090 ();
 sg13g2_decap_8 FILLER_20_1097 ();
 sg13g2_decap_8 FILLER_20_1104 ();
 sg13g2_decap_8 FILLER_20_1111 ();
 sg13g2_decap_8 FILLER_20_1118 ();
 sg13g2_decap_8 FILLER_20_1125 ();
 sg13g2_decap_8 FILLER_20_1132 ();
 sg13g2_decap_8 FILLER_20_1139 ();
 sg13g2_decap_8 FILLER_20_1146 ();
 sg13g2_decap_8 FILLER_20_1153 ();
 sg13g2_decap_8 FILLER_20_1160 ();
 sg13g2_decap_8 FILLER_20_1167 ();
 sg13g2_decap_8 FILLER_20_1174 ();
 sg13g2_decap_8 FILLER_20_1181 ();
 sg13g2_decap_8 FILLER_20_1188 ();
 sg13g2_decap_8 FILLER_20_1195 ();
 sg13g2_decap_8 FILLER_20_1202 ();
 sg13g2_decap_8 FILLER_20_1209 ();
 sg13g2_decap_8 FILLER_20_1216 ();
 sg13g2_decap_8 FILLER_20_1223 ();
 sg13g2_decap_8 FILLER_20_1230 ();
 sg13g2_decap_8 FILLER_20_1237 ();
 sg13g2_decap_8 FILLER_20_1244 ();
 sg13g2_decap_8 FILLER_20_1251 ();
 sg13g2_decap_8 FILLER_20_1258 ();
 sg13g2_decap_8 FILLER_20_1265 ();
 sg13g2_decap_8 FILLER_20_1272 ();
 sg13g2_decap_8 FILLER_20_1279 ();
 sg13g2_decap_8 FILLER_20_1286 ();
 sg13g2_decap_8 FILLER_20_1293 ();
 sg13g2_decap_8 FILLER_20_1300 ();
 sg13g2_decap_8 FILLER_20_1307 ();
 sg13g2_fill_1 FILLER_20_1314 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_117 ();
 sg13g2_fill_2 FILLER_21_149 ();
 sg13g2_fill_1 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_decap_4 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_fill_2 FILLER_21_234 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_350 ();
 sg13g2_fill_2 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_fill_2 FILLER_21_397 ();
 sg13g2_fill_1 FILLER_21_399 ();
 sg13g2_fill_1 FILLER_21_439 ();
 sg13g2_fill_1 FILLER_21_458 ();
 sg13g2_fill_1 FILLER_21_498 ();
 sg13g2_fill_1 FILLER_21_508 ();
 sg13g2_fill_1 FILLER_21_544 ();
 sg13g2_fill_2 FILLER_21_562 ();
 sg13g2_decap_4 FILLER_21_590 ();
 sg13g2_fill_2 FILLER_21_594 ();
 sg13g2_decap_8 FILLER_21_626 ();
 sg13g2_fill_1 FILLER_21_633 ();
 sg13g2_decap_4 FILLER_21_687 ();
 sg13g2_fill_1 FILLER_21_691 ();
 sg13g2_fill_2 FILLER_21_696 ();
 sg13g2_decap_4 FILLER_21_703 ();
 sg13g2_fill_2 FILLER_21_707 ();
 sg13g2_fill_2 FILLER_21_734 ();
 sg13g2_fill_2 FILLER_21_746 ();
 sg13g2_decap_8 FILLER_21_768 ();
 sg13g2_fill_1 FILLER_21_775 ();
 sg13g2_decap_4 FILLER_21_789 ();
 sg13g2_fill_1 FILLER_21_797 ();
 sg13g2_decap_8 FILLER_21_802 ();
 sg13g2_fill_2 FILLER_21_817 ();
 sg13g2_fill_1 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_838 ();
 sg13g2_fill_2 FILLER_21_845 ();
 sg13g2_decap_4 FILLER_21_851 ();
 sg13g2_fill_2 FILLER_21_855 ();
 sg13g2_decap_4 FILLER_21_869 ();
 sg13g2_decap_4 FILLER_21_888 ();
 sg13g2_fill_2 FILLER_21_892 ();
 sg13g2_fill_2 FILLER_21_899 ();
 sg13g2_fill_1 FILLER_21_901 ();
 sg13g2_fill_2 FILLER_21_907 ();
 sg13g2_fill_1 FILLER_21_909 ();
 sg13g2_fill_2 FILLER_21_931 ();
 sg13g2_fill_1 FILLER_21_933 ();
 sg13g2_decap_8 FILLER_21_952 ();
 sg13g2_decap_8 FILLER_21_959 ();
 sg13g2_fill_2 FILLER_21_966 ();
 sg13g2_fill_2 FILLER_21_1007 ();
 sg13g2_decap_8 FILLER_21_1031 ();
 sg13g2_decap_8 FILLER_21_1038 ();
 sg13g2_decap_8 FILLER_21_1045 ();
 sg13g2_decap_8 FILLER_21_1052 ();
 sg13g2_decap_8 FILLER_21_1059 ();
 sg13g2_decap_8 FILLER_21_1066 ();
 sg13g2_decap_8 FILLER_21_1073 ();
 sg13g2_decap_8 FILLER_21_1080 ();
 sg13g2_decap_8 FILLER_21_1087 ();
 sg13g2_decap_8 FILLER_21_1094 ();
 sg13g2_decap_8 FILLER_21_1101 ();
 sg13g2_decap_8 FILLER_21_1108 ();
 sg13g2_decap_8 FILLER_21_1115 ();
 sg13g2_decap_8 FILLER_21_1122 ();
 sg13g2_decap_8 FILLER_21_1129 ();
 sg13g2_decap_8 FILLER_21_1136 ();
 sg13g2_decap_8 FILLER_21_1143 ();
 sg13g2_decap_8 FILLER_21_1150 ();
 sg13g2_decap_8 FILLER_21_1157 ();
 sg13g2_decap_8 FILLER_21_1164 ();
 sg13g2_decap_8 FILLER_21_1171 ();
 sg13g2_decap_8 FILLER_21_1178 ();
 sg13g2_decap_8 FILLER_21_1185 ();
 sg13g2_decap_8 FILLER_21_1192 ();
 sg13g2_decap_8 FILLER_21_1199 ();
 sg13g2_decap_8 FILLER_21_1206 ();
 sg13g2_decap_8 FILLER_21_1213 ();
 sg13g2_decap_8 FILLER_21_1220 ();
 sg13g2_decap_8 FILLER_21_1227 ();
 sg13g2_decap_8 FILLER_21_1234 ();
 sg13g2_decap_8 FILLER_21_1241 ();
 sg13g2_decap_8 FILLER_21_1248 ();
 sg13g2_decap_8 FILLER_21_1255 ();
 sg13g2_decap_8 FILLER_21_1262 ();
 sg13g2_decap_8 FILLER_21_1269 ();
 sg13g2_decap_8 FILLER_21_1276 ();
 sg13g2_decap_8 FILLER_21_1283 ();
 sg13g2_decap_8 FILLER_21_1290 ();
 sg13g2_decap_8 FILLER_21_1297 ();
 sg13g2_decap_8 FILLER_21_1304 ();
 sg13g2_decap_4 FILLER_21_1311 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_135 ();
 sg13g2_fill_2 FILLER_22_167 ();
 sg13g2_fill_1 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_217 ();
 sg13g2_fill_2 FILLER_22_222 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_fill_2 FILLER_22_321 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_fill_1 FILLER_22_342 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_424 ();
 sg13g2_fill_1 FILLER_22_460 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_fill_2 FILLER_22_480 ();
 sg13g2_fill_1 FILLER_22_482 ();
 sg13g2_fill_2 FILLER_22_487 ();
 sg13g2_fill_1 FILLER_22_520 ();
 sg13g2_fill_2 FILLER_22_531 ();
 sg13g2_decap_8 FILLER_22_587 ();
 sg13g2_fill_1 FILLER_22_594 ();
 sg13g2_decap_8 FILLER_22_599 ();
 sg13g2_fill_2 FILLER_22_606 ();
 sg13g2_decap_4 FILLER_22_642 ();
 sg13g2_fill_2 FILLER_22_646 ();
 sg13g2_decap_8 FILLER_22_660 ();
 sg13g2_decap_8 FILLER_22_667 ();
 sg13g2_fill_1 FILLER_22_674 ();
 sg13g2_fill_2 FILLER_22_683 ();
 sg13g2_fill_1 FILLER_22_685 ();
 sg13g2_fill_1 FILLER_22_705 ();
 sg13g2_decap_8 FILLER_22_716 ();
 sg13g2_decap_8 FILLER_22_723 ();
 sg13g2_fill_2 FILLER_22_730 ();
 sg13g2_decap_4 FILLER_22_742 ();
 sg13g2_fill_2 FILLER_22_755 ();
 sg13g2_fill_1 FILLER_22_757 ();
 sg13g2_decap_4 FILLER_22_766 ();
 sg13g2_fill_1 FILLER_22_770 ();
 sg13g2_fill_1 FILLER_22_801 ();
 sg13g2_fill_2 FILLER_22_816 ();
 sg13g2_fill_1 FILLER_22_818 ();
 sg13g2_fill_1 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_879 ();
 sg13g2_fill_2 FILLER_22_909 ();
 sg13g2_fill_2 FILLER_22_932 ();
 sg13g2_fill_1 FILLER_22_934 ();
 sg13g2_decap_8 FILLER_22_945 ();
 sg13g2_decap_8 FILLER_22_952 ();
 sg13g2_decap_8 FILLER_22_959 ();
 sg13g2_decap_4 FILLER_22_966 ();
 sg13g2_fill_2 FILLER_22_970 ();
 sg13g2_fill_2 FILLER_22_985 ();
 sg13g2_fill_1 FILLER_22_987 ();
 sg13g2_decap_8 FILLER_22_1045 ();
 sg13g2_decap_8 FILLER_22_1052 ();
 sg13g2_decap_8 FILLER_22_1059 ();
 sg13g2_decap_8 FILLER_22_1066 ();
 sg13g2_decap_8 FILLER_22_1073 ();
 sg13g2_decap_8 FILLER_22_1080 ();
 sg13g2_decap_8 FILLER_22_1087 ();
 sg13g2_decap_8 FILLER_22_1094 ();
 sg13g2_decap_8 FILLER_22_1101 ();
 sg13g2_decap_8 FILLER_22_1108 ();
 sg13g2_decap_8 FILLER_22_1115 ();
 sg13g2_decap_8 FILLER_22_1122 ();
 sg13g2_decap_8 FILLER_22_1129 ();
 sg13g2_decap_8 FILLER_22_1136 ();
 sg13g2_decap_8 FILLER_22_1143 ();
 sg13g2_decap_8 FILLER_22_1150 ();
 sg13g2_decap_8 FILLER_22_1157 ();
 sg13g2_decap_8 FILLER_22_1164 ();
 sg13g2_decap_8 FILLER_22_1171 ();
 sg13g2_decap_8 FILLER_22_1178 ();
 sg13g2_decap_8 FILLER_22_1185 ();
 sg13g2_decap_8 FILLER_22_1192 ();
 sg13g2_decap_8 FILLER_22_1199 ();
 sg13g2_decap_8 FILLER_22_1206 ();
 sg13g2_decap_8 FILLER_22_1213 ();
 sg13g2_decap_8 FILLER_22_1220 ();
 sg13g2_decap_8 FILLER_22_1227 ();
 sg13g2_decap_8 FILLER_22_1234 ();
 sg13g2_decap_8 FILLER_22_1241 ();
 sg13g2_decap_8 FILLER_22_1248 ();
 sg13g2_decap_8 FILLER_22_1255 ();
 sg13g2_decap_8 FILLER_22_1262 ();
 sg13g2_decap_8 FILLER_22_1269 ();
 sg13g2_decap_8 FILLER_22_1276 ();
 sg13g2_decap_8 FILLER_22_1283 ();
 sg13g2_decap_8 FILLER_22_1290 ();
 sg13g2_decap_8 FILLER_22_1297 ();
 sg13g2_decap_8 FILLER_22_1304 ();
 sg13g2_decap_4 FILLER_22_1311 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_decap_4 FILLER_23_122 ();
 sg13g2_fill_2 FILLER_23_126 ();
 sg13g2_decap_4 FILLER_23_142 ();
 sg13g2_fill_2 FILLER_23_146 ();
 sg13g2_fill_1 FILLER_23_152 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_fill_2 FILLER_23_178 ();
 sg13g2_fill_1 FILLER_23_202 ();
 sg13g2_fill_2 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_241 ();
 sg13g2_decap_4 FILLER_23_256 ();
 sg13g2_fill_2 FILLER_23_260 ();
 sg13g2_fill_2 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_374 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_4 FILLER_23_393 ();
 sg13g2_fill_2 FILLER_23_397 ();
 sg13g2_fill_2 FILLER_23_420 ();
 sg13g2_fill_2 FILLER_23_452 ();
 sg13g2_fill_2 FILLER_23_468 ();
 sg13g2_fill_1 FILLER_23_470 ();
 sg13g2_decap_4 FILLER_23_502 ();
 sg13g2_fill_1 FILLER_23_506 ();
 sg13g2_fill_1 FILLER_23_523 ();
 sg13g2_fill_2 FILLER_23_539 ();
 sg13g2_fill_1 FILLER_23_541 ();
 sg13g2_decap_4 FILLER_23_581 ();
 sg13g2_fill_1 FILLER_23_594 ();
 sg13g2_decap_4 FILLER_23_621 ();
 sg13g2_decap_4 FILLER_23_632 ();
 sg13g2_fill_2 FILLER_23_636 ();
 sg13g2_decap_8 FILLER_23_654 ();
 sg13g2_fill_2 FILLER_23_669 ();
 sg13g2_decap_4 FILLER_23_679 ();
 sg13g2_fill_2 FILLER_23_688 ();
 sg13g2_fill_1 FILLER_23_690 ();
 sg13g2_decap_4 FILLER_23_704 ();
 sg13g2_fill_1 FILLER_23_708 ();
 sg13g2_decap_4 FILLER_23_724 ();
 sg13g2_fill_2 FILLER_23_728 ();
 sg13g2_decap_4 FILLER_23_751 ();
 sg13g2_fill_2 FILLER_23_768 ();
 sg13g2_fill_2 FILLER_23_777 ();
 sg13g2_fill_2 FILLER_23_783 ();
 sg13g2_fill_1 FILLER_23_793 ();
 sg13g2_decap_8 FILLER_23_815 ();
 sg13g2_decap_8 FILLER_23_822 ();
 sg13g2_fill_1 FILLER_23_829 ();
 sg13g2_fill_2 FILLER_23_840 ();
 sg13g2_decap_4 FILLER_23_848 ();
 sg13g2_fill_2 FILLER_23_862 ();
 sg13g2_fill_1 FILLER_23_864 ();
 sg13g2_fill_1 FILLER_23_879 ();
 sg13g2_decap_8 FILLER_23_897 ();
 sg13g2_fill_2 FILLER_23_904 ();
 sg13g2_decap_4 FILLER_23_921 ();
 sg13g2_decap_4 FILLER_23_944 ();
 sg13g2_fill_2 FILLER_23_948 ();
 sg13g2_decap_8 FILLER_23_1028 ();
 sg13g2_decap_8 FILLER_23_1035 ();
 sg13g2_decap_8 FILLER_23_1042 ();
 sg13g2_decap_8 FILLER_23_1049 ();
 sg13g2_decap_8 FILLER_23_1056 ();
 sg13g2_decap_8 FILLER_23_1063 ();
 sg13g2_decap_8 FILLER_23_1070 ();
 sg13g2_decap_8 FILLER_23_1077 ();
 sg13g2_decap_8 FILLER_23_1084 ();
 sg13g2_decap_8 FILLER_23_1091 ();
 sg13g2_decap_8 FILLER_23_1098 ();
 sg13g2_decap_8 FILLER_23_1105 ();
 sg13g2_decap_8 FILLER_23_1112 ();
 sg13g2_decap_8 FILLER_23_1119 ();
 sg13g2_decap_8 FILLER_23_1126 ();
 sg13g2_decap_8 FILLER_23_1133 ();
 sg13g2_decap_8 FILLER_23_1140 ();
 sg13g2_decap_8 FILLER_23_1147 ();
 sg13g2_decap_8 FILLER_23_1154 ();
 sg13g2_decap_8 FILLER_23_1161 ();
 sg13g2_decap_8 FILLER_23_1168 ();
 sg13g2_decap_8 FILLER_23_1175 ();
 sg13g2_decap_8 FILLER_23_1182 ();
 sg13g2_decap_8 FILLER_23_1189 ();
 sg13g2_decap_8 FILLER_23_1196 ();
 sg13g2_decap_8 FILLER_23_1203 ();
 sg13g2_decap_8 FILLER_23_1210 ();
 sg13g2_decap_8 FILLER_23_1217 ();
 sg13g2_decap_8 FILLER_23_1224 ();
 sg13g2_decap_8 FILLER_23_1231 ();
 sg13g2_decap_8 FILLER_23_1238 ();
 sg13g2_decap_8 FILLER_23_1245 ();
 sg13g2_decap_8 FILLER_23_1252 ();
 sg13g2_decap_8 FILLER_23_1259 ();
 sg13g2_decap_8 FILLER_23_1266 ();
 sg13g2_decap_8 FILLER_23_1273 ();
 sg13g2_decap_8 FILLER_23_1280 ();
 sg13g2_decap_8 FILLER_23_1287 ();
 sg13g2_decap_8 FILLER_23_1294 ();
 sg13g2_decap_8 FILLER_23_1301 ();
 sg13g2_decap_8 FILLER_23_1308 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_fill_2 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_decap_8 FILLER_24_190 ();
 sg13g2_decap_4 FILLER_24_197 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_232 ();
 sg13g2_fill_1 FILLER_24_280 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_323 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_fill_2 FILLER_24_345 ();
 sg13g2_fill_1 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_fill_2 FILLER_24_438 ();
 sg13g2_fill_1 FILLER_24_440 ();
 sg13g2_fill_2 FILLER_24_450 ();
 sg13g2_fill_2 FILLER_24_460 ();
 sg13g2_fill_1 FILLER_24_462 ();
 sg13g2_fill_1 FILLER_24_468 ();
 sg13g2_fill_2 FILLER_24_484 ();
 sg13g2_fill_1 FILLER_24_512 ();
 sg13g2_decap_8 FILLER_24_544 ();
 sg13g2_decap_4 FILLER_24_551 ();
 sg13g2_decap_4 FILLER_24_585 ();
 sg13g2_fill_2 FILLER_24_589 ();
 sg13g2_decap_4 FILLER_24_644 ();
 sg13g2_decap_4 FILLER_24_660 ();
 sg13g2_fill_2 FILLER_24_692 ();
 sg13g2_fill_1 FILLER_24_694 ();
 sg13g2_decap_4 FILLER_24_707 ();
 sg13g2_fill_2 FILLER_24_721 ();
 sg13g2_fill_1 FILLER_24_731 ();
 sg13g2_fill_1 FILLER_24_736 ();
 sg13g2_fill_2 FILLER_24_759 ();
 sg13g2_fill_1 FILLER_24_779 ();
 sg13g2_decap_4 FILLER_24_791 ();
 sg13g2_fill_2 FILLER_24_795 ();
 sg13g2_fill_1 FILLER_24_802 ();
 sg13g2_fill_2 FILLER_24_813 ();
 sg13g2_fill_1 FILLER_24_815 ();
 sg13g2_fill_2 FILLER_24_824 ();
 sg13g2_fill_2 FILLER_24_840 ();
 sg13g2_fill_1 FILLER_24_842 ();
 sg13g2_decap_8 FILLER_24_863 ();
 sg13g2_fill_2 FILLER_24_870 ();
 sg13g2_fill_1 FILLER_24_872 ();
 sg13g2_fill_2 FILLER_24_884 ();
 sg13g2_fill_1 FILLER_24_886 ();
 sg13g2_fill_1 FILLER_24_894 ();
 sg13g2_decap_4 FILLER_24_929 ();
 sg13g2_fill_2 FILLER_24_933 ();
 sg13g2_decap_8 FILLER_24_945 ();
 sg13g2_decap_4 FILLER_24_952 ();
 sg13g2_fill_2 FILLER_24_956 ();
 sg13g2_fill_2 FILLER_24_971 ();
 sg13g2_fill_1 FILLER_24_987 ();
 sg13g2_fill_1 FILLER_24_1002 ();
 sg13g2_decap_8 FILLER_24_1020 ();
 sg13g2_decap_8 FILLER_24_1027 ();
 sg13g2_decap_8 FILLER_24_1034 ();
 sg13g2_decap_8 FILLER_24_1041 ();
 sg13g2_decap_8 FILLER_24_1048 ();
 sg13g2_decap_8 FILLER_24_1055 ();
 sg13g2_decap_8 FILLER_24_1062 ();
 sg13g2_decap_8 FILLER_24_1069 ();
 sg13g2_decap_8 FILLER_24_1076 ();
 sg13g2_decap_8 FILLER_24_1083 ();
 sg13g2_decap_8 FILLER_24_1090 ();
 sg13g2_decap_8 FILLER_24_1097 ();
 sg13g2_decap_8 FILLER_24_1104 ();
 sg13g2_decap_8 FILLER_24_1111 ();
 sg13g2_decap_8 FILLER_24_1118 ();
 sg13g2_decap_8 FILLER_24_1125 ();
 sg13g2_decap_8 FILLER_24_1132 ();
 sg13g2_decap_8 FILLER_24_1139 ();
 sg13g2_decap_8 FILLER_24_1146 ();
 sg13g2_decap_8 FILLER_24_1153 ();
 sg13g2_decap_8 FILLER_24_1160 ();
 sg13g2_decap_8 FILLER_24_1167 ();
 sg13g2_decap_8 FILLER_24_1174 ();
 sg13g2_decap_8 FILLER_24_1181 ();
 sg13g2_decap_8 FILLER_24_1188 ();
 sg13g2_decap_8 FILLER_24_1195 ();
 sg13g2_decap_8 FILLER_24_1202 ();
 sg13g2_decap_8 FILLER_24_1209 ();
 sg13g2_decap_8 FILLER_24_1216 ();
 sg13g2_decap_8 FILLER_24_1223 ();
 sg13g2_decap_8 FILLER_24_1230 ();
 sg13g2_decap_8 FILLER_24_1237 ();
 sg13g2_decap_8 FILLER_24_1244 ();
 sg13g2_decap_8 FILLER_24_1251 ();
 sg13g2_decap_8 FILLER_24_1258 ();
 sg13g2_decap_8 FILLER_24_1265 ();
 sg13g2_decap_8 FILLER_24_1272 ();
 sg13g2_decap_8 FILLER_24_1279 ();
 sg13g2_decap_8 FILLER_24_1286 ();
 sg13g2_decap_8 FILLER_24_1293 ();
 sg13g2_decap_8 FILLER_24_1300 ();
 sg13g2_decap_8 FILLER_24_1307 ();
 sg13g2_fill_1 FILLER_24_1314 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_146 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_fill_2 FILLER_25_330 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_fill_1 FILLER_25_396 ();
 sg13g2_fill_1 FILLER_25_409 ();
 sg13g2_decap_4 FILLER_25_414 ();
 sg13g2_fill_2 FILLER_25_418 ();
 sg13g2_decap_4 FILLER_25_472 ();
 sg13g2_fill_2 FILLER_25_481 ();
 sg13g2_fill_1 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_492 ();
 sg13g2_fill_2 FILLER_25_499 ();
 sg13g2_decap_4 FILLER_25_562 ();
 sg13g2_fill_2 FILLER_25_566 ();
 sg13g2_decap_4 FILLER_25_571 ();
 sg13g2_fill_1 FILLER_25_589 ();
 sg13g2_fill_2 FILLER_25_595 ();
 sg13g2_fill_1 FILLER_25_597 ();
 sg13g2_fill_1 FILLER_25_611 ();
 sg13g2_fill_2 FILLER_25_628 ();
 sg13g2_fill_2 FILLER_25_641 ();
 sg13g2_fill_2 FILLER_25_656 ();
 sg13g2_decap_4 FILLER_25_666 ();
 sg13g2_fill_1 FILLER_25_670 ();
 sg13g2_decap_8 FILLER_25_677 ();
 sg13g2_decap_4 FILLER_25_684 ();
 sg13g2_decap_4 FILLER_25_696 ();
 sg13g2_fill_1 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_723 ();
 sg13g2_decap_4 FILLER_25_730 ();
 sg13g2_decap_4 FILLER_25_739 ();
 sg13g2_fill_1 FILLER_25_743 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_4 FILLER_25_756 ();
 sg13g2_fill_2 FILLER_25_769 ();
 sg13g2_fill_1 FILLER_25_771 ();
 sg13g2_fill_2 FILLER_25_788 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_4 FILLER_25_826 ();
 sg13g2_fill_2 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_4 FILLER_25_894 ();
 sg13g2_fill_1 FILLER_25_910 ();
 sg13g2_fill_2 FILLER_25_922 ();
 sg13g2_fill_1 FILLER_25_924 ();
 sg13g2_fill_2 FILLER_25_954 ();
 sg13g2_fill_2 FILLER_25_960 ();
 sg13g2_fill_2 FILLER_25_966 ();
 sg13g2_decap_8 FILLER_25_1036 ();
 sg13g2_decap_8 FILLER_25_1043 ();
 sg13g2_decap_8 FILLER_25_1050 ();
 sg13g2_decap_8 FILLER_25_1057 ();
 sg13g2_decap_8 FILLER_25_1064 ();
 sg13g2_decap_8 FILLER_25_1071 ();
 sg13g2_decap_8 FILLER_25_1078 ();
 sg13g2_decap_8 FILLER_25_1085 ();
 sg13g2_decap_8 FILLER_25_1092 ();
 sg13g2_decap_8 FILLER_25_1099 ();
 sg13g2_decap_8 FILLER_25_1106 ();
 sg13g2_decap_8 FILLER_25_1113 ();
 sg13g2_decap_8 FILLER_25_1120 ();
 sg13g2_decap_8 FILLER_25_1127 ();
 sg13g2_decap_8 FILLER_25_1134 ();
 sg13g2_decap_8 FILLER_25_1141 ();
 sg13g2_decap_8 FILLER_25_1148 ();
 sg13g2_decap_8 FILLER_25_1155 ();
 sg13g2_decap_8 FILLER_25_1162 ();
 sg13g2_decap_8 FILLER_25_1169 ();
 sg13g2_decap_8 FILLER_25_1176 ();
 sg13g2_decap_8 FILLER_25_1183 ();
 sg13g2_decap_8 FILLER_25_1190 ();
 sg13g2_decap_8 FILLER_25_1197 ();
 sg13g2_decap_8 FILLER_25_1204 ();
 sg13g2_decap_8 FILLER_25_1211 ();
 sg13g2_decap_8 FILLER_25_1218 ();
 sg13g2_decap_8 FILLER_25_1225 ();
 sg13g2_decap_8 FILLER_25_1232 ();
 sg13g2_decap_8 FILLER_25_1239 ();
 sg13g2_decap_8 FILLER_25_1246 ();
 sg13g2_decap_8 FILLER_25_1253 ();
 sg13g2_decap_8 FILLER_25_1260 ();
 sg13g2_decap_8 FILLER_25_1267 ();
 sg13g2_decap_8 FILLER_25_1274 ();
 sg13g2_decap_8 FILLER_25_1281 ();
 sg13g2_decap_8 FILLER_25_1288 ();
 sg13g2_decap_8 FILLER_25_1295 ();
 sg13g2_decap_8 FILLER_25_1302 ();
 sg13g2_decap_4 FILLER_25_1309 ();
 sg13g2_fill_2 FILLER_25_1313 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_decap_8 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_fill_2 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_327 ();
 sg13g2_fill_1 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_348 ();
 sg13g2_fill_1 FILLER_26_357 ();
 sg13g2_fill_2 FILLER_26_379 ();
 sg13g2_fill_1 FILLER_26_407 ();
 sg13g2_fill_2 FILLER_26_466 ();
 sg13g2_fill_1 FILLER_26_508 ();
 sg13g2_fill_2 FILLER_26_519 ();
 sg13g2_fill_2 FILLER_26_603 ();
 sg13g2_fill_1 FILLER_26_605 ();
 sg13g2_decap_4 FILLER_26_610 ();
 sg13g2_fill_1 FILLER_26_614 ();
 sg13g2_fill_1 FILLER_26_619 ();
 sg13g2_fill_2 FILLER_26_629 ();
 sg13g2_fill_1 FILLER_26_631 ();
 sg13g2_fill_2 FILLER_26_682 ();
 sg13g2_fill_1 FILLER_26_684 ();
 sg13g2_decap_8 FILLER_26_699 ();
 sg13g2_fill_1 FILLER_26_706 ();
 sg13g2_fill_2 FILLER_26_720 ();
 sg13g2_decap_4 FILLER_26_730 ();
 sg13g2_fill_1 FILLER_26_734 ();
 sg13g2_decap_4 FILLER_26_739 ();
 sg13g2_fill_2 FILLER_26_743 ();
 sg13g2_fill_2 FILLER_26_760 ();
 sg13g2_fill_1 FILLER_26_762 ();
 sg13g2_fill_1 FILLER_26_768 ();
 sg13g2_decap_4 FILLER_26_774 ();
 sg13g2_fill_1 FILLER_26_778 ();
 sg13g2_fill_2 FILLER_26_789 ();
 sg13g2_fill_1 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_811 ();
 sg13g2_decap_4 FILLER_26_818 ();
 sg13g2_fill_1 FILLER_26_837 ();
 sg13g2_decap_8 FILLER_26_842 ();
 sg13g2_fill_2 FILLER_26_866 ();
 sg13g2_fill_1 FILLER_26_868 ();
 sg13g2_fill_1 FILLER_26_878 ();
 sg13g2_decap_8 FILLER_26_884 ();
 sg13g2_decap_8 FILLER_26_891 ();
 sg13g2_decap_8 FILLER_26_898 ();
 sg13g2_decap_8 FILLER_26_910 ();
 sg13g2_fill_2 FILLER_26_917 ();
 sg13g2_fill_1 FILLER_26_919 ();
 sg13g2_decap_4 FILLER_26_931 ();
 sg13g2_fill_2 FILLER_26_935 ();
 sg13g2_decap_4 FILLER_26_947 ();
 sg13g2_decap_8 FILLER_26_1026 ();
 sg13g2_decap_8 FILLER_26_1033 ();
 sg13g2_decap_8 FILLER_26_1040 ();
 sg13g2_decap_8 FILLER_26_1047 ();
 sg13g2_decap_8 FILLER_26_1054 ();
 sg13g2_decap_8 FILLER_26_1061 ();
 sg13g2_decap_8 FILLER_26_1068 ();
 sg13g2_decap_8 FILLER_26_1075 ();
 sg13g2_decap_8 FILLER_26_1082 ();
 sg13g2_decap_8 FILLER_26_1089 ();
 sg13g2_decap_8 FILLER_26_1096 ();
 sg13g2_decap_8 FILLER_26_1103 ();
 sg13g2_decap_8 FILLER_26_1110 ();
 sg13g2_decap_8 FILLER_26_1117 ();
 sg13g2_decap_8 FILLER_26_1124 ();
 sg13g2_decap_8 FILLER_26_1131 ();
 sg13g2_decap_8 FILLER_26_1138 ();
 sg13g2_decap_8 FILLER_26_1145 ();
 sg13g2_decap_8 FILLER_26_1152 ();
 sg13g2_decap_8 FILLER_26_1159 ();
 sg13g2_decap_8 FILLER_26_1166 ();
 sg13g2_decap_8 FILLER_26_1173 ();
 sg13g2_decap_8 FILLER_26_1180 ();
 sg13g2_decap_8 FILLER_26_1187 ();
 sg13g2_decap_8 FILLER_26_1194 ();
 sg13g2_decap_8 FILLER_26_1201 ();
 sg13g2_decap_8 FILLER_26_1208 ();
 sg13g2_decap_8 FILLER_26_1215 ();
 sg13g2_decap_8 FILLER_26_1222 ();
 sg13g2_decap_8 FILLER_26_1229 ();
 sg13g2_decap_8 FILLER_26_1236 ();
 sg13g2_decap_8 FILLER_26_1243 ();
 sg13g2_decap_8 FILLER_26_1250 ();
 sg13g2_decap_8 FILLER_26_1257 ();
 sg13g2_decap_8 FILLER_26_1264 ();
 sg13g2_decap_8 FILLER_26_1271 ();
 sg13g2_decap_8 FILLER_26_1278 ();
 sg13g2_decap_8 FILLER_26_1285 ();
 sg13g2_decap_8 FILLER_26_1292 ();
 sg13g2_decap_8 FILLER_26_1299 ();
 sg13g2_decap_8 FILLER_26_1306 ();
 sg13g2_fill_2 FILLER_26_1313 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_fill_1 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_217 ();
 sg13g2_fill_1 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_decap_4 FILLER_27_271 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_320 ();
 sg13g2_decap_4 FILLER_27_365 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_decap_4 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_411 ();
 sg13g2_fill_1 FILLER_27_413 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_fill_2 FILLER_27_476 ();
 sg13g2_fill_1 FILLER_27_478 ();
 sg13g2_fill_2 FILLER_27_551 ();
 sg13g2_decap_8 FILLER_27_557 ();
 sg13g2_decap_8 FILLER_27_564 ();
 sg13g2_fill_1 FILLER_27_571 ();
 sg13g2_decap_8 FILLER_27_576 ();
 sg13g2_decap_8 FILLER_27_583 ();
 sg13g2_decap_8 FILLER_27_590 ();
 sg13g2_decap_4 FILLER_27_597 ();
 sg13g2_decap_8 FILLER_27_631 ();
 sg13g2_fill_2 FILLER_27_638 ();
 sg13g2_decap_4 FILLER_27_662 ();
 sg13g2_fill_1 FILLER_27_666 ();
 sg13g2_fill_1 FILLER_27_683 ();
 sg13g2_fill_1 FILLER_27_694 ();
 sg13g2_fill_2 FILLER_27_708 ();
 sg13g2_fill_1 FILLER_27_730 ();
 sg13g2_fill_2 FILLER_27_742 ();
 sg13g2_fill_1 FILLER_27_744 ();
 sg13g2_fill_2 FILLER_27_759 ();
 sg13g2_decap_4 FILLER_27_783 ();
 sg13g2_fill_1 FILLER_27_797 ();
 sg13g2_fill_2 FILLER_27_814 ();
 sg13g2_fill_2 FILLER_27_829 ();
 sg13g2_fill_1 FILLER_27_831 ();
 sg13g2_fill_1 FILLER_27_867 ();
 sg13g2_fill_2 FILLER_27_873 ();
 sg13g2_decap_4 FILLER_27_890 ();
 sg13g2_fill_1 FILLER_27_894 ();
 sg13g2_fill_1 FILLER_27_916 ();
 sg13g2_fill_1 FILLER_27_933 ();
 sg13g2_decap_8 FILLER_27_939 ();
 sg13g2_decap_4 FILLER_27_946 ();
 sg13g2_fill_2 FILLER_27_950 ();
 sg13g2_fill_2 FILLER_27_965 ();
 sg13g2_fill_1 FILLER_27_967 ();
 sg13g2_decap_8 FILLER_27_1031 ();
 sg13g2_decap_8 FILLER_27_1038 ();
 sg13g2_decap_8 FILLER_27_1045 ();
 sg13g2_decap_8 FILLER_27_1052 ();
 sg13g2_decap_8 FILLER_27_1059 ();
 sg13g2_decap_8 FILLER_27_1066 ();
 sg13g2_decap_8 FILLER_27_1073 ();
 sg13g2_decap_8 FILLER_27_1080 ();
 sg13g2_decap_8 FILLER_27_1087 ();
 sg13g2_decap_8 FILLER_27_1094 ();
 sg13g2_decap_8 FILLER_27_1101 ();
 sg13g2_decap_8 FILLER_27_1108 ();
 sg13g2_decap_8 FILLER_27_1115 ();
 sg13g2_decap_8 FILLER_27_1122 ();
 sg13g2_decap_8 FILLER_27_1129 ();
 sg13g2_decap_8 FILLER_27_1136 ();
 sg13g2_decap_8 FILLER_27_1143 ();
 sg13g2_decap_8 FILLER_27_1150 ();
 sg13g2_decap_8 FILLER_27_1157 ();
 sg13g2_decap_8 FILLER_27_1164 ();
 sg13g2_decap_8 FILLER_27_1171 ();
 sg13g2_decap_8 FILLER_27_1178 ();
 sg13g2_decap_8 FILLER_27_1185 ();
 sg13g2_decap_8 FILLER_27_1192 ();
 sg13g2_decap_8 FILLER_27_1199 ();
 sg13g2_decap_8 FILLER_27_1206 ();
 sg13g2_decap_8 FILLER_27_1213 ();
 sg13g2_decap_8 FILLER_27_1220 ();
 sg13g2_decap_8 FILLER_27_1227 ();
 sg13g2_decap_8 FILLER_27_1234 ();
 sg13g2_decap_8 FILLER_27_1241 ();
 sg13g2_decap_8 FILLER_27_1248 ();
 sg13g2_decap_8 FILLER_27_1255 ();
 sg13g2_decap_8 FILLER_27_1262 ();
 sg13g2_decap_8 FILLER_27_1269 ();
 sg13g2_decap_8 FILLER_27_1276 ();
 sg13g2_decap_8 FILLER_27_1283 ();
 sg13g2_decap_8 FILLER_27_1290 ();
 sg13g2_decap_8 FILLER_27_1297 ();
 sg13g2_decap_8 FILLER_27_1304 ();
 sg13g2_decap_4 FILLER_27_1311 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_107 ();
 sg13g2_fill_2 FILLER_28_138 ();
 sg13g2_fill_1 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_154 ();
 sg13g2_fill_1 FILLER_28_184 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_367 ();
 sg13g2_fill_1 FILLER_28_394 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_28_440 ();
 sg13g2_decap_4 FILLER_28_503 ();
 sg13g2_fill_1 FILLER_28_507 ();
 sg13g2_fill_2 FILLER_28_586 ();
 sg13g2_fill_1 FILLER_28_588 ();
 sg13g2_fill_1 FILLER_28_626 ();
 sg13g2_fill_2 FILLER_28_637 ();
 sg13g2_fill_1 FILLER_28_639 ();
 sg13g2_fill_1 FILLER_28_649 ();
 sg13g2_decap_4 FILLER_28_656 ();
 sg13g2_fill_2 FILLER_28_660 ();
 sg13g2_decap_8 FILLER_28_693 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_4 FILLER_28_720 ();
 sg13g2_decap_8 FILLER_28_738 ();
 sg13g2_fill_1 FILLER_28_754 ();
 sg13g2_decap_8 FILLER_28_771 ();
 sg13g2_fill_2 FILLER_28_778 ();
 sg13g2_decap_8 FILLER_28_801 ();
 sg13g2_fill_1 FILLER_28_808 ();
 sg13g2_decap_8 FILLER_28_835 ();
 sg13g2_decap_8 FILLER_28_842 ();
 sg13g2_fill_2 FILLER_28_849 ();
 sg13g2_decap_4 FILLER_28_861 ();
 sg13g2_fill_1 FILLER_28_865 ();
 sg13g2_fill_2 FILLER_28_871 ();
 sg13g2_fill_1 FILLER_28_882 ();
 sg13g2_fill_1 FILLER_28_887 ();
 sg13g2_decap_4 FILLER_28_913 ();
 sg13g2_decap_4 FILLER_28_931 ();
 sg13g2_decap_4 FILLER_28_947 ();
 sg13g2_decap_8 FILLER_28_955 ();
 sg13g2_fill_1 FILLER_28_962 ();
 sg13g2_fill_2 FILLER_28_1009 ();
 sg13g2_fill_1 FILLER_28_1011 ();
 sg13g2_decap_8 FILLER_28_1028 ();
 sg13g2_decap_8 FILLER_28_1035 ();
 sg13g2_decap_8 FILLER_28_1042 ();
 sg13g2_decap_8 FILLER_28_1049 ();
 sg13g2_decap_8 FILLER_28_1056 ();
 sg13g2_decap_8 FILLER_28_1063 ();
 sg13g2_decap_8 FILLER_28_1070 ();
 sg13g2_decap_8 FILLER_28_1077 ();
 sg13g2_decap_8 FILLER_28_1084 ();
 sg13g2_decap_8 FILLER_28_1091 ();
 sg13g2_decap_8 FILLER_28_1098 ();
 sg13g2_decap_8 FILLER_28_1105 ();
 sg13g2_decap_8 FILLER_28_1112 ();
 sg13g2_decap_8 FILLER_28_1119 ();
 sg13g2_decap_8 FILLER_28_1126 ();
 sg13g2_decap_8 FILLER_28_1133 ();
 sg13g2_decap_8 FILLER_28_1140 ();
 sg13g2_decap_8 FILLER_28_1147 ();
 sg13g2_decap_8 FILLER_28_1154 ();
 sg13g2_decap_8 FILLER_28_1161 ();
 sg13g2_decap_8 FILLER_28_1168 ();
 sg13g2_decap_8 FILLER_28_1175 ();
 sg13g2_decap_8 FILLER_28_1182 ();
 sg13g2_decap_8 FILLER_28_1189 ();
 sg13g2_decap_8 FILLER_28_1196 ();
 sg13g2_decap_8 FILLER_28_1203 ();
 sg13g2_decap_8 FILLER_28_1210 ();
 sg13g2_decap_8 FILLER_28_1217 ();
 sg13g2_decap_8 FILLER_28_1224 ();
 sg13g2_decap_8 FILLER_28_1231 ();
 sg13g2_decap_8 FILLER_28_1238 ();
 sg13g2_decap_8 FILLER_28_1245 ();
 sg13g2_decap_8 FILLER_28_1252 ();
 sg13g2_decap_8 FILLER_28_1259 ();
 sg13g2_decap_8 FILLER_28_1266 ();
 sg13g2_decap_8 FILLER_28_1273 ();
 sg13g2_decap_8 FILLER_28_1280 ();
 sg13g2_decap_8 FILLER_28_1287 ();
 sg13g2_decap_8 FILLER_28_1294 ();
 sg13g2_decap_8 FILLER_28_1301 ();
 sg13g2_decap_8 FILLER_28_1308 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_96 ();
 sg13g2_fill_2 FILLER_29_160 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_decap_4 FILLER_29_188 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_207 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_244 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_262 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_373 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_2 FILLER_29_474 ();
 sg13g2_fill_1 FILLER_29_476 ();
 sg13g2_fill_1 FILLER_29_486 ();
 sg13g2_decap_8 FILLER_29_495 ();
 sg13g2_decap_4 FILLER_29_502 ();
 sg13g2_fill_2 FILLER_29_536 ();
 sg13g2_decap_8 FILLER_29_543 ();
 sg13g2_fill_1 FILLER_29_550 ();
 sg13g2_decap_8 FILLER_29_555 ();
 sg13g2_decap_8 FILLER_29_562 ();
 sg13g2_fill_1 FILLER_29_569 ();
 sg13g2_decap_4 FILLER_29_574 ();
 sg13g2_fill_2 FILLER_29_578 ();
 sg13g2_fill_2 FILLER_29_588 ();
 sg13g2_decap_4 FILLER_29_609 ();
 sg13g2_decap_4 FILLER_29_621 ();
 sg13g2_fill_2 FILLER_29_643 ();
 sg13g2_fill_1 FILLER_29_652 ();
 sg13g2_fill_2 FILLER_29_667 ();
 sg13g2_fill_1 FILLER_29_669 ();
 sg13g2_fill_1 FILLER_29_678 ();
 sg13g2_fill_2 FILLER_29_695 ();
 sg13g2_fill_1 FILLER_29_697 ();
 sg13g2_fill_2 FILLER_29_720 ();
 sg13g2_fill_1 FILLER_29_722 ();
 sg13g2_fill_2 FILLER_29_738 ();
 sg13g2_fill_1 FILLER_29_740 ();
 sg13g2_fill_2 FILLER_29_751 ();
 sg13g2_fill_1 FILLER_29_753 ();
 sg13g2_fill_2 FILLER_29_760 ();
 sg13g2_fill_2 FILLER_29_771 ();
 sg13g2_decap_8 FILLER_29_788 ();
 sg13g2_fill_1 FILLER_29_805 ();
 sg13g2_decap_4 FILLER_29_810 ();
 sg13g2_fill_1 FILLER_29_814 ();
 sg13g2_fill_2 FILLER_29_829 ();
 sg13g2_fill_2 FILLER_29_861 ();
 sg13g2_fill_1 FILLER_29_863 ();
 sg13g2_fill_2 FILLER_29_894 ();
 sg13g2_decap_4 FILLER_29_913 ();
 sg13g2_decap_8 FILLER_29_927 ();
 sg13g2_fill_1 FILLER_29_934 ();
 sg13g2_fill_1 FILLER_29_939 ();
 sg13g2_fill_2 FILLER_29_966 ();
 sg13g2_fill_1 FILLER_29_979 ();
 sg13g2_fill_1 FILLER_29_998 ();
 sg13g2_fill_1 FILLER_29_1016 ();
 sg13g2_decap_8 FILLER_29_1043 ();
 sg13g2_decap_8 FILLER_29_1050 ();
 sg13g2_decap_8 FILLER_29_1057 ();
 sg13g2_decap_8 FILLER_29_1064 ();
 sg13g2_decap_8 FILLER_29_1071 ();
 sg13g2_decap_8 FILLER_29_1078 ();
 sg13g2_decap_8 FILLER_29_1085 ();
 sg13g2_decap_8 FILLER_29_1092 ();
 sg13g2_decap_8 FILLER_29_1099 ();
 sg13g2_decap_8 FILLER_29_1106 ();
 sg13g2_decap_8 FILLER_29_1113 ();
 sg13g2_decap_8 FILLER_29_1120 ();
 sg13g2_decap_8 FILLER_29_1127 ();
 sg13g2_decap_8 FILLER_29_1134 ();
 sg13g2_decap_8 FILLER_29_1141 ();
 sg13g2_decap_8 FILLER_29_1148 ();
 sg13g2_decap_8 FILLER_29_1155 ();
 sg13g2_decap_8 FILLER_29_1162 ();
 sg13g2_decap_8 FILLER_29_1169 ();
 sg13g2_decap_8 FILLER_29_1176 ();
 sg13g2_decap_8 FILLER_29_1183 ();
 sg13g2_decap_8 FILLER_29_1190 ();
 sg13g2_decap_8 FILLER_29_1197 ();
 sg13g2_decap_8 FILLER_29_1204 ();
 sg13g2_decap_8 FILLER_29_1211 ();
 sg13g2_decap_8 FILLER_29_1218 ();
 sg13g2_decap_8 FILLER_29_1225 ();
 sg13g2_decap_8 FILLER_29_1232 ();
 sg13g2_decap_8 FILLER_29_1239 ();
 sg13g2_decap_8 FILLER_29_1246 ();
 sg13g2_decap_8 FILLER_29_1253 ();
 sg13g2_decap_8 FILLER_29_1260 ();
 sg13g2_decap_8 FILLER_29_1267 ();
 sg13g2_decap_8 FILLER_29_1274 ();
 sg13g2_decap_8 FILLER_29_1281 ();
 sg13g2_decap_8 FILLER_29_1288 ();
 sg13g2_decap_8 FILLER_29_1295 ();
 sg13g2_decap_8 FILLER_29_1302 ();
 sg13g2_decap_4 FILLER_29_1309 ();
 sg13g2_fill_2 FILLER_29_1313 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_4 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_227 ();
 sg13g2_fill_2 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_decap_4 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_307 ();
 sg13g2_decap_8 FILLER_30_330 ();
 sg13g2_decap_4 FILLER_30_337 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_8 FILLER_30_404 ();
 sg13g2_fill_2 FILLER_30_411 ();
 sg13g2_decap_4 FILLER_30_446 ();
 sg13g2_fill_1 FILLER_30_450 ();
 sg13g2_fill_1 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_534 ();
 sg13g2_decap_4 FILLER_30_541 ();
 sg13g2_fill_2 FILLER_30_545 ();
 sg13g2_fill_2 FILLER_30_577 ();
 sg13g2_fill_2 FILLER_30_586 ();
 sg13g2_fill_1 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_610 ();
 sg13g2_fill_2 FILLER_30_617 ();
 sg13g2_fill_1 FILLER_30_634 ();
 sg13g2_fill_2 FILLER_30_653 ();
 sg13g2_fill_1 FILLER_30_655 ();
 sg13g2_fill_2 FILLER_30_668 ();
 sg13g2_fill_1 FILLER_30_670 ();
 sg13g2_fill_2 FILLER_30_675 ();
 sg13g2_fill_1 FILLER_30_677 ();
 sg13g2_decap_8 FILLER_30_684 ();
 sg13g2_fill_1 FILLER_30_691 ();
 sg13g2_decap_4 FILLER_30_700 ();
 sg13g2_fill_2 FILLER_30_712 ();
 sg13g2_fill_1 FILLER_30_720 ();
 sg13g2_decap_4 FILLER_30_731 ();
 sg13g2_fill_1 FILLER_30_735 ();
 sg13g2_fill_1 FILLER_30_741 ();
 sg13g2_fill_2 FILLER_30_755 ();
 sg13g2_decap_4 FILLER_30_789 ();
 sg13g2_decap_8 FILLER_30_806 ();
 sg13g2_decap_8 FILLER_30_813 ();
 sg13g2_fill_1 FILLER_30_820 ();
 sg13g2_decap_8 FILLER_30_827 ();
 sg13g2_fill_2 FILLER_30_834 ();
 sg13g2_decap_8 FILLER_30_845 ();
 sg13g2_fill_2 FILLER_30_856 ();
 sg13g2_decap_8 FILLER_30_863 ();
 sg13g2_decap_8 FILLER_30_870 ();
 sg13g2_decap_4 FILLER_30_882 ();
 sg13g2_fill_2 FILLER_30_895 ();
 sg13g2_fill_1 FILLER_30_897 ();
 sg13g2_fill_2 FILLER_30_902 ();
 sg13g2_fill_1 FILLER_30_904 ();
 sg13g2_fill_2 FILLER_30_922 ();
 sg13g2_fill_2 FILLER_30_950 ();
 sg13g2_fill_2 FILLER_30_960 ();
 sg13g2_fill_2 FILLER_30_970 ();
 sg13g2_fill_1 FILLER_30_972 ();
 sg13g2_fill_1 FILLER_30_1025 ();
 sg13g2_decap_8 FILLER_30_1034 ();
 sg13g2_decap_8 FILLER_30_1041 ();
 sg13g2_decap_8 FILLER_30_1048 ();
 sg13g2_decap_8 FILLER_30_1055 ();
 sg13g2_decap_8 FILLER_30_1062 ();
 sg13g2_decap_8 FILLER_30_1069 ();
 sg13g2_decap_8 FILLER_30_1076 ();
 sg13g2_decap_8 FILLER_30_1083 ();
 sg13g2_decap_8 FILLER_30_1090 ();
 sg13g2_decap_8 FILLER_30_1097 ();
 sg13g2_decap_8 FILLER_30_1104 ();
 sg13g2_decap_8 FILLER_30_1111 ();
 sg13g2_decap_8 FILLER_30_1118 ();
 sg13g2_decap_8 FILLER_30_1125 ();
 sg13g2_decap_8 FILLER_30_1132 ();
 sg13g2_decap_8 FILLER_30_1139 ();
 sg13g2_decap_8 FILLER_30_1146 ();
 sg13g2_decap_8 FILLER_30_1153 ();
 sg13g2_decap_8 FILLER_30_1160 ();
 sg13g2_decap_8 FILLER_30_1167 ();
 sg13g2_decap_8 FILLER_30_1174 ();
 sg13g2_decap_8 FILLER_30_1181 ();
 sg13g2_decap_8 FILLER_30_1188 ();
 sg13g2_decap_8 FILLER_30_1195 ();
 sg13g2_decap_8 FILLER_30_1202 ();
 sg13g2_decap_8 FILLER_30_1209 ();
 sg13g2_decap_8 FILLER_30_1216 ();
 sg13g2_decap_8 FILLER_30_1223 ();
 sg13g2_decap_8 FILLER_30_1230 ();
 sg13g2_decap_8 FILLER_30_1237 ();
 sg13g2_decap_8 FILLER_30_1244 ();
 sg13g2_decap_8 FILLER_30_1251 ();
 sg13g2_decap_8 FILLER_30_1258 ();
 sg13g2_decap_8 FILLER_30_1265 ();
 sg13g2_decap_8 FILLER_30_1272 ();
 sg13g2_decap_8 FILLER_30_1279 ();
 sg13g2_decap_8 FILLER_30_1286 ();
 sg13g2_decap_8 FILLER_30_1293 ();
 sg13g2_decap_8 FILLER_30_1300 ();
 sg13g2_decap_8 FILLER_30_1307 ();
 sg13g2_fill_1 FILLER_30_1314 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_137 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_197 ();
 sg13g2_decap_4 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_decap_4 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_fill_2 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_2 FILLER_31_409 ();
 sg13g2_decap_4 FILLER_31_416 ();
 sg13g2_fill_1 FILLER_31_425 ();
 sg13g2_decap_4 FILLER_31_438 ();
 sg13g2_fill_1 FILLER_31_442 ();
 sg13g2_decap_4 FILLER_31_448 ();
 sg13g2_fill_2 FILLER_31_490 ();
 sg13g2_fill_2 FILLER_31_501 ();
 sg13g2_fill_1 FILLER_31_503 ();
 sg13g2_fill_2 FILLER_31_529 ();
 sg13g2_fill_1 FILLER_31_531 ();
 sg13g2_fill_1 FILLER_31_566 ();
 sg13g2_decap_4 FILLER_31_597 ();
 sg13g2_fill_2 FILLER_31_601 ();
 sg13g2_fill_1 FILLER_31_626 ();
 sg13g2_decap_4 FILLER_31_640 ();
 sg13g2_fill_2 FILLER_31_680 ();
 sg13g2_fill_2 FILLER_31_707 ();
 sg13g2_fill_2 FILLER_31_714 ();
 sg13g2_fill_1 FILLER_31_716 ();
 sg13g2_decap_4 FILLER_31_741 ();
 sg13g2_decap_4 FILLER_31_748 ();
 sg13g2_fill_1 FILLER_31_752 ();
 sg13g2_decap_8 FILLER_31_761 ();
 sg13g2_decap_4 FILLER_31_768 ();
 sg13g2_fill_1 FILLER_31_772 ();
 sg13g2_decap_8 FILLER_31_778 ();
 sg13g2_fill_2 FILLER_31_785 ();
 sg13g2_decap_4 FILLER_31_795 ();
 sg13g2_decap_8 FILLER_31_804 ();
 sg13g2_fill_2 FILLER_31_828 ();
 sg13g2_fill_1 FILLER_31_843 ();
 sg13g2_fill_2 FILLER_31_867 ();
 sg13g2_fill_2 FILLER_31_886 ();
 sg13g2_fill_2 FILLER_31_909 ();
 sg13g2_fill_2 FILLER_31_921 ();
 sg13g2_fill_1 FILLER_31_923 ();
 sg13g2_decap_4 FILLER_31_928 ();
 sg13g2_fill_2 FILLER_31_932 ();
 sg13g2_fill_2 FILLER_31_948 ();
 sg13g2_fill_2 FILLER_31_1005 ();
 sg13g2_fill_1 FILLER_31_1007 ();
 sg13g2_decap_8 FILLER_31_1062 ();
 sg13g2_decap_8 FILLER_31_1069 ();
 sg13g2_decap_8 FILLER_31_1076 ();
 sg13g2_decap_8 FILLER_31_1083 ();
 sg13g2_decap_8 FILLER_31_1090 ();
 sg13g2_decap_8 FILLER_31_1097 ();
 sg13g2_decap_8 FILLER_31_1104 ();
 sg13g2_decap_8 FILLER_31_1111 ();
 sg13g2_decap_8 FILLER_31_1118 ();
 sg13g2_decap_8 FILLER_31_1125 ();
 sg13g2_decap_8 FILLER_31_1132 ();
 sg13g2_decap_8 FILLER_31_1139 ();
 sg13g2_decap_8 FILLER_31_1146 ();
 sg13g2_decap_8 FILLER_31_1153 ();
 sg13g2_decap_8 FILLER_31_1160 ();
 sg13g2_decap_8 FILLER_31_1167 ();
 sg13g2_decap_8 FILLER_31_1174 ();
 sg13g2_decap_8 FILLER_31_1181 ();
 sg13g2_decap_8 FILLER_31_1188 ();
 sg13g2_decap_8 FILLER_31_1195 ();
 sg13g2_decap_8 FILLER_31_1202 ();
 sg13g2_decap_8 FILLER_31_1209 ();
 sg13g2_decap_8 FILLER_31_1216 ();
 sg13g2_decap_8 FILLER_31_1223 ();
 sg13g2_decap_8 FILLER_31_1230 ();
 sg13g2_decap_8 FILLER_31_1237 ();
 sg13g2_decap_8 FILLER_31_1244 ();
 sg13g2_decap_8 FILLER_31_1251 ();
 sg13g2_decap_8 FILLER_31_1258 ();
 sg13g2_decap_8 FILLER_31_1265 ();
 sg13g2_decap_8 FILLER_31_1272 ();
 sg13g2_decap_8 FILLER_31_1279 ();
 sg13g2_decap_8 FILLER_31_1286 ();
 sg13g2_decap_8 FILLER_31_1293 ();
 sg13g2_decap_8 FILLER_31_1300 ();
 sg13g2_decap_8 FILLER_31_1307 ();
 sg13g2_fill_1 FILLER_31_1314 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_135 ();
 sg13g2_decap_8 FILLER_32_146 ();
 sg13g2_fill_2 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_164 ();
 sg13g2_decap_8 FILLER_32_178 ();
 sg13g2_fill_2 FILLER_32_194 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_decap_4 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_320 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_32_402 ();
 sg13g2_fill_1 FILLER_32_404 ();
 sg13g2_decap_4 FILLER_32_431 ();
 sg13g2_fill_2 FILLER_32_461 ();
 sg13g2_fill_1 FILLER_32_463 ();
 sg13g2_fill_2 FILLER_32_498 ();
 sg13g2_fill_1 FILLER_32_500 ();
 sg13g2_fill_2 FILLER_32_509 ();
 sg13g2_decap_4 FILLER_32_524 ();
 sg13g2_fill_2 FILLER_32_532 ();
 sg13g2_fill_1 FILLER_32_534 ();
 sg13g2_fill_2 FILLER_32_545 ();
 sg13g2_fill_2 FILLER_32_577 ();
 sg13g2_decap_8 FILLER_32_584 ();
 sg13g2_decap_4 FILLER_32_595 ();
 sg13g2_fill_1 FILLER_32_599 ();
 sg13g2_decap_8 FILLER_32_607 ();
 sg13g2_decap_8 FILLER_32_633 ();
 sg13g2_decap_8 FILLER_32_640 ();
 sg13g2_fill_1 FILLER_32_647 ();
 sg13g2_decap_8 FILLER_32_657 ();
 sg13g2_fill_2 FILLER_32_664 ();
 sg13g2_fill_1 FILLER_32_666 ();
 sg13g2_decap_8 FILLER_32_672 ();
 sg13g2_fill_2 FILLER_32_679 ();
 sg13g2_fill_1 FILLER_32_681 ();
 sg13g2_fill_2 FILLER_32_690 ();
 sg13g2_fill_2 FILLER_32_703 ();
 sg13g2_fill_2 FILLER_32_725 ();
 sg13g2_fill_1 FILLER_32_727 ();
 sg13g2_fill_1 FILLER_32_763 ();
 sg13g2_fill_2 FILLER_32_768 ();
 sg13g2_fill_1 FILLER_32_775 ();
 sg13g2_fill_1 FILLER_32_791 ();
 sg13g2_decap_4 FILLER_32_802 ();
 sg13g2_decap_8 FILLER_32_810 ();
 sg13g2_fill_1 FILLER_32_832 ();
 sg13g2_fill_2 FILLER_32_853 ();
 sg13g2_fill_1 FILLER_32_855 ();
 sg13g2_decap_4 FILLER_32_876 ();
 sg13g2_fill_1 FILLER_32_880 ();
 sg13g2_decap_4 FILLER_32_886 ();
 sg13g2_fill_1 FILLER_32_890 ();
 sg13g2_fill_2 FILLER_32_895 ();
 sg13g2_fill_2 FILLER_32_919 ();
 sg13g2_fill_2 FILLER_32_931 ();
 sg13g2_fill_1 FILLER_32_933 ();
 sg13g2_fill_2 FILLER_32_953 ();
 sg13g2_fill_2 FILLER_32_970 ();
 sg13g2_fill_1 FILLER_32_972 ();
 sg13g2_decap_8 FILLER_32_1061 ();
 sg13g2_decap_8 FILLER_32_1068 ();
 sg13g2_decap_8 FILLER_32_1075 ();
 sg13g2_decap_8 FILLER_32_1082 ();
 sg13g2_decap_8 FILLER_32_1089 ();
 sg13g2_decap_8 FILLER_32_1096 ();
 sg13g2_decap_8 FILLER_32_1103 ();
 sg13g2_decap_8 FILLER_32_1110 ();
 sg13g2_decap_8 FILLER_32_1117 ();
 sg13g2_decap_8 FILLER_32_1124 ();
 sg13g2_decap_8 FILLER_32_1131 ();
 sg13g2_decap_8 FILLER_32_1138 ();
 sg13g2_decap_8 FILLER_32_1145 ();
 sg13g2_decap_8 FILLER_32_1152 ();
 sg13g2_decap_8 FILLER_32_1159 ();
 sg13g2_decap_8 FILLER_32_1166 ();
 sg13g2_decap_8 FILLER_32_1173 ();
 sg13g2_decap_8 FILLER_32_1180 ();
 sg13g2_decap_8 FILLER_32_1187 ();
 sg13g2_decap_8 FILLER_32_1194 ();
 sg13g2_decap_8 FILLER_32_1201 ();
 sg13g2_decap_8 FILLER_32_1208 ();
 sg13g2_decap_8 FILLER_32_1215 ();
 sg13g2_decap_8 FILLER_32_1222 ();
 sg13g2_decap_8 FILLER_32_1229 ();
 sg13g2_decap_8 FILLER_32_1236 ();
 sg13g2_decap_8 FILLER_32_1243 ();
 sg13g2_decap_8 FILLER_32_1250 ();
 sg13g2_decap_8 FILLER_32_1257 ();
 sg13g2_decap_8 FILLER_32_1264 ();
 sg13g2_decap_8 FILLER_32_1271 ();
 sg13g2_decap_8 FILLER_32_1278 ();
 sg13g2_decap_8 FILLER_32_1285 ();
 sg13g2_decap_8 FILLER_32_1292 ();
 sg13g2_decap_8 FILLER_32_1299 ();
 sg13g2_decap_8 FILLER_32_1306 ();
 sg13g2_fill_2 FILLER_32_1313 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_1 FILLER_33_100 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_143 ();
 sg13g2_fill_1 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_256 ();
 sg13g2_decap_4 FILLER_33_261 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_decap_4 FILLER_33_314 ();
 sg13g2_decap_4 FILLER_33_331 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_4 FILLER_33_380 ();
 sg13g2_fill_2 FILLER_33_384 ();
 sg13g2_fill_2 FILLER_33_403 ();
 sg13g2_fill_1 FILLER_33_405 ();
 sg13g2_fill_1 FILLER_33_443 ();
 sg13g2_decap_4 FILLER_33_469 ();
 sg13g2_fill_1 FILLER_33_498 ();
 sg13g2_fill_2 FILLER_33_535 ();
 sg13g2_decap_8 FILLER_33_554 ();
 sg13g2_decap_4 FILLER_33_561 ();
 sg13g2_fill_2 FILLER_33_565 ();
 sg13g2_fill_1 FILLER_33_619 ();
 sg13g2_decap_4 FILLER_33_642 ();
 sg13g2_decap_8 FILLER_33_680 ();
 sg13g2_fill_1 FILLER_33_687 ();
 sg13g2_fill_2 FILLER_33_693 ();
 sg13g2_fill_2 FILLER_33_701 ();
 sg13g2_fill_2 FILLER_33_709 ();
 sg13g2_fill_2 FILLER_33_731 ();
 sg13g2_fill_1 FILLER_33_733 ();
 sg13g2_decap_4 FILLER_33_739 ();
 sg13g2_fill_1 FILLER_33_743 ();
 sg13g2_fill_1 FILLER_33_747 ();
 sg13g2_fill_1 FILLER_33_758 ();
 sg13g2_fill_1 FILLER_33_786 ();
 sg13g2_fill_2 FILLER_33_792 ();
 sg13g2_fill_2 FILLER_33_808 ();
 sg13g2_fill_2 FILLER_33_818 ();
 sg13g2_decap_4 FILLER_33_828 ();
 sg13g2_fill_2 FILLER_33_832 ();
 sg13g2_fill_2 FILLER_33_843 ();
 sg13g2_decap_4 FILLER_33_855 ();
 sg13g2_fill_2 FILLER_33_859 ();
 sg13g2_fill_2 FILLER_33_878 ();
 sg13g2_decap_4 FILLER_33_897 ();
 sg13g2_fill_2 FILLER_33_901 ();
 sg13g2_fill_1 FILLER_33_911 ();
 sg13g2_decap_8 FILLER_33_934 ();
 sg13g2_fill_2 FILLER_33_950 ();
 sg13g2_fill_2 FILLER_33_965 ();
 sg13g2_fill_1 FILLER_33_967 ();
 sg13g2_decap_4 FILLER_33_973 ();
 sg13g2_fill_2 FILLER_33_985 ();
 sg13g2_fill_1 FILLER_33_987 ();
 sg13g2_decap_8 FILLER_33_1028 ();
 sg13g2_decap_4 FILLER_33_1035 ();
 sg13g2_decap_8 FILLER_33_1043 ();
 sg13g2_decap_8 FILLER_33_1050 ();
 sg13g2_decap_8 FILLER_33_1057 ();
 sg13g2_decap_8 FILLER_33_1064 ();
 sg13g2_decap_8 FILLER_33_1071 ();
 sg13g2_decap_8 FILLER_33_1078 ();
 sg13g2_decap_8 FILLER_33_1085 ();
 sg13g2_decap_8 FILLER_33_1092 ();
 sg13g2_decap_8 FILLER_33_1099 ();
 sg13g2_decap_8 FILLER_33_1106 ();
 sg13g2_decap_8 FILLER_33_1113 ();
 sg13g2_decap_8 FILLER_33_1120 ();
 sg13g2_decap_8 FILLER_33_1127 ();
 sg13g2_decap_8 FILLER_33_1134 ();
 sg13g2_decap_8 FILLER_33_1141 ();
 sg13g2_decap_8 FILLER_33_1148 ();
 sg13g2_decap_8 FILLER_33_1155 ();
 sg13g2_decap_8 FILLER_33_1162 ();
 sg13g2_decap_8 FILLER_33_1169 ();
 sg13g2_decap_8 FILLER_33_1176 ();
 sg13g2_decap_8 FILLER_33_1183 ();
 sg13g2_decap_8 FILLER_33_1190 ();
 sg13g2_decap_8 FILLER_33_1197 ();
 sg13g2_decap_8 FILLER_33_1204 ();
 sg13g2_decap_8 FILLER_33_1211 ();
 sg13g2_decap_8 FILLER_33_1218 ();
 sg13g2_decap_8 FILLER_33_1225 ();
 sg13g2_decap_8 FILLER_33_1232 ();
 sg13g2_decap_8 FILLER_33_1239 ();
 sg13g2_decap_8 FILLER_33_1246 ();
 sg13g2_decap_8 FILLER_33_1253 ();
 sg13g2_decap_8 FILLER_33_1260 ();
 sg13g2_decap_8 FILLER_33_1267 ();
 sg13g2_decap_8 FILLER_33_1274 ();
 sg13g2_decap_8 FILLER_33_1281 ();
 sg13g2_decap_8 FILLER_33_1288 ();
 sg13g2_decap_8 FILLER_33_1295 ();
 sg13g2_decap_8 FILLER_33_1302 ();
 sg13g2_decap_4 FILLER_33_1309 ();
 sg13g2_fill_2 FILLER_33_1313 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_100 ();
 sg13g2_fill_2 FILLER_34_136 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_fill_2 FILLER_34_152 ();
 sg13g2_fill_1 FILLER_34_154 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_227 ();
 sg13g2_decap_4 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_267 ();
 sg13g2_fill_2 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_290 ();
 sg13g2_decap_8 FILLER_34_309 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_decap_4 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_fill_2 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_fill_2 FILLER_34_394 ();
 sg13g2_fill_1 FILLER_34_396 ();
 sg13g2_fill_2 FILLER_34_432 ();
 sg13g2_fill_1 FILLER_34_442 ();
 sg13g2_decap_8 FILLER_34_479 ();
 sg13g2_decap_8 FILLER_34_486 ();
 sg13g2_fill_2 FILLER_34_493 ();
 sg13g2_decap_4 FILLER_34_504 ();
 sg13g2_fill_2 FILLER_34_508 ();
 sg13g2_decap_4 FILLER_34_521 ();
 sg13g2_decap_4 FILLER_34_534 ();
 sg13g2_fill_1 FILLER_34_538 ();
 sg13g2_decap_8 FILLER_34_551 ();
 sg13g2_decap_8 FILLER_34_570 ();
 sg13g2_fill_1 FILLER_34_577 ();
 sg13g2_decap_4 FILLER_34_582 ();
 sg13g2_fill_2 FILLER_34_586 ();
 sg13g2_fill_2 FILLER_34_601 ();
 sg13g2_fill_1 FILLER_34_603 ();
 sg13g2_fill_1 FILLER_34_608 ();
 sg13g2_decap_8 FILLER_34_619 ();
 sg13g2_decap_8 FILLER_34_626 ();
 sg13g2_decap_4 FILLER_34_633 ();
 sg13g2_fill_2 FILLER_34_637 ();
 sg13g2_decap_4 FILLER_34_655 ();
 sg13g2_fill_2 FILLER_34_659 ();
 sg13g2_fill_2 FILLER_34_712 ();
 sg13g2_fill_1 FILLER_34_714 ();
 sg13g2_fill_2 FILLER_34_723 ();
 sg13g2_fill_1 FILLER_34_725 ();
 sg13g2_decap_4 FILLER_34_738 ();
 sg13g2_fill_1 FILLER_34_742 ();
 sg13g2_fill_1 FILLER_34_768 ();
 sg13g2_fill_1 FILLER_34_786 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_4 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_807 ();
 sg13g2_fill_2 FILLER_34_832 ();
 sg13g2_fill_2 FILLER_34_852 ();
 sg13g2_fill_1 FILLER_34_854 ();
 sg13g2_fill_2 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_34_875 ();
 sg13g2_decap_8 FILLER_34_890 ();
 sg13g2_fill_2 FILLER_34_897 ();
 sg13g2_fill_1 FILLER_34_909 ();
 sg13g2_decap_8 FILLER_34_915 ();
 sg13g2_fill_2 FILLER_34_927 ();
 sg13g2_fill_1 FILLER_34_929 ();
 sg13g2_fill_1 FILLER_34_939 ();
 sg13g2_fill_1 FILLER_34_950 ();
 sg13g2_fill_1 FILLER_34_969 ();
 sg13g2_decap_8 FILLER_34_1054 ();
 sg13g2_decap_8 FILLER_34_1061 ();
 sg13g2_decap_8 FILLER_34_1068 ();
 sg13g2_decap_8 FILLER_34_1075 ();
 sg13g2_decap_8 FILLER_34_1082 ();
 sg13g2_decap_8 FILLER_34_1089 ();
 sg13g2_decap_8 FILLER_34_1096 ();
 sg13g2_decap_8 FILLER_34_1103 ();
 sg13g2_decap_8 FILLER_34_1110 ();
 sg13g2_decap_8 FILLER_34_1117 ();
 sg13g2_decap_8 FILLER_34_1124 ();
 sg13g2_decap_8 FILLER_34_1131 ();
 sg13g2_decap_8 FILLER_34_1138 ();
 sg13g2_decap_8 FILLER_34_1145 ();
 sg13g2_decap_8 FILLER_34_1152 ();
 sg13g2_decap_8 FILLER_34_1159 ();
 sg13g2_decap_8 FILLER_34_1166 ();
 sg13g2_decap_8 FILLER_34_1173 ();
 sg13g2_decap_8 FILLER_34_1180 ();
 sg13g2_decap_8 FILLER_34_1187 ();
 sg13g2_decap_8 FILLER_34_1194 ();
 sg13g2_decap_8 FILLER_34_1201 ();
 sg13g2_decap_8 FILLER_34_1208 ();
 sg13g2_decap_8 FILLER_34_1215 ();
 sg13g2_decap_8 FILLER_34_1222 ();
 sg13g2_decap_8 FILLER_34_1229 ();
 sg13g2_decap_8 FILLER_34_1236 ();
 sg13g2_decap_8 FILLER_34_1243 ();
 sg13g2_decap_8 FILLER_34_1250 ();
 sg13g2_decap_8 FILLER_34_1257 ();
 sg13g2_decap_8 FILLER_34_1264 ();
 sg13g2_decap_8 FILLER_34_1271 ();
 sg13g2_decap_8 FILLER_34_1278 ();
 sg13g2_decap_8 FILLER_34_1285 ();
 sg13g2_decap_8 FILLER_34_1292 ();
 sg13g2_decap_8 FILLER_34_1299 ();
 sg13g2_decap_8 FILLER_34_1306 ();
 sg13g2_fill_2 FILLER_34_1313 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_fill_1 FILLER_35_127 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_146 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_decap_4 FILLER_35_159 ();
 sg13g2_fill_1 FILLER_35_163 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_fill_2 FILLER_35_174 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_fill_1 FILLER_35_247 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_1 FILLER_35_262 ();
 sg13g2_decap_8 FILLER_35_267 ();
 sg13g2_fill_1 FILLER_35_274 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_fill_1 FILLER_35_312 ();
 sg13g2_fill_2 FILLER_35_339 ();
 sg13g2_fill_1 FILLER_35_341 ();
 sg13g2_decap_4 FILLER_35_352 ();
 sg13g2_fill_2 FILLER_35_356 ();
 sg13g2_decap_4 FILLER_35_362 ();
 sg13g2_fill_1 FILLER_35_366 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_fill_2 FILLER_35_429 ();
 sg13g2_fill_1 FILLER_35_435 ();
 sg13g2_fill_1 FILLER_35_459 ();
 sg13g2_decap_8 FILLER_35_481 ();
 sg13g2_fill_2 FILLER_35_488 ();
 sg13g2_decap_4 FILLER_35_529 ();
 sg13g2_fill_2 FILLER_35_569 ();
 sg13g2_fill_1 FILLER_35_579 ();
 sg13g2_fill_2 FILLER_35_606 ();
 sg13g2_fill_1 FILLER_35_608 ();
 sg13g2_fill_1 FILLER_35_613 ();
 sg13g2_decap_8 FILLER_35_633 ();
 sg13g2_decap_8 FILLER_35_640 ();
 sg13g2_decap_8 FILLER_35_647 ();
 sg13g2_fill_2 FILLER_35_654 ();
 sg13g2_decap_8 FILLER_35_664 ();
 sg13g2_decap_8 FILLER_35_682 ();
 sg13g2_decap_4 FILLER_35_697 ();
 sg13g2_decap_8 FILLER_35_712 ();
 sg13g2_decap_8 FILLER_35_719 ();
 sg13g2_fill_2 FILLER_35_726 ();
 sg13g2_fill_1 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_738 ();
 sg13g2_fill_2 FILLER_35_745 ();
 sg13g2_fill_1 FILLER_35_747 ();
 sg13g2_decap_8 FILLER_35_757 ();
 sg13g2_fill_1 FILLER_35_764 ();
 sg13g2_decap_8 FILLER_35_785 ();
 sg13g2_fill_1 FILLER_35_810 ();
 sg13g2_decap_4 FILLER_35_816 ();
 sg13g2_fill_2 FILLER_35_820 ();
 sg13g2_decap_8 FILLER_35_834 ();
 sg13g2_decap_4 FILLER_35_841 ();
 sg13g2_fill_1 FILLER_35_845 ();
 sg13g2_decap_8 FILLER_35_850 ();
 sg13g2_decap_4 FILLER_35_857 ();
 sg13g2_fill_2 FILLER_35_861 ();
 sg13g2_fill_2 FILLER_35_867 ();
 sg13g2_fill_1 FILLER_35_869 ();
 sg13g2_decap_8 FILLER_35_925 ();
 sg13g2_fill_2 FILLER_35_947 ();
 sg13g2_decap_8 FILLER_35_967 ();
 sg13g2_decap_8 FILLER_35_974 ();
 sg13g2_decap_8 FILLER_35_981 ();
 sg13g2_fill_2 FILLER_35_993 ();
 sg13g2_fill_1 FILLER_35_995 ();
 sg13g2_fill_2 FILLER_35_1001 ();
 sg13g2_fill_2 FILLER_35_1029 ();
 sg13g2_fill_1 FILLER_35_1031 ();
 sg13g2_decap_8 FILLER_35_1058 ();
 sg13g2_decap_8 FILLER_35_1065 ();
 sg13g2_decap_8 FILLER_35_1072 ();
 sg13g2_decap_8 FILLER_35_1079 ();
 sg13g2_decap_8 FILLER_35_1086 ();
 sg13g2_decap_8 FILLER_35_1093 ();
 sg13g2_decap_8 FILLER_35_1100 ();
 sg13g2_decap_8 FILLER_35_1107 ();
 sg13g2_decap_8 FILLER_35_1114 ();
 sg13g2_decap_8 FILLER_35_1121 ();
 sg13g2_decap_8 FILLER_35_1128 ();
 sg13g2_decap_8 FILLER_35_1135 ();
 sg13g2_decap_8 FILLER_35_1142 ();
 sg13g2_decap_8 FILLER_35_1149 ();
 sg13g2_decap_8 FILLER_35_1156 ();
 sg13g2_decap_8 FILLER_35_1163 ();
 sg13g2_decap_8 FILLER_35_1170 ();
 sg13g2_decap_8 FILLER_35_1177 ();
 sg13g2_decap_8 FILLER_35_1184 ();
 sg13g2_decap_8 FILLER_35_1191 ();
 sg13g2_decap_8 FILLER_35_1198 ();
 sg13g2_decap_8 FILLER_35_1205 ();
 sg13g2_decap_8 FILLER_35_1212 ();
 sg13g2_decap_8 FILLER_35_1219 ();
 sg13g2_decap_8 FILLER_35_1226 ();
 sg13g2_decap_8 FILLER_35_1233 ();
 sg13g2_decap_8 FILLER_35_1240 ();
 sg13g2_decap_8 FILLER_35_1247 ();
 sg13g2_decap_8 FILLER_35_1254 ();
 sg13g2_decap_8 FILLER_35_1261 ();
 sg13g2_decap_8 FILLER_35_1268 ();
 sg13g2_decap_8 FILLER_35_1275 ();
 sg13g2_decap_8 FILLER_35_1282 ();
 sg13g2_decap_8 FILLER_35_1289 ();
 sg13g2_decap_8 FILLER_35_1296 ();
 sg13g2_decap_8 FILLER_35_1303 ();
 sg13g2_decap_4 FILLER_35_1310 ();
 sg13g2_fill_1 FILLER_35_1314 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_103 ();
 sg13g2_fill_1 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_155 ();
 sg13g2_fill_2 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_decap_4 FILLER_36_193 ();
 sg13g2_decap_4 FILLER_36_201 ();
 sg13g2_decap_4 FILLER_36_213 ();
 sg13g2_fill_2 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_243 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_fill_1 FILLER_36_389 ();
 sg13g2_decap_4 FILLER_36_394 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_fill_1 FILLER_36_425 ();
 sg13g2_fill_2 FILLER_36_461 ();
 sg13g2_fill_1 FILLER_36_463 ();
 sg13g2_fill_1 FILLER_36_490 ();
 sg13g2_decap_4 FILLER_36_495 ();
 sg13g2_fill_1 FILLER_36_499 ();
 sg13g2_decap_8 FILLER_36_505 ();
 sg13g2_fill_2 FILLER_36_512 ();
 sg13g2_decap_4 FILLER_36_518 ();
 sg13g2_fill_2 FILLER_36_522 ();
 sg13g2_fill_2 FILLER_36_532 ();
 sg13g2_fill_1 FILLER_36_534 ();
 sg13g2_fill_2 FILLER_36_539 ();
 sg13g2_fill_2 FILLER_36_545 ();
 sg13g2_decap_4 FILLER_36_555 ();
 sg13g2_fill_2 FILLER_36_559 ();
 sg13g2_fill_2 FILLER_36_587 ();
 sg13g2_fill_2 FILLER_36_598 ();
 sg13g2_fill_1 FILLER_36_600 ();
 sg13g2_fill_2 FILLER_36_645 ();
 sg13g2_decap_4 FILLER_36_660 ();
 sg13g2_fill_1 FILLER_36_664 ();
 sg13g2_fill_2 FILLER_36_681 ();
 sg13g2_fill_1 FILLER_36_683 ();
 sg13g2_fill_2 FILLER_36_688 ();
 sg13g2_fill_2 FILLER_36_695 ();
 sg13g2_decap_8 FILLER_36_706 ();
 sg13g2_decap_8 FILLER_36_713 ();
 sg13g2_fill_2 FILLER_36_730 ();
 sg13g2_fill_1 FILLER_36_740 ();
 sg13g2_fill_2 FILLER_36_758 ();
 sg13g2_fill_1 FILLER_36_765 ();
 sg13g2_fill_2 FILLER_36_771 ();
 sg13g2_fill_1 FILLER_36_773 ();
 sg13g2_decap_8 FILLER_36_778 ();
 sg13g2_decap_4 FILLER_36_790 ();
 sg13g2_decap_4 FILLER_36_818 ();
 sg13g2_decap_4 FILLER_36_831 ();
 sg13g2_fill_2 FILLER_36_845 ();
 sg13g2_decap_4 FILLER_36_869 ();
 sg13g2_decap_8 FILLER_36_886 ();
 sg13g2_decap_4 FILLER_36_893 ();
 sg13g2_fill_1 FILLER_36_897 ();
 sg13g2_decap_4 FILLER_36_902 ();
 sg13g2_fill_1 FILLER_36_930 ();
 sg13g2_fill_1 FILLER_36_954 ();
 sg13g2_decap_4 FILLER_36_962 ();
 sg13g2_decap_8 FILLER_36_1052 ();
 sg13g2_decap_8 FILLER_36_1059 ();
 sg13g2_decap_8 FILLER_36_1066 ();
 sg13g2_decap_8 FILLER_36_1073 ();
 sg13g2_decap_8 FILLER_36_1080 ();
 sg13g2_decap_8 FILLER_36_1087 ();
 sg13g2_decap_8 FILLER_36_1094 ();
 sg13g2_decap_8 FILLER_36_1101 ();
 sg13g2_decap_8 FILLER_36_1108 ();
 sg13g2_decap_8 FILLER_36_1115 ();
 sg13g2_decap_8 FILLER_36_1122 ();
 sg13g2_decap_8 FILLER_36_1129 ();
 sg13g2_decap_8 FILLER_36_1136 ();
 sg13g2_decap_8 FILLER_36_1143 ();
 sg13g2_decap_8 FILLER_36_1150 ();
 sg13g2_decap_8 FILLER_36_1157 ();
 sg13g2_decap_8 FILLER_36_1164 ();
 sg13g2_decap_8 FILLER_36_1171 ();
 sg13g2_decap_8 FILLER_36_1178 ();
 sg13g2_decap_8 FILLER_36_1185 ();
 sg13g2_decap_8 FILLER_36_1192 ();
 sg13g2_decap_8 FILLER_36_1199 ();
 sg13g2_decap_8 FILLER_36_1206 ();
 sg13g2_decap_8 FILLER_36_1213 ();
 sg13g2_decap_8 FILLER_36_1220 ();
 sg13g2_decap_8 FILLER_36_1227 ();
 sg13g2_decap_8 FILLER_36_1234 ();
 sg13g2_decap_8 FILLER_36_1241 ();
 sg13g2_decap_8 FILLER_36_1248 ();
 sg13g2_decap_8 FILLER_36_1255 ();
 sg13g2_decap_8 FILLER_36_1262 ();
 sg13g2_decap_8 FILLER_36_1269 ();
 sg13g2_decap_8 FILLER_36_1276 ();
 sg13g2_decap_8 FILLER_36_1283 ();
 sg13g2_decap_8 FILLER_36_1290 ();
 sg13g2_decap_8 FILLER_36_1297 ();
 sg13g2_decap_8 FILLER_36_1304 ();
 sg13g2_decap_4 FILLER_36_1311 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_114 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_121 ();
 sg13g2_fill_1 FILLER_37_140 ();
 sg13g2_fill_1 FILLER_37_198 ();
 sg13g2_fill_2 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_fill_2 FILLER_37_259 ();
 sg13g2_fill_1 FILLER_37_261 ();
 sg13g2_fill_2 FILLER_37_266 ();
 sg13g2_decap_4 FILLER_37_317 ();
 sg13g2_fill_1 FILLER_37_321 ();
 sg13g2_fill_2 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_345 ();
 sg13g2_decap_4 FILLER_37_350 ();
 sg13g2_fill_2 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_decap_8 FILLER_37_431 ();
 sg13g2_decap_8 FILLER_37_442 ();
 sg13g2_decap_8 FILLER_37_449 ();
 sg13g2_fill_1 FILLER_37_468 ();
 sg13g2_fill_1 FILLER_37_474 ();
 sg13g2_fill_1 FILLER_37_479 ();
 sg13g2_fill_2 FILLER_37_515 ();
 sg13g2_fill_1 FILLER_37_517 ();
 sg13g2_fill_1 FILLER_37_523 ();
 sg13g2_fill_2 FILLER_37_534 ();
 sg13g2_fill_1 FILLER_37_562 ();
 sg13g2_decap_8 FILLER_37_568 ();
 sg13g2_fill_1 FILLER_37_586 ();
 sg13g2_decap_4 FILLER_37_616 ();
 sg13g2_fill_2 FILLER_37_632 ();
 sg13g2_fill_2 FILLER_37_642 ();
 sg13g2_fill_1 FILLER_37_644 ();
 sg13g2_fill_2 FILLER_37_670 ();
 sg13g2_fill_1 FILLER_37_691 ();
 sg13g2_fill_2 FILLER_37_709 ();
 sg13g2_fill_2 FILLER_37_721 ();
 sg13g2_fill_1 FILLER_37_723 ();
 sg13g2_decap_8 FILLER_37_748 ();
 sg13g2_fill_2 FILLER_37_755 ();
 sg13g2_fill_2 FILLER_37_772 ();
 sg13g2_fill_1 FILLER_37_774 ();
 sg13g2_decap_4 FILLER_37_789 ();
 sg13g2_fill_2 FILLER_37_800 ();
 sg13g2_decap_8 FILLER_37_806 ();
 sg13g2_decap_4 FILLER_37_813 ();
 sg13g2_fill_1 FILLER_37_817 ();
 sg13g2_fill_2 FILLER_37_835 ();
 sg13g2_fill_1 FILLER_37_848 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_fill_2 FILLER_37_919 ();
 sg13g2_decap_8 FILLER_37_928 ();
 sg13g2_fill_2 FILLER_37_935 ();
 sg13g2_decap_8 FILLER_37_944 ();
 sg13g2_fill_1 FILLER_37_951 ();
 sg13g2_decap_8 FILLER_37_968 ();
 sg13g2_fill_2 FILLER_37_975 ();
 sg13g2_decap_8 FILLER_37_1059 ();
 sg13g2_decap_8 FILLER_37_1066 ();
 sg13g2_decap_8 FILLER_37_1073 ();
 sg13g2_decap_8 FILLER_37_1080 ();
 sg13g2_decap_8 FILLER_37_1087 ();
 sg13g2_decap_8 FILLER_37_1094 ();
 sg13g2_decap_8 FILLER_37_1101 ();
 sg13g2_decap_8 FILLER_37_1108 ();
 sg13g2_decap_8 FILLER_37_1115 ();
 sg13g2_decap_8 FILLER_37_1122 ();
 sg13g2_decap_8 FILLER_37_1129 ();
 sg13g2_decap_8 FILLER_37_1136 ();
 sg13g2_decap_8 FILLER_37_1143 ();
 sg13g2_decap_8 FILLER_37_1150 ();
 sg13g2_decap_8 FILLER_37_1157 ();
 sg13g2_decap_8 FILLER_37_1164 ();
 sg13g2_decap_8 FILLER_37_1171 ();
 sg13g2_decap_8 FILLER_37_1178 ();
 sg13g2_decap_8 FILLER_37_1185 ();
 sg13g2_decap_8 FILLER_37_1192 ();
 sg13g2_decap_8 FILLER_37_1199 ();
 sg13g2_decap_8 FILLER_37_1206 ();
 sg13g2_decap_8 FILLER_37_1213 ();
 sg13g2_decap_8 FILLER_37_1220 ();
 sg13g2_decap_8 FILLER_37_1227 ();
 sg13g2_decap_8 FILLER_37_1234 ();
 sg13g2_decap_8 FILLER_37_1241 ();
 sg13g2_decap_8 FILLER_37_1248 ();
 sg13g2_decap_8 FILLER_37_1255 ();
 sg13g2_decap_8 FILLER_37_1262 ();
 sg13g2_decap_8 FILLER_37_1269 ();
 sg13g2_decap_8 FILLER_37_1276 ();
 sg13g2_decap_8 FILLER_37_1283 ();
 sg13g2_decap_8 FILLER_37_1290 ();
 sg13g2_decap_8 FILLER_37_1297 ();
 sg13g2_decap_8 FILLER_37_1304 ();
 sg13g2_decap_4 FILLER_37_1311 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_91 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_2 FILLER_38_145 ();
 sg13g2_fill_2 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_235 ();
 sg13g2_fill_1 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_decap_4 FILLER_38_337 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_2 FILLER_38_347 ();
 sg13g2_fill_1 FILLER_38_349 ();
 sg13g2_decap_4 FILLER_38_355 ();
 sg13g2_fill_2 FILLER_38_393 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_fill_1 FILLER_38_410 ();
 sg13g2_fill_2 FILLER_38_415 ();
 sg13g2_fill_1 FILLER_38_417 ();
 sg13g2_fill_2 FILLER_38_458 ();
 sg13g2_fill_2 FILLER_38_481 ();
 sg13g2_fill_1 FILLER_38_492 ();
 sg13g2_decap_4 FILLER_38_497 ();
 sg13g2_fill_2 FILLER_38_511 ();
 sg13g2_fill_2 FILLER_38_529 ();
 sg13g2_decap_8 FILLER_38_563 ();
 sg13g2_decap_8 FILLER_38_570 ();
 sg13g2_fill_1 FILLER_38_577 ();
 sg13g2_decap_4 FILLER_38_594 ();
 sg13g2_fill_2 FILLER_38_598 ();
 sg13g2_fill_1 FILLER_38_610 ();
 sg13g2_fill_2 FILLER_38_618 ();
 sg13g2_decap_8 FILLER_38_651 ();
 sg13g2_fill_2 FILLER_38_658 ();
 sg13g2_fill_1 FILLER_38_660 ();
 sg13g2_decap_8 FILLER_38_668 ();
 sg13g2_decap_8 FILLER_38_675 ();
 sg13g2_decap_8 FILLER_38_682 ();
 sg13g2_fill_2 FILLER_38_702 ();
 sg13g2_fill_1 FILLER_38_708 ();
 sg13g2_decap_4 FILLER_38_713 ();
 sg13g2_fill_2 FILLER_38_717 ();
 sg13g2_fill_1 FILLER_38_729 ();
 sg13g2_fill_1 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_fill_2 FILLER_38_756 ();
 sg13g2_fill_1 FILLER_38_758 ();
 sg13g2_fill_1 FILLER_38_768 ();
 sg13g2_fill_1 FILLER_38_777 ();
 sg13g2_fill_2 FILLER_38_815 ();
 sg13g2_fill_1 FILLER_38_835 ();
 sg13g2_decap_4 FILLER_38_850 ();
 sg13g2_fill_2 FILLER_38_854 ();
 sg13g2_fill_2 FILLER_38_886 ();
 sg13g2_fill_1 FILLER_38_888 ();
 sg13g2_fill_2 FILLER_38_910 ();
 sg13g2_fill_1 FILLER_38_912 ();
 sg13g2_fill_1 FILLER_38_918 ();
 sg13g2_fill_2 FILLER_38_936 ();
 sg13g2_decap_4 FILLER_38_973 ();
 sg13g2_fill_1 FILLER_38_981 ();
 sg13g2_fill_2 FILLER_38_1012 ();
 sg13g2_decap_8 FILLER_38_1066 ();
 sg13g2_decap_8 FILLER_38_1073 ();
 sg13g2_decap_8 FILLER_38_1080 ();
 sg13g2_decap_8 FILLER_38_1087 ();
 sg13g2_decap_8 FILLER_38_1094 ();
 sg13g2_decap_8 FILLER_38_1101 ();
 sg13g2_decap_8 FILLER_38_1108 ();
 sg13g2_decap_8 FILLER_38_1115 ();
 sg13g2_decap_8 FILLER_38_1122 ();
 sg13g2_decap_8 FILLER_38_1129 ();
 sg13g2_decap_8 FILLER_38_1136 ();
 sg13g2_decap_8 FILLER_38_1143 ();
 sg13g2_decap_8 FILLER_38_1150 ();
 sg13g2_decap_8 FILLER_38_1157 ();
 sg13g2_decap_8 FILLER_38_1164 ();
 sg13g2_decap_8 FILLER_38_1171 ();
 sg13g2_decap_8 FILLER_38_1178 ();
 sg13g2_decap_8 FILLER_38_1185 ();
 sg13g2_decap_8 FILLER_38_1192 ();
 sg13g2_decap_8 FILLER_38_1199 ();
 sg13g2_decap_8 FILLER_38_1206 ();
 sg13g2_decap_8 FILLER_38_1213 ();
 sg13g2_decap_8 FILLER_38_1220 ();
 sg13g2_decap_8 FILLER_38_1227 ();
 sg13g2_decap_8 FILLER_38_1234 ();
 sg13g2_decap_8 FILLER_38_1241 ();
 sg13g2_decap_8 FILLER_38_1248 ();
 sg13g2_decap_8 FILLER_38_1255 ();
 sg13g2_decap_8 FILLER_38_1262 ();
 sg13g2_decap_8 FILLER_38_1269 ();
 sg13g2_decap_8 FILLER_38_1276 ();
 sg13g2_decap_8 FILLER_38_1283 ();
 sg13g2_decap_8 FILLER_38_1290 ();
 sg13g2_decap_8 FILLER_38_1297 ();
 sg13g2_decap_8 FILLER_38_1304 ();
 sg13g2_decap_4 FILLER_38_1311 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_fill_2 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_183 ();
 sg13g2_fill_2 FILLER_39_206 ();
 sg13g2_fill_1 FILLER_39_208 ();
 sg13g2_fill_2 FILLER_39_235 ();
 sg13g2_fill_1 FILLER_39_237 ();
 sg13g2_decap_4 FILLER_39_243 ();
 sg13g2_fill_1 FILLER_39_247 ();
 sg13g2_decap_8 FILLER_39_305 ();
 sg13g2_fill_2 FILLER_39_325 ();
 sg13g2_fill_2 FILLER_39_360 ();
 sg13g2_fill_1 FILLER_39_362 ();
 sg13g2_decap_4 FILLER_39_368 ();
 sg13g2_fill_2 FILLER_39_372 ();
 sg13g2_decap_4 FILLER_39_378 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_decap_8 FILLER_39_391 ();
 sg13g2_fill_2 FILLER_39_398 ();
 sg13g2_decap_8 FILLER_39_407 ();
 sg13g2_fill_1 FILLER_39_422 ();
 sg13g2_decap_8 FILLER_39_466 ();
 sg13g2_fill_2 FILLER_39_473 ();
 sg13g2_fill_1 FILLER_39_475 ();
 sg13g2_fill_1 FILLER_39_515 ();
 sg13g2_fill_2 FILLER_39_522 ();
 sg13g2_fill_2 FILLER_39_552 ();
 sg13g2_fill_1 FILLER_39_599 ();
 sg13g2_decap_8 FILLER_39_605 ();
 sg13g2_fill_2 FILLER_39_617 ();
 sg13g2_fill_2 FILLER_39_644 ();
 sg13g2_fill_2 FILLER_39_650 ();
 sg13g2_fill_2 FILLER_39_710 ();
 sg13g2_fill_1 FILLER_39_728 ();
 sg13g2_decap_4 FILLER_39_733 ();
 sg13g2_fill_1 FILLER_39_737 ();
 sg13g2_decap_4 FILLER_39_753 ();
 sg13g2_fill_2 FILLER_39_757 ();
 sg13g2_decap_4 FILLER_39_769 ();
 sg13g2_fill_1 FILLER_39_773 ();
 sg13g2_decap_4 FILLER_39_778 ();
 sg13g2_fill_1 FILLER_39_782 ();
 sg13g2_decap_4 FILLER_39_798 ();
 sg13g2_fill_2 FILLER_39_802 ();
 sg13g2_fill_2 FILLER_39_808 ();
 sg13g2_fill_1 FILLER_39_810 ();
 sg13g2_fill_2 FILLER_39_821 ();
 sg13g2_fill_1 FILLER_39_823 ();
 sg13g2_decap_8 FILLER_39_829 ();
 sg13g2_fill_2 FILLER_39_836 ();
 sg13g2_decap_8 FILLER_39_872 ();
 sg13g2_decap_4 FILLER_39_879 ();
 sg13g2_fill_1 FILLER_39_883 ();
 sg13g2_decap_8 FILLER_39_892 ();
 sg13g2_decap_4 FILLER_39_899 ();
 sg13g2_fill_1 FILLER_39_903 ();
 sg13g2_fill_2 FILLER_39_926 ();
 sg13g2_fill_1 FILLER_39_928 ();
 sg13g2_fill_2 FILLER_39_963 ();
 sg13g2_fill_1 FILLER_39_965 ();
 sg13g2_fill_2 FILLER_39_1023 ();
 sg13g2_decap_8 FILLER_39_1051 ();
 sg13g2_decap_8 FILLER_39_1058 ();
 sg13g2_decap_8 FILLER_39_1065 ();
 sg13g2_decap_8 FILLER_39_1072 ();
 sg13g2_decap_8 FILLER_39_1079 ();
 sg13g2_decap_8 FILLER_39_1086 ();
 sg13g2_decap_8 FILLER_39_1093 ();
 sg13g2_decap_8 FILLER_39_1100 ();
 sg13g2_decap_8 FILLER_39_1107 ();
 sg13g2_decap_8 FILLER_39_1114 ();
 sg13g2_decap_8 FILLER_39_1121 ();
 sg13g2_decap_8 FILLER_39_1128 ();
 sg13g2_decap_8 FILLER_39_1135 ();
 sg13g2_decap_8 FILLER_39_1142 ();
 sg13g2_decap_8 FILLER_39_1149 ();
 sg13g2_decap_8 FILLER_39_1156 ();
 sg13g2_decap_8 FILLER_39_1163 ();
 sg13g2_decap_8 FILLER_39_1170 ();
 sg13g2_decap_8 FILLER_39_1177 ();
 sg13g2_decap_8 FILLER_39_1184 ();
 sg13g2_decap_8 FILLER_39_1191 ();
 sg13g2_decap_8 FILLER_39_1198 ();
 sg13g2_decap_8 FILLER_39_1205 ();
 sg13g2_decap_8 FILLER_39_1212 ();
 sg13g2_decap_8 FILLER_39_1219 ();
 sg13g2_decap_8 FILLER_39_1226 ();
 sg13g2_decap_8 FILLER_39_1233 ();
 sg13g2_decap_8 FILLER_39_1240 ();
 sg13g2_decap_8 FILLER_39_1247 ();
 sg13g2_decap_8 FILLER_39_1254 ();
 sg13g2_decap_8 FILLER_39_1261 ();
 sg13g2_decap_8 FILLER_39_1268 ();
 sg13g2_decap_8 FILLER_39_1275 ();
 sg13g2_decap_8 FILLER_39_1282 ();
 sg13g2_decap_8 FILLER_39_1289 ();
 sg13g2_decap_8 FILLER_39_1296 ();
 sg13g2_decap_8 FILLER_39_1303 ();
 sg13g2_decap_4 FILLER_39_1310 ();
 sg13g2_fill_1 FILLER_39_1314 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_fill_1 FILLER_40_126 ();
 sg13g2_decap_4 FILLER_40_145 ();
 sg13g2_fill_2 FILLER_40_149 ();
 sg13g2_decap_4 FILLER_40_155 ();
 sg13g2_decap_8 FILLER_40_163 ();
 sg13g2_fill_2 FILLER_40_170 ();
 sg13g2_fill_1 FILLER_40_212 ();
 sg13g2_fill_2 FILLER_40_226 ();
 sg13g2_fill_1 FILLER_40_228 ();
 sg13g2_decap_8 FILLER_40_264 ();
 sg13g2_fill_2 FILLER_40_271 ();
 sg13g2_decap_8 FILLER_40_330 ();
 sg13g2_decap_8 FILLER_40_341 ();
 sg13g2_decap_8 FILLER_40_348 ();
 sg13g2_fill_2 FILLER_40_355 ();
 sg13g2_fill_1 FILLER_40_362 ();
 sg13g2_fill_2 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_fill_2 FILLER_40_385 ();
 sg13g2_fill_1 FILLER_40_387 ();
 sg13g2_decap_4 FILLER_40_414 ();
 sg13g2_fill_2 FILLER_40_418 ();
 sg13g2_decap_4 FILLER_40_446 ();
 sg13g2_fill_1 FILLER_40_450 ();
 sg13g2_decap_4 FILLER_40_455 ();
 sg13g2_fill_2 FILLER_40_459 ();
 sg13g2_fill_1 FILLER_40_491 ();
 sg13g2_decap_8 FILLER_40_499 ();
 sg13g2_fill_2 FILLER_40_506 ();
 sg13g2_fill_1 FILLER_40_508 ();
 sg13g2_fill_1 FILLER_40_531 ();
 sg13g2_decap_8 FILLER_40_558 ();
 sg13g2_fill_2 FILLER_40_569 ();
 sg13g2_fill_1 FILLER_40_571 ();
 sg13g2_decap_8 FILLER_40_576 ();
 sg13g2_decap_4 FILLER_40_583 ();
 sg13g2_fill_1 FILLER_40_587 ();
 sg13g2_fill_1 FILLER_40_614 ();
 sg13g2_decap_4 FILLER_40_620 ();
 sg13g2_fill_2 FILLER_40_629 ();
 sg13g2_decap_8 FILLER_40_663 ();
 sg13g2_decap_8 FILLER_40_670 ();
 sg13g2_fill_2 FILLER_40_677 ();
 sg13g2_decap_4 FILLER_40_691 ();
 sg13g2_fill_2 FILLER_40_695 ();
 sg13g2_decap_4 FILLER_40_718 ();
 sg13g2_fill_1 FILLER_40_722 ();
 sg13g2_decap_4 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_745 ();
 sg13g2_fill_2 FILLER_40_767 ();
 sg13g2_fill_1 FILLER_40_769 ();
 sg13g2_decap_8 FILLER_40_853 ();
 sg13g2_decap_4 FILLER_40_909 ();
 sg13g2_fill_1 FILLER_40_913 ();
 sg13g2_fill_2 FILLER_40_919 ();
 sg13g2_fill_2 FILLER_40_930 ();
 sg13g2_fill_1 FILLER_40_932 ();
 sg13g2_decap_8 FILLER_40_941 ();
 sg13g2_fill_1 FILLER_40_948 ();
 sg13g2_decap_4 FILLER_40_957 ();
 sg13g2_fill_1 FILLER_40_987 ();
 sg13g2_fill_1 FILLER_40_1010 ();
 sg13g2_fill_1 FILLER_40_1031 ();
 sg13g2_decap_8 FILLER_40_1063 ();
 sg13g2_decap_8 FILLER_40_1070 ();
 sg13g2_decap_8 FILLER_40_1077 ();
 sg13g2_decap_8 FILLER_40_1084 ();
 sg13g2_decap_8 FILLER_40_1091 ();
 sg13g2_decap_8 FILLER_40_1098 ();
 sg13g2_decap_8 FILLER_40_1105 ();
 sg13g2_decap_8 FILLER_40_1112 ();
 sg13g2_decap_8 FILLER_40_1119 ();
 sg13g2_decap_8 FILLER_40_1126 ();
 sg13g2_decap_8 FILLER_40_1133 ();
 sg13g2_decap_8 FILLER_40_1140 ();
 sg13g2_decap_8 FILLER_40_1147 ();
 sg13g2_decap_8 FILLER_40_1154 ();
 sg13g2_decap_8 FILLER_40_1161 ();
 sg13g2_decap_8 FILLER_40_1168 ();
 sg13g2_decap_8 FILLER_40_1175 ();
 sg13g2_decap_8 FILLER_40_1182 ();
 sg13g2_decap_8 FILLER_40_1189 ();
 sg13g2_decap_8 FILLER_40_1196 ();
 sg13g2_decap_8 FILLER_40_1203 ();
 sg13g2_decap_8 FILLER_40_1210 ();
 sg13g2_decap_8 FILLER_40_1217 ();
 sg13g2_decap_8 FILLER_40_1224 ();
 sg13g2_decap_8 FILLER_40_1231 ();
 sg13g2_decap_8 FILLER_40_1238 ();
 sg13g2_decap_8 FILLER_40_1245 ();
 sg13g2_decap_8 FILLER_40_1252 ();
 sg13g2_decap_8 FILLER_40_1259 ();
 sg13g2_decap_8 FILLER_40_1266 ();
 sg13g2_decap_8 FILLER_40_1273 ();
 sg13g2_decap_8 FILLER_40_1280 ();
 sg13g2_decap_8 FILLER_40_1287 ();
 sg13g2_decap_8 FILLER_40_1294 ();
 sg13g2_decap_8 FILLER_40_1301 ();
 sg13g2_decap_8 FILLER_40_1308 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_fill_1 FILLER_41_133 ();
 sg13g2_fill_1 FILLER_41_199 ();
 sg13g2_fill_1 FILLER_41_205 ();
 sg13g2_fill_2 FILLER_41_241 ();
 sg13g2_fill_1 FILLER_41_256 ();
 sg13g2_fill_2 FILLER_41_270 ();
 sg13g2_fill_1 FILLER_41_272 ();
 sg13g2_decap_4 FILLER_41_292 ();
 sg13g2_fill_1 FILLER_41_296 ();
 sg13g2_fill_2 FILLER_41_313 ();
 sg13g2_fill_2 FILLER_41_319 ();
 sg13g2_fill_1 FILLER_41_321 ();
 sg13g2_fill_1 FILLER_41_379 ();
 sg13g2_decap_8 FILLER_41_388 ();
 sg13g2_decap_8 FILLER_41_403 ();
 sg13g2_decap_8 FILLER_41_410 ();
 sg13g2_fill_1 FILLER_41_417 ();
 sg13g2_fill_1 FILLER_41_430 ();
 sg13g2_fill_1 FILLER_41_435 ();
 sg13g2_fill_2 FILLER_41_479 ();
 sg13g2_fill_1 FILLER_41_481 ();
 sg13g2_fill_2 FILLER_41_489 ();
 sg13g2_decap_8 FILLER_41_495 ();
 sg13g2_fill_1 FILLER_41_502 ();
 sg13g2_decap_4 FILLER_41_506 ();
 sg13g2_fill_2 FILLER_41_510 ();
 sg13g2_fill_2 FILLER_41_523 ();
 sg13g2_fill_1 FILLER_41_525 ();
 sg13g2_decap_8 FILLER_41_530 ();
 sg13g2_fill_2 FILLER_41_537 ();
 sg13g2_decap_8 FILLER_41_547 ();
 sg13g2_fill_2 FILLER_41_554 ();
 sg13g2_fill_1 FILLER_41_556 ();
 sg13g2_decap_4 FILLER_41_583 ();
 sg13g2_fill_2 FILLER_41_587 ();
 sg13g2_fill_2 FILLER_41_597 ();
 sg13g2_decap_8 FILLER_41_603 ();
 sg13g2_decap_4 FILLER_41_610 ();
 sg13g2_decap_8 FILLER_41_634 ();
 sg13g2_decap_8 FILLER_41_649 ();
 sg13g2_fill_2 FILLER_41_669 ();
 sg13g2_fill_2 FILLER_41_679 ();
 sg13g2_fill_1 FILLER_41_696 ();
 sg13g2_fill_2 FILLER_41_702 ();
 sg13g2_fill_1 FILLER_41_704 ();
 sg13g2_fill_2 FILLER_41_712 ();
 sg13g2_fill_2 FILLER_41_727 ();
 sg13g2_fill_1 FILLER_41_729 ();
 sg13g2_fill_2 FILLER_41_755 ();
 sg13g2_fill_1 FILLER_41_757 ();
 sg13g2_fill_2 FILLER_41_777 ();
 sg13g2_fill_2 FILLER_41_783 ();
 sg13g2_fill_1 FILLER_41_785 ();
 sg13g2_decap_8 FILLER_41_810 ();
 sg13g2_fill_2 FILLER_41_817 ();
 sg13g2_fill_2 FILLER_41_823 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_fill_2 FILLER_41_836 ();
 sg13g2_decap_4 FILLER_41_843 ();
 sg13g2_fill_2 FILLER_41_847 ();
 sg13g2_decap_4 FILLER_41_870 ();
 sg13g2_fill_2 FILLER_41_874 ();
 sg13g2_fill_1 FILLER_41_880 ();
 sg13g2_decap_4 FILLER_41_891 ();
 sg13g2_fill_2 FILLER_41_903 ();
 sg13g2_fill_1 FILLER_41_905 ();
 sg13g2_fill_1 FILLER_41_929 ();
 sg13g2_fill_1 FILLER_41_987 ();
 sg13g2_decap_8 FILLER_41_1053 ();
 sg13g2_decap_8 FILLER_41_1060 ();
 sg13g2_decap_8 FILLER_41_1067 ();
 sg13g2_decap_8 FILLER_41_1074 ();
 sg13g2_decap_8 FILLER_41_1081 ();
 sg13g2_decap_8 FILLER_41_1088 ();
 sg13g2_decap_8 FILLER_41_1095 ();
 sg13g2_decap_8 FILLER_41_1102 ();
 sg13g2_decap_8 FILLER_41_1109 ();
 sg13g2_decap_8 FILLER_41_1116 ();
 sg13g2_decap_8 FILLER_41_1123 ();
 sg13g2_decap_8 FILLER_41_1130 ();
 sg13g2_decap_8 FILLER_41_1137 ();
 sg13g2_decap_8 FILLER_41_1144 ();
 sg13g2_decap_8 FILLER_41_1151 ();
 sg13g2_decap_8 FILLER_41_1158 ();
 sg13g2_decap_8 FILLER_41_1165 ();
 sg13g2_decap_8 FILLER_41_1172 ();
 sg13g2_decap_8 FILLER_41_1179 ();
 sg13g2_decap_8 FILLER_41_1186 ();
 sg13g2_decap_8 FILLER_41_1193 ();
 sg13g2_decap_8 FILLER_41_1200 ();
 sg13g2_decap_8 FILLER_41_1207 ();
 sg13g2_decap_8 FILLER_41_1214 ();
 sg13g2_decap_8 FILLER_41_1221 ();
 sg13g2_decap_8 FILLER_41_1228 ();
 sg13g2_decap_8 FILLER_41_1235 ();
 sg13g2_decap_8 FILLER_41_1242 ();
 sg13g2_decap_8 FILLER_41_1249 ();
 sg13g2_decap_8 FILLER_41_1256 ();
 sg13g2_decap_8 FILLER_41_1263 ();
 sg13g2_decap_8 FILLER_41_1270 ();
 sg13g2_decap_8 FILLER_41_1277 ();
 sg13g2_decap_8 FILLER_41_1284 ();
 sg13g2_decap_8 FILLER_41_1291 ();
 sg13g2_decap_8 FILLER_41_1298 ();
 sg13g2_decap_8 FILLER_41_1305 ();
 sg13g2_fill_2 FILLER_41_1312 ();
 sg13g2_fill_1 FILLER_41_1314 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_fill_1 FILLER_42_149 ();
 sg13g2_fill_1 FILLER_42_159 ();
 sg13g2_fill_2 FILLER_42_174 ();
 sg13g2_fill_1 FILLER_42_176 ();
 sg13g2_fill_1 FILLER_42_199 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_fill_1 FILLER_42_224 ();
 sg13g2_decap_4 FILLER_42_251 ();
 sg13g2_fill_2 FILLER_42_281 ();
 sg13g2_decap_8 FILLER_42_309 ();
 sg13g2_fill_2 FILLER_42_316 ();
 sg13g2_fill_1 FILLER_42_318 ();
 sg13g2_fill_2 FILLER_42_349 ();
 sg13g2_fill_1 FILLER_42_351 ();
 sg13g2_decap_8 FILLER_42_356 ();
 sg13g2_fill_1 FILLER_42_363 ();
 sg13g2_decap_8 FILLER_42_368 ();
 sg13g2_fill_2 FILLER_42_444 ();
 sg13g2_fill_1 FILLER_42_446 ();
 sg13g2_fill_2 FILLER_42_451 ();
 sg13g2_fill_1 FILLER_42_453 ();
 sg13g2_fill_2 FILLER_42_526 ();
 sg13g2_decap_8 FILLER_42_558 ();
 sg13g2_fill_2 FILLER_42_565 ();
 sg13g2_fill_1 FILLER_42_567 ();
 sg13g2_fill_2 FILLER_42_572 ();
 sg13g2_fill_1 FILLER_42_574 ();
 sg13g2_fill_2 FILLER_42_583 ();
 sg13g2_fill_1 FILLER_42_606 ();
 sg13g2_fill_2 FILLER_42_635 ();
 sg13g2_fill_1 FILLER_42_637 ();
 sg13g2_decap_4 FILLER_42_675 ();
 sg13g2_fill_2 FILLER_42_688 ();
 sg13g2_fill_1 FILLER_42_695 ();
 sg13g2_fill_1 FILLER_42_723 ();
 sg13g2_fill_2 FILLER_42_729 ();
 sg13g2_fill_2 FILLER_42_784 ();
 sg13g2_decap_4 FILLER_42_809 ();
 sg13g2_fill_2 FILLER_42_813 ();
 sg13g2_decap_8 FILLER_42_841 ();
 sg13g2_decap_4 FILLER_42_848 ();
 sg13g2_fill_1 FILLER_42_852 ();
 sg13g2_decap_8 FILLER_42_861 ();
 sg13g2_fill_2 FILLER_42_868 ();
 sg13g2_decap_8 FILLER_42_885 ();
 sg13g2_fill_2 FILLER_42_892 ();
 sg13g2_decap_4 FILLER_42_908 ();
 sg13g2_fill_2 FILLER_42_912 ();
 sg13g2_decap_4 FILLER_42_924 ();
 sg13g2_fill_2 FILLER_42_928 ();
 sg13g2_fill_2 FILLER_42_939 ();
 sg13g2_fill_1 FILLER_42_941 ();
 sg13g2_decap_4 FILLER_42_967 ();
 sg13g2_fill_1 FILLER_42_988 ();
 sg13g2_fill_1 FILLER_42_1003 ();
 sg13g2_fill_2 FILLER_42_1030 ();
 sg13g2_fill_1 FILLER_42_1032 ();
 sg13g2_decap_8 FILLER_42_1059 ();
 sg13g2_decap_8 FILLER_42_1066 ();
 sg13g2_decap_8 FILLER_42_1073 ();
 sg13g2_decap_8 FILLER_42_1080 ();
 sg13g2_decap_8 FILLER_42_1087 ();
 sg13g2_decap_8 FILLER_42_1094 ();
 sg13g2_decap_8 FILLER_42_1101 ();
 sg13g2_decap_8 FILLER_42_1108 ();
 sg13g2_decap_8 FILLER_42_1115 ();
 sg13g2_decap_8 FILLER_42_1122 ();
 sg13g2_decap_8 FILLER_42_1129 ();
 sg13g2_decap_8 FILLER_42_1136 ();
 sg13g2_decap_8 FILLER_42_1143 ();
 sg13g2_decap_8 FILLER_42_1150 ();
 sg13g2_decap_8 FILLER_42_1157 ();
 sg13g2_decap_8 FILLER_42_1164 ();
 sg13g2_decap_8 FILLER_42_1171 ();
 sg13g2_decap_8 FILLER_42_1178 ();
 sg13g2_decap_8 FILLER_42_1185 ();
 sg13g2_decap_8 FILLER_42_1192 ();
 sg13g2_decap_8 FILLER_42_1199 ();
 sg13g2_decap_8 FILLER_42_1206 ();
 sg13g2_decap_8 FILLER_42_1213 ();
 sg13g2_decap_8 FILLER_42_1220 ();
 sg13g2_decap_8 FILLER_42_1227 ();
 sg13g2_decap_8 FILLER_42_1234 ();
 sg13g2_decap_8 FILLER_42_1241 ();
 sg13g2_decap_8 FILLER_42_1248 ();
 sg13g2_decap_8 FILLER_42_1255 ();
 sg13g2_decap_8 FILLER_42_1262 ();
 sg13g2_decap_8 FILLER_42_1269 ();
 sg13g2_decap_8 FILLER_42_1276 ();
 sg13g2_decap_8 FILLER_42_1283 ();
 sg13g2_decap_8 FILLER_42_1290 ();
 sg13g2_decap_8 FILLER_42_1297 ();
 sg13g2_decap_8 FILLER_42_1304 ();
 sg13g2_decap_4 FILLER_42_1311 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_4 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_121 ();
 sg13g2_fill_2 FILLER_43_127 ();
 sg13g2_fill_1 FILLER_43_129 ();
 sg13g2_fill_2 FILLER_43_148 ();
 sg13g2_fill_1 FILLER_43_150 ();
 sg13g2_fill_1 FILLER_43_187 ();
 sg13g2_decap_4 FILLER_43_224 ();
 sg13g2_fill_1 FILLER_43_228 ();
 sg13g2_fill_2 FILLER_43_234 ();
 sg13g2_fill_1 FILLER_43_244 ();
 sg13g2_fill_1 FILLER_43_271 ();
 sg13g2_fill_2 FILLER_43_289 ();
 sg13g2_fill_1 FILLER_43_321 ();
 sg13g2_fill_2 FILLER_43_327 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_fill_2 FILLER_43_334 ();
 sg13g2_fill_1 FILLER_43_388 ();
 sg13g2_fill_1 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_422 ();
 sg13g2_fill_2 FILLER_43_445 ();
 sg13g2_fill_1 FILLER_43_447 ();
 sg13g2_decap_4 FILLER_43_461 ();
 sg13g2_fill_1 FILLER_43_465 ();
 sg13g2_decap_4 FILLER_43_473 ();
 sg13g2_fill_2 FILLER_43_477 ();
 sg13g2_fill_2 FILLER_43_484 ();
 sg13g2_decap_4 FILLER_43_493 ();
 sg13g2_fill_1 FILLER_43_497 ();
 sg13g2_decap_4 FILLER_43_506 ();
 sg13g2_fill_2 FILLER_43_528 ();
 sg13g2_fill_1 FILLER_43_530 ();
 sg13g2_fill_1 FILLER_43_536 ();
 sg13g2_fill_1 FILLER_43_541 ();
 sg13g2_fill_2 FILLER_43_598 ();
 sg13g2_fill_1 FILLER_43_600 ();
 sg13g2_decap_4 FILLER_43_609 ();
 sg13g2_fill_2 FILLER_43_618 ();
 sg13g2_fill_1 FILLER_43_620 ();
 sg13g2_decap_8 FILLER_43_647 ();
 sg13g2_decap_8 FILLER_43_654 ();
 sg13g2_fill_2 FILLER_43_661 ();
 sg13g2_fill_1 FILLER_43_663 ();
 sg13g2_decap_8 FILLER_43_668 ();
 sg13g2_fill_1 FILLER_43_680 ();
 sg13g2_decap_8 FILLER_43_685 ();
 sg13g2_decap_8 FILLER_43_692 ();
 sg13g2_fill_2 FILLER_43_699 ();
 sg13g2_fill_1 FILLER_43_705 ();
 sg13g2_decap_8 FILLER_43_710 ();
 sg13g2_decap_4 FILLER_43_717 ();
 sg13g2_fill_2 FILLER_43_721 ();
 sg13g2_decap_4 FILLER_43_727 ();
 sg13g2_fill_2 FILLER_43_740 ();
 sg13g2_fill_1 FILLER_43_747 ();
 sg13g2_decap_8 FILLER_43_762 ();
 sg13g2_decap_8 FILLER_43_779 ();
 sg13g2_fill_2 FILLER_43_791 ();
 sg13g2_decap_4 FILLER_43_803 ();
 sg13g2_fill_1 FILLER_43_822 ();
 sg13g2_decap_4 FILLER_43_840 ();
 sg13g2_fill_2 FILLER_43_865 ();
 sg13g2_fill_1 FILLER_43_867 ();
 sg13g2_fill_1 FILLER_43_908 ();
 sg13g2_decap_4 FILLER_43_972 ();
 sg13g2_fill_1 FILLER_43_976 ();
 sg13g2_fill_2 FILLER_43_1011 ();
 sg13g2_fill_1 FILLER_43_1013 ();
 sg13g2_fill_2 FILLER_43_1023 ();
 sg13g2_decap_8 FILLER_43_1066 ();
 sg13g2_decap_8 FILLER_43_1073 ();
 sg13g2_decap_8 FILLER_43_1080 ();
 sg13g2_decap_8 FILLER_43_1087 ();
 sg13g2_decap_8 FILLER_43_1094 ();
 sg13g2_decap_8 FILLER_43_1101 ();
 sg13g2_decap_8 FILLER_43_1108 ();
 sg13g2_decap_8 FILLER_43_1115 ();
 sg13g2_decap_8 FILLER_43_1122 ();
 sg13g2_decap_8 FILLER_43_1129 ();
 sg13g2_decap_8 FILLER_43_1136 ();
 sg13g2_decap_8 FILLER_43_1143 ();
 sg13g2_decap_8 FILLER_43_1150 ();
 sg13g2_decap_8 FILLER_43_1157 ();
 sg13g2_decap_8 FILLER_43_1164 ();
 sg13g2_decap_8 FILLER_43_1171 ();
 sg13g2_decap_8 FILLER_43_1178 ();
 sg13g2_decap_8 FILLER_43_1185 ();
 sg13g2_decap_8 FILLER_43_1192 ();
 sg13g2_decap_8 FILLER_43_1199 ();
 sg13g2_decap_8 FILLER_43_1206 ();
 sg13g2_decap_8 FILLER_43_1213 ();
 sg13g2_decap_8 FILLER_43_1220 ();
 sg13g2_decap_8 FILLER_43_1227 ();
 sg13g2_decap_8 FILLER_43_1234 ();
 sg13g2_decap_8 FILLER_43_1241 ();
 sg13g2_decap_8 FILLER_43_1248 ();
 sg13g2_decap_8 FILLER_43_1255 ();
 sg13g2_decap_8 FILLER_43_1262 ();
 sg13g2_decap_8 FILLER_43_1269 ();
 sg13g2_decap_8 FILLER_43_1276 ();
 sg13g2_decap_8 FILLER_43_1283 ();
 sg13g2_decap_8 FILLER_43_1290 ();
 sg13g2_decap_8 FILLER_43_1297 ();
 sg13g2_decap_8 FILLER_43_1304 ();
 sg13g2_decap_4 FILLER_43_1311 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_fill_2 FILLER_44_162 ();
 sg13g2_fill_1 FILLER_44_178 ();
 sg13g2_fill_2 FILLER_44_183 ();
 sg13g2_fill_1 FILLER_44_185 ();
 sg13g2_decap_4 FILLER_44_209 ();
 sg13g2_fill_2 FILLER_44_243 ();
 sg13g2_fill_1 FILLER_44_259 ();
 sg13g2_fill_2 FILLER_44_286 ();
 sg13g2_fill_2 FILLER_44_292 ();
 sg13g2_decap_4 FILLER_44_311 ();
 sg13g2_fill_2 FILLER_44_315 ();
 sg13g2_decap_4 FILLER_44_330 ();
 sg13g2_fill_2 FILLER_44_334 ();
 sg13g2_fill_2 FILLER_44_350 ();
 sg13g2_fill_1 FILLER_44_352 ();
 sg13g2_decap_8 FILLER_44_362 ();
 sg13g2_fill_2 FILLER_44_369 ();
 sg13g2_fill_1 FILLER_44_384 ();
 sg13g2_fill_2 FILLER_44_463 ();
 sg13g2_fill_1 FILLER_44_465 ();
 sg13g2_decap_8 FILLER_44_492 ();
 sg13g2_fill_1 FILLER_44_499 ();
 sg13g2_decap_4 FILLER_44_533 ();
 sg13g2_fill_1 FILLER_44_537 ();
 sg13g2_decap_8 FILLER_44_542 ();
 sg13g2_fill_1 FILLER_44_549 ();
 sg13g2_decap_8 FILLER_44_576 ();
 sg13g2_decap_4 FILLER_44_587 ();
 sg13g2_fill_2 FILLER_44_602 ();
 sg13g2_fill_1 FILLER_44_614 ();
 sg13g2_decap_4 FILLER_44_623 ();
 sg13g2_fill_1 FILLER_44_684 ();
 sg13g2_fill_1 FILLER_44_716 ();
 sg13g2_decap_8 FILLER_44_743 ();
 sg13g2_decap_4 FILLER_44_750 ();
 sg13g2_fill_1 FILLER_44_754 ();
 sg13g2_decap_8 FILLER_44_764 ();
 sg13g2_decap_4 FILLER_44_771 ();
 sg13g2_decap_8 FILLER_44_779 ();
 sg13g2_fill_2 FILLER_44_786 ();
 sg13g2_decap_8 FILLER_44_796 ();
 sg13g2_fill_1 FILLER_44_803 ();
 sg13g2_fill_2 FILLER_44_814 ();
 sg13g2_fill_1 FILLER_44_816 ();
 sg13g2_fill_1 FILLER_44_841 ();
 sg13g2_fill_2 FILLER_44_866 ();
 sg13g2_decap_8 FILLER_44_882 ();
 sg13g2_fill_2 FILLER_44_889 ();
 sg13g2_fill_1 FILLER_44_891 ();
 sg13g2_decap_8 FILLER_44_907 ();
 sg13g2_decap_4 FILLER_44_914 ();
 sg13g2_fill_1 FILLER_44_918 ();
 sg13g2_decap_4 FILLER_44_935 ();
 sg13g2_fill_2 FILLER_44_939 ();
 sg13g2_fill_2 FILLER_44_946 ();
 sg13g2_decap_4 FILLER_44_978 ();
 sg13g2_fill_2 FILLER_44_992 ();
 sg13g2_fill_1 FILLER_44_994 ();
 sg13g2_fill_2 FILLER_44_999 ();
 sg13g2_fill_1 FILLER_44_1001 ();
 sg13g2_fill_2 FILLER_44_1037 ();
 sg13g2_fill_1 FILLER_44_1039 ();
 sg13g2_decap_8 FILLER_44_1066 ();
 sg13g2_decap_8 FILLER_44_1073 ();
 sg13g2_decap_8 FILLER_44_1080 ();
 sg13g2_decap_8 FILLER_44_1087 ();
 sg13g2_decap_8 FILLER_44_1094 ();
 sg13g2_decap_8 FILLER_44_1101 ();
 sg13g2_decap_8 FILLER_44_1108 ();
 sg13g2_decap_8 FILLER_44_1115 ();
 sg13g2_decap_8 FILLER_44_1122 ();
 sg13g2_decap_8 FILLER_44_1129 ();
 sg13g2_decap_8 FILLER_44_1136 ();
 sg13g2_decap_8 FILLER_44_1143 ();
 sg13g2_decap_8 FILLER_44_1150 ();
 sg13g2_decap_8 FILLER_44_1157 ();
 sg13g2_decap_8 FILLER_44_1164 ();
 sg13g2_decap_8 FILLER_44_1171 ();
 sg13g2_decap_8 FILLER_44_1178 ();
 sg13g2_decap_8 FILLER_44_1185 ();
 sg13g2_decap_8 FILLER_44_1192 ();
 sg13g2_decap_8 FILLER_44_1199 ();
 sg13g2_decap_8 FILLER_44_1206 ();
 sg13g2_decap_8 FILLER_44_1213 ();
 sg13g2_decap_8 FILLER_44_1220 ();
 sg13g2_decap_8 FILLER_44_1227 ();
 sg13g2_decap_8 FILLER_44_1234 ();
 sg13g2_decap_8 FILLER_44_1241 ();
 sg13g2_decap_8 FILLER_44_1248 ();
 sg13g2_decap_8 FILLER_44_1255 ();
 sg13g2_decap_8 FILLER_44_1262 ();
 sg13g2_decap_8 FILLER_44_1269 ();
 sg13g2_decap_8 FILLER_44_1276 ();
 sg13g2_decap_8 FILLER_44_1283 ();
 sg13g2_decap_8 FILLER_44_1290 ();
 sg13g2_decap_8 FILLER_44_1297 ();
 sg13g2_decap_8 FILLER_44_1304 ();
 sg13g2_decap_4 FILLER_44_1311 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_fill_2 FILLER_45_110 ();
 sg13g2_fill_1 FILLER_45_112 ();
 sg13g2_decap_4 FILLER_45_127 ();
 sg13g2_fill_2 FILLER_45_135 ();
 sg13g2_fill_2 FILLER_45_142 ();
 sg13g2_fill_1 FILLER_45_144 ();
 sg13g2_fill_2 FILLER_45_205 ();
 sg13g2_fill_1 FILLER_45_218 ();
 sg13g2_fill_2 FILLER_45_228 ();
 sg13g2_fill_2 FILLER_45_235 ();
 sg13g2_fill_1 FILLER_45_237 ();
 sg13g2_fill_2 FILLER_45_264 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_fill_2 FILLER_45_318 ();
 sg13g2_fill_1 FILLER_45_351 ();
 sg13g2_fill_2 FILLER_45_383 ();
 sg13g2_decap_8 FILLER_45_390 ();
 sg13g2_fill_1 FILLER_45_397 ();
 sg13g2_fill_2 FILLER_45_402 ();
 sg13g2_fill_1 FILLER_45_404 ();
 sg13g2_decap_4 FILLER_45_414 ();
 sg13g2_fill_2 FILLER_45_418 ();
 sg13g2_decap_8 FILLER_45_433 ();
 sg13g2_fill_2 FILLER_45_461 ();
 sg13g2_fill_1 FILLER_45_463 ();
 sg13g2_decap_8 FILLER_45_485 ();
 sg13g2_fill_2 FILLER_45_492 ();
 sg13g2_decap_8 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_518 ();
 sg13g2_fill_2 FILLER_45_525 ();
 sg13g2_fill_1 FILLER_45_527 ();
 sg13g2_decap_4 FILLER_45_554 ();
 sg13g2_fill_2 FILLER_45_567 ();
 sg13g2_fill_1 FILLER_45_569 ();
 sg13g2_fill_2 FILLER_45_609 ();
 sg13g2_fill_1 FILLER_45_611 ();
 sg13g2_decap_8 FILLER_45_620 ();
 sg13g2_fill_1 FILLER_45_631 ();
 sg13g2_fill_2 FILLER_45_666 ();
 sg13g2_fill_1 FILLER_45_668 ();
 sg13g2_decap_8 FILLER_45_699 ();
 sg13g2_fill_1 FILLER_45_706 ();
 sg13g2_decap_8 FILLER_45_718 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_4 FILLER_45_732 ();
 sg13g2_fill_1 FILLER_45_736 ();
 sg13g2_fill_2 FILLER_45_756 ();
 sg13g2_fill_2 FILLER_45_762 ();
 sg13g2_fill_1 FILLER_45_764 ();
 sg13g2_fill_1 FILLER_45_796 ();
 sg13g2_decap_8 FILLER_45_817 ();
 sg13g2_fill_1 FILLER_45_824 ();
 sg13g2_decap_8 FILLER_45_830 ();
 sg13g2_fill_2 FILLER_45_837 ();
 sg13g2_fill_1 FILLER_45_839 ();
 sg13g2_decap_4 FILLER_45_860 ();
 sg13g2_fill_1 FILLER_45_864 ();
 sg13g2_fill_1 FILLER_45_884 ();
 sg13g2_decap_4 FILLER_45_890 ();
 sg13g2_decap_8 FILLER_45_908 ();
 sg13g2_decap_4 FILLER_45_915 ();
 sg13g2_fill_1 FILLER_45_923 ();
 sg13g2_fill_1 FILLER_45_934 ();
 sg13g2_fill_2 FILLER_45_943 ();
 sg13g2_fill_1 FILLER_45_945 ();
 sg13g2_fill_1 FILLER_45_954 ();
 sg13g2_fill_2 FILLER_45_973 ();
 sg13g2_fill_2 FILLER_45_980 ();
 sg13g2_decap_8 FILLER_45_1065 ();
 sg13g2_decap_8 FILLER_45_1072 ();
 sg13g2_decap_8 FILLER_45_1079 ();
 sg13g2_decap_8 FILLER_45_1086 ();
 sg13g2_decap_8 FILLER_45_1093 ();
 sg13g2_decap_8 FILLER_45_1100 ();
 sg13g2_decap_8 FILLER_45_1107 ();
 sg13g2_decap_8 FILLER_45_1114 ();
 sg13g2_decap_8 FILLER_45_1121 ();
 sg13g2_decap_8 FILLER_45_1128 ();
 sg13g2_decap_8 FILLER_45_1135 ();
 sg13g2_decap_8 FILLER_45_1142 ();
 sg13g2_decap_8 FILLER_45_1149 ();
 sg13g2_decap_8 FILLER_45_1156 ();
 sg13g2_decap_8 FILLER_45_1163 ();
 sg13g2_decap_8 FILLER_45_1170 ();
 sg13g2_decap_8 FILLER_45_1177 ();
 sg13g2_decap_8 FILLER_45_1184 ();
 sg13g2_decap_8 FILLER_45_1191 ();
 sg13g2_decap_8 FILLER_45_1198 ();
 sg13g2_decap_8 FILLER_45_1205 ();
 sg13g2_decap_8 FILLER_45_1212 ();
 sg13g2_decap_8 FILLER_45_1219 ();
 sg13g2_decap_8 FILLER_45_1226 ();
 sg13g2_decap_8 FILLER_45_1233 ();
 sg13g2_decap_8 FILLER_45_1240 ();
 sg13g2_decap_8 FILLER_45_1247 ();
 sg13g2_decap_8 FILLER_45_1254 ();
 sg13g2_decap_8 FILLER_45_1261 ();
 sg13g2_decap_8 FILLER_45_1268 ();
 sg13g2_decap_8 FILLER_45_1275 ();
 sg13g2_decap_8 FILLER_45_1282 ();
 sg13g2_decap_8 FILLER_45_1289 ();
 sg13g2_decap_8 FILLER_45_1296 ();
 sg13g2_decap_8 FILLER_45_1303 ();
 sg13g2_decap_4 FILLER_45_1310 ();
 sg13g2_fill_1 FILLER_45_1314 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_4 FILLER_46_175 ();
 sg13g2_fill_1 FILLER_46_179 ();
 sg13g2_fill_1 FILLER_46_184 ();
 sg13g2_fill_2 FILLER_46_230 ();
 sg13g2_fill_1 FILLER_46_232 ();
 sg13g2_fill_2 FILLER_46_260 ();
 sg13g2_decap_8 FILLER_46_288 ();
 sg13g2_decap_8 FILLER_46_295 ();
 sg13g2_fill_1 FILLER_46_302 ();
 sg13g2_fill_2 FILLER_46_337 ();
 sg13g2_fill_2 FILLER_46_361 ();
 sg13g2_fill_2 FILLER_46_371 ();
 sg13g2_fill_1 FILLER_46_373 ();
 sg13g2_fill_2 FILLER_46_379 ();
 sg13g2_fill_1 FILLER_46_381 ();
 sg13g2_fill_1 FILLER_46_453 ();
 sg13g2_fill_1 FILLER_46_490 ();
 sg13g2_decap_4 FILLER_46_516 ();
 sg13g2_decap_4 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_544 ();
 sg13g2_fill_2 FILLER_46_551 ();
 sg13g2_fill_1 FILLER_46_553 ();
 sg13g2_fill_2 FILLER_46_580 ();
 sg13g2_fill_1 FILLER_46_582 ();
 sg13g2_decap_8 FILLER_46_591 ();
 sg13g2_fill_2 FILLER_46_613 ();
 sg13g2_fill_1 FILLER_46_615 ();
 sg13g2_fill_1 FILLER_46_642 ();
 sg13g2_decap_8 FILLER_46_647 ();
 sg13g2_fill_1 FILLER_46_680 ();
 sg13g2_fill_2 FILLER_46_686 ();
 sg13g2_fill_1 FILLER_46_688 ();
 sg13g2_decap_4 FILLER_46_741 ();
 sg13g2_fill_1 FILLER_46_745 ();
 sg13g2_decap_4 FILLER_46_754 ();
 sg13g2_fill_2 FILLER_46_763 ();
 sg13g2_decap_8 FILLER_46_770 ();
 sg13g2_fill_1 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_782 ();
 sg13g2_decap_4 FILLER_46_819 ();
 sg13g2_fill_2 FILLER_46_823 ();
 sg13g2_fill_2 FILLER_46_828 ();
 sg13g2_fill_1 FILLER_46_830 ();
 sg13g2_fill_2 FILLER_46_847 ();
 sg13g2_fill_1 FILLER_46_849 ();
 sg13g2_decap_4 FILLER_46_862 ();
 sg13g2_fill_1 FILLER_46_889 ();
 sg13g2_fill_2 FILLER_46_906 ();
 sg13g2_fill_2 FILLER_46_995 ();
 sg13g2_fill_1 FILLER_46_997 ();
 sg13g2_fill_2 FILLER_46_1002 ();
 sg13g2_fill_2 FILLER_46_1026 ();
 sg13g2_fill_2 FILLER_46_1047 ();
 sg13g2_fill_1 FILLER_46_1049 ();
 sg13g2_decap_8 FILLER_46_1054 ();
 sg13g2_decap_8 FILLER_46_1061 ();
 sg13g2_decap_8 FILLER_46_1068 ();
 sg13g2_decap_8 FILLER_46_1075 ();
 sg13g2_decap_8 FILLER_46_1082 ();
 sg13g2_decap_8 FILLER_46_1089 ();
 sg13g2_decap_8 FILLER_46_1096 ();
 sg13g2_decap_8 FILLER_46_1103 ();
 sg13g2_decap_8 FILLER_46_1110 ();
 sg13g2_decap_8 FILLER_46_1117 ();
 sg13g2_decap_8 FILLER_46_1124 ();
 sg13g2_decap_8 FILLER_46_1131 ();
 sg13g2_decap_8 FILLER_46_1138 ();
 sg13g2_decap_8 FILLER_46_1145 ();
 sg13g2_decap_8 FILLER_46_1152 ();
 sg13g2_decap_8 FILLER_46_1159 ();
 sg13g2_decap_8 FILLER_46_1166 ();
 sg13g2_decap_8 FILLER_46_1173 ();
 sg13g2_decap_8 FILLER_46_1180 ();
 sg13g2_decap_8 FILLER_46_1187 ();
 sg13g2_decap_8 FILLER_46_1194 ();
 sg13g2_decap_8 FILLER_46_1201 ();
 sg13g2_decap_8 FILLER_46_1208 ();
 sg13g2_decap_8 FILLER_46_1215 ();
 sg13g2_decap_8 FILLER_46_1222 ();
 sg13g2_decap_8 FILLER_46_1229 ();
 sg13g2_decap_8 FILLER_46_1236 ();
 sg13g2_decap_8 FILLER_46_1243 ();
 sg13g2_decap_8 FILLER_46_1250 ();
 sg13g2_decap_8 FILLER_46_1257 ();
 sg13g2_decap_8 FILLER_46_1264 ();
 sg13g2_decap_8 FILLER_46_1271 ();
 sg13g2_decap_8 FILLER_46_1278 ();
 sg13g2_decap_8 FILLER_46_1285 ();
 sg13g2_decap_8 FILLER_46_1292 ();
 sg13g2_decap_8 FILLER_46_1299 ();
 sg13g2_decap_8 FILLER_46_1306 ();
 sg13g2_fill_2 FILLER_46_1313 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_4 FILLER_47_77 ();
 sg13g2_fill_1 FILLER_47_81 ();
 sg13g2_fill_2 FILLER_47_117 ();
 sg13g2_fill_1 FILLER_47_119 ();
 sg13g2_fill_2 FILLER_47_130 ();
 sg13g2_fill_2 FILLER_47_137 ();
 sg13g2_fill_1 FILLER_47_139 ();
 sg13g2_fill_1 FILLER_47_153 ();
 sg13g2_decap_8 FILLER_47_208 ();
 sg13g2_fill_1 FILLER_47_219 ();
 sg13g2_fill_2 FILLER_47_229 ();
 sg13g2_fill_2 FILLER_47_255 ();
 sg13g2_fill_1 FILLER_47_257 ();
 sg13g2_fill_2 FILLER_47_266 ();
 sg13g2_fill_1 FILLER_47_268 ();
 sg13g2_fill_2 FILLER_47_277 ();
 sg13g2_decap_4 FILLER_47_296 ();
 sg13g2_fill_1 FILLER_47_300 ();
 sg13g2_fill_2 FILLER_47_322 ();
 sg13g2_fill_2 FILLER_47_332 ();
 sg13g2_fill_1 FILLER_47_334 ();
 sg13g2_fill_1 FILLER_47_340 ();
 sg13g2_fill_2 FILLER_47_374 ();
 sg13g2_decap_4 FILLER_47_380 ();
 sg13g2_fill_2 FILLER_47_384 ();
 sg13g2_fill_2 FILLER_47_391 ();
 sg13g2_decap_4 FILLER_47_397 ();
 sg13g2_fill_1 FILLER_47_401 ();
 sg13g2_decap_4 FILLER_47_419 ();
 sg13g2_fill_2 FILLER_47_423 ();
 sg13g2_fill_1 FILLER_47_438 ();
 sg13g2_decap_4 FILLER_47_464 ();
 sg13g2_fill_2 FILLER_47_472 ();
 sg13g2_fill_1 FILLER_47_474 ();
 sg13g2_decap_4 FILLER_47_480 ();
 sg13g2_fill_2 FILLER_47_484 ();
 sg13g2_decap_8 FILLER_47_491 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_fill_1 FILLER_47_518 ();
 sg13g2_fill_2 FILLER_47_527 ();
 sg13g2_fill_2 FILLER_47_546 ();
 sg13g2_fill_1 FILLER_47_564 ();
 sg13g2_decap_8 FILLER_47_573 ();
 sg13g2_fill_2 FILLER_47_632 ();
 sg13g2_fill_1 FILLER_47_634 ();
 sg13g2_decap_4 FILLER_47_643 ();
 sg13g2_fill_2 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_657 ();
 sg13g2_fill_1 FILLER_47_664 ();
 sg13g2_fill_2 FILLER_47_669 ();
 sg13g2_decap_8 FILLER_47_710 ();
 sg13g2_fill_1 FILLER_47_717 ();
 sg13g2_decap_8 FILLER_47_804 ();
 sg13g2_fill_2 FILLER_47_811 ();
 sg13g2_decap_8 FILLER_47_836 ();
 sg13g2_fill_2 FILLER_47_843 ();
 sg13g2_fill_2 FILLER_47_862 ();
 sg13g2_fill_1 FILLER_47_880 ();
 sg13g2_fill_2 FILLER_47_896 ();
 sg13g2_decap_4 FILLER_47_902 ();
 sg13g2_fill_1 FILLER_47_906 ();
 sg13g2_decap_8 FILLER_47_915 ();
 sg13g2_decap_8 FILLER_47_922 ();
 sg13g2_decap_4 FILLER_47_929 ();
 sg13g2_fill_2 FILLER_47_933 ();
 sg13g2_fill_2 FILLER_47_940 ();
 sg13g2_decap_4 FILLER_47_952 ();
 sg13g2_fill_1 FILLER_47_956 ();
 sg13g2_fill_2 FILLER_47_974 ();
 sg13g2_decap_8 FILLER_47_1057 ();
 sg13g2_decap_8 FILLER_47_1064 ();
 sg13g2_decap_8 FILLER_47_1071 ();
 sg13g2_decap_8 FILLER_47_1078 ();
 sg13g2_decap_8 FILLER_47_1085 ();
 sg13g2_decap_8 FILLER_47_1092 ();
 sg13g2_decap_8 FILLER_47_1099 ();
 sg13g2_decap_8 FILLER_47_1106 ();
 sg13g2_decap_8 FILLER_47_1113 ();
 sg13g2_decap_8 FILLER_47_1120 ();
 sg13g2_decap_8 FILLER_47_1127 ();
 sg13g2_decap_8 FILLER_47_1134 ();
 sg13g2_decap_8 FILLER_47_1141 ();
 sg13g2_decap_8 FILLER_47_1148 ();
 sg13g2_decap_8 FILLER_47_1155 ();
 sg13g2_decap_8 FILLER_47_1162 ();
 sg13g2_decap_8 FILLER_47_1169 ();
 sg13g2_decap_8 FILLER_47_1176 ();
 sg13g2_decap_8 FILLER_47_1183 ();
 sg13g2_decap_8 FILLER_47_1190 ();
 sg13g2_decap_8 FILLER_47_1197 ();
 sg13g2_decap_8 FILLER_47_1204 ();
 sg13g2_decap_8 FILLER_47_1211 ();
 sg13g2_decap_8 FILLER_47_1218 ();
 sg13g2_decap_8 FILLER_47_1225 ();
 sg13g2_decap_8 FILLER_47_1232 ();
 sg13g2_decap_8 FILLER_47_1239 ();
 sg13g2_decap_8 FILLER_47_1246 ();
 sg13g2_decap_8 FILLER_47_1253 ();
 sg13g2_decap_8 FILLER_47_1260 ();
 sg13g2_decap_8 FILLER_47_1267 ();
 sg13g2_decap_8 FILLER_47_1274 ();
 sg13g2_decap_8 FILLER_47_1281 ();
 sg13g2_decap_8 FILLER_47_1288 ();
 sg13g2_decap_8 FILLER_47_1295 ();
 sg13g2_decap_8 FILLER_47_1302 ();
 sg13g2_decap_4 FILLER_47_1309 ();
 sg13g2_fill_2 FILLER_47_1313 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_4 FILLER_48_84 ();
 sg13g2_fill_1 FILLER_48_88 ();
 sg13g2_decap_4 FILLER_48_125 ();
 sg13g2_fill_2 FILLER_48_129 ();
 sg13g2_fill_2 FILLER_48_175 ();
 sg13g2_fill_2 FILLER_48_190 ();
 sg13g2_fill_2 FILLER_48_201 ();
 sg13g2_fill_1 FILLER_48_229 ();
 sg13g2_fill_1 FILLER_48_239 ();
 sg13g2_decap_4 FILLER_48_263 ();
 sg13g2_fill_2 FILLER_48_267 ();
 sg13g2_fill_2 FILLER_48_409 ();
 sg13g2_decap_8 FILLER_48_437 ();
 sg13g2_fill_2 FILLER_48_444 ();
 sg13g2_fill_2 FILLER_48_454 ();
 sg13g2_fill_1 FILLER_48_456 ();
 sg13g2_decap_8 FILLER_48_503 ();
 sg13g2_decap_4 FILLER_48_538 ();
 sg13g2_decap_8 FILLER_48_549 ();
 sg13g2_decap_4 FILLER_48_556 ();
 sg13g2_fill_1 FILLER_48_560 ();
 sg13g2_decap_4 FILLER_48_584 ();
 sg13g2_fill_2 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_594 ();
 sg13g2_decap_8 FILLER_48_601 ();
 sg13g2_decap_4 FILLER_48_608 ();
 sg13g2_fill_2 FILLER_48_621 ();
 sg13g2_decap_8 FILLER_48_649 ();
 sg13g2_decap_4 FILLER_48_671 ();
 sg13g2_fill_2 FILLER_48_684 ();
 sg13g2_fill_1 FILLER_48_686 ();
 sg13g2_decap_4 FILLER_48_691 ();
 sg13g2_fill_2 FILLER_48_695 ();
 sg13g2_fill_2 FILLER_48_707 ();
 sg13g2_fill_2 FILLER_48_739 ();
 sg13g2_fill_1 FILLER_48_741 ();
 sg13g2_decap_4 FILLER_48_747 ();
 sg13g2_fill_1 FILLER_48_751 ();
 sg13g2_fill_2 FILLER_48_756 ();
 sg13g2_fill_1 FILLER_48_758 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_fill_2 FILLER_48_777 ();
 sg13g2_fill_1 FILLER_48_779 ();
 sg13g2_decap_4 FILLER_48_805 ();
 sg13g2_fill_1 FILLER_48_809 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_fill_2 FILLER_48_822 ();
 sg13g2_fill_2 FILLER_48_829 ();
 sg13g2_fill_1 FILLER_48_831 ();
 sg13g2_fill_1 FILLER_48_836 ();
 sg13g2_fill_2 FILLER_48_844 ();
 sg13g2_fill_1 FILLER_48_846 ();
 sg13g2_decap_8 FILLER_48_856 ();
 sg13g2_decap_8 FILLER_48_863 ();
 sg13g2_fill_2 FILLER_48_882 ();
 sg13g2_fill_2 FILLER_48_904 ();
 sg13g2_fill_1 FILLER_48_906 ();
 sg13g2_decap_4 FILLER_48_925 ();
 sg13g2_decap_8 FILLER_48_933 ();
 sg13g2_decap_8 FILLER_48_944 ();
 sg13g2_fill_2 FILLER_48_951 ();
 sg13g2_fill_2 FILLER_48_984 ();
 sg13g2_fill_1 FILLER_48_986 ();
 sg13g2_fill_2 FILLER_48_1027 ();
 sg13g2_fill_1 FILLER_48_1029 ();
 sg13g2_decap_8 FILLER_48_1057 ();
 sg13g2_decap_8 FILLER_48_1064 ();
 sg13g2_decap_8 FILLER_48_1071 ();
 sg13g2_decap_8 FILLER_48_1078 ();
 sg13g2_decap_8 FILLER_48_1085 ();
 sg13g2_decap_8 FILLER_48_1092 ();
 sg13g2_decap_8 FILLER_48_1099 ();
 sg13g2_decap_8 FILLER_48_1106 ();
 sg13g2_decap_8 FILLER_48_1113 ();
 sg13g2_decap_8 FILLER_48_1120 ();
 sg13g2_decap_8 FILLER_48_1127 ();
 sg13g2_decap_8 FILLER_48_1134 ();
 sg13g2_decap_8 FILLER_48_1141 ();
 sg13g2_decap_8 FILLER_48_1148 ();
 sg13g2_decap_8 FILLER_48_1155 ();
 sg13g2_decap_8 FILLER_48_1162 ();
 sg13g2_decap_8 FILLER_48_1169 ();
 sg13g2_decap_8 FILLER_48_1176 ();
 sg13g2_decap_8 FILLER_48_1183 ();
 sg13g2_decap_8 FILLER_48_1190 ();
 sg13g2_decap_8 FILLER_48_1197 ();
 sg13g2_decap_8 FILLER_48_1204 ();
 sg13g2_decap_8 FILLER_48_1211 ();
 sg13g2_decap_8 FILLER_48_1218 ();
 sg13g2_decap_8 FILLER_48_1225 ();
 sg13g2_decap_8 FILLER_48_1232 ();
 sg13g2_decap_8 FILLER_48_1239 ();
 sg13g2_decap_8 FILLER_48_1246 ();
 sg13g2_decap_8 FILLER_48_1253 ();
 sg13g2_decap_8 FILLER_48_1260 ();
 sg13g2_decap_8 FILLER_48_1267 ();
 sg13g2_decap_8 FILLER_48_1274 ();
 sg13g2_decap_8 FILLER_48_1281 ();
 sg13g2_decap_8 FILLER_48_1288 ();
 sg13g2_decap_8 FILLER_48_1295 ();
 sg13g2_decap_8 FILLER_48_1302 ();
 sg13g2_decap_4 FILLER_48_1309 ();
 sg13g2_fill_2 FILLER_48_1313 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_4 FILLER_49_84 ();
 sg13g2_fill_1 FILLER_49_88 ();
 sg13g2_fill_2 FILLER_49_97 ();
 sg13g2_fill_2 FILLER_49_112 ();
 sg13g2_fill_1 FILLER_49_114 ();
 sg13g2_decap_4 FILLER_49_128 ();
 sg13g2_fill_1 FILLER_49_132 ();
 sg13g2_fill_1 FILLER_49_142 ();
 sg13g2_fill_2 FILLER_49_211 ();
 sg13g2_fill_1 FILLER_49_213 ();
 sg13g2_fill_1 FILLER_49_218 ();
 sg13g2_fill_1 FILLER_49_234 ();
 sg13g2_fill_2 FILLER_49_261 ();
 sg13g2_fill_2 FILLER_49_294 ();
 sg13g2_fill_1 FILLER_49_296 ();
 sg13g2_fill_1 FILLER_49_319 ();
 sg13g2_decap_8 FILLER_49_328 ();
 sg13g2_fill_2 FILLER_49_335 ();
 sg13g2_fill_2 FILLER_49_349 ();
 sg13g2_fill_1 FILLER_49_402 ();
 sg13g2_decap_8 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_49_414 ();
 sg13g2_decap_8 FILLER_49_421 ();
 sg13g2_decap_8 FILLER_49_428 ();
 sg13g2_fill_2 FILLER_49_435 ();
 sg13g2_fill_2 FILLER_49_473 ();
 sg13g2_fill_2 FILLER_49_483 ();
 sg13g2_fill_1 FILLER_49_485 ();
 sg13g2_fill_2 FILLER_49_515 ();
 sg13g2_fill_1 FILLER_49_517 ();
 sg13g2_fill_2 FILLER_49_531 ();
 sg13g2_decap_4 FILLER_49_611 ();
 sg13g2_fill_1 FILLER_49_625 ();
 sg13g2_fill_2 FILLER_49_691 ();
 sg13g2_decap_8 FILLER_49_736 ();
 sg13g2_decap_8 FILLER_49_748 ();
 sg13g2_fill_1 FILLER_49_755 ();
 sg13g2_fill_1 FILLER_49_766 ();
 sg13g2_fill_1 FILLER_49_791 ();
 sg13g2_decap_4 FILLER_49_797 ();
 sg13g2_fill_1 FILLER_49_841 ();
 sg13g2_fill_1 FILLER_49_864 ();
 sg13g2_decap_8 FILLER_49_873 ();
 sg13g2_fill_1 FILLER_49_880 ();
 sg13g2_fill_2 FILLER_49_885 ();
 sg13g2_fill_2 FILLER_49_900 ();
 sg13g2_fill_2 FILLER_49_955 ();
 sg13g2_fill_2 FILLER_49_976 ();
 sg13g2_fill_1 FILLER_49_978 ();
 sg13g2_fill_2 FILLER_49_1001 ();
 sg13g2_fill_1 FILLER_49_1003 ();
 sg13g2_decap_8 FILLER_49_1060 ();
 sg13g2_decap_8 FILLER_49_1067 ();
 sg13g2_decap_8 FILLER_49_1074 ();
 sg13g2_decap_8 FILLER_49_1081 ();
 sg13g2_decap_8 FILLER_49_1088 ();
 sg13g2_decap_8 FILLER_49_1095 ();
 sg13g2_decap_8 FILLER_49_1102 ();
 sg13g2_decap_8 FILLER_49_1109 ();
 sg13g2_decap_8 FILLER_49_1116 ();
 sg13g2_decap_8 FILLER_49_1123 ();
 sg13g2_decap_8 FILLER_49_1130 ();
 sg13g2_decap_8 FILLER_49_1137 ();
 sg13g2_decap_8 FILLER_49_1144 ();
 sg13g2_decap_8 FILLER_49_1151 ();
 sg13g2_decap_8 FILLER_49_1158 ();
 sg13g2_decap_8 FILLER_49_1165 ();
 sg13g2_decap_8 FILLER_49_1172 ();
 sg13g2_decap_8 FILLER_49_1179 ();
 sg13g2_decap_8 FILLER_49_1186 ();
 sg13g2_decap_8 FILLER_49_1193 ();
 sg13g2_decap_8 FILLER_49_1200 ();
 sg13g2_decap_8 FILLER_49_1207 ();
 sg13g2_decap_8 FILLER_49_1214 ();
 sg13g2_decap_8 FILLER_49_1221 ();
 sg13g2_decap_8 FILLER_49_1228 ();
 sg13g2_decap_8 FILLER_49_1235 ();
 sg13g2_decap_8 FILLER_49_1242 ();
 sg13g2_decap_8 FILLER_49_1249 ();
 sg13g2_decap_8 FILLER_49_1256 ();
 sg13g2_decap_8 FILLER_49_1263 ();
 sg13g2_decap_8 FILLER_49_1270 ();
 sg13g2_decap_8 FILLER_49_1277 ();
 sg13g2_decap_8 FILLER_49_1284 ();
 sg13g2_decap_8 FILLER_49_1291 ();
 sg13g2_decap_8 FILLER_49_1298 ();
 sg13g2_decap_8 FILLER_49_1305 ();
 sg13g2_fill_2 FILLER_49_1312 ();
 sg13g2_fill_1 FILLER_49_1314 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_4 FILLER_50_77 ();
 sg13g2_fill_2 FILLER_50_81 ();
 sg13g2_fill_1 FILLER_50_109 ();
 sg13g2_fill_1 FILLER_50_150 ();
 sg13g2_fill_2 FILLER_50_165 ();
 sg13g2_fill_1 FILLER_50_180 ();
 sg13g2_fill_1 FILLER_50_206 ();
 sg13g2_fill_2 FILLER_50_221 ();
 sg13g2_decap_8 FILLER_50_228 ();
 sg13g2_fill_1 FILLER_50_235 ();
 sg13g2_decap_4 FILLER_50_241 ();
 sg13g2_fill_1 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_250 ();
 sg13g2_decap_4 FILLER_50_257 ();
 sg13g2_fill_2 FILLER_50_270 ();
 sg13g2_fill_1 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_321 ();
 sg13g2_fill_1 FILLER_50_327 ();
 sg13g2_decap_8 FILLER_50_332 ();
 sg13g2_decap_4 FILLER_50_339 ();
 sg13g2_decap_4 FILLER_50_389 ();
 sg13g2_fill_1 FILLER_50_436 ();
 sg13g2_fill_2 FILLER_50_450 ();
 sg13g2_fill_2 FILLER_50_476 ();
 sg13g2_fill_2 FILLER_50_488 ();
 sg13g2_fill_1 FILLER_50_490 ();
 sg13g2_decap_4 FILLER_50_511 ();
 sg13g2_fill_2 FILLER_50_515 ();
 sg13g2_fill_2 FILLER_50_522 ();
 sg13g2_decap_4 FILLER_50_532 ();
 sg13g2_decap_8 FILLER_50_553 ();
 sg13g2_decap_4 FILLER_50_565 ();
 sg13g2_fill_1 FILLER_50_569 ();
 sg13g2_fill_1 FILLER_50_583 ();
 sg13g2_decap_4 FILLER_50_633 ();
 sg13g2_fill_2 FILLER_50_637 ();
 sg13g2_fill_1 FILLER_50_653 ();
 sg13g2_decap_8 FILLER_50_667 ();
 sg13g2_fill_2 FILLER_50_674 ();
 sg13g2_decap_4 FILLER_50_680 ();
 sg13g2_decap_8 FILLER_50_694 ();
 sg13g2_fill_2 FILLER_50_701 ();
 sg13g2_decap_4 FILLER_50_716 ();
 sg13g2_fill_1 FILLER_50_720 ();
 sg13g2_fill_2 FILLER_50_736 ();
 sg13g2_fill_1 FILLER_50_738 ();
 sg13g2_fill_2 FILLER_50_754 ();
 sg13g2_fill_1 FILLER_50_756 ();
 sg13g2_fill_2 FILLER_50_777 ();
 sg13g2_decap_8 FILLER_50_783 ();
 sg13g2_decap_8 FILLER_50_790 ();
 sg13g2_decap_4 FILLER_50_818 ();
 sg13g2_fill_2 FILLER_50_831 ();
 sg13g2_decap_4 FILLER_50_838 ();
 sg13g2_fill_1 FILLER_50_842 ();
 sg13g2_decap_4 FILLER_50_852 ();
 sg13g2_fill_2 FILLER_50_861 ();
 sg13g2_fill_2 FILLER_50_886 ();
 sg13g2_fill_1 FILLER_50_888 ();
 sg13g2_decap_8 FILLER_50_899 ();
 sg13g2_fill_1 FILLER_50_906 ();
 sg13g2_decap_8 FILLER_50_922 ();
 sg13g2_decap_8 FILLER_50_929 ();
 sg13g2_decap_4 FILLER_50_936 ();
 sg13g2_fill_1 FILLER_50_940 ();
 sg13g2_decap_8 FILLER_50_945 ();
 sg13g2_decap_4 FILLER_50_952 ();
 sg13g2_fill_1 FILLER_50_956 ();
 sg13g2_fill_1 FILLER_50_995 ();
 sg13g2_fill_2 FILLER_50_1013 ();
 sg13g2_fill_1 FILLER_50_1019 ();
 sg13g2_decap_8 FILLER_50_1050 ();
 sg13g2_decap_8 FILLER_50_1057 ();
 sg13g2_decap_8 FILLER_50_1064 ();
 sg13g2_decap_8 FILLER_50_1071 ();
 sg13g2_decap_8 FILLER_50_1078 ();
 sg13g2_decap_8 FILLER_50_1085 ();
 sg13g2_decap_8 FILLER_50_1092 ();
 sg13g2_decap_8 FILLER_50_1099 ();
 sg13g2_decap_8 FILLER_50_1106 ();
 sg13g2_decap_8 FILLER_50_1113 ();
 sg13g2_decap_8 FILLER_50_1120 ();
 sg13g2_decap_8 FILLER_50_1127 ();
 sg13g2_decap_8 FILLER_50_1134 ();
 sg13g2_decap_8 FILLER_50_1141 ();
 sg13g2_decap_8 FILLER_50_1148 ();
 sg13g2_decap_8 FILLER_50_1155 ();
 sg13g2_decap_8 FILLER_50_1162 ();
 sg13g2_decap_8 FILLER_50_1169 ();
 sg13g2_decap_8 FILLER_50_1176 ();
 sg13g2_decap_8 FILLER_50_1183 ();
 sg13g2_decap_8 FILLER_50_1190 ();
 sg13g2_decap_8 FILLER_50_1197 ();
 sg13g2_decap_8 FILLER_50_1204 ();
 sg13g2_decap_8 FILLER_50_1211 ();
 sg13g2_decap_8 FILLER_50_1218 ();
 sg13g2_decap_8 FILLER_50_1225 ();
 sg13g2_decap_8 FILLER_50_1232 ();
 sg13g2_decap_8 FILLER_50_1239 ();
 sg13g2_decap_8 FILLER_50_1246 ();
 sg13g2_decap_8 FILLER_50_1253 ();
 sg13g2_decap_8 FILLER_50_1260 ();
 sg13g2_decap_8 FILLER_50_1267 ();
 sg13g2_decap_8 FILLER_50_1274 ();
 sg13g2_decap_8 FILLER_50_1281 ();
 sg13g2_decap_8 FILLER_50_1288 ();
 sg13g2_decap_8 FILLER_50_1295 ();
 sg13g2_decap_8 FILLER_50_1302 ();
 sg13g2_decap_4 FILLER_50_1309 ();
 sg13g2_fill_2 FILLER_50_1313 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_fill_2 FILLER_51_115 ();
 sg13g2_fill_2 FILLER_51_132 ();
 sg13g2_fill_1 FILLER_51_134 ();
 sg13g2_fill_2 FILLER_51_201 ();
 sg13g2_fill_1 FILLER_51_203 ();
 sg13g2_fill_1 FILLER_51_266 ();
 sg13g2_fill_2 FILLER_51_292 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_325 ();
 sg13g2_fill_1 FILLER_51_332 ();
 sg13g2_decap_8 FILLER_51_346 ();
 sg13g2_fill_2 FILLER_51_353 ();
 sg13g2_decap_4 FILLER_51_363 ();
 sg13g2_fill_2 FILLER_51_381 ();
 sg13g2_fill_2 FILLER_51_388 ();
 sg13g2_fill_1 FILLER_51_390 ();
 sg13g2_fill_2 FILLER_51_399 ();
 sg13g2_fill_1 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_426 ();
 sg13g2_fill_2 FILLER_51_432 ();
 sg13g2_fill_1 FILLER_51_444 ();
 sg13g2_fill_2 FILLER_51_480 ();
 sg13g2_fill_1 FILLER_51_494 ();
 sg13g2_decap_4 FILLER_51_499 ();
 sg13g2_fill_2 FILLER_51_537 ();
 sg13g2_fill_1 FILLER_51_539 ();
 sg13g2_fill_2 FILLER_51_591 ();
 sg13g2_fill_1 FILLER_51_593 ();
 sg13g2_fill_1 FILLER_51_611 ();
 sg13g2_fill_1 FILLER_51_630 ();
 sg13g2_fill_2 FILLER_51_635 ();
 sg13g2_fill_2 FILLER_51_673 ();
 sg13g2_fill_1 FILLER_51_688 ();
 sg13g2_fill_2 FILLER_51_729 ();
 sg13g2_fill_1 FILLER_51_731 ();
 sg13g2_decap_4 FILLER_51_750 ();
 sg13g2_fill_2 FILLER_51_754 ();
 sg13g2_decap_8 FILLER_51_764 ();
 sg13g2_fill_1 FILLER_51_771 ();
 sg13g2_decap_4 FILLER_51_787 ();
 sg13g2_fill_1 FILLER_51_791 ();
 sg13g2_decap_4 FILLER_51_804 ();
 sg13g2_decap_4 FILLER_51_830 ();
 sg13g2_decap_4 FILLER_51_846 ();
 sg13g2_fill_2 FILLER_51_850 ();
 sg13g2_decap_8 FILLER_51_860 ();
 sg13g2_fill_2 FILLER_51_867 ();
 sg13g2_fill_1 FILLER_51_869 ();
 sg13g2_fill_1 FILLER_51_922 ();
 sg13g2_fill_1 FILLER_51_956 ();
 sg13g2_decap_4 FILLER_51_969 ();
 sg13g2_decap_4 FILLER_51_986 ();
 sg13g2_fill_1 FILLER_51_1016 ();
 sg13g2_decap_8 FILLER_51_1040 ();
 sg13g2_decap_8 FILLER_51_1047 ();
 sg13g2_decap_8 FILLER_51_1054 ();
 sg13g2_decap_8 FILLER_51_1061 ();
 sg13g2_decap_8 FILLER_51_1068 ();
 sg13g2_decap_8 FILLER_51_1075 ();
 sg13g2_decap_8 FILLER_51_1082 ();
 sg13g2_decap_8 FILLER_51_1089 ();
 sg13g2_decap_8 FILLER_51_1096 ();
 sg13g2_decap_8 FILLER_51_1103 ();
 sg13g2_decap_8 FILLER_51_1110 ();
 sg13g2_decap_8 FILLER_51_1117 ();
 sg13g2_decap_8 FILLER_51_1124 ();
 sg13g2_decap_8 FILLER_51_1131 ();
 sg13g2_decap_8 FILLER_51_1138 ();
 sg13g2_decap_8 FILLER_51_1145 ();
 sg13g2_decap_8 FILLER_51_1152 ();
 sg13g2_decap_8 FILLER_51_1159 ();
 sg13g2_decap_8 FILLER_51_1166 ();
 sg13g2_decap_8 FILLER_51_1173 ();
 sg13g2_decap_8 FILLER_51_1180 ();
 sg13g2_decap_8 FILLER_51_1187 ();
 sg13g2_decap_8 FILLER_51_1194 ();
 sg13g2_decap_8 FILLER_51_1201 ();
 sg13g2_decap_8 FILLER_51_1208 ();
 sg13g2_decap_8 FILLER_51_1215 ();
 sg13g2_decap_8 FILLER_51_1222 ();
 sg13g2_decap_8 FILLER_51_1229 ();
 sg13g2_decap_8 FILLER_51_1236 ();
 sg13g2_decap_8 FILLER_51_1243 ();
 sg13g2_decap_8 FILLER_51_1250 ();
 sg13g2_decap_8 FILLER_51_1257 ();
 sg13g2_decap_8 FILLER_51_1264 ();
 sg13g2_decap_8 FILLER_51_1271 ();
 sg13g2_decap_8 FILLER_51_1278 ();
 sg13g2_decap_8 FILLER_51_1285 ();
 sg13g2_decap_8 FILLER_51_1292 ();
 sg13g2_decap_8 FILLER_51_1299 ();
 sg13g2_decap_8 FILLER_51_1306 ();
 sg13g2_fill_2 FILLER_51_1313 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_fill_2 FILLER_52_91 ();
 sg13g2_fill_1 FILLER_52_93 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_fill_2 FILLER_52_105 ();
 sg13g2_fill_2 FILLER_52_120 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_fill_1 FILLER_52_165 ();
 sg13g2_decap_4 FILLER_52_170 ();
 sg13g2_fill_1 FILLER_52_218 ();
 sg13g2_decap_4 FILLER_52_234 ();
 sg13g2_fill_1 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_261 ();
 sg13g2_fill_1 FILLER_52_263 ();
 sg13g2_fill_2 FILLER_52_333 ();
 sg13g2_fill_2 FILLER_52_344 ();
 sg13g2_decap_4 FILLER_52_359 ();
 sg13g2_fill_2 FILLER_52_373 ();
 sg13g2_fill_1 FILLER_52_375 ();
 sg13g2_decap_4 FILLER_52_414 ();
 sg13g2_fill_1 FILLER_52_423 ();
 sg13g2_fill_2 FILLER_52_450 ();
 sg13g2_fill_1 FILLER_52_452 ();
 sg13g2_fill_1 FILLER_52_458 ();
 sg13g2_fill_1 FILLER_52_464 ();
 sg13g2_decap_8 FILLER_52_473 ();
 sg13g2_fill_2 FILLER_52_480 ();
 sg13g2_fill_2 FILLER_52_487 ();
 sg13g2_fill_1 FILLER_52_489 ();
 sg13g2_fill_2 FILLER_52_519 ();
 sg13g2_fill_1 FILLER_52_521 ();
 sg13g2_decap_8 FILLER_52_526 ();
 sg13g2_decap_8 FILLER_52_533 ();
 sg13g2_decap_4 FILLER_52_540 ();
 sg13g2_fill_2 FILLER_52_544 ();
 sg13g2_fill_1 FILLER_52_550 ();
 sg13g2_fill_2 FILLER_52_564 ();
 sg13g2_fill_1 FILLER_52_579 ();
 sg13g2_decap_8 FILLER_52_695 ();
 sg13g2_decap_8 FILLER_52_702 ();
 sg13g2_fill_2 FILLER_52_722 ();
 sg13g2_fill_1 FILLER_52_724 ();
 sg13g2_decap_8 FILLER_52_729 ();
 sg13g2_fill_2 FILLER_52_736 ();
 sg13g2_fill_2 FILLER_52_759 ();
 sg13g2_fill_1 FILLER_52_775 ();
 sg13g2_decap_8 FILLER_52_793 ();
 sg13g2_fill_1 FILLER_52_811 ();
 sg13g2_decap_4 FILLER_52_816 ();
 sg13g2_decap_4 FILLER_52_825 ();
 sg13g2_fill_1 FILLER_52_829 ();
 sg13g2_fill_1 FILLER_52_835 ();
 sg13g2_decap_4 FILLER_52_841 ();
 sg13g2_fill_2 FILLER_52_845 ();
 sg13g2_decap_4 FILLER_52_867 ();
 sg13g2_fill_1 FILLER_52_871 ();
 sg13g2_decap_8 FILLER_52_927 ();
 sg13g2_decap_4 FILLER_52_934 ();
 sg13g2_fill_1 FILLER_52_938 ();
 sg13g2_fill_2 FILLER_52_951 ();
 sg13g2_fill_1 FILLER_52_953 ();
 sg13g2_fill_2 FILLER_52_959 ();
 sg13g2_fill_1 FILLER_52_961 ();
 sg13g2_fill_2 FILLER_52_967 ();
 sg13g2_fill_1 FILLER_52_969 ();
 sg13g2_decap_4 FILLER_52_1022 ();
 sg13g2_decap_8 FILLER_52_1052 ();
 sg13g2_decap_8 FILLER_52_1059 ();
 sg13g2_decap_8 FILLER_52_1066 ();
 sg13g2_decap_8 FILLER_52_1073 ();
 sg13g2_decap_8 FILLER_52_1080 ();
 sg13g2_decap_8 FILLER_52_1087 ();
 sg13g2_decap_8 FILLER_52_1094 ();
 sg13g2_decap_8 FILLER_52_1101 ();
 sg13g2_decap_8 FILLER_52_1108 ();
 sg13g2_decap_8 FILLER_52_1115 ();
 sg13g2_decap_8 FILLER_52_1122 ();
 sg13g2_decap_8 FILLER_52_1129 ();
 sg13g2_decap_8 FILLER_52_1136 ();
 sg13g2_decap_8 FILLER_52_1143 ();
 sg13g2_decap_8 FILLER_52_1150 ();
 sg13g2_decap_8 FILLER_52_1157 ();
 sg13g2_decap_8 FILLER_52_1164 ();
 sg13g2_decap_8 FILLER_52_1171 ();
 sg13g2_decap_8 FILLER_52_1178 ();
 sg13g2_decap_8 FILLER_52_1185 ();
 sg13g2_decap_8 FILLER_52_1192 ();
 sg13g2_decap_8 FILLER_52_1199 ();
 sg13g2_decap_8 FILLER_52_1206 ();
 sg13g2_decap_8 FILLER_52_1213 ();
 sg13g2_decap_8 FILLER_52_1220 ();
 sg13g2_decap_8 FILLER_52_1227 ();
 sg13g2_decap_8 FILLER_52_1234 ();
 sg13g2_decap_8 FILLER_52_1241 ();
 sg13g2_decap_8 FILLER_52_1248 ();
 sg13g2_decap_8 FILLER_52_1255 ();
 sg13g2_decap_8 FILLER_52_1262 ();
 sg13g2_decap_8 FILLER_52_1269 ();
 sg13g2_decap_8 FILLER_52_1276 ();
 sg13g2_decap_8 FILLER_52_1283 ();
 sg13g2_decap_8 FILLER_52_1290 ();
 sg13g2_decap_8 FILLER_52_1297 ();
 sg13g2_decap_8 FILLER_52_1304 ();
 sg13g2_decap_4 FILLER_52_1311 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_4 FILLER_53_84 ();
 sg13g2_fill_2 FILLER_53_114 ();
 sg13g2_fill_1 FILLER_53_121 ();
 sg13g2_fill_1 FILLER_53_148 ();
 sg13g2_fill_2 FILLER_53_167 ();
 sg13g2_fill_2 FILLER_53_204 ();
 sg13g2_fill_2 FILLER_53_215 ();
 sg13g2_fill_1 FILLER_53_217 ();
 sg13g2_fill_1 FILLER_53_222 ();
 sg13g2_decap_8 FILLER_53_227 ();
 sg13g2_fill_2 FILLER_53_234 ();
 sg13g2_fill_2 FILLER_53_241 ();
 sg13g2_fill_1 FILLER_53_243 ();
 sg13g2_fill_2 FILLER_53_274 ();
 sg13g2_fill_1 FILLER_53_276 ();
 sg13g2_fill_2 FILLER_53_282 ();
 sg13g2_fill_1 FILLER_53_284 ();
 sg13g2_fill_1 FILLER_53_302 ();
 sg13g2_fill_1 FILLER_53_337 ();
 sg13g2_decap_8 FILLER_53_346 ();
 sg13g2_fill_1 FILLER_53_353 ();
 sg13g2_fill_1 FILLER_53_375 ();
 sg13g2_fill_2 FILLER_53_385 ();
 sg13g2_fill_2 FILLER_53_404 ();
 sg13g2_fill_1 FILLER_53_406 ();
 sg13g2_fill_2 FILLER_53_450 ();
 sg13g2_fill_1 FILLER_53_452 ();
 sg13g2_decap_8 FILLER_53_492 ();
 sg13g2_decap_8 FILLER_53_499 ();
 sg13g2_fill_1 FILLER_53_506 ();
 sg13g2_fill_1 FILLER_53_510 ();
 sg13g2_fill_1 FILLER_53_543 ();
 sg13g2_fill_1 FILLER_53_591 ();
 sg13g2_decap_4 FILLER_53_597 ();
 sg13g2_decap_8 FILLER_53_613 ();
 sg13g2_fill_2 FILLER_53_620 ();
 sg13g2_fill_1 FILLER_53_622 ();
 sg13g2_fill_2 FILLER_53_645 ();
 sg13g2_decap_8 FILLER_53_681 ();
 sg13g2_fill_2 FILLER_53_688 ();
 sg13g2_decap_8 FILLER_53_738 ();
 sg13g2_fill_2 FILLER_53_745 ();
 sg13g2_fill_1 FILLER_53_747 ();
 sg13g2_fill_1 FILLER_53_757 ();
 sg13g2_fill_2 FILLER_53_784 ();
 sg13g2_fill_2 FILLER_53_795 ();
 sg13g2_fill_1 FILLER_53_797 ();
 sg13g2_decap_8 FILLER_53_808 ();
 sg13g2_decap_8 FILLER_53_815 ();
 sg13g2_fill_1 FILLER_53_822 ();
 sg13g2_fill_1 FILLER_53_844 ();
 sg13g2_decap_8 FILLER_53_849 ();
 sg13g2_fill_1 FILLER_53_856 ();
 sg13g2_decap_8 FILLER_53_861 ();
 sg13g2_decap_4 FILLER_53_873 ();
 sg13g2_fill_1 FILLER_53_877 ();
 sg13g2_decap_8 FILLER_53_888 ();
 sg13g2_fill_1 FILLER_53_895 ();
 sg13g2_decap_8 FILLER_53_900 ();
 sg13g2_fill_2 FILLER_53_907 ();
 sg13g2_fill_1 FILLER_53_909 ();
 sg13g2_decap_4 FILLER_53_937 ();
 sg13g2_fill_2 FILLER_53_941 ();
 sg13g2_decap_4 FILLER_53_957 ();
 sg13g2_fill_2 FILLER_53_971 ();
 sg13g2_fill_1 FILLER_53_973 ();
 sg13g2_decap_8 FILLER_53_1045 ();
 sg13g2_decap_8 FILLER_53_1052 ();
 sg13g2_decap_8 FILLER_53_1059 ();
 sg13g2_decap_8 FILLER_53_1066 ();
 sg13g2_decap_8 FILLER_53_1073 ();
 sg13g2_decap_8 FILLER_53_1080 ();
 sg13g2_decap_8 FILLER_53_1087 ();
 sg13g2_decap_8 FILLER_53_1094 ();
 sg13g2_decap_8 FILLER_53_1101 ();
 sg13g2_decap_8 FILLER_53_1108 ();
 sg13g2_decap_8 FILLER_53_1115 ();
 sg13g2_decap_8 FILLER_53_1122 ();
 sg13g2_decap_8 FILLER_53_1129 ();
 sg13g2_decap_8 FILLER_53_1136 ();
 sg13g2_decap_8 FILLER_53_1143 ();
 sg13g2_decap_8 FILLER_53_1150 ();
 sg13g2_decap_8 FILLER_53_1157 ();
 sg13g2_decap_8 FILLER_53_1164 ();
 sg13g2_decap_8 FILLER_53_1171 ();
 sg13g2_decap_8 FILLER_53_1178 ();
 sg13g2_decap_8 FILLER_53_1185 ();
 sg13g2_decap_8 FILLER_53_1192 ();
 sg13g2_decap_8 FILLER_53_1199 ();
 sg13g2_decap_8 FILLER_53_1206 ();
 sg13g2_decap_8 FILLER_53_1213 ();
 sg13g2_decap_8 FILLER_53_1220 ();
 sg13g2_decap_8 FILLER_53_1227 ();
 sg13g2_decap_8 FILLER_53_1234 ();
 sg13g2_decap_8 FILLER_53_1241 ();
 sg13g2_decap_8 FILLER_53_1248 ();
 sg13g2_decap_8 FILLER_53_1255 ();
 sg13g2_decap_8 FILLER_53_1262 ();
 sg13g2_decap_8 FILLER_53_1269 ();
 sg13g2_decap_8 FILLER_53_1276 ();
 sg13g2_decap_8 FILLER_53_1283 ();
 sg13g2_decap_8 FILLER_53_1290 ();
 sg13g2_decap_8 FILLER_53_1297 ();
 sg13g2_decap_8 FILLER_53_1304 ();
 sg13g2_decap_4 FILLER_53_1311 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_fill_1 FILLER_54_91 ();
 sg13g2_fill_1 FILLER_54_113 ();
 sg13g2_fill_2 FILLER_54_124 ();
 sg13g2_fill_1 FILLER_54_126 ();
 sg13g2_fill_2 FILLER_54_131 ();
 sg13g2_fill_1 FILLER_54_141 ();
 sg13g2_fill_1 FILLER_54_181 ();
 sg13g2_fill_2 FILLER_54_243 ();
 sg13g2_fill_1 FILLER_54_245 ();
 sg13g2_fill_2 FILLER_54_274 ();
 sg13g2_fill_1 FILLER_54_276 ();
 sg13g2_fill_2 FILLER_54_281 ();
 sg13g2_fill_2 FILLER_54_288 ();
 sg13g2_fill_2 FILLER_54_298 ();
 sg13g2_fill_1 FILLER_54_338 ();
 sg13g2_decap_4 FILLER_54_344 ();
 sg13g2_fill_2 FILLER_54_348 ();
 sg13g2_decap_8 FILLER_54_363 ();
 sg13g2_decap_4 FILLER_54_370 ();
 sg13g2_fill_2 FILLER_54_374 ();
 sg13g2_fill_2 FILLER_54_380 ();
 sg13g2_fill_1 FILLER_54_382 ();
 sg13g2_fill_1 FILLER_54_401 ();
 sg13g2_fill_1 FILLER_54_412 ();
 sg13g2_fill_2 FILLER_54_421 ();
 sg13g2_fill_1 FILLER_54_423 ();
 sg13g2_fill_1 FILLER_54_433 ();
 sg13g2_decap_4 FILLER_54_462 ();
 sg13g2_fill_2 FILLER_54_466 ();
 sg13g2_fill_1 FILLER_54_481 ();
 sg13g2_fill_2 FILLER_54_493 ();
 sg13g2_fill_2 FILLER_54_503 ();
 sg13g2_fill_1 FILLER_54_505 ();
 sg13g2_fill_2 FILLER_54_519 ();
 sg13g2_fill_1 FILLER_54_521 ();
 sg13g2_decap_4 FILLER_54_530 ();
 sg13g2_fill_2 FILLER_54_534 ();
 sg13g2_fill_2 FILLER_54_593 ();
 sg13g2_fill_1 FILLER_54_617 ();
 sg13g2_fill_1 FILLER_54_623 ();
 sg13g2_fill_1 FILLER_54_632 ();
 sg13g2_fill_1 FILLER_54_641 ();
 sg13g2_fill_1 FILLER_54_730 ();
 sg13g2_decap_4 FILLER_54_754 ();
 sg13g2_fill_1 FILLER_54_772 ();
 sg13g2_fill_2 FILLER_54_777 ();
 sg13g2_fill_1 FILLER_54_779 ();
 sg13g2_fill_2 FILLER_54_790 ();
 sg13g2_fill_1 FILLER_54_792 ();
 sg13g2_decap_4 FILLER_54_801 ();
 sg13g2_fill_2 FILLER_54_812 ();
 sg13g2_fill_1 FILLER_54_833 ();
 sg13g2_fill_2 FILLER_54_843 ();
 sg13g2_fill_1 FILLER_54_845 ();
 sg13g2_fill_2 FILLER_54_872 ();
 sg13g2_fill_1 FILLER_54_874 ();
 sg13g2_decap_4 FILLER_54_886 ();
 sg13g2_fill_2 FILLER_54_901 ();
 sg13g2_fill_2 FILLER_54_912 ();
 sg13g2_decap_4 FILLER_54_922 ();
 sg13g2_fill_2 FILLER_54_926 ();
 sg13g2_fill_1 FILLER_54_959 ();
 sg13g2_fill_2 FILLER_54_984 ();
 sg13g2_fill_1 FILLER_54_1000 ();
 sg13g2_decap_8 FILLER_54_1053 ();
 sg13g2_decap_8 FILLER_54_1060 ();
 sg13g2_decap_8 FILLER_54_1067 ();
 sg13g2_decap_8 FILLER_54_1074 ();
 sg13g2_decap_8 FILLER_54_1081 ();
 sg13g2_decap_8 FILLER_54_1088 ();
 sg13g2_decap_8 FILLER_54_1095 ();
 sg13g2_decap_8 FILLER_54_1102 ();
 sg13g2_decap_8 FILLER_54_1109 ();
 sg13g2_decap_8 FILLER_54_1116 ();
 sg13g2_decap_8 FILLER_54_1123 ();
 sg13g2_decap_8 FILLER_54_1130 ();
 sg13g2_decap_8 FILLER_54_1137 ();
 sg13g2_decap_8 FILLER_54_1144 ();
 sg13g2_decap_8 FILLER_54_1151 ();
 sg13g2_decap_8 FILLER_54_1158 ();
 sg13g2_decap_8 FILLER_54_1165 ();
 sg13g2_decap_8 FILLER_54_1172 ();
 sg13g2_decap_8 FILLER_54_1179 ();
 sg13g2_decap_8 FILLER_54_1186 ();
 sg13g2_decap_8 FILLER_54_1193 ();
 sg13g2_decap_8 FILLER_54_1200 ();
 sg13g2_decap_8 FILLER_54_1207 ();
 sg13g2_decap_8 FILLER_54_1214 ();
 sg13g2_decap_8 FILLER_54_1221 ();
 sg13g2_decap_8 FILLER_54_1228 ();
 sg13g2_decap_8 FILLER_54_1235 ();
 sg13g2_decap_8 FILLER_54_1242 ();
 sg13g2_decap_8 FILLER_54_1249 ();
 sg13g2_decap_8 FILLER_54_1256 ();
 sg13g2_decap_8 FILLER_54_1263 ();
 sg13g2_decap_8 FILLER_54_1270 ();
 sg13g2_decap_8 FILLER_54_1277 ();
 sg13g2_decap_8 FILLER_54_1284 ();
 sg13g2_decap_8 FILLER_54_1291 ();
 sg13g2_decap_8 FILLER_54_1298 ();
 sg13g2_decap_8 FILLER_54_1305 ();
 sg13g2_fill_2 FILLER_54_1312 ();
 sg13g2_fill_1 FILLER_54_1314 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_4 FILLER_55_91 ();
 sg13g2_fill_2 FILLER_55_121 ();
 sg13g2_fill_2 FILLER_55_167 ();
 sg13g2_fill_1 FILLER_55_207 ();
 sg13g2_decap_4 FILLER_55_221 ();
 sg13g2_decap_4 FILLER_55_234 ();
 sg13g2_fill_2 FILLER_55_269 ();
 sg13g2_fill_2 FILLER_55_276 ();
 sg13g2_decap_4 FILLER_55_342 ();
 sg13g2_fill_2 FILLER_55_346 ();
 sg13g2_decap_8 FILLER_55_356 ();
 sg13g2_fill_2 FILLER_55_363 ();
 sg13g2_fill_1 FILLER_55_388 ();
 sg13g2_decap_8 FILLER_55_412 ();
 sg13g2_fill_2 FILLER_55_419 ();
 sg13g2_fill_1 FILLER_55_455 ();
 sg13g2_decap_4 FILLER_55_461 ();
 sg13g2_fill_1 FILLER_55_465 ();
 sg13g2_decap_8 FILLER_55_487 ();
 sg13g2_decap_8 FILLER_55_494 ();
 sg13g2_decap_4 FILLER_55_501 ();
 sg13g2_fill_2 FILLER_55_505 ();
 sg13g2_decap_4 FILLER_55_538 ();
 sg13g2_fill_1 FILLER_55_542 ();
 sg13g2_decap_4 FILLER_55_553 ();
 sg13g2_fill_1 FILLER_55_584 ();
 sg13g2_decap_4 FILLER_55_625 ();
 sg13g2_fill_2 FILLER_55_629 ();
 sg13g2_fill_2 FILLER_55_637 ();
 sg13g2_fill_1 FILLER_55_647 ();
 sg13g2_decap_8 FILLER_55_654 ();
 sg13g2_fill_2 FILLER_55_661 ();
 sg13g2_fill_1 FILLER_55_663 ();
 sg13g2_decap_4 FILLER_55_687 ();
 sg13g2_fill_1 FILLER_55_691 ();
 sg13g2_fill_2 FILLER_55_733 ();
 sg13g2_fill_2 FILLER_55_757 ();
 sg13g2_fill_1 FILLER_55_765 ();
 sg13g2_fill_1 FILLER_55_772 ();
 sg13g2_fill_2 FILLER_55_787 ();
 sg13g2_fill_1 FILLER_55_789 ();
 sg13g2_decap_8 FILLER_55_800 ();
 sg13g2_fill_2 FILLER_55_807 ();
 sg13g2_fill_1 FILLER_55_809 ();
 sg13g2_decap_4 FILLER_55_814 ();
 sg13g2_fill_1 FILLER_55_818 ();
 sg13g2_fill_2 FILLER_55_836 ();
 sg13g2_fill_2 FILLER_55_843 ();
 sg13g2_decap_8 FILLER_55_869 ();
 sg13g2_fill_1 FILLER_55_876 ();
 sg13g2_fill_2 FILLER_55_889 ();
 sg13g2_decap_4 FILLER_55_928 ();
 sg13g2_fill_2 FILLER_55_932 ();
 sg13g2_decap_4 FILLER_55_938 ();
 sg13g2_fill_1 FILLER_55_942 ();
 sg13g2_fill_2 FILLER_55_948 ();
 sg13g2_fill_1 FILLER_55_950 ();
 sg13g2_decap_4 FILLER_55_955 ();
 sg13g2_fill_1 FILLER_55_959 ();
 sg13g2_fill_1 FILLER_55_1020 ();
 sg13g2_fill_2 FILLER_55_1035 ();
 sg13g2_decap_8 FILLER_55_1041 ();
 sg13g2_decap_8 FILLER_55_1048 ();
 sg13g2_decap_8 FILLER_55_1055 ();
 sg13g2_decap_8 FILLER_55_1062 ();
 sg13g2_decap_8 FILLER_55_1069 ();
 sg13g2_decap_8 FILLER_55_1076 ();
 sg13g2_decap_8 FILLER_55_1083 ();
 sg13g2_decap_8 FILLER_55_1090 ();
 sg13g2_decap_8 FILLER_55_1097 ();
 sg13g2_decap_8 FILLER_55_1104 ();
 sg13g2_decap_8 FILLER_55_1111 ();
 sg13g2_decap_8 FILLER_55_1118 ();
 sg13g2_decap_8 FILLER_55_1125 ();
 sg13g2_decap_8 FILLER_55_1132 ();
 sg13g2_decap_8 FILLER_55_1139 ();
 sg13g2_decap_8 FILLER_55_1146 ();
 sg13g2_decap_8 FILLER_55_1153 ();
 sg13g2_decap_8 FILLER_55_1160 ();
 sg13g2_decap_8 FILLER_55_1167 ();
 sg13g2_decap_8 FILLER_55_1174 ();
 sg13g2_decap_8 FILLER_55_1181 ();
 sg13g2_decap_8 FILLER_55_1188 ();
 sg13g2_decap_8 FILLER_55_1195 ();
 sg13g2_decap_8 FILLER_55_1202 ();
 sg13g2_decap_8 FILLER_55_1209 ();
 sg13g2_decap_8 FILLER_55_1216 ();
 sg13g2_decap_8 FILLER_55_1223 ();
 sg13g2_decap_8 FILLER_55_1230 ();
 sg13g2_decap_8 FILLER_55_1237 ();
 sg13g2_decap_8 FILLER_55_1244 ();
 sg13g2_decap_8 FILLER_55_1251 ();
 sg13g2_decap_8 FILLER_55_1258 ();
 sg13g2_decap_8 FILLER_55_1265 ();
 sg13g2_decap_8 FILLER_55_1272 ();
 sg13g2_decap_8 FILLER_55_1279 ();
 sg13g2_decap_8 FILLER_55_1286 ();
 sg13g2_decap_8 FILLER_55_1293 ();
 sg13g2_decap_8 FILLER_55_1300 ();
 sg13g2_decap_8 FILLER_55_1307 ();
 sg13g2_fill_1 FILLER_55_1314 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_fill_1 FILLER_56_105 ();
 sg13g2_fill_2 FILLER_56_119 ();
 sg13g2_fill_1 FILLER_56_121 ();
 sg13g2_decap_8 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_163 ();
 sg13g2_fill_2 FILLER_56_216 ();
 sg13g2_fill_1 FILLER_56_218 ();
 sg13g2_decap_4 FILLER_56_268 ();
 sg13g2_fill_2 FILLER_56_282 ();
 sg13g2_fill_1 FILLER_56_297 ();
 sg13g2_fill_2 FILLER_56_413 ();
 sg13g2_fill_1 FILLER_56_434 ();
 sg13g2_fill_1 FILLER_56_440 ();
 sg13g2_fill_1 FILLER_56_464 ();
 sg13g2_decap_4 FILLER_56_483 ();
 sg13g2_fill_1 FILLER_56_497 ();
 sg13g2_fill_2 FILLER_56_506 ();
 sg13g2_fill_1 FILLER_56_508 ();
 sg13g2_decap_4 FILLER_56_535 ();
 sg13g2_fill_2 FILLER_56_539 ();
 sg13g2_decap_4 FILLER_56_546 ();
 sg13g2_fill_1 FILLER_56_580 ();
 sg13g2_decap_4 FILLER_56_603 ();
 sg13g2_decap_4 FILLER_56_629 ();
 sg13g2_fill_1 FILLER_56_639 ();
 sg13g2_decap_4 FILLER_56_707 ();
 sg13g2_fill_1 FILLER_56_711 ();
 sg13g2_fill_2 FILLER_56_725 ();
 sg13g2_fill_1 FILLER_56_727 ();
 sg13g2_fill_1 FILLER_56_738 ();
 sg13g2_fill_2 FILLER_56_744 ();
 sg13g2_fill_1 FILLER_56_746 ();
 sg13g2_decap_4 FILLER_56_752 ();
 sg13g2_fill_2 FILLER_56_756 ();
 sg13g2_fill_1 FILLER_56_769 ();
 sg13g2_fill_1 FILLER_56_776 ();
 sg13g2_fill_1 FILLER_56_802 ();
 sg13g2_fill_2 FILLER_56_824 ();
 sg13g2_fill_1 FILLER_56_826 ();
 sg13g2_fill_1 FILLER_56_875 ();
 sg13g2_decap_4 FILLER_56_890 ();
 sg13g2_fill_1 FILLER_56_894 ();
 sg13g2_fill_2 FILLER_56_913 ();
 sg13g2_fill_1 FILLER_56_915 ();
 sg13g2_fill_2 FILLER_56_921 ();
 sg13g2_fill_1 FILLER_56_923 ();
 sg13g2_fill_2 FILLER_56_968 ();
 sg13g2_fill_1 FILLER_56_970 ();
 sg13g2_fill_1 FILLER_56_989 ();
 sg13g2_fill_2 FILLER_56_998 ();
 sg13g2_fill_1 FILLER_56_1000 ();
 sg13g2_decap_8 FILLER_56_1005 ();
 sg13g2_decap_8 FILLER_56_1012 ();
 sg13g2_decap_8 FILLER_56_1019 ();
 sg13g2_decap_8 FILLER_56_1026 ();
 sg13g2_decap_8 FILLER_56_1033 ();
 sg13g2_decap_8 FILLER_56_1040 ();
 sg13g2_decap_8 FILLER_56_1047 ();
 sg13g2_decap_8 FILLER_56_1054 ();
 sg13g2_decap_8 FILLER_56_1061 ();
 sg13g2_decap_8 FILLER_56_1068 ();
 sg13g2_decap_8 FILLER_56_1075 ();
 sg13g2_decap_8 FILLER_56_1082 ();
 sg13g2_decap_8 FILLER_56_1089 ();
 sg13g2_decap_8 FILLER_56_1096 ();
 sg13g2_decap_8 FILLER_56_1103 ();
 sg13g2_decap_8 FILLER_56_1110 ();
 sg13g2_decap_8 FILLER_56_1117 ();
 sg13g2_decap_8 FILLER_56_1124 ();
 sg13g2_decap_8 FILLER_56_1131 ();
 sg13g2_decap_8 FILLER_56_1138 ();
 sg13g2_decap_8 FILLER_56_1145 ();
 sg13g2_decap_8 FILLER_56_1152 ();
 sg13g2_decap_8 FILLER_56_1159 ();
 sg13g2_decap_8 FILLER_56_1166 ();
 sg13g2_decap_8 FILLER_56_1173 ();
 sg13g2_decap_8 FILLER_56_1180 ();
 sg13g2_decap_8 FILLER_56_1187 ();
 sg13g2_decap_8 FILLER_56_1194 ();
 sg13g2_decap_8 FILLER_56_1201 ();
 sg13g2_decap_8 FILLER_56_1208 ();
 sg13g2_decap_8 FILLER_56_1215 ();
 sg13g2_decap_8 FILLER_56_1222 ();
 sg13g2_decap_8 FILLER_56_1229 ();
 sg13g2_decap_8 FILLER_56_1236 ();
 sg13g2_decap_8 FILLER_56_1243 ();
 sg13g2_decap_8 FILLER_56_1250 ();
 sg13g2_decap_8 FILLER_56_1257 ();
 sg13g2_decap_8 FILLER_56_1264 ();
 sg13g2_decap_8 FILLER_56_1271 ();
 sg13g2_decap_8 FILLER_56_1278 ();
 sg13g2_decap_8 FILLER_56_1285 ();
 sg13g2_decap_8 FILLER_56_1292 ();
 sg13g2_decap_8 FILLER_56_1299 ();
 sg13g2_decap_8 FILLER_56_1306 ();
 sg13g2_fill_2 FILLER_56_1313 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_4 FILLER_57_91 ();
 sg13g2_fill_2 FILLER_57_95 ();
 sg13g2_fill_1 FILLER_57_132 ();
 sg13g2_fill_2 FILLER_57_159 ();
 sg13g2_fill_2 FILLER_57_179 ();
 sg13g2_fill_1 FILLER_57_181 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_fill_1 FILLER_57_224 ();
 sg13g2_decap_4 FILLER_57_233 ();
 sg13g2_fill_1 FILLER_57_237 ();
 sg13g2_fill_2 FILLER_57_252 ();
 sg13g2_fill_1 FILLER_57_254 ();
 sg13g2_fill_1 FILLER_57_259 ();
 sg13g2_fill_2 FILLER_57_264 ();
 sg13g2_fill_1 FILLER_57_324 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_fill_2 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_348 ();
 sg13g2_fill_2 FILLER_57_367 ();
 sg13g2_decap_8 FILLER_57_381 ();
 sg13g2_fill_1 FILLER_57_388 ();
 sg13g2_decap_4 FILLER_57_393 ();
 sg13g2_fill_1 FILLER_57_397 ();
 sg13g2_decap_8 FILLER_57_403 ();
 sg13g2_decap_4 FILLER_57_410 ();
 sg13g2_fill_1 FILLER_57_414 ();
 sg13g2_decap_8 FILLER_57_419 ();
 sg13g2_fill_2 FILLER_57_426 ();
 sg13g2_fill_1 FILLER_57_436 ();
 sg13g2_fill_1 FILLER_57_442 ();
 sg13g2_decap_4 FILLER_57_447 ();
 sg13g2_fill_1 FILLER_57_451 ();
 sg13g2_fill_1 FILLER_57_509 ();
 sg13g2_decap_8 FILLER_57_536 ();
 sg13g2_fill_2 FILLER_57_557 ();
 sg13g2_fill_2 FILLER_57_564 ();
 sg13g2_decap_4 FILLER_57_612 ();
 sg13g2_decap_8 FILLER_57_620 ();
 sg13g2_fill_2 FILLER_57_627 ();
 sg13g2_decap_4 FILLER_57_634 ();
 sg13g2_fill_2 FILLER_57_638 ();
 sg13g2_decap_8 FILLER_57_651 ();
 sg13g2_fill_2 FILLER_57_658 ();
 sg13g2_decap_4 FILLER_57_683 ();
 sg13g2_decap_8 FILLER_57_705 ();
 sg13g2_decap_4 FILLER_57_725 ();
 sg13g2_fill_1 FILLER_57_729 ();
 sg13g2_fill_2 FILLER_57_740 ();
 sg13g2_fill_1 FILLER_57_742 ();
 sg13g2_decap_8 FILLER_57_747 ();
 sg13g2_fill_1 FILLER_57_754 ();
 sg13g2_fill_2 FILLER_57_776 ();
 sg13g2_fill_1 FILLER_57_778 ();
 sg13g2_fill_1 FILLER_57_790 ();
 sg13g2_decap_8 FILLER_57_800 ();
 sg13g2_fill_2 FILLER_57_807 ();
 sg13g2_decap_8 FILLER_57_814 ();
 sg13g2_fill_2 FILLER_57_821 ();
 sg13g2_decap_4 FILLER_57_836 ();
 sg13g2_fill_2 FILLER_57_845 ();
 sg13g2_fill_2 FILLER_57_857 ();
 sg13g2_decap_8 FILLER_57_863 ();
 sg13g2_decap_4 FILLER_57_870 ();
 sg13g2_fill_2 FILLER_57_874 ();
 sg13g2_fill_1 FILLER_57_893 ();
 sg13g2_decap_8 FILLER_57_907 ();
 sg13g2_decap_4 FILLER_57_914 ();
 sg13g2_fill_2 FILLER_57_918 ();
 sg13g2_fill_2 FILLER_57_929 ();
 sg13g2_fill_1 FILLER_57_931 ();
 sg13g2_fill_2 FILLER_57_976 ();
 sg13g2_decap_8 FILLER_57_1004 ();
 sg13g2_decap_8 FILLER_57_1011 ();
 sg13g2_decap_8 FILLER_57_1018 ();
 sg13g2_decap_8 FILLER_57_1025 ();
 sg13g2_decap_8 FILLER_57_1032 ();
 sg13g2_decap_8 FILLER_57_1039 ();
 sg13g2_decap_8 FILLER_57_1046 ();
 sg13g2_decap_8 FILLER_57_1053 ();
 sg13g2_decap_8 FILLER_57_1060 ();
 sg13g2_decap_8 FILLER_57_1067 ();
 sg13g2_decap_8 FILLER_57_1074 ();
 sg13g2_decap_8 FILLER_57_1081 ();
 sg13g2_decap_8 FILLER_57_1088 ();
 sg13g2_decap_8 FILLER_57_1095 ();
 sg13g2_decap_8 FILLER_57_1102 ();
 sg13g2_decap_8 FILLER_57_1109 ();
 sg13g2_decap_8 FILLER_57_1116 ();
 sg13g2_decap_8 FILLER_57_1123 ();
 sg13g2_decap_8 FILLER_57_1130 ();
 sg13g2_decap_8 FILLER_57_1137 ();
 sg13g2_decap_8 FILLER_57_1144 ();
 sg13g2_decap_8 FILLER_57_1151 ();
 sg13g2_decap_8 FILLER_57_1158 ();
 sg13g2_decap_8 FILLER_57_1165 ();
 sg13g2_decap_8 FILLER_57_1172 ();
 sg13g2_decap_8 FILLER_57_1179 ();
 sg13g2_decap_8 FILLER_57_1186 ();
 sg13g2_decap_8 FILLER_57_1193 ();
 sg13g2_decap_8 FILLER_57_1200 ();
 sg13g2_decap_8 FILLER_57_1207 ();
 sg13g2_decap_8 FILLER_57_1214 ();
 sg13g2_decap_8 FILLER_57_1221 ();
 sg13g2_decap_8 FILLER_57_1228 ();
 sg13g2_decap_8 FILLER_57_1235 ();
 sg13g2_decap_8 FILLER_57_1242 ();
 sg13g2_decap_8 FILLER_57_1249 ();
 sg13g2_decap_8 FILLER_57_1256 ();
 sg13g2_decap_8 FILLER_57_1263 ();
 sg13g2_decap_8 FILLER_57_1270 ();
 sg13g2_decap_8 FILLER_57_1277 ();
 sg13g2_decap_8 FILLER_57_1284 ();
 sg13g2_decap_8 FILLER_57_1291 ();
 sg13g2_decap_8 FILLER_57_1298 ();
 sg13g2_decap_8 FILLER_57_1305 ();
 sg13g2_fill_2 FILLER_57_1312 ();
 sg13g2_fill_1 FILLER_57_1314 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_91 ();
 sg13g2_fill_1 FILLER_58_128 ();
 sg13g2_fill_2 FILLER_58_155 ();
 sg13g2_fill_1 FILLER_58_157 ();
 sg13g2_decap_8 FILLER_58_162 ();
 sg13g2_fill_2 FILLER_58_169 ();
 sg13g2_decap_8 FILLER_58_176 ();
 sg13g2_fill_2 FILLER_58_183 ();
 sg13g2_fill_1 FILLER_58_185 ();
 sg13g2_fill_2 FILLER_58_240 ();
 sg13g2_fill_2 FILLER_58_282 ();
 sg13g2_decap_4 FILLER_58_297 ();
 sg13g2_fill_2 FILLER_58_301 ();
 sg13g2_fill_1 FILLER_58_307 ();
 sg13g2_fill_2 FILLER_58_312 ();
 sg13g2_fill_1 FILLER_58_342 ();
 sg13g2_fill_2 FILLER_58_347 ();
 sg13g2_fill_2 FILLER_58_359 ();
 sg13g2_fill_1 FILLER_58_361 ();
 sg13g2_decap_4 FILLER_58_371 ();
 sg13g2_fill_2 FILLER_58_375 ();
 sg13g2_decap_4 FILLER_58_390 ();
 sg13g2_fill_1 FILLER_58_394 ();
 sg13g2_fill_2 FILLER_58_422 ();
 sg13g2_decap_4 FILLER_58_459 ();
 sg13g2_decap_8 FILLER_58_467 ();
 sg13g2_fill_2 FILLER_58_474 ();
 sg13g2_fill_1 FILLER_58_494 ();
 sg13g2_decap_4 FILLER_58_500 ();
 sg13g2_fill_1 FILLER_58_504 ();
 sg13g2_decap_4 FILLER_58_512 ();
 sg13g2_decap_8 FILLER_58_528 ();
 sg13g2_fill_2 FILLER_58_535 ();
 sg13g2_fill_1 FILLER_58_537 ();
 sg13g2_fill_2 FILLER_58_543 ();
 sg13g2_fill_2 FILLER_58_557 ();
 sg13g2_fill_1 FILLER_58_559 ();
 sg13g2_decap_4 FILLER_58_595 ();
 sg13g2_fill_1 FILLER_58_599 ();
 sg13g2_fill_1 FILLER_58_621 ();
 sg13g2_fill_2 FILLER_58_643 ();
 sg13g2_fill_1 FILLER_58_681 ();
 sg13g2_fill_2 FILLER_58_730 ();
 sg13g2_fill_1 FILLER_58_732 ();
 sg13g2_fill_1 FILLER_58_769 ();
 sg13g2_fill_2 FILLER_58_791 ();
 sg13g2_fill_1 FILLER_58_805 ();
 sg13g2_decap_4 FILLER_58_825 ();
 sg13g2_fill_2 FILLER_58_829 ();
 sg13g2_fill_2 FILLER_58_836 ();
 sg13g2_decap_4 FILLER_58_843 ();
 sg13g2_fill_1 FILLER_58_847 ();
 sg13g2_fill_2 FILLER_58_907 ();
 sg13g2_fill_1 FILLER_58_909 ();
 sg13g2_fill_2 FILLER_58_936 ();
 sg13g2_fill_2 FILLER_58_973 ();
 sg13g2_fill_1 FILLER_58_975 ();
 sg13g2_decap_8 FILLER_58_1002 ();
 sg13g2_decap_8 FILLER_58_1009 ();
 sg13g2_decap_8 FILLER_58_1016 ();
 sg13g2_decap_8 FILLER_58_1023 ();
 sg13g2_decap_8 FILLER_58_1030 ();
 sg13g2_decap_8 FILLER_58_1037 ();
 sg13g2_decap_8 FILLER_58_1044 ();
 sg13g2_decap_8 FILLER_58_1051 ();
 sg13g2_decap_8 FILLER_58_1058 ();
 sg13g2_decap_8 FILLER_58_1065 ();
 sg13g2_decap_8 FILLER_58_1072 ();
 sg13g2_decap_8 FILLER_58_1079 ();
 sg13g2_decap_8 FILLER_58_1086 ();
 sg13g2_decap_8 FILLER_58_1093 ();
 sg13g2_decap_8 FILLER_58_1100 ();
 sg13g2_decap_8 FILLER_58_1107 ();
 sg13g2_decap_8 FILLER_58_1114 ();
 sg13g2_decap_8 FILLER_58_1121 ();
 sg13g2_decap_8 FILLER_58_1128 ();
 sg13g2_decap_8 FILLER_58_1135 ();
 sg13g2_decap_8 FILLER_58_1142 ();
 sg13g2_decap_8 FILLER_58_1149 ();
 sg13g2_decap_8 FILLER_58_1156 ();
 sg13g2_decap_8 FILLER_58_1163 ();
 sg13g2_decap_8 FILLER_58_1170 ();
 sg13g2_decap_8 FILLER_58_1177 ();
 sg13g2_decap_8 FILLER_58_1184 ();
 sg13g2_decap_8 FILLER_58_1191 ();
 sg13g2_decap_8 FILLER_58_1198 ();
 sg13g2_decap_8 FILLER_58_1205 ();
 sg13g2_decap_8 FILLER_58_1212 ();
 sg13g2_decap_8 FILLER_58_1219 ();
 sg13g2_decap_8 FILLER_58_1226 ();
 sg13g2_decap_8 FILLER_58_1233 ();
 sg13g2_decap_8 FILLER_58_1240 ();
 sg13g2_decap_8 FILLER_58_1247 ();
 sg13g2_decap_8 FILLER_58_1254 ();
 sg13g2_decap_8 FILLER_58_1261 ();
 sg13g2_decap_8 FILLER_58_1268 ();
 sg13g2_decap_8 FILLER_58_1275 ();
 sg13g2_decap_8 FILLER_58_1282 ();
 sg13g2_decap_8 FILLER_58_1289 ();
 sg13g2_decap_8 FILLER_58_1296 ();
 sg13g2_decap_8 FILLER_58_1303 ();
 sg13g2_decap_4 FILLER_58_1310 ();
 sg13g2_fill_1 FILLER_58_1314 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_fill_1 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_54 ();
 sg13g2_decap_8 FILLER_59_61 ();
 sg13g2_decap_8 FILLER_59_68 ();
 sg13g2_decap_8 FILLER_59_75 ();
 sg13g2_decap_8 FILLER_59_82 ();
 sg13g2_decap_8 FILLER_59_89 ();
 sg13g2_fill_1 FILLER_59_124 ();
 sg13g2_fill_2 FILLER_59_130 ();
 sg13g2_decap_8 FILLER_59_142 ();
 sg13g2_fill_2 FILLER_59_149 ();
 sg13g2_fill_1 FILLER_59_172 ();
 sg13g2_fill_2 FILLER_59_181 ();
 sg13g2_fill_1 FILLER_59_196 ();
 sg13g2_fill_2 FILLER_59_202 ();
 sg13g2_fill_1 FILLER_59_204 ();
 sg13g2_fill_2 FILLER_59_218 ();
 sg13g2_decap_4 FILLER_59_239 ();
 sg13g2_fill_1 FILLER_59_255 ();
 sg13g2_decap_4 FILLER_59_264 ();
 sg13g2_fill_1 FILLER_59_278 ();
 sg13g2_decap_8 FILLER_59_305 ();
 sg13g2_decap_4 FILLER_59_312 ();
 sg13g2_fill_2 FILLER_59_316 ();
 sg13g2_fill_2 FILLER_59_323 ();
 sg13g2_fill_1 FILLER_59_325 ();
 sg13g2_fill_1 FILLER_59_361 ();
 sg13g2_decap_4 FILLER_59_428 ();
 sg13g2_fill_2 FILLER_59_444 ();
 sg13g2_fill_2 FILLER_59_451 ();
 sg13g2_fill_1 FILLER_59_453 ();
 sg13g2_fill_2 FILLER_59_463 ();
 sg13g2_fill_1 FILLER_59_465 ();
 sg13g2_fill_2 FILLER_59_479 ();
 sg13g2_fill_1 FILLER_59_481 ();
 sg13g2_decap_4 FILLER_59_502 ();
 sg13g2_fill_2 FILLER_59_540 ();
 sg13g2_decap_8 FILLER_59_570 ();
 sg13g2_fill_2 FILLER_59_577 ();
 sg13g2_fill_1 FILLER_59_579 ();
 sg13g2_fill_2 FILLER_59_584 ();
 sg13g2_fill_2 FILLER_59_591 ();
 sg13g2_fill_1 FILLER_59_593 ();
 sg13g2_fill_2 FILLER_59_604 ();
 sg13g2_decap_8 FILLER_59_616 ();
 sg13g2_decap_4 FILLER_59_623 ();
 sg13g2_decap_8 FILLER_59_631 ();
 sg13g2_fill_2 FILLER_59_659 ();
 sg13g2_decap_8 FILLER_59_683 ();
 sg13g2_fill_2 FILLER_59_690 ();
 sg13g2_fill_2 FILLER_59_705 ();
 sg13g2_decap_8 FILLER_59_776 ();
 sg13g2_fill_2 FILLER_59_783 ();
 sg13g2_fill_1 FILLER_59_785 ();
 sg13g2_fill_2 FILLER_59_805 ();
 sg13g2_decap_4 FILLER_59_817 ();
 sg13g2_fill_2 FILLER_59_827 ();
 sg13g2_fill_2 FILLER_59_851 ();
 sg13g2_decap_4 FILLER_59_861 ();
 sg13g2_fill_1 FILLER_59_865 ();
 sg13g2_fill_2 FILLER_59_874 ();
 sg13g2_fill_1 FILLER_59_876 ();
 sg13g2_fill_2 FILLER_59_895 ();
 sg13g2_fill_1 FILLER_59_897 ();
 sg13g2_fill_2 FILLER_59_903 ();
 sg13g2_fill_1 FILLER_59_905 ();
 sg13g2_decap_8 FILLER_59_911 ();
 sg13g2_decap_8 FILLER_59_918 ();
 sg13g2_fill_2 FILLER_59_925 ();
 sg13g2_decap_4 FILLER_59_947 ();
 sg13g2_fill_2 FILLER_59_951 ();
 sg13g2_fill_2 FILLER_59_966 ();
 sg13g2_fill_1 FILLER_59_987 ();
 sg13g2_decap_8 FILLER_59_1006 ();
 sg13g2_decap_8 FILLER_59_1013 ();
 sg13g2_decap_8 FILLER_59_1020 ();
 sg13g2_decap_8 FILLER_59_1027 ();
 sg13g2_decap_8 FILLER_59_1034 ();
 sg13g2_decap_8 FILLER_59_1041 ();
 sg13g2_decap_8 FILLER_59_1048 ();
 sg13g2_decap_8 FILLER_59_1055 ();
 sg13g2_decap_8 FILLER_59_1062 ();
 sg13g2_decap_8 FILLER_59_1069 ();
 sg13g2_decap_8 FILLER_59_1076 ();
 sg13g2_decap_8 FILLER_59_1083 ();
 sg13g2_decap_8 FILLER_59_1090 ();
 sg13g2_decap_8 FILLER_59_1097 ();
 sg13g2_decap_8 FILLER_59_1104 ();
 sg13g2_decap_8 FILLER_59_1111 ();
 sg13g2_decap_8 FILLER_59_1118 ();
 sg13g2_decap_8 FILLER_59_1125 ();
 sg13g2_decap_8 FILLER_59_1132 ();
 sg13g2_decap_8 FILLER_59_1139 ();
 sg13g2_decap_8 FILLER_59_1146 ();
 sg13g2_decap_8 FILLER_59_1153 ();
 sg13g2_decap_8 FILLER_59_1160 ();
 sg13g2_decap_8 FILLER_59_1167 ();
 sg13g2_decap_8 FILLER_59_1174 ();
 sg13g2_decap_8 FILLER_59_1181 ();
 sg13g2_decap_8 FILLER_59_1188 ();
 sg13g2_decap_8 FILLER_59_1195 ();
 sg13g2_decap_8 FILLER_59_1202 ();
 sg13g2_decap_8 FILLER_59_1209 ();
 sg13g2_decap_8 FILLER_59_1216 ();
 sg13g2_decap_8 FILLER_59_1223 ();
 sg13g2_decap_8 FILLER_59_1230 ();
 sg13g2_decap_8 FILLER_59_1237 ();
 sg13g2_decap_8 FILLER_59_1244 ();
 sg13g2_decap_8 FILLER_59_1251 ();
 sg13g2_decap_8 FILLER_59_1258 ();
 sg13g2_decap_8 FILLER_59_1265 ();
 sg13g2_decap_8 FILLER_59_1272 ();
 sg13g2_decap_8 FILLER_59_1279 ();
 sg13g2_decap_8 FILLER_59_1286 ();
 sg13g2_decap_8 FILLER_59_1293 ();
 sg13g2_decap_8 FILLER_59_1300 ();
 sg13g2_decap_8 FILLER_59_1307 ();
 sg13g2_fill_1 FILLER_59_1314 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_14 ();
 sg13g2_fill_2 FILLER_60_52 ();
 sg13g2_decap_8 FILLER_60_80 ();
 sg13g2_decap_4 FILLER_60_87 ();
 sg13g2_fill_1 FILLER_60_91 ();
 sg13g2_fill_2 FILLER_60_118 ();
 sg13g2_fill_2 FILLER_60_125 ();
 sg13g2_fill_2 FILLER_60_144 ();
 sg13g2_fill_1 FILLER_60_146 ();
 sg13g2_fill_1 FILLER_60_168 ();
 sg13g2_fill_1 FILLER_60_195 ();
 sg13g2_fill_2 FILLER_60_210 ();
 sg13g2_fill_1 FILLER_60_212 ();
 sg13g2_fill_2 FILLER_60_241 ();
 sg13g2_fill_1 FILLER_60_251 ();
 sg13g2_fill_1 FILLER_60_266 ();
 sg13g2_fill_2 FILLER_60_272 ();
 sg13g2_fill_1 FILLER_60_274 ();
 sg13g2_fill_2 FILLER_60_279 ();
 sg13g2_fill_2 FILLER_60_285 ();
 sg13g2_fill_1 FILLER_60_287 ();
 sg13g2_fill_2 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_60_324 ();
 sg13g2_fill_1 FILLER_60_337 ();
 sg13g2_fill_2 FILLER_60_362 ();
 sg13g2_fill_1 FILLER_60_364 ();
 sg13g2_fill_1 FILLER_60_379 ();
 sg13g2_decap_4 FILLER_60_392 ();
 sg13g2_fill_2 FILLER_60_396 ();
 sg13g2_decap_8 FILLER_60_403 ();
 sg13g2_decap_4 FILLER_60_410 ();
 sg13g2_fill_2 FILLER_60_414 ();
 sg13g2_decap_4 FILLER_60_434 ();
 sg13g2_fill_2 FILLER_60_446 ();
 sg13g2_fill_2 FILLER_60_452 ();
 sg13g2_decap_4 FILLER_60_488 ();
 sg13g2_decap_8 FILLER_60_528 ();
 sg13g2_fill_2 FILLER_60_535 ();
 sg13g2_fill_2 FILLER_60_555 ();
 sg13g2_fill_2 FILLER_60_565 ();
 sg13g2_fill_1 FILLER_60_567 ();
 sg13g2_fill_2 FILLER_60_650 ();
 sg13g2_fill_1 FILLER_60_688 ();
 sg13g2_decap_4 FILLER_60_693 ();
 sg13g2_fill_1 FILLER_60_697 ();
 sg13g2_fill_2 FILLER_60_715 ();
 sg13g2_fill_1 FILLER_60_717 ();
 sg13g2_decap_8 FILLER_60_722 ();
 sg13g2_fill_2 FILLER_60_729 ();
 sg13g2_fill_1 FILLER_60_745 ();
 sg13g2_fill_1 FILLER_60_766 ();
 sg13g2_decap_4 FILLER_60_774 ();
 sg13g2_decap_4 FILLER_60_783 ();
 sg13g2_fill_1 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_793 ();
 sg13g2_decap_4 FILLER_60_800 ();
 sg13g2_decap_4 FILLER_60_824 ();
 sg13g2_fill_2 FILLER_60_828 ();
 sg13g2_decap_4 FILLER_60_842 ();
 sg13g2_decap_4 FILLER_60_857 ();
 sg13g2_fill_2 FILLER_60_884 ();
 sg13g2_fill_2 FILLER_60_894 ();
 sg13g2_fill_1 FILLER_60_896 ();
 sg13g2_fill_2 FILLER_60_937 ();
 sg13g2_decap_8 FILLER_60_1017 ();
 sg13g2_decap_8 FILLER_60_1024 ();
 sg13g2_decap_8 FILLER_60_1031 ();
 sg13g2_decap_8 FILLER_60_1038 ();
 sg13g2_decap_8 FILLER_60_1045 ();
 sg13g2_decap_8 FILLER_60_1052 ();
 sg13g2_decap_8 FILLER_60_1059 ();
 sg13g2_decap_8 FILLER_60_1066 ();
 sg13g2_decap_8 FILLER_60_1073 ();
 sg13g2_decap_8 FILLER_60_1080 ();
 sg13g2_decap_8 FILLER_60_1087 ();
 sg13g2_decap_8 FILLER_60_1094 ();
 sg13g2_decap_8 FILLER_60_1101 ();
 sg13g2_decap_8 FILLER_60_1108 ();
 sg13g2_decap_8 FILLER_60_1115 ();
 sg13g2_decap_8 FILLER_60_1122 ();
 sg13g2_decap_8 FILLER_60_1129 ();
 sg13g2_decap_8 FILLER_60_1136 ();
 sg13g2_decap_8 FILLER_60_1143 ();
 sg13g2_decap_8 FILLER_60_1150 ();
 sg13g2_decap_8 FILLER_60_1157 ();
 sg13g2_decap_8 FILLER_60_1164 ();
 sg13g2_decap_8 FILLER_60_1171 ();
 sg13g2_decap_8 FILLER_60_1178 ();
 sg13g2_decap_8 FILLER_60_1185 ();
 sg13g2_decap_8 FILLER_60_1192 ();
 sg13g2_decap_8 FILLER_60_1199 ();
 sg13g2_decap_8 FILLER_60_1206 ();
 sg13g2_decap_8 FILLER_60_1213 ();
 sg13g2_decap_8 FILLER_60_1220 ();
 sg13g2_decap_8 FILLER_60_1227 ();
 sg13g2_decap_8 FILLER_60_1234 ();
 sg13g2_decap_8 FILLER_60_1241 ();
 sg13g2_decap_8 FILLER_60_1248 ();
 sg13g2_decap_8 FILLER_60_1255 ();
 sg13g2_decap_8 FILLER_60_1262 ();
 sg13g2_decap_8 FILLER_60_1269 ();
 sg13g2_decap_8 FILLER_60_1276 ();
 sg13g2_decap_8 FILLER_60_1283 ();
 sg13g2_decap_8 FILLER_60_1290 ();
 sg13g2_decap_8 FILLER_60_1297 ();
 sg13g2_decap_8 FILLER_60_1304 ();
 sg13g2_decap_4 FILLER_60_1311 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_4 FILLER_61_21 ();
 sg13g2_fill_1 FILLER_61_25 ();
 sg13g2_fill_2 FILLER_61_43 ();
 sg13g2_decap_8 FILLER_61_75 ();
 sg13g2_decap_8 FILLER_61_82 ();
 sg13g2_decap_8 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_96 ();
 sg13g2_fill_2 FILLER_61_115 ();
 sg13g2_fill_1 FILLER_61_117 ();
 sg13g2_fill_2 FILLER_61_127 ();
 sg13g2_fill_2 FILLER_61_177 ();
 sg13g2_fill_1 FILLER_61_179 ();
 sg13g2_fill_2 FILLER_61_189 ();
 sg13g2_fill_1 FILLER_61_191 ();
 sg13g2_fill_2 FILLER_61_205 ();
 sg13g2_fill_1 FILLER_61_207 ();
 sg13g2_fill_2 FILLER_61_234 ();
 sg13g2_fill_1 FILLER_61_292 ();
 sg13g2_decap_4 FILLER_61_297 ();
 sg13g2_fill_1 FILLER_61_301 ();
 sg13g2_fill_2 FILLER_61_323 ();
 sg13g2_fill_1 FILLER_61_329 ();
 sg13g2_fill_1 FILLER_61_391 ();
 sg13g2_fill_1 FILLER_61_422 ();
 sg13g2_decap_4 FILLER_61_459 ();
 sg13g2_fill_2 FILLER_61_463 ();
 sg13g2_fill_1 FILLER_61_469 ();
 sg13g2_decap_8 FILLER_61_478 ();
 sg13g2_decap_4 FILLER_61_485 ();
 sg13g2_fill_1 FILLER_61_489 ();
 sg13g2_decap_4 FILLER_61_504 ();
 sg13g2_decap_8 FILLER_61_548 ();
 sg13g2_decap_8 FILLER_61_555 ();
 sg13g2_fill_2 FILLER_61_562 ();
 sg13g2_decap_8 FILLER_61_574 ();
 sg13g2_fill_2 FILLER_61_581 ();
 sg13g2_fill_1 FILLER_61_583 ();
 sg13g2_decap_8 FILLER_61_588 ();
 sg13g2_decap_8 FILLER_61_595 ();
 sg13g2_decap_8 FILLER_61_602 ();
 sg13g2_fill_1 FILLER_61_609 ();
 sg13g2_fill_2 FILLER_61_646 ();
 sg13g2_fill_2 FILLER_61_653 ();
 sg13g2_fill_1 FILLER_61_677 ();
 sg13g2_fill_2 FILLER_61_730 ();
 sg13g2_fill_1 FILLER_61_732 ();
 sg13g2_fill_2 FILLER_61_753 ();
 sg13g2_fill_2 FILLER_61_763 ();
 sg13g2_fill_1 FILLER_61_765 ();
 sg13g2_decap_4 FILLER_61_774 ();
 sg13g2_decap_4 FILLER_61_801 ();
 sg13g2_fill_1 FILLER_61_827 ();
 sg13g2_fill_2 FILLER_61_851 ();
 sg13g2_decap_8 FILLER_61_858 ();
 sg13g2_decap_4 FILLER_61_865 ();
 sg13g2_fill_1 FILLER_61_869 ();
 sg13g2_fill_2 FILLER_61_893 ();
 sg13g2_fill_1 FILLER_61_921 ();
 sg13g2_fill_1 FILLER_61_953 ();
 sg13g2_fill_2 FILLER_61_963 ();
 sg13g2_decap_8 FILLER_61_987 ();
 sg13g2_decap_8 FILLER_61_998 ();
 sg13g2_decap_8 FILLER_61_1005 ();
 sg13g2_decap_8 FILLER_61_1012 ();
 sg13g2_decap_8 FILLER_61_1019 ();
 sg13g2_decap_8 FILLER_61_1026 ();
 sg13g2_decap_8 FILLER_61_1033 ();
 sg13g2_decap_8 FILLER_61_1040 ();
 sg13g2_decap_8 FILLER_61_1047 ();
 sg13g2_decap_8 FILLER_61_1054 ();
 sg13g2_decap_8 FILLER_61_1061 ();
 sg13g2_decap_8 FILLER_61_1068 ();
 sg13g2_decap_8 FILLER_61_1075 ();
 sg13g2_decap_8 FILLER_61_1082 ();
 sg13g2_decap_8 FILLER_61_1089 ();
 sg13g2_decap_8 FILLER_61_1096 ();
 sg13g2_decap_8 FILLER_61_1103 ();
 sg13g2_decap_8 FILLER_61_1110 ();
 sg13g2_decap_8 FILLER_61_1117 ();
 sg13g2_decap_8 FILLER_61_1124 ();
 sg13g2_decap_8 FILLER_61_1131 ();
 sg13g2_decap_8 FILLER_61_1138 ();
 sg13g2_decap_8 FILLER_61_1145 ();
 sg13g2_decap_8 FILLER_61_1152 ();
 sg13g2_decap_8 FILLER_61_1159 ();
 sg13g2_decap_8 FILLER_61_1166 ();
 sg13g2_decap_8 FILLER_61_1173 ();
 sg13g2_decap_8 FILLER_61_1180 ();
 sg13g2_decap_8 FILLER_61_1187 ();
 sg13g2_decap_8 FILLER_61_1194 ();
 sg13g2_decap_8 FILLER_61_1201 ();
 sg13g2_decap_8 FILLER_61_1208 ();
 sg13g2_decap_8 FILLER_61_1215 ();
 sg13g2_decap_8 FILLER_61_1222 ();
 sg13g2_decap_8 FILLER_61_1229 ();
 sg13g2_decap_8 FILLER_61_1236 ();
 sg13g2_decap_8 FILLER_61_1243 ();
 sg13g2_decap_8 FILLER_61_1250 ();
 sg13g2_decap_8 FILLER_61_1257 ();
 sg13g2_decap_8 FILLER_61_1264 ();
 sg13g2_decap_8 FILLER_61_1271 ();
 sg13g2_decap_8 FILLER_61_1278 ();
 sg13g2_decap_8 FILLER_61_1285 ();
 sg13g2_decap_8 FILLER_61_1292 ();
 sg13g2_decap_8 FILLER_61_1299 ();
 sg13g2_decap_8 FILLER_61_1306 ();
 sg13g2_fill_2 FILLER_61_1313 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_fill_2 FILLER_62_21 ();
 sg13g2_fill_1 FILLER_62_23 ();
 sg13g2_decap_4 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_80 ();
 sg13g2_decap_8 FILLER_62_87 ();
 sg13g2_decap_4 FILLER_62_94 ();
 sg13g2_fill_2 FILLER_62_98 ();
 sg13g2_fill_2 FILLER_62_126 ();
 sg13g2_fill_1 FILLER_62_128 ();
 sg13g2_fill_1 FILLER_62_143 ();
 sg13g2_decap_8 FILLER_62_200 ();
 sg13g2_decap_4 FILLER_62_207 ();
 sg13g2_decap_4 FILLER_62_215 ();
 sg13g2_fill_2 FILLER_62_223 ();
 sg13g2_fill_1 FILLER_62_225 ();
 sg13g2_decap_4 FILLER_62_231 ();
 sg13g2_decap_4 FILLER_62_240 ();
 sg13g2_fill_2 FILLER_62_244 ();
 sg13g2_decap_4 FILLER_62_264 ();
 sg13g2_fill_1 FILLER_62_268 ();
 sg13g2_decap_4 FILLER_62_333 ();
 sg13g2_fill_1 FILLER_62_337 ();
 sg13g2_decap_8 FILLER_62_342 ();
 sg13g2_fill_2 FILLER_62_349 ();
 sg13g2_fill_1 FILLER_62_351 ();
 sg13g2_fill_2 FILLER_62_357 ();
 sg13g2_fill_1 FILLER_62_359 ();
 sg13g2_fill_2 FILLER_62_401 ();
 sg13g2_fill_1 FILLER_62_407 ();
 sg13g2_fill_2 FILLER_62_412 ();
 sg13g2_fill_1 FILLER_62_414 ();
 sg13g2_fill_2 FILLER_62_452 ();
 sg13g2_fill_1 FILLER_62_454 ();
 sg13g2_fill_2 FILLER_62_474 ();
 sg13g2_decap_4 FILLER_62_480 ();
 sg13g2_fill_2 FILLER_62_484 ();
 sg13g2_decap_8 FILLER_62_507 ();
 sg13g2_decap_8 FILLER_62_514 ();
 sg13g2_decap_8 FILLER_62_521 ();
 sg13g2_decap_8 FILLER_62_597 ();
 sg13g2_fill_2 FILLER_62_604 ();
 sg13g2_fill_1 FILLER_62_611 ();
 sg13g2_fill_2 FILLER_62_628 ();
 sg13g2_decap_8 FILLER_62_636 ();
 sg13g2_decap_8 FILLER_62_643 ();
 sg13g2_fill_2 FILLER_62_650 ();
 sg13g2_fill_1 FILLER_62_652 ();
 sg13g2_fill_2 FILLER_62_666 ();
 sg13g2_decap_8 FILLER_62_672 ();
 sg13g2_fill_1 FILLER_62_679 ();
 sg13g2_decap_8 FILLER_62_684 ();
 sg13g2_fill_2 FILLER_62_691 ();
 sg13g2_fill_1 FILLER_62_693 ();
 sg13g2_decap_4 FILLER_62_709 ();
 sg13g2_fill_2 FILLER_62_713 ();
 sg13g2_fill_2 FILLER_62_745 ();
 sg13g2_decap_8 FILLER_62_769 ();
 sg13g2_fill_2 FILLER_62_776 ();
 sg13g2_fill_1 FILLER_62_787 ();
 sg13g2_decap_8 FILLER_62_793 ();
 sg13g2_decap_4 FILLER_62_800 ();
 sg13g2_decap_8 FILLER_62_822 ();
 sg13g2_decap_4 FILLER_62_834 ();
 sg13g2_fill_1 FILLER_62_838 ();
 sg13g2_decap_4 FILLER_62_850 ();
 sg13g2_fill_2 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_901 ();
 sg13g2_fill_2 FILLER_62_919 ();
 sg13g2_fill_1 FILLER_62_921 ();
 sg13g2_fill_2 FILLER_62_992 ();
 sg13g2_decap_8 FILLER_62_998 ();
 sg13g2_decap_8 FILLER_62_1005 ();
 sg13g2_decap_8 FILLER_62_1012 ();
 sg13g2_decap_8 FILLER_62_1019 ();
 sg13g2_decap_8 FILLER_62_1026 ();
 sg13g2_decap_8 FILLER_62_1033 ();
 sg13g2_decap_8 FILLER_62_1040 ();
 sg13g2_decap_8 FILLER_62_1047 ();
 sg13g2_decap_8 FILLER_62_1054 ();
 sg13g2_decap_8 FILLER_62_1061 ();
 sg13g2_decap_8 FILLER_62_1068 ();
 sg13g2_decap_8 FILLER_62_1075 ();
 sg13g2_decap_8 FILLER_62_1082 ();
 sg13g2_decap_8 FILLER_62_1089 ();
 sg13g2_decap_8 FILLER_62_1096 ();
 sg13g2_decap_8 FILLER_62_1103 ();
 sg13g2_decap_8 FILLER_62_1110 ();
 sg13g2_decap_8 FILLER_62_1117 ();
 sg13g2_decap_8 FILLER_62_1124 ();
 sg13g2_decap_8 FILLER_62_1131 ();
 sg13g2_decap_8 FILLER_62_1138 ();
 sg13g2_decap_8 FILLER_62_1145 ();
 sg13g2_decap_8 FILLER_62_1152 ();
 sg13g2_decap_8 FILLER_62_1159 ();
 sg13g2_decap_8 FILLER_62_1166 ();
 sg13g2_decap_8 FILLER_62_1173 ();
 sg13g2_decap_8 FILLER_62_1180 ();
 sg13g2_decap_8 FILLER_62_1187 ();
 sg13g2_decap_8 FILLER_62_1194 ();
 sg13g2_decap_8 FILLER_62_1201 ();
 sg13g2_decap_8 FILLER_62_1208 ();
 sg13g2_decap_8 FILLER_62_1215 ();
 sg13g2_decap_8 FILLER_62_1222 ();
 sg13g2_decap_8 FILLER_62_1229 ();
 sg13g2_decap_8 FILLER_62_1236 ();
 sg13g2_decap_8 FILLER_62_1243 ();
 sg13g2_decap_8 FILLER_62_1250 ();
 sg13g2_decap_8 FILLER_62_1257 ();
 sg13g2_decap_8 FILLER_62_1264 ();
 sg13g2_decap_8 FILLER_62_1271 ();
 sg13g2_decap_8 FILLER_62_1278 ();
 sg13g2_decap_8 FILLER_62_1285 ();
 sg13g2_decap_8 FILLER_62_1292 ();
 sg13g2_decap_8 FILLER_62_1299 ();
 sg13g2_decap_8 FILLER_62_1306 ();
 sg13g2_fill_2 FILLER_62_1313 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_fill_2 FILLER_63_11 ();
 sg13g2_fill_2 FILLER_63_39 ();
 sg13g2_fill_1 FILLER_63_66 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_fill_1 FILLER_63_155 ();
 sg13g2_fill_1 FILLER_63_161 ();
 sg13g2_fill_2 FILLER_63_179 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_fill_2 FILLER_63_231 ();
 sg13g2_fill_1 FILLER_63_233 ();
 sg13g2_decap_8 FILLER_63_244 ();
 sg13g2_fill_2 FILLER_63_251 ();
 sg13g2_fill_2 FILLER_63_258 ();
 sg13g2_fill_2 FILLER_63_273 ();
 sg13g2_fill_2 FILLER_63_294 ();
 sg13g2_fill_2 FILLER_63_305 ();
 sg13g2_fill_2 FILLER_63_325 ();
 sg13g2_fill_2 FILLER_63_340 ();
 sg13g2_fill_1 FILLER_63_342 ();
 sg13g2_fill_2 FILLER_63_356 ();
 sg13g2_fill_2 FILLER_63_380 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_fill_1 FILLER_63_388 ();
 sg13g2_fill_2 FILLER_63_467 ();
 sg13g2_fill_2 FILLER_63_474 ();
 sg13g2_fill_1 FILLER_63_476 ();
 sg13g2_fill_1 FILLER_63_485 ();
 sg13g2_decap_8 FILLER_63_491 ();
 sg13g2_decap_8 FILLER_63_498 ();
 sg13g2_decap_4 FILLER_63_512 ();
 sg13g2_fill_2 FILLER_63_516 ();
 sg13g2_decap_8 FILLER_63_534 ();
 sg13g2_fill_1 FILLER_63_541 ();
 sg13g2_decap_4 FILLER_63_557 ();
 sg13g2_decap_8 FILLER_63_565 ();
 sg13g2_decap_4 FILLER_63_572 ();
 sg13g2_fill_2 FILLER_63_576 ();
 sg13g2_fill_1 FILLER_63_586 ();
 sg13g2_decap_4 FILLER_63_609 ();
 sg13g2_fill_1 FILLER_63_642 ();
 sg13g2_fill_1 FILLER_63_695 ();
 sg13g2_fill_2 FILLER_63_706 ();
 sg13g2_fill_1 FILLER_63_708 ();
 sg13g2_decap_8 FILLER_63_739 ();
 sg13g2_decap_8 FILLER_63_746 ();
 sg13g2_fill_1 FILLER_63_753 ();
 sg13g2_decap_8 FILLER_63_759 ();
 sg13g2_fill_2 FILLER_63_766 ();
 sg13g2_fill_1 FILLER_63_768 ();
 sg13g2_decap_4 FILLER_63_789 ();
 sg13g2_fill_2 FILLER_63_814 ();
 sg13g2_fill_2 FILLER_63_824 ();
 sg13g2_decap_4 FILLER_63_855 ();
 sg13g2_fill_1 FILLER_63_859 ();
 sg13g2_fill_2 FILLER_63_870 ();
 sg13g2_decap_4 FILLER_63_877 ();
 sg13g2_fill_2 FILLER_63_881 ();
 sg13g2_fill_1 FILLER_63_891 ();
 sg13g2_decap_4 FILLER_63_899 ();
 sg13g2_fill_2 FILLER_63_903 ();
 sg13g2_decap_4 FILLER_63_909 ();
 sg13g2_fill_2 FILLER_63_913 ();
 sg13g2_decap_4 FILLER_63_957 ();
 sg13g2_decap_8 FILLER_63_1009 ();
 sg13g2_decap_8 FILLER_63_1016 ();
 sg13g2_decap_8 FILLER_63_1023 ();
 sg13g2_decap_8 FILLER_63_1030 ();
 sg13g2_decap_8 FILLER_63_1037 ();
 sg13g2_decap_8 FILLER_63_1044 ();
 sg13g2_decap_8 FILLER_63_1051 ();
 sg13g2_decap_8 FILLER_63_1058 ();
 sg13g2_decap_8 FILLER_63_1065 ();
 sg13g2_decap_8 FILLER_63_1072 ();
 sg13g2_decap_8 FILLER_63_1079 ();
 sg13g2_decap_8 FILLER_63_1086 ();
 sg13g2_decap_8 FILLER_63_1093 ();
 sg13g2_decap_8 FILLER_63_1100 ();
 sg13g2_decap_8 FILLER_63_1107 ();
 sg13g2_decap_8 FILLER_63_1114 ();
 sg13g2_decap_8 FILLER_63_1121 ();
 sg13g2_decap_8 FILLER_63_1128 ();
 sg13g2_decap_8 FILLER_63_1135 ();
 sg13g2_decap_8 FILLER_63_1142 ();
 sg13g2_decap_8 FILLER_63_1149 ();
 sg13g2_decap_8 FILLER_63_1156 ();
 sg13g2_decap_8 FILLER_63_1163 ();
 sg13g2_decap_8 FILLER_63_1170 ();
 sg13g2_decap_8 FILLER_63_1177 ();
 sg13g2_decap_8 FILLER_63_1184 ();
 sg13g2_decap_8 FILLER_63_1191 ();
 sg13g2_decap_8 FILLER_63_1198 ();
 sg13g2_decap_8 FILLER_63_1205 ();
 sg13g2_decap_8 FILLER_63_1212 ();
 sg13g2_decap_8 FILLER_63_1219 ();
 sg13g2_decap_8 FILLER_63_1226 ();
 sg13g2_decap_8 FILLER_63_1233 ();
 sg13g2_decap_8 FILLER_63_1240 ();
 sg13g2_decap_8 FILLER_63_1247 ();
 sg13g2_decap_8 FILLER_63_1254 ();
 sg13g2_decap_8 FILLER_63_1261 ();
 sg13g2_decap_8 FILLER_63_1268 ();
 sg13g2_decap_8 FILLER_63_1275 ();
 sg13g2_decap_8 FILLER_63_1282 ();
 sg13g2_decap_8 FILLER_63_1289 ();
 sg13g2_decap_8 FILLER_63_1296 ();
 sg13g2_decap_8 FILLER_63_1303 ();
 sg13g2_decap_4 FILLER_63_1310 ();
 sg13g2_fill_1 FILLER_63_1314 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_16 ();
 sg13g2_fill_1 FILLER_64_46 ();
 sg13g2_fill_1 FILLER_64_61 ();
 sg13g2_decap_8 FILLER_64_85 ();
 sg13g2_decap_4 FILLER_64_92 ();
 sg13g2_fill_2 FILLER_64_96 ();
 sg13g2_fill_2 FILLER_64_132 ();
 sg13g2_fill_2 FILLER_64_160 ();
 sg13g2_fill_1 FILLER_64_162 ();
 sg13g2_fill_1 FILLER_64_168 ();
 sg13g2_fill_2 FILLER_64_200 ();
 sg13g2_fill_1 FILLER_64_202 ();
 sg13g2_fill_2 FILLER_64_230 ();
 sg13g2_fill_1 FILLER_64_232 ();
 sg13g2_fill_2 FILLER_64_326 ();
 sg13g2_fill_1 FILLER_64_328 ();
 sg13g2_fill_2 FILLER_64_334 ();
 sg13g2_fill_1 FILLER_64_336 ();
 sg13g2_fill_2 FILLER_64_354 ();
 sg13g2_fill_2 FILLER_64_396 ();
 sg13g2_fill_1 FILLER_64_398 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_2 FILLER_64_414 ();
 sg13g2_fill_1 FILLER_64_430 ();
 sg13g2_fill_2 FILLER_64_435 ();
 sg13g2_fill_1 FILLER_64_437 ();
 sg13g2_fill_2 FILLER_64_447 ();
 sg13g2_fill_1 FILLER_64_458 ();
 sg13g2_decap_4 FILLER_64_463 ();
 sg13g2_fill_1 FILLER_64_471 ();
 sg13g2_fill_2 FILLER_64_525 ();
 sg13g2_fill_2 FILLER_64_534 ();
 sg13g2_fill_1 FILLER_64_542 ();
 sg13g2_decap_8 FILLER_64_601 ();
 sg13g2_fill_1 FILLER_64_608 ();
 sg13g2_fill_2 FILLER_64_614 ();
 sg13g2_fill_1 FILLER_64_616 ();
 sg13g2_fill_1 FILLER_64_630 ();
 sg13g2_decap_8 FILLER_64_636 ();
 sg13g2_fill_1 FILLER_64_646 ();
 sg13g2_decap_8 FILLER_64_668 ();
 sg13g2_decap_8 FILLER_64_675 ();
 sg13g2_decap_4 FILLER_64_682 ();
 sg13g2_decap_8 FILLER_64_710 ();
 sg13g2_fill_2 FILLER_64_717 ();
 sg13g2_fill_1 FILLER_64_719 ();
 sg13g2_decap_8 FILLER_64_724 ();
 sg13g2_decap_8 FILLER_64_731 ();
 sg13g2_decap_4 FILLER_64_738 ();
 sg13g2_fill_2 FILLER_64_742 ();
 sg13g2_fill_1 FILLER_64_791 ();
 sg13g2_decap_8 FILLER_64_800 ();
 sg13g2_fill_2 FILLER_64_807 ();
 sg13g2_fill_1 FILLER_64_809 ();
 sg13g2_fill_2 FILLER_64_817 ();
 sg13g2_decap_4 FILLER_64_837 ();
 sg13g2_fill_2 FILLER_64_841 ();
 sg13g2_fill_1 FILLER_64_851 ();
 sg13g2_decap_4 FILLER_64_881 ();
 sg13g2_fill_1 FILLER_64_894 ();
 sg13g2_fill_1 FILLER_64_921 ();
 sg13g2_fill_1 FILLER_64_958 ();
 sg13g2_decap_8 FILLER_64_994 ();
 sg13g2_decap_8 FILLER_64_1001 ();
 sg13g2_decap_8 FILLER_64_1008 ();
 sg13g2_decap_8 FILLER_64_1015 ();
 sg13g2_decap_8 FILLER_64_1022 ();
 sg13g2_decap_8 FILLER_64_1029 ();
 sg13g2_decap_8 FILLER_64_1036 ();
 sg13g2_decap_8 FILLER_64_1043 ();
 sg13g2_decap_8 FILLER_64_1050 ();
 sg13g2_decap_8 FILLER_64_1057 ();
 sg13g2_decap_8 FILLER_64_1064 ();
 sg13g2_decap_8 FILLER_64_1071 ();
 sg13g2_decap_8 FILLER_64_1078 ();
 sg13g2_decap_8 FILLER_64_1085 ();
 sg13g2_decap_8 FILLER_64_1092 ();
 sg13g2_decap_8 FILLER_64_1099 ();
 sg13g2_decap_8 FILLER_64_1106 ();
 sg13g2_decap_8 FILLER_64_1113 ();
 sg13g2_decap_8 FILLER_64_1120 ();
 sg13g2_decap_8 FILLER_64_1127 ();
 sg13g2_decap_8 FILLER_64_1134 ();
 sg13g2_decap_8 FILLER_64_1141 ();
 sg13g2_decap_8 FILLER_64_1148 ();
 sg13g2_decap_8 FILLER_64_1155 ();
 sg13g2_decap_8 FILLER_64_1162 ();
 sg13g2_decap_8 FILLER_64_1169 ();
 sg13g2_decap_8 FILLER_64_1176 ();
 sg13g2_decap_8 FILLER_64_1183 ();
 sg13g2_decap_8 FILLER_64_1190 ();
 sg13g2_decap_8 FILLER_64_1197 ();
 sg13g2_decap_8 FILLER_64_1204 ();
 sg13g2_decap_8 FILLER_64_1211 ();
 sg13g2_decap_8 FILLER_64_1218 ();
 sg13g2_decap_8 FILLER_64_1225 ();
 sg13g2_decap_8 FILLER_64_1232 ();
 sg13g2_decap_8 FILLER_64_1239 ();
 sg13g2_decap_8 FILLER_64_1246 ();
 sg13g2_decap_8 FILLER_64_1253 ();
 sg13g2_decap_8 FILLER_64_1260 ();
 sg13g2_decap_8 FILLER_64_1267 ();
 sg13g2_decap_8 FILLER_64_1274 ();
 sg13g2_decap_8 FILLER_64_1281 ();
 sg13g2_decap_8 FILLER_64_1288 ();
 sg13g2_decap_8 FILLER_64_1295 ();
 sg13g2_decap_8 FILLER_64_1302 ();
 sg13g2_decap_4 FILLER_64_1309 ();
 sg13g2_fill_2 FILLER_64_1313 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_78 ();
 sg13g2_fill_1 FILLER_65_80 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_4 FILLER_65_91 ();
 sg13g2_fill_2 FILLER_65_95 ();
 sg13g2_fill_2 FILLER_65_120 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_fill_2 FILLER_65_171 ();
 sg13g2_decap_8 FILLER_65_191 ();
 sg13g2_decap_4 FILLER_65_198 ();
 sg13g2_fill_2 FILLER_65_202 ();
 sg13g2_fill_2 FILLER_65_208 ();
 sg13g2_fill_1 FILLER_65_210 ();
 sg13g2_decap_4 FILLER_65_217 ();
 sg13g2_fill_2 FILLER_65_261 ();
 sg13g2_fill_2 FILLER_65_295 ();
 sg13g2_fill_2 FILLER_65_314 ();
 sg13g2_fill_2 FILLER_65_348 ();
 sg13g2_fill_1 FILLER_65_350 ();
 sg13g2_fill_1 FILLER_65_364 ();
 sg13g2_fill_2 FILLER_65_455 ();
 sg13g2_fill_1 FILLER_65_471 ();
 sg13g2_fill_2 FILLER_65_493 ();
 sg13g2_fill_2 FILLER_65_512 ();
 sg13g2_fill_2 FILLER_65_518 ();
 sg13g2_fill_1 FILLER_65_520 ();
 sg13g2_fill_2 FILLER_65_526 ();
 sg13g2_decap_4 FILLER_65_535 ();
 sg13g2_fill_2 FILLER_65_586 ();
 sg13g2_fill_1 FILLER_65_588 ();
 sg13g2_fill_2 FILLER_65_647 ();
 sg13g2_decap_8 FILLER_65_663 ();
 sg13g2_decap_4 FILLER_65_670 ();
 sg13g2_fill_2 FILLER_65_674 ();
 sg13g2_fill_1 FILLER_65_766 ();
 sg13g2_fill_2 FILLER_65_778 ();
 sg13g2_fill_1 FILLER_65_780 ();
 sg13g2_decap_4 FILLER_65_798 ();
 sg13g2_fill_2 FILLER_65_815 ();
 sg13g2_decap_8 FILLER_65_827 ();
 sg13g2_fill_2 FILLER_65_834 ();
 sg13g2_fill_1 FILLER_65_836 ();
 sg13g2_decap_4 FILLER_65_842 ();
 sg13g2_fill_1 FILLER_65_854 ();
 sg13g2_fill_2 FILLER_65_869 ();
 sg13g2_fill_1 FILLER_65_871 ();
 sg13g2_fill_2 FILLER_65_885 ();
 sg13g2_fill_1 FILLER_65_898 ();
 sg13g2_decap_8 FILLER_65_912 ();
 sg13g2_fill_2 FILLER_65_957 ();
 sg13g2_fill_1 FILLER_65_968 ();
 sg13g2_decap_8 FILLER_65_1000 ();
 sg13g2_decap_8 FILLER_65_1007 ();
 sg13g2_decap_8 FILLER_65_1014 ();
 sg13g2_decap_8 FILLER_65_1021 ();
 sg13g2_decap_8 FILLER_65_1028 ();
 sg13g2_decap_8 FILLER_65_1035 ();
 sg13g2_decap_8 FILLER_65_1042 ();
 sg13g2_decap_8 FILLER_65_1049 ();
 sg13g2_decap_8 FILLER_65_1056 ();
 sg13g2_decap_8 FILLER_65_1063 ();
 sg13g2_decap_8 FILLER_65_1070 ();
 sg13g2_decap_8 FILLER_65_1077 ();
 sg13g2_decap_8 FILLER_65_1084 ();
 sg13g2_decap_8 FILLER_65_1091 ();
 sg13g2_decap_8 FILLER_65_1098 ();
 sg13g2_decap_8 FILLER_65_1105 ();
 sg13g2_decap_8 FILLER_65_1112 ();
 sg13g2_decap_8 FILLER_65_1119 ();
 sg13g2_decap_8 FILLER_65_1126 ();
 sg13g2_decap_8 FILLER_65_1133 ();
 sg13g2_decap_8 FILLER_65_1140 ();
 sg13g2_decap_8 FILLER_65_1147 ();
 sg13g2_decap_8 FILLER_65_1154 ();
 sg13g2_decap_8 FILLER_65_1161 ();
 sg13g2_decap_8 FILLER_65_1168 ();
 sg13g2_decap_8 FILLER_65_1175 ();
 sg13g2_decap_8 FILLER_65_1182 ();
 sg13g2_decap_8 FILLER_65_1189 ();
 sg13g2_decap_8 FILLER_65_1196 ();
 sg13g2_decap_8 FILLER_65_1203 ();
 sg13g2_decap_8 FILLER_65_1210 ();
 sg13g2_decap_8 FILLER_65_1217 ();
 sg13g2_decap_8 FILLER_65_1224 ();
 sg13g2_decap_8 FILLER_65_1231 ();
 sg13g2_decap_8 FILLER_65_1238 ();
 sg13g2_decap_8 FILLER_65_1245 ();
 sg13g2_decap_8 FILLER_65_1252 ();
 sg13g2_decap_8 FILLER_65_1259 ();
 sg13g2_decap_8 FILLER_65_1266 ();
 sg13g2_decap_8 FILLER_65_1273 ();
 sg13g2_decap_8 FILLER_65_1280 ();
 sg13g2_decap_8 FILLER_65_1287 ();
 sg13g2_decap_8 FILLER_65_1294 ();
 sg13g2_decap_8 FILLER_65_1301 ();
 sg13g2_decap_8 FILLER_65_1308 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_21 ();
 sg13g2_fill_2 FILLER_66_74 ();
 sg13g2_fill_1 FILLER_66_76 ();
 sg13g2_fill_2 FILLER_66_150 ();
 sg13g2_fill_1 FILLER_66_152 ();
 sg13g2_fill_2 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_247 ();
 sg13g2_fill_2 FILLER_66_282 ();
 sg13g2_fill_2 FILLER_66_289 ();
 sg13g2_fill_1 FILLER_66_291 ();
 sg13g2_decap_4 FILLER_66_391 ();
 sg13g2_fill_2 FILLER_66_395 ();
 sg13g2_fill_1 FILLER_66_405 ();
 sg13g2_decap_8 FILLER_66_466 ();
 sg13g2_fill_1 FILLER_66_473 ();
 sg13g2_fill_1 FILLER_66_478 ();
 sg13g2_decap_8 FILLER_66_483 ();
 sg13g2_decap_4 FILLER_66_490 ();
 sg13g2_fill_2 FILLER_66_494 ();
 sg13g2_fill_1 FILLER_66_543 ();
 sg13g2_fill_1 FILLER_66_580 ();
 sg13g2_decap_8 FILLER_66_594 ();
 sg13g2_decap_8 FILLER_66_601 ();
 sg13g2_fill_2 FILLER_66_626 ();
 sg13g2_fill_1 FILLER_66_633 ();
 sg13g2_fill_2 FILLER_66_659 ();
 sg13g2_fill_1 FILLER_66_692 ();
 sg13g2_fill_1 FILLER_66_726 ();
 sg13g2_fill_1 FILLER_66_757 ();
 sg13g2_fill_1 FILLER_66_777 ();
 sg13g2_fill_1 FILLER_66_797 ();
 sg13g2_decap_4 FILLER_66_841 ();
 sg13g2_fill_2 FILLER_66_863 ();
 sg13g2_fill_1 FILLER_66_865 ();
 sg13g2_fill_2 FILLER_66_940 ();
 sg13g2_fill_1 FILLER_66_942 ();
 sg13g2_decap_8 FILLER_66_996 ();
 sg13g2_decap_8 FILLER_66_1003 ();
 sg13g2_decap_8 FILLER_66_1010 ();
 sg13g2_decap_8 FILLER_66_1017 ();
 sg13g2_decap_8 FILLER_66_1024 ();
 sg13g2_decap_8 FILLER_66_1031 ();
 sg13g2_decap_8 FILLER_66_1038 ();
 sg13g2_decap_8 FILLER_66_1045 ();
 sg13g2_decap_8 FILLER_66_1052 ();
 sg13g2_decap_8 FILLER_66_1059 ();
 sg13g2_decap_8 FILLER_66_1066 ();
 sg13g2_decap_8 FILLER_66_1073 ();
 sg13g2_decap_8 FILLER_66_1080 ();
 sg13g2_decap_8 FILLER_66_1087 ();
 sg13g2_decap_8 FILLER_66_1094 ();
 sg13g2_decap_8 FILLER_66_1101 ();
 sg13g2_decap_8 FILLER_66_1108 ();
 sg13g2_decap_8 FILLER_66_1115 ();
 sg13g2_decap_8 FILLER_66_1122 ();
 sg13g2_decap_8 FILLER_66_1129 ();
 sg13g2_decap_8 FILLER_66_1136 ();
 sg13g2_decap_8 FILLER_66_1143 ();
 sg13g2_decap_8 FILLER_66_1150 ();
 sg13g2_decap_8 FILLER_66_1157 ();
 sg13g2_decap_8 FILLER_66_1164 ();
 sg13g2_decap_8 FILLER_66_1171 ();
 sg13g2_decap_8 FILLER_66_1178 ();
 sg13g2_decap_8 FILLER_66_1185 ();
 sg13g2_decap_8 FILLER_66_1192 ();
 sg13g2_decap_8 FILLER_66_1199 ();
 sg13g2_decap_8 FILLER_66_1206 ();
 sg13g2_decap_8 FILLER_66_1213 ();
 sg13g2_decap_8 FILLER_66_1220 ();
 sg13g2_decap_8 FILLER_66_1227 ();
 sg13g2_decap_8 FILLER_66_1234 ();
 sg13g2_decap_8 FILLER_66_1241 ();
 sg13g2_decap_8 FILLER_66_1248 ();
 sg13g2_decap_8 FILLER_66_1255 ();
 sg13g2_decap_8 FILLER_66_1262 ();
 sg13g2_decap_8 FILLER_66_1269 ();
 sg13g2_decap_8 FILLER_66_1276 ();
 sg13g2_decap_8 FILLER_66_1283 ();
 sg13g2_decap_8 FILLER_66_1290 ();
 sg13g2_decap_8 FILLER_66_1297 ();
 sg13g2_decap_8 FILLER_66_1304 ();
 sg13g2_decap_4 FILLER_66_1311 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_fill_2 FILLER_67_53 ();
 sg13g2_fill_2 FILLER_67_81 ();
 sg13g2_fill_2 FILLER_67_118 ();
 sg13g2_fill_1 FILLER_67_138 ();
 sg13g2_fill_1 FILLER_67_143 ();
 sg13g2_fill_1 FILLER_67_187 ();
 sg13g2_fill_1 FILLER_67_193 ();
 sg13g2_fill_2 FILLER_67_198 ();
 sg13g2_fill_1 FILLER_67_200 ();
 sg13g2_decap_8 FILLER_67_306 ();
 sg13g2_fill_1 FILLER_67_339 ();
 sg13g2_fill_2 FILLER_67_371 ();
 sg13g2_fill_1 FILLER_67_373 ();
 sg13g2_decap_8 FILLER_67_391 ();
 sg13g2_fill_2 FILLER_67_398 ();
 sg13g2_fill_2 FILLER_67_412 ();
 sg13g2_fill_2 FILLER_67_423 ();
 sg13g2_fill_1 FILLER_67_439 ();
 sg13g2_fill_1 FILLER_67_448 ();
 sg13g2_fill_1 FILLER_67_457 ();
 sg13g2_decap_8 FILLER_67_494 ();
 sg13g2_decap_4 FILLER_67_501 ();
 sg13g2_fill_2 FILLER_67_512 ();
 sg13g2_fill_1 FILLER_67_514 ();
 sg13g2_decap_8 FILLER_67_526 ();
 sg13g2_fill_2 FILLER_67_537 ();
 sg13g2_fill_1 FILLER_67_628 ();
 sg13g2_fill_2 FILLER_67_651 ();
 sg13g2_fill_1 FILLER_67_653 ();
 sg13g2_fill_2 FILLER_67_660 ();
 sg13g2_fill_1 FILLER_67_662 ();
 sg13g2_fill_2 FILLER_67_682 ();
 sg13g2_fill_1 FILLER_67_684 ();
 sg13g2_fill_1 FILLER_67_746 ();
 sg13g2_decap_4 FILLER_67_773 ();
 sg13g2_fill_2 FILLER_67_807 ();
 sg13g2_fill_1 FILLER_67_809 ();
 sg13g2_decap_4 FILLER_67_830 ();
 sg13g2_decap_8 FILLER_67_866 ();
 sg13g2_fill_2 FILLER_67_873 ();
 sg13g2_fill_1 FILLER_67_875 ();
 sg13g2_fill_2 FILLER_67_887 ();
 sg13g2_fill_2 FILLER_67_897 ();
 sg13g2_fill_1 FILLER_67_918 ();
 sg13g2_fill_1 FILLER_67_940 ();
 sg13g2_fill_2 FILLER_67_980 ();
 sg13g2_decap_8 FILLER_67_986 ();
 sg13g2_decap_8 FILLER_67_993 ();
 sg13g2_decap_8 FILLER_67_1000 ();
 sg13g2_decap_8 FILLER_67_1007 ();
 sg13g2_decap_8 FILLER_67_1014 ();
 sg13g2_decap_8 FILLER_67_1021 ();
 sg13g2_decap_8 FILLER_67_1028 ();
 sg13g2_decap_8 FILLER_67_1035 ();
 sg13g2_decap_8 FILLER_67_1042 ();
 sg13g2_decap_8 FILLER_67_1049 ();
 sg13g2_decap_8 FILLER_67_1056 ();
 sg13g2_decap_8 FILLER_67_1063 ();
 sg13g2_decap_8 FILLER_67_1070 ();
 sg13g2_decap_8 FILLER_67_1077 ();
 sg13g2_decap_8 FILLER_67_1084 ();
 sg13g2_decap_8 FILLER_67_1091 ();
 sg13g2_decap_8 FILLER_67_1098 ();
 sg13g2_decap_8 FILLER_67_1105 ();
 sg13g2_decap_8 FILLER_67_1112 ();
 sg13g2_decap_8 FILLER_67_1119 ();
 sg13g2_decap_8 FILLER_67_1126 ();
 sg13g2_decap_8 FILLER_67_1133 ();
 sg13g2_decap_8 FILLER_67_1140 ();
 sg13g2_decap_8 FILLER_67_1147 ();
 sg13g2_decap_8 FILLER_67_1154 ();
 sg13g2_decap_8 FILLER_67_1161 ();
 sg13g2_decap_8 FILLER_67_1168 ();
 sg13g2_decap_8 FILLER_67_1175 ();
 sg13g2_decap_8 FILLER_67_1182 ();
 sg13g2_decap_8 FILLER_67_1189 ();
 sg13g2_decap_8 FILLER_67_1196 ();
 sg13g2_decap_8 FILLER_67_1203 ();
 sg13g2_decap_8 FILLER_67_1210 ();
 sg13g2_decap_8 FILLER_67_1217 ();
 sg13g2_decap_8 FILLER_67_1224 ();
 sg13g2_decap_8 FILLER_67_1231 ();
 sg13g2_decap_8 FILLER_67_1238 ();
 sg13g2_decap_8 FILLER_67_1245 ();
 sg13g2_decap_8 FILLER_67_1252 ();
 sg13g2_decap_8 FILLER_67_1259 ();
 sg13g2_decap_8 FILLER_67_1266 ();
 sg13g2_decap_8 FILLER_67_1273 ();
 sg13g2_decap_8 FILLER_67_1280 ();
 sg13g2_decap_8 FILLER_67_1287 ();
 sg13g2_decap_8 FILLER_67_1294 ();
 sg13g2_decap_8 FILLER_67_1301 ();
 sg13g2_decap_8 FILLER_67_1308 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_4 ();
 sg13g2_fill_2 FILLER_68_96 ();
 sg13g2_fill_1 FILLER_68_98 ();
 sg13g2_fill_2 FILLER_68_143 ();
 sg13g2_fill_1 FILLER_68_145 ();
 sg13g2_fill_2 FILLER_68_171 ();
 sg13g2_fill_1 FILLER_68_173 ();
 sg13g2_fill_2 FILLER_68_191 ();
 sg13g2_decap_4 FILLER_68_240 ();
 sg13g2_fill_2 FILLER_68_253 ();
 sg13g2_decap_4 FILLER_68_297 ();
 sg13g2_decap_8 FILLER_68_335 ();
 sg13g2_decap_8 FILLER_68_342 ();
 sg13g2_decap_4 FILLER_68_366 ();
 sg13g2_fill_2 FILLER_68_370 ();
 sg13g2_fill_2 FILLER_68_403 ();
 sg13g2_fill_2 FILLER_68_441 ();
 sg13g2_fill_2 FILLER_68_451 ();
 sg13g2_fill_2 FILLER_68_462 ();
 sg13g2_decap_8 FILLER_68_485 ();
 sg13g2_fill_2 FILLER_68_492 ();
 sg13g2_fill_1 FILLER_68_494 ();
 sg13g2_fill_2 FILLER_68_548 ();
 sg13g2_fill_1 FILLER_68_550 ();
 sg13g2_fill_2 FILLER_68_577 ();
 sg13g2_fill_1 FILLER_68_579 ();
 sg13g2_decap_4 FILLER_68_598 ();
 sg13g2_fill_2 FILLER_68_602 ();
 sg13g2_decap_4 FILLER_68_608 ();
 sg13g2_fill_1 FILLER_68_623 ();
 sg13g2_fill_1 FILLER_68_639 ();
 sg13g2_fill_1 FILLER_68_668 ();
 sg13g2_fill_2 FILLER_68_676 ();
 sg13g2_fill_1 FILLER_68_678 ();
 sg13g2_fill_1 FILLER_68_695 ();
 sg13g2_decap_4 FILLER_68_701 ();
 sg13g2_fill_2 FILLER_68_705 ();
 sg13g2_decap_4 FILLER_68_715 ();
 sg13g2_fill_1 FILLER_68_719 ();
 sg13g2_decap_8 FILLER_68_724 ();
 sg13g2_fill_2 FILLER_68_731 ();
 sg13g2_decap_4 FILLER_68_750 ();
 sg13g2_fill_1 FILLER_68_754 ();
 sg13g2_fill_2 FILLER_68_776 ();
 sg13g2_decap_4 FILLER_68_792 ();
 sg13g2_fill_2 FILLER_68_796 ();
 sg13g2_decap_8 FILLER_68_803 ();
 sg13g2_decap_8 FILLER_68_844 ();
 sg13g2_decap_8 FILLER_68_851 ();
 sg13g2_decap_4 FILLER_68_858 ();
 sg13g2_fill_1 FILLER_68_871 ();
 sg13g2_decap_4 FILLER_68_881 ();
 sg13g2_fill_1 FILLER_68_944 ();
 sg13g2_fill_2 FILLER_68_954 ();
 sg13g2_fill_1 FILLER_68_956 ();
 sg13g2_fill_1 FILLER_68_988 ();
 sg13g2_decap_4 FILLER_68_993 ();
 sg13g2_fill_1 FILLER_68_1001 ();
 sg13g2_decap_4 FILLER_68_1006 ();
 sg13g2_decap_8 FILLER_68_1014 ();
 sg13g2_decap_8 FILLER_68_1021 ();
 sg13g2_decap_8 FILLER_68_1028 ();
 sg13g2_decap_8 FILLER_68_1035 ();
 sg13g2_decap_8 FILLER_68_1042 ();
 sg13g2_decap_8 FILLER_68_1049 ();
 sg13g2_decap_8 FILLER_68_1056 ();
 sg13g2_decap_8 FILLER_68_1063 ();
 sg13g2_decap_8 FILLER_68_1070 ();
 sg13g2_decap_8 FILLER_68_1077 ();
 sg13g2_decap_8 FILLER_68_1084 ();
 sg13g2_decap_8 FILLER_68_1091 ();
 sg13g2_decap_8 FILLER_68_1098 ();
 sg13g2_decap_8 FILLER_68_1105 ();
 sg13g2_decap_8 FILLER_68_1112 ();
 sg13g2_decap_8 FILLER_68_1119 ();
 sg13g2_decap_8 FILLER_68_1126 ();
 sg13g2_decap_8 FILLER_68_1133 ();
 sg13g2_decap_8 FILLER_68_1140 ();
 sg13g2_decap_8 FILLER_68_1147 ();
 sg13g2_decap_8 FILLER_68_1154 ();
 sg13g2_decap_8 FILLER_68_1161 ();
 sg13g2_decap_8 FILLER_68_1168 ();
 sg13g2_decap_8 FILLER_68_1175 ();
 sg13g2_decap_8 FILLER_68_1182 ();
 sg13g2_decap_8 FILLER_68_1189 ();
 sg13g2_decap_8 FILLER_68_1196 ();
 sg13g2_decap_8 FILLER_68_1203 ();
 sg13g2_decap_8 FILLER_68_1210 ();
 sg13g2_decap_8 FILLER_68_1217 ();
 sg13g2_decap_8 FILLER_68_1224 ();
 sg13g2_decap_8 FILLER_68_1231 ();
 sg13g2_decap_8 FILLER_68_1238 ();
 sg13g2_decap_8 FILLER_68_1245 ();
 sg13g2_decap_8 FILLER_68_1252 ();
 sg13g2_decap_8 FILLER_68_1259 ();
 sg13g2_decap_8 FILLER_68_1266 ();
 sg13g2_decap_8 FILLER_68_1273 ();
 sg13g2_decap_8 FILLER_68_1280 ();
 sg13g2_decap_8 FILLER_68_1287 ();
 sg13g2_decap_8 FILLER_68_1294 ();
 sg13g2_decap_8 FILLER_68_1301 ();
 sg13g2_decap_8 FILLER_68_1308 ();
 sg13g2_fill_2 FILLER_69_77 ();
 sg13g2_fill_1 FILLER_69_124 ();
 sg13g2_fill_1 FILLER_69_168 ();
 sg13g2_fill_1 FILLER_69_200 ();
 sg13g2_fill_1 FILLER_69_211 ();
 sg13g2_decap_8 FILLER_69_221 ();
 sg13g2_fill_1 FILLER_69_233 ();
 sg13g2_fill_2 FILLER_69_274 ();
 sg13g2_fill_1 FILLER_69_323 ();
 sg13g2_fill_2 FILLER_69_328 ();
 sg13g2_fill_1 FILLER_69_330 ();
 sg13g2_decap_4 FILLER_69_379 ();
 sg13g2_fill_2 FILLER_69_419 ();
 sg13g2_decap_4 FILLER_69_425 ();
 sg13g2_decap_4 FILLER_69_433 ();
 sg13g2_fill_1 FILLER_69_437 ();
 sg13g2_decap_4 FILLER_69_447 ();
 sg13g2_fill_1 FILLER_69_451 ();
 sg13g2_fill_2 FILLER_69_460 ();
 sg13g2_fill_2 FILLER_69_517 ();
 sg13g2_decap_4 FILLER_69_566 ();
 sg13g2_decap_8 FILLER_69_609 ();
 sg13g2_fill_2 FILLER_69_616 ();
 sg13g2_fill_1 FILLER_69_618 ();
 sg13g2_fill_2 FILLER_69_654 ();
 sg13g2_fill_1 FILLER_69_662 ();
 sg13g2_fill_2 FILLER_69_688 ();
 sg13g2_fill_2 FILLER_69_699 ();
 sg13g2_decap_4 FILLER_69_731 ();
 sg13g2_fill_2 FILLER_69_735 ();
 sg13g2_decap_4 FILLER_69_742 ();
 sg13g2_fill_1 FILLER_69_746 ();
 sg13g2_fill_1 FILLER_69_778 ();
 sg13g2_fill_2 FILLER_69_784 ();
 sg13g2_decap_4 FILLER_69_795 ();
 sg13g2_fill_2 FILLER_69_799 ();
 sg13g2_decap_4 FILLER_69_822 ();
 sg13g2_fill_2 FILLER_69_894 ();
 sg13g2_fill_2 FILLER_69_909 ();
 sg13g2_fill_2 FILLER_69_924 ();
 sg13g2_decap_8 FILLER_69_1027 ();
 sg13g2_decap_8 FILLER_69_1034 ();
 sg13g2_decap_8 FILLER_69_1041 ();
 sg13g2_decap_8 FILLER_69_1048 ();
 sg13g2_decap_8 FILLER_69_1055 ();
 sg13g2_decap_8 FILLER_69_1062 ();
 sg13g2_decap_8 FILLER_69_1069 ();
 sg13g2_decap_8 FILLER_69_1076 ();
 sg13g2_decap_8 FILLER_69_1083 ();
 sg13g2_decap_8 FILLER_69_1090 ();
 sg13g2_decap_8 FILLER_69_1097 ();
 sg13g2_decap_8 FILLER_69_1104 ();
 sg13g2_decap_8 FILLER_69_1111 ();
 sg13g2_decap_8 FILLER_69_1118 ();
 sg13g2_decap_8 FILLER_69_1125 ();
 sg13g2_decap_8 FILLER_69_1132 ();
 sg13g2_decap_8 FILLER_69_1139 ();
 sg13g2_decap_8 FILLER_69_1146 ();
 sg13g2_decap_8 FILLER_69_1153 ();
 sg13g2_decap_8 FILLER_69_1160 ();
 sg13g2_decap_8 FILLER_69_1167 ();
 sg13g2_decap_8 FILLER_69_1174 ();
 sg13g2_decap_8 FILLER_69_1181 ();
 sg13g2_decap_8 FILLER_69_1188 ();
 sg13g2_decap_8 FILLER_69_1195 ();
 sg13g2_decap_8 FILLER_69_1202 ();
 sg13g2_decap_8 FILLER_69_1209 ();
 sg13g2_decap_8 FILLER_69_1216 ();
 sg13g2_decap_8 FILLER_69_1223 ();
 sg13g2_decap_8 FILLER_69_1230 ();
 sg13g2_decap_8 FILLER_69_1237 ();
 sg13g2_decap_8 FILLER_69_1244 ();
 sg13g2_decap_8 FILLER_69_1251 ();
 sg13g2_decap_8 FILLER_69_1258 ();
 sg13g2_decap_8 FILLER_69_1265 ();
 sg13g2_decap_8 FILLER_69_1272 ();
 sg13g2_decap_8 FILLER_69_1279 ();
 sg13g2_decap_8 FILLER_69_1286 ();
 sg13g2_decap_8 FILLER_69_1293 ();
 sg13g2_decap_8 FILLER_69_1300 ();
 sg13g2_decap_8 FILLER_69_1307 ();
 sg13g2_fill_1 FILLER_69_1314 ();
 sg13g2_fill_1 FILLER_70_54 ();
 sg13g2_fill_2 FILLER_70_81 ();
 sg13g2_fill_1 FILLER_70_145 ();
 sg13g2_fill_1 FILLER_70_151 ();
 sg13g2_fill_2 FILLER_70_161 ();
 sg13g2_fill_1 FILLER_70_163 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_4 FILLER_70_189 ();
 sg13g2_fill_1 FILLER_70_193 ();
 sg13g2_fill_1 FILLER_70_199 ();
 sg13g2_decap_4 FILLER_70_235 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_decap_4 FILLER_70_301 ();
 sg13g2_fill_2 FILLER_70_310 ();
 sg13g2_decap_4 FILLER_70_320 ();
 sg13g2_fill_2 FILLER_70_324 ();
 sg13g2_decap_8 FILLER_70_334 ();
 sg13g2_fill_2 FILLER_70_341 ();
 sg13g2_fill_2 FILLER_70_348 ();
 sg13g2_fill_1 FILLER_70_355 ();
 sg13g2_fill_2 FILLER_70_405 ();
 sg13g2_fill_1 FILLER_70_501 ();
 sg13g2_fill_2 FILLER_70_541 ();
 sg13g2_fill_1 FILLER_70_605 ();
 sg13g2_fill_2 FILLER_70_665 ();
 sg13g2_fill_1 FILLER_70_681 ();
 sg13g2_decap_4 FILLER_70_746 ();
 sg13g2_fill_2 FILLER_70_750 ();
 sg13g2_fill_2 FILLER_70_756 ();
 sg13g2_decap_8 FILLER_70_762 ();
 sg13g2_decap_4 FILLER_70_769 ();
 sg13g2_fill_2 FILLER_70_773 ();
 sg13g2_decap_4 FILLER_70_806 ();
 sg13g2_fill_1 FILLER_70_815 ();
 sg13g2_fill_1 FILLER_70_829 ();
 sg13g2_fill_1 FILLER_70_854 ();
 sg13g2_fill_2 FILLER_70_873 ();
 sg13g2_fill_1 FILLER_70_875 ();
 sg13g2_fill_2 FILLER_70_902 ();
 sg13g2_fill_2 FILLER_70_974 ();
 sg13g2_fill_1 FILLER_70_976 ();
 sg13g2_fill_2 FILLER_70_999 ();
 sg13g2_decap_8 FILLER_70_1033 ();
 sg13g2_decap_8 FILLER_70_1040 ();
 sg13g2_decap_8 FILLER_70_1047 ();
 sg13g2_decap_8 FILLER_70_1054 ();
 sg13g2_decap_8 FILLER_70_1061 ();
 sg13g2_decap_8 FILLER_70_1068 ();
 sg13g2_decap_8 FILLER_70_1075 ();
 sg13g2_decap_8 FILLER_70_1082 ();
 sg13g2_decap_8 FILLER_70_1089 ();
 sg13g2_decap_8 FILLER_70_1096 ();
 sg13g2_decap_8 FILLER_70_1103 ();
 sg13g2_decap_8 FILLER_70_1110 ();
 sg13g2_decap_8 FILLER_70_1117 ();
 sg13g2_decap_8 FILLER_70_1124 ();
 sg13g2_decap_8 FILLER_70_1131 ();
 sg13g2_decap_8 FILLER_70_1138 ();
 sg13g2_decap_8 FILLER_70_1145 ();
 sg13g2_decap_8 FILLER_70_1152 ();
 sg13g2_decap_8 FILLER_70_1159 ();
 sg13g2_decap_8 FILLER_70_1166 ();
 sg13g2_decap_8 FILLER_70_1173 ();
 sg13g2_decap_8 FILLER_70_1180 ();
 sg13g2_decap_8 FILLER_70_1187 ();
 sg13g2_decap_8 FILLER_70_1194 ();
 sg13g2_decap_8 FILLER_70_1201 ();
 sg13g2_decap_8 FILLER_70_1208 ();
 sg13g2_decap_8 FILLER_70_1215 ();
 sg13g2_decap_8 FILLER_70_1222 ();
 sg13g2_decap_8 FILLER_70_1229 ();
 sg13g2_decap_8 FILLER_70_1236 ();
 sg13g2_decap_8 FILLER_70_1243 ();
 sg13g2_decap_8 FILLER_70_1250 ();
 sg13g2_decap_8 FILLER_70_1257 ();
 sg13g2_decap_8 FILLER_70_1264 ();
 sg13g2_decap_8 FILLER_70_1271 ();
 sg13g2_decap_8 FILLER_70_1278 ();
 sg13g2_decap_8 FILLER_70_1285 ();
 sg13g2_decap_8 FILLER_70_1292 ();
 sg13g2_decap_8 FILLER_70_1299 ();
 sg13g2_decap_8 FILLER_70_1306 ();
 sg13g2_fill_2 FILLER_70_1313 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_2 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_44 ();
 sg13g2_fill_2 FILLER_71_54 ();
 sg13g2_fill_1 FILLER_71_75 ();
 sg13g2_fill_2 FILLER_71_106 ();
 sg13g2_fill_1 FILLER_71_108 ();
 sg13g2_fill_2 FILLER_71_166 ();
 sg13g2_fill_2 FILLER_71_203 ();
 sg13g2_fill_2 FILLER_71_271 ();
 sg13g2_fill_1 FILLER_71_273 ();
 sg13g2_fill_2 FILLER_71_352 ();
 sg13g2_fill_2 FILLER_71_385 ();
 sg13g2_fill_1 FILLER_71_387 ();
 sg13g2_fill_1 FILLER_71_401 ();
 sg13g2_fill_1 FILLER_71_412 ();
 sg13g2_decap_8 FILLER_71_430 ();
 sg13g2_fill_1 FILLER_71_437 ();
 sg13g2_fill_1 FILLER_71_460 ();
 sg13g2_fill_1 FILLER_71_479 ();
 sg13g2_fill_2 FILLER_71_498 ();
 sg13g2_fill_1 FILLER_71_500 ();
 sg13g2_fill_2 FILLER_71_509 ();
 sg13g2_fill_1 FILLER_71_511 ();
 sg13g2_decap_4 FILLER_71_573 ();
 sg13g2_fill_1 FILLER_71_577 ();
 sg13g2_fill_1 FILLER_71_621 ();
 sg13g2_fill_2 FILLER_71_692 ();
 sg13g2_fill_2 FILLER_71_717 ();
 sg13g2_decap_4 FILLER_71_772 ();
 sg13g2_fill_1 FILLER_71_776 ();
 sg13g2_fill_2 FILLER_71_785 ();
 sg13g2_fill_1 FILLER_71_787 ();
 sg13g2_fill_2 FILLER_71_793 ();
 sg13g2_fill_1 FILLER_71_827 ();
 sg13g2_fill_2 FILLER_71_885 ();
 sg13g2_fill_2 FILLER_71_891 ();
 sg13g2_fill_1 FILLER_71_915 ();
 sg13g2_fill_1 FILLER_71_1023 ();
 sg13g2_decap_8 FILLER_71_1045 ();
 sg13g2_decap_8 FILLER_71_1052 ();
 sg13g2_decap_8 FILLER_71_1059 ();
 sg13g2_decap_8 FILLER_71_1066 ();
 sg13g2_decap_8 FILLER_71_1073 ();
 sg13g2_decap_8 FILLER_71_1080 ();
 sg13g2_decap_8 FILLER_71_1087 ();
 sg13g2_decap_8 FILLER_71_1094 ();
 sg13g2_decap_8 FILLER_71_1101 ();
 sg13g2_decap_8 FILLER_71_1108 ();
 sg13g2_decap_8 FILLER_71_1115 ();
 sg13g2_decap_8 FILLER_71_1122 ();
 sg13g2_decap_8 FILLER_71_1129 ();
 sg13g2_decap_8 FILLER_71_1136 ();
 sg13g2_decap_8 FILLER_71_1143 ();
 sg13g2_decap_8 FILLER_71_1150 ();
 sg13g2_decap_8 FILLER_71_1157 ();
 sg13g2_decap_8 FILLER_71_1164 ();
 sg13g2_decap_8 FILLER_71_1171 ();
 sg13g2_decap_8 FILLER_71_1178 ();
 sg13g2_decap_8 FILLER_71_1185 ();
 sg13g2_decap_8 FILLER_71_1192 ();
 sg13g2_decap_8 FILLER_71_1199 ();
 sg13g2_decap_8 FILLER_71_1206 ();
 sg13g2_decap_8 FILLER_71_1213 ();
 sg13g2_decap_8 FILLER_71_1220 ();
 sg13g2_decap_8 FILLER_71_1227 ();
 sg13g2_decap_8 FILLER_71_1234 ();
 sg13g2_decap_8 FILLER_71_1241 ();
 sg13g2_decap_8 FILLER_71_1248 ();
 sg13g2_decap_8 FILLER_71_1255 ();
 sg13g2_decap_8 FILLER_71_1262 ();
 sg13g2_decap_8 FILLER_71_1269 ();
 sg13g2_decap_8 FILLER_71_1276 ();
 sg13g2_decap_8 FILLER_71_1283 ();
 sg13g2_decap_8 FILLER_71_1290 ();
 sg13g2_decap_8 FILLER_71_1297 ();
 sg13g2_decap_8 FILLER_71_1304 ();
 sg13g2_decap_4 FILLER_71_1311 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_2 ();
 sg13g2_fill_2 FILLER_72_38 ();
 sg13g2_fill_1 FILLER_72_40 ();
 sg13g2_fill_2 FILLER_72_50 ();
 sg13g2_fill_1 FILLER_72_88 ();
 sg13g2_fill_1 FILLER_72_141 ();
 sg13g2_fill_2 FILLER_72_146 ();
 sg13g2_fill_1 FILLER_72_148 ();
 sg13g2_decap_4 FILLER_72_171 ();
 sg13g2_fill_2 FILLER_72_189 ();
 sg13g2_fill_1 FILLER_72_191 ();
 sg13g2_fill_1 FILLER_72_212 ();
 sg13g2_fill_1 FILLER_72_225 ();
 sg13g2_decap_4 FILLER_72_231 ();
 sg13g2_fill_2 FILLER_72_235 ();
 sg13g2_decap_4 FILLER_72_241 ();
 sg13g2_fill_2 FILLER_72_245 ();
 sg13g2_fill_1 FILLER_72_255 ();
 sg13g2_fill_2 FILLER_72_287 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_fill_1 FILLER_72_307 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_fill_1 FILLER_72_317 ();
 sg13g2_decap_4 FILLER_72_327 ();
 sg13g2_fill_1 FILLER_72_331 ();
 sg13g2_fill_1 FILLER_72_358 ();
 sg13g2_fill_2 FILLER_72_371 ();
 sg13g2_fill_1 FILLER_72_373 ();
 sg13g2_fill_1 FILLER_72_413 ();
 sg13g2_fill_2 FILLER_72_426 ();
 sg13g2_fill_1 FILLER_72_437 ();
 sg13g2_fill_2 FILLER_72_442 ();
 sg13g2_fill_2 FILLER_72_453 ();
 sg13g2_fill_1 FILLER_72_455 ();
 sg13g2_fill_1 FILLER_72_522 ();
 sg13g2_fill_2 FILLER_72_532 ();
 sg13g2_fill_1 FILLER_72_534 ();
 sg13g2_fill_2 FILLER_72_565 ();
 sg13g2_fill_2 FILLER_72_711 ();
 sg13g2_fill_2 FILLER_72_747 ();
 sg13g2_fill_1 FILLER_72_749 ();
 sg13g2_decap_4 FILLER_72_762 ();
 sg13g2_fill_1 FILLER_72_807 ();
 sg13g2_fill_1 FILLER_72_853 ();
 sg13g2_fill_1 FILLER_72_871 ();
 sg13g2_fill_1 FILLER_72_894 ();
 sg13g2_fill_2 FILLER_72_903 ();
 sg13g2_fill_1 FILLER_72_917 ();
 sg13g2_fill_2 FILLER_72_984 ();
 sg13g2_decap_8 FILLER_72_1047 ();
 sg13g2_decap_8 FILLER_72_1054 ();
 sg13g2_decap_8 FILLER_72_1061 ();
 sg13g2_decap_8 FILLER_72_1068 ();
 sg13g2_decap_8 FILLER_72_1075 ();
 sg13g2_decap_8 FILLER_72_1082 ();
 sg13g2_decap_8 FILLER_72_1089 ();
 sg13g2_decap_8 FILLER_72_1096 ();
 sg13g2_decap_8 FILLER_72_1103 ();
 sg13g2_decap_8 FILLER_72_1110 ();
 sg13g2_decap_8 FILLER_72_1117 ();
 sg13g2_decap_8 FILLER_72_1124 ();
 sg13g2_decap_8 FILLER_72_1131 ();
 sg13g2_decap_8 FILLER_72_1138 ();
 sg13g2_decap_8 FILLER_72_1145 ();
 sg13g2_decap_8 FILLER_72_1152 ();
 sg13g2_decap_8 FILLER_72_1159 ();
 sg13g2_decap_8 FILLER_72_1166 ();
 sg13g2_decap_8 FILLER_72_1173 ();
 sg13g2_decap_8 FILLER_72_1180 ();
 sg13g2_decap_8 FILLER_72_1187 ();
 sg13g2_decap_8 FILLER_72_1194 ();
 sg13g2_decap_8 FILLER_72_1201 ();
 sg13g2_decap_8 FILLER_72_1208 ();
 sg13g2_decap_8 FILLER_72_1215 ();
 sg13g2_decap_8 FILLER_72_1222 ();
 sg13g2_decap_8 FILLER_72_1229 ();
 sg13g2_decap_8 FILLER_72_1236 ();
 sg13g2_decap_8 FILLER_72_1243 ();
 sg13g2_decap_8 FILLER_72_1250 ();
 sg13g2_decap_8 FILLER_72_1257 ();
 sg13g2_decap_8 FILLER_72_1264 ();
 sg13g2_decap_8 FILLER_72_1271 ();
 sg13g2_decap_8 FILLER_72_1278 ();
 sg13g2_decap_8 FILLER_72_1285 ();
 sg13g2_decap_8 FILLER_72_1292 ();
 sg13g2_decap_8 FILLER_72_1299 ();
 sg13g2_decap_8 FILLER_72_1306 ();
 sg13g2_fill_2 FILLER_72_1313 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_87 ();
 sg13g2_fill_1 FILLER_73_89 ();
 sg13g2_fill_2 FILLER_73_164 ();
 sg13g2_decap_4 FILLER_73_248 ();
 sg13g2_fill_2 FILLER_73_252 ();
 sg13g2_fill_1 FILLER_73_303 ();
 sg13g2_fill_2 FILLER_73_312 ();
 sg13g2_fill_2 FILLER_73_332 ();
 sg13g2_fill_2 FILLER_73_360 ();
 sg13g2_fill_2 FILLER_73_367 ();
 sg13g2_fill_2 FILLER_73_374 ();
 sg13g2_fill_1 FILLER_73_389 ();
 sg13g2_fill_2 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_421 ();
 sg13g2_fill_2 FILLER_73_425 ();
 sg13g2_fill_2 FILLER_73_458 ();
 sg13g2_fill_1 FILLER_73_460 ();
 sg13g2_decap_4 FILLER_73_486 ();
 sg13g2_fill_1 FILLER_73_490 ();
 sg13g2_decap_4 FILLER_73_496 ();
 sg13g2_fill_1 FILLER_73_500 ();
 sg13g2_fill_2 FILLER_73_505 ();
 sg13g2_decap_4 FILLER_73_511 ();
 sg13g2_fill_1 FILLER_73_557 ();
 sg13g2_fill_1 FILLER_73_596 ();
 sg13g2_decap_4 FILLER_73_606 ();
 sg13g2_fill_1 FILLER_73_610 ();
 sg13g2_decap_8 FILLER_73_633 ();
 sg13g2_fill_1 FILLER_73_640 ();
 sg13g2_fill_2 FILLER_73_649 ();
 sg13g2_fill_2 FILLER_73_655 ();
 sg13g2_fill_2 FILLER_73_693 ();
 sg13g2_fill_1 FILLER_73_704 ();
 sg13g2_fill_1 FILLER_73_710 ();
 sg13g2_fill_2 FILLER_73_725 ();
 sg13g2_fill_1 FILLER_73_760 ();
 sg13g2_decap_8 FILLER_73_783 ();
 sg13g2_fill_1 FILLER_73_790 ();
 sg13g2_fill_2 FILLER_73_809 ();
 sg13g2_fill_1 FILLER_73_837 ();
 sg13g2_fill_1 FILLER_73_843 ();
 sg13g2_fill_2 FILLER_73_870 ();
 sg13g2_fill_1 FILLER_73_872 ();
 sg13g2_fill_2 FILLER_73_954 ();
 sg13g2_fill_2 FILLER_73_972 ();
 sg13g2_fill_1 FILLER_73_974 ();
 sg13g2_fill_2 FILLER_73_992 ();
 sg13g2_decap_8 FILLER_73_1038 ();
 sg13g2_decap_8 FILLER_73_1045 ();
 sg13g2_decap_8 FILLER_73_1052 ();
 sg13g2_decap_8 FILLER_73_1059 ();
 sg13g2_decap_8 FILLER_73_1066 ();
 sg13g2_decap_8 FILLER_73_1073 ();
 sg13g2_decap_8 FILLER_73_1080 ();
 sg13g2_decap_8 FILLER_73_1087 ();
 sg13g2_decap_8 FILLER_73_1094 ();
 sg13g2_decap_8 FILLER_73_1101 ();
 sg13g2_decap_8 FILLER_73_1108 ();
 sg13g2_decap_8 FILLER_73_1115 ();
 sg13g2_decap_8 FILLER_73_1122 ();
 sg13g2_decap_8 FILLER_73_1129 ();
 sg13g2_decap_8 FILLER_73_1136 ();
 sg13g2_decap_8 FILLER_73_1143 ();
 sg13g2_decap_8 FILLER_73_1150 ();
 sg13g2_decap_8 FILLER_73_1157 ();
 sg13g2_decap_8 FILLER_73_1164 ();
 sg13g2_decap_8 FILLER_73_1171 ();
 sg13g2_decap_8 FILLER_73_1178 ();
 sg13g2_decap_8 FILLER_73_1185 ();
 sg13g2_decap_8 FILLER_73_1192 ();
 sg13g2_decap_8 FILLER_73_1199 ();
 sg13g2_decap_8 FILLER_73_1206 ();
 sg13g2_decap_8 FILLER_73_1213 ();
 sg13g2_decap_8 FILLER_73_1220 ();
 sg13g2_decap_8 FILLER_73_1227 ();
 sg13g2_decap_8 FILLER_73_1234 ();
 sg13g2_decap_8 FILLER_73_1241 ();
 sg13g2_decap_8 FILLER_73_1248 ();
 sg13g2_decap_8 FILLER_73_1255 ();
 sg13g2_decap_8 FILLER_73_1262 ();
 sg13g2_decap_8 FILLER_73_1269 ();
 sg13g2_decap_8 FILLER_73_1276 ();
 sg13g2_decap_8 FILLER_73_1283 ();
 sg13g2_decap_8 FILLER_73_1290 ();
 sg13g2_decap_8 FILLER_73_1297 ();
 sg13g2_decap_8 FILLER_73_1304 ();
 sg13g2_decap_4 FILLER_73_1311 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_2 ();
 sg13g2_fill_1 FILLER_74_42 ();
 sg13g2_fill_1 FILLER_74_56 ();
 sg13g2_fill_2 FILLER_74_62 ();
 sg13g2_fill_1 FILLER_74_64 ();
 sg13g2_fill_1 FILLER_74_115 ();
 sg13g2_fill_2 FILLER_74_135 ();
 sg13g2_decap_8 FILLER_74_153 ();
 sg13g2_decap_8 FILLER_74_160 ();
 sg13g2_decap_8 FILLER_74_167 ();
 sg13g2_fill_2 FILLER_74_174 ();
 sg13g2_fill_2 FILLER_74_202 ();
 sg13g2_fill_2 FILLER_74_208 ();
 sg13g2_fill_1 FILLER_74_229 ();
 sg13g2_decap_4 FILLER_74_243 ();
 sg13g2_fill_1 FILLER_74_247 ();
 sg13g2_decap_8 FILLER_74_274 ();
 sg13g2_fill_2 FILLER_74_281 ();
 sg13g2_fill_2 FILLER_74_313 ();
 sg13g2_fill_2 FILLER_74_341 ();
 sg13g2_fill_2 FILLER_74_376 ();
 sg13g2_fill_1 FILLER_74_378 ();
 sg13g2_fill_2 FILLER_74_426 ();
 sg13g2_fill_1 FILLER_74_428 ();
 sg13g2_fill_2 FILLER_74_434 ();
 sg13g2_fill_1 FILLER_74_436 ();
 sg13g2_fill_2 FILLER_74_488 ();
 sg13g2_decap_8 FILLER_74_516 ();
 sg13g2_decap_4 FILLER_74_523 ();
 sg13g2_fill_1 FILLER_74_527 ();
 sg13g2_decap_8 FILLER_74_532 ();
 sg13g2_decap_4 FILLER_74_539 ();
 sg13g2_fill_2 FILLER_74_543 ();
 sg13g2_fill_1 FILLER_74_576 ();
 sg13g2_fill_1 FILLER_74_608 ();
 sg13g2_decap_4 FILLER_74_629 ();
 sg13g2_fill_1 FILLER_74_633 ();
 sg13g2_fill_2 FILLER_74_660 ();
 sg13g2_fill_1 FILLER_74_676 ();
 sg13g2_fill_1 FILLER_74_760 ();
 sg13g2_fill_1 FILLER_74_840 ();
 sg13g2_decap_4 FILLER_74_853 ();
 sg13g2_fill_1 FILLER_74_857 ();
 sg13g2_fill_2 FILLER_74_875 ();
 sg13g2_fill_1 FILLER_74_877 ();
 sg13g2_fill_1 FILLER_74_922 ();
 sg13g2_fill_1 FILLER_74_935 ();
 sg13g2_decap_8 FILLER_74_1049 ();
 sg13g2_decap_8 FILLER_74_1056 ();
 sg13g2_decap_8 FILLER_74_1063 ();
 sg13g2_decap_8 FILLER_74_1070 ();
 sg13g2_decap_8 FILLER_74_1077 ();
 sg13g2_decap_8 FILLER_74_1084 ();
 sg13g2_decap_8 FILLER_74_1091 ();
 sg13g2_decap_8 FILLER_74_1098 ();
 sg13g2_decap_8 FILLER_74_1105 ();
 sg13g2_decap_8 FILLER_74_1112 ();
 sg13g2_decap_8 FILLER_74_1119 ();
 sg13g2_decap_8 FILLER_74_1126 ();
 sg13g2_decap_8 FILLER_74_1133 ();
 sg13g2_decap_8 FILLER_74_1140 ();
 sg13g2_decap_8 FILLER_74_1147 ();
 sg13g2_decap_8 FILLER_74_1154 ();
 sg13g2_decap_8 FILLER_74_1161 ();
 sg13g2_decap_8 FILLER_74_1168 ();
 sg13g2_decap_8 FILLER_74_1175 ();
 sg13g2_decap_8 FILLER_74_1182 ();
 sg13g2_decap_8 FILLER_74_1189 ();
 sg13g2_decap_8 FILLER_74_1196 ();
 sg13g2_decap_8 FILLER_74_1203 ();
 sg13g2_decap_8 FILLER_74_1210 ();
 sg13g2_decap_8 FILLER_74_1217 ();
 sg13g2_decap_8 FILLER_74_1224 ();
 sg13g2_decap_8 FILLER_74_1231 ();
 sg13g2_decap_8 FILLER_74_1238 ();
 sg13g2_decap_8 FILLER_74_1245 ();
 sg13g2_decap_8 FILLER_74_1252 ();
 sg13g2_decap_8 FILLER_74_1259 ();
 sg13g2_decap_8 FILLER_74_1266 ();
 sg13g2_decap_8 FILLER_74_1273 ();
 sg13g2_decap_8 FILLER_74_1280 ();
 sg13g2_decap_8 FILLER_74_1287 ();
 sg13g2_decap_8 FILLER_74_1294 ();
 sg13g2_decap_8 FILLER_74_1301 ();
 sg13g2_decap_8 FILLER_74_1308 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_7 ();
 sg13g2_fill_1 FILLER_75_9 ();
 sg13g2_fill_1 FILLER_75_49 ();
 sg13g2_fill_2 FILLER_75_59 ();
 sg13g2_fill_1 FILLER_75_66 ();
 sg13g2_fill_2 FILLER_75_107 ();
 sg13g2_decap_8 FILLER_75_149 ();
 sg13g2_decap_8 FILLER_75_156 ();
 sg13g2_fill_1 FILLER_75_163 ();
 sg13g2_decap_8 FILLER_75_169 ();
 sg13g2_decap_4 FILLER_75_176 ();
 sg13g2_fill_2 FILLER_75_180 ();
 sg13g2_fill_2 FILLER_75_208 ();
 sg13g2_decap_8 FILLER_75_251 ();
 sg13g2_fill_1 FILLER_75_258 ();
 sg13g2_fill_2 FILLER_75_263 ();
 sg13g2_fill_1 FILLER_75_342 ();
 sg13g2_fill_1 FILLER_75_352 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_decap_8 FILLER_75_372 ();
 sg13g2_fill_2 FILLER_75_387 ();
 sg13g2_fill_1 FILLER_75_389 ();
 sg13g2_fill_1 FILLER_75_394 ();
 sg13g2_decap_8 FILLER_75_413 ();
 sg13g2_fill_1 FILLER_75_420 ();
 sg13g2_fill_1 FILLER_75_426 ();
 sg13g2_fill_2 FILLER_75_478 ();
 sg13g2_fill_2 FILLER_75_489 ();
 sg13g2_fill_1 FILLER_75_491 ();
 sg13g2_decap_8 FILLER_75_549 ();
 sg13g2_fill_1 FILLER_75_556 ();
 sg13g2_fill_2 FILLER_75_587 ();
 sg13g2_fill_1 FILLER_75_626 ();
 sg13g2_decap_4 FILLER_75_653 ();
 sg13g2_fill_1 FILLER_75_742 ();
 sg13g2_decap_8 FILLER_75_762 ();
 sg13g2_fill_2 FILLER_75_818 ();
 sg13g2_fill_1 FILLER_75_945 ();
 sg13g2_fill_2 FILLER_75_1012 ();
 sg13g2_decap_8 FILLER_75_1044 ();
 sg13g2_decap_8 FILLER_75_1051 ();
 sg13g2_decap_8 FILLER_75_1058 ();
 sg13g2_decap_8 FILLER_75_1065 ();
 sg13g2_decap_8 FILLER_75_1072 ();
 sg13g2_decap_8 FILLER_75_1079 ();
 sg13g2_decap_8 FILLER_75_1086 ();
 sg13g2_decap_8 FILLER_75_1093 ();
 sg13g2_decap_8 FILLER_75_1100 ();
 sg13g2_decap_8 FILLER_75_1107 ();
 sg13g2_decap_8 FILLER_75_1114 ();
 sg13g2_decap_8 FILLER_75_1121 ();
 sg13g2_decap_8 FILLER_75_1128 ();
 sg13g2_decap_8 FILLER_75_1135 ();
 sg13g2_decap_8 FILLER_75_1142 ();
 sg13g2_decap_8 FILLER_75_1149 ();
 sg13g2_decap_8 FILLER_75_1156 ();
 sg13g2_decap_8 FILLER_75_1163 ();
 sg13g2_decap_8 FILLER_75_1170 ();
 sg13g2_decap_8 FILLER_75_1177 ();
 sg13g2_decap_8 FILLER_75_1184 ();
 sg13g2_decap_8 FILLER_75_1191 ();
 sg13g2_decap_8 FILLER_75_1198 ();
 sg13g2_decap_8 FILLER_75_1205 ();
 sg13g2_decap_8 FILLER_75_1212 ();
 sg13g2_decap_8 FILLER_75_1219 ();
 sg13g2_decap_8 FILLER_75_1226 ();
 sg13g2_decap_8 FILLER_75_1233 ();
 sg13g2_decap_8 FILLER_75_1240 ();
 sg13g2_decap_8 FILLER_75_1247 ();
 sg13g2_decap_8 FILLER_75_1254 ();
 sg13g2_decap_8 FILLER_75_1261 ();
 sg13g2_decap_8 FILLER_75_1268 ();
 sg13g2_decap_8 FILLER_75_1275 ();
 sg13g2_decap_8 FILLER_75_1282 ();
 sg13g2_decap_8 FILLER_75_1289 ();
 sg13g2_decap_8 FILLER_75_1296 ();
 sg13g2_decap_8 FILLER_75_1303 ();
 sg13g2_decap_4 FILLER_75_1310 ();
 sg13g2_fill_1 FILLER_75_1314 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_41 ();
 sg13g2_fill_1 FILLER_76_57 ();
 sg13g2_fill_2 FILLER_76_99 ();
 sg13g2_fill_1 FILLER_76_115 ();
 sg13g2_decap_8 FILLER_76_149 ();
 sg13g2_decap_8 FILLER_76_156 ();
 sg13g2_decap_8 FILLER_76_163 ();
 sg13g2_decap_4 FILLER_76_170 ();
 sg13g2_fill_2 FILLER_76_209 ();
 sg13g2_fill_2 FILLER_76_285 ();
 sg13g2_fill_2 FILLER_76_309 ();
 sg13g2_fill_2 FILLER_76_334 ();
 sg13g2_decap_4 FILLER_76_362 ();
 sg13g2_decap_4 FILLER_76_384 ();
 sg13g2_fill_1 FILLER_76_388 ();
 sg13g2_fill_1 FILLER_76_419 ();
 sg13g2_fill_1 FILLER_76_446 ();
 sg13g2_fill_2 FILLER_76_451 ();
 sg13g2_fill_1 FILLER_76_457 ();
 sg13g2_fill_1 FILLER_76_505 ();
 sg13g2_decap_8 FILLER_76_510 ();
 sg13g2_fill_2 FILLER_76_517 ();
 sg13g2_fill_1 FILLER_76_519 ();
 sg13g2_fill_2 FILLER_76_528 ();
 sg13g2_fill_2 FILLER_76_535 ();
 sg13g2_fill_1 FILLER_76_537 ();
 sg13g2_decap_4 FILLER_76_571 ();
 sg13g2_fill_1 FILLER_76_580 ();
 sg13g2_fill_2 FILLER_76_587 ();
 sg13g2_fill_1 FILLER_76_612 ();
 sg13g2_decap_8 FILLER_76_627 ();
 sg13g2_decap_4 FILLER_76_634 ();
 sg13g2_fill_2 FILLER_76_646 ();
 sg13g2_fill_1 FILLER_76_665 ();
 sg13g2_fill_2 FILLER_76_682 ();
 sg13g2_fill_1 FILLER_76_697 ();
 sg13g2_fill_2 FILLER_76_724 ();
 sg13g2_fill_1 FILLER_76_755 ();
 sg13g2_fill_1 FILLER_76_779 ();
 sg13g2_decap_4 FILLER_76_784 ();
 sg13g2_fill_1 FILLER_76_788 ();
 sg13g2_fill_1 FILLER_76_863 ();
 sg13g2_decap_8 FILLER_76_867 ();
 sg13g2_fill_1 FILLER_76_964 ();
 sg13g2_fill_2 FILLER_76_1020 ();
 sg13g2_fill_1 FILLER_76_1022 ();
 sg13g2_decap_8 FILLER_76_1040 ();
 sg13g2_decap_8 FILLER_76_1047 ();
 sg13g2_decap_8 FILLER_76_1054 ();
 sg13g2_decap_8 FILLER_76_1061 ();
 sg13g2_decap_8 FILLER_76_1068 ();
 sg13g2_decap_8 FILLER_76_1075 ();
 sg13g2_decap_8 FILLER_76_1082 ();
 sg13g2_decap_8 FILLER_76_1089 ();
 sg13g2_decap_8 FILLER_76_1096 ();
 sg13g2_decap_8 FILLER_76_1103 ();
 sg13g2_decap_8 FILLER_76_1110 ();
 sg13g2_decap_8 FILLER_76_1117 ();
 sg13g2_decap_8 FILLER_76_1124 ();
 sg13g2_decap_8 FILLER_76_1131 ();
 sg13g2_decap_8 FILLER_76_1138 ();
 sg13g2_decap_8 FILLER_76_1145 ();
 sg13g2_decap_8 FILLER_76_1152 ();
 sg13g2_decap_8 FILLER_76_1159 ();
 sg13g2_decap_8 FILLER_76_1166 ();
 sg13g2_decap_8 FILLER_76_1173 ();
 sg13g2_decap_8 FILLER_76_1180 ();
 sg13g2_decap_8 FILLER_76_1187 ();
 sg13g2_decap_8 FILLER_76_1194 ();
 sg13g2_decap_8 FILLER_76_1201 ();
 sg13g2_decap_8 FILLER_76_1208 ();
 sg13g2_decap_8 FILLER_76_1215 ();
 sg13g2_decap_8 FILLER_76_1222 ();
 sg13g2_decap_8 FILLER_76_1229 ();
 sg13g2_decap_8 FILLER_76_1236 ();
 sg13g2_decap_8 FILLER_76_1243 ();
 sg13g2_decap_8 FILLER_76_1250 ();
 sg13g2_decap_8 FILLER_76_1257 ();
 sg13g2_decap_8 FILLER_76_1264 ();
 sg13g2_decap_8 FILLER_76_1271 ();
 sg13g2_decap_8 FILLER_76_1278 ();
 sg13g2_decap_8 FILLER_76_1285 ();
 sg13g2_decap_8 FILLER_76_1292 ();
 sg13g2_decap_8 FILLER_76_1299 ();
 sg13g2_decap_8 FILLER_76_1306 ();
 sg13g2_fill_2 FILLER_76_1313 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_14 ();
 sg13g2_fill_1 FILLER_77_16 ();
 sg13g2_fill_1 FILLER_77_52 ();
 sg13g2_fill_2 FILLER_77_58 ();
 sg13g2_fill_2 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_152 ();
 sg13g2_decap_8 FILLER_77_159 ();
 sg13g2_decap_8 FILLER_77_166 ();
 sg13g2_decap_8 FILLER_77_173 ();
 sg13g2_decap_4 FILLER_77_180 ();
 sg13g2_fill_1 FILLER_77_184 ();
 sg13g2_fill_2 FILLER_77_189 ();
 sg13g2_fill_1 FILLER_77_221 ();
 sg13g2_fill_1 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_250 ();
 sg13g2_fill_2 FILLER_77_257 ();
 sg13g2_fill_1 FILLER_77_259 ();
 sg13g2_decap_4 FILLER_77_278 ();
 sg13g2_fill_2 FILLER_77_282 ();
 sg13g2_decap_8 FILLER_77_289 ();
 sg13g2_fill_1 FILLER_77_296 ();
 sg13g2_fill_2 FILLER_77_328 ();
 sg13g2_fill_1 FILLER_77_330 ();
 sg13g2_fill_2 FILLER_77_348 ();
 sg13g2_fill_1 FILLER_77_398 ();
 sg13g2_fill_2 FILLER_77_434 ();
 sg13g2_fill_2 FILLER_77_450 ();
 sg13g2_fill_2 FILLER_77_457 ();
 sg13g2_fill_2 FILLER_77_482 ();
 sg13g2_fill_1 FILLER_77_484 ();
 sg13g2_decap_4 FILLER_77_498 ();
 sg13g2_fill_2 FILLER_77_502 ();
 sg13g2_fill_1 FILLER_77_560 ();
 sg13g2_fill_2 FILLER_77_593 ();
 sg13g2_fill_1 FILLER_77_595 ();
 sg13g2_fill_2 FILLER_77_623 ();
 sg13g2_fill_1 FILLER_77_625 ();
 sg13g2_fill_2 FILLER_77_652 ();
 sg13g2_fill_2 FILLER_77_711 ();
 sg13g2_fill_1 FILLER_77_713 ();
 sg13g2_fill_2 FILLER_77_800 ();
 sg13g2_fill_1 FILLER_77_807 ();
 sg13g2_fill_2 FILLER_77_822 ();
 sg13g2_fill_1 FILLER_77_829 ();
 sg13g2_fill_1 FILLER_77_887 ();
 sg13g2_fill_1 FILLER_77_949 ();
 sg13g2_decap_8 FILLER_77_1040 ();
 sg13g2_decap_8 FILLER_77_1047 ();
 sg13g2_decap_8 FILLER_77_1054 ();
 sg13g2_decap_8 FILLER_77_1061 ();
 sg13g2_decap_8 FILLER_77_1068 ();
 sg13g2_decap_8 FILLER_77_1075 ();
 sg13g2_decap_8 FILLER_77_1082 ();
 sg13g2_decap_8 FILLER_77_1089 ();
 sg13g2_decap_8 FILLER_77_1096 ();
 sg13g2_decap_8 FILLER_77_1103 ();
 sg13g2_decap_8 FILLER_77_1110 ();
 sg13g2_decap_8 FILLER_77_1117 ();
 sg13g2_decap_8 FILLER_77_1124 ();
 sg13g2_decap_8 FILLER_77_1131 ();
 sg13g2_decap_8 FILLER_77_1138 ();
 sg13g2_decap_8 FILLER_77_1145 ();
 sg13g2_decap_8 FILLER_77_1152 ();
 sg13g2_decap_8 FILLER_77_1159 ();
 sg13g2_decap_8 FILLER_77_1166 ();
 sg13g2_decap_8 FILLER_77_1173 ();
 sg13g2_decap_8 FILLER_77_1180 ();
 sg13g2_decap_8 FILLER_77_1187 ();
 sg13g2_decap_8 FILLER_77_1194 ();
 sg13g2_decap_8 FILLER_77_1201 ();
 sg13g2_decap_8 FILLER_77_1208 ();
 sg13g2_decap_8 FILLER_77_1215 ();
 sg13g2_decap_8 FILLER_77_1222 ();
 sg13g2_decap_8 FILLER_77_1229 ();
 sg13g2_decap_8 FILLER_77_1236 ();
 sg13g2_decap_8 FILLER_77_1243 ();
 sg13g2_decap_8 FILLER_77_1250 ();
 sg13g2_decap_8 FILLER_77_1257 ();
 sg13g2_decap_8 FILLER_77_1264 ();
 sg13g2_decap_8 FILLER_77_1271 ();
 sg13g2_decap_8 FILLER_77_1278 ();
 sg13g2_decap_8 FILLER_77_1285 ();
 sg13g2_decap_8 FILLER_77_1292 ();
 sg13g2_decap_8 FILLER_77_1299 ();
 sg13g2_decap_8 FILLER_77_1306 ();
 sg13g2_fill_2 FILLER_77_1313 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_fill_2 FILLER_78_32 ();
 sg13g2_fill_1 FILLER_78_114 ();
 sg13g2_decap_8 FILLER_78_151 ();
 sg13g2_decap_8 FILLER_78_158 ();
 sg13g2_decap_8 FILLER_78_165 ();
 sg13g2_fill_2 FILLER_78_236 ();
 sg13g2_decap_8 FILLER_78_264 ();
 sg13g2_decap_4 FILLER_78_271 ();
 sg13g2_fill_2 FILLER_78_275 ();
 sg13g2_decap_8 FILLER_78_306 ();
 sg13g2_fill_2 FILLER_78_313 ();
 sg13g2_fill_2 FILLER_78_341 ();
 sg13g2_fill_1 FILLER_78_343 ();
 sg13g2_decap_4 FILLER_78_375 ();
 sg13g2_fill_1 FILLER_78_405 ();
 sg13g2_decap_8 FILLER_78_521 ();
 sg13g2_decap_8 FILLER_78_528 ();
 sg13g2_decap_8 FILLER_78_535 ();
 sg13g2_fill_2 FILLER_78_542 ();
 sg13g2_fill_1 FILLER_78_544 ();
 sg13g2_decap_8 FILLER_78_549 ();
 sg13g2_fill_2 FILLER_78_564 ();
 sg13g2_fill_1 FILLER_78_566 ();
 sg13g2_fill_2 FILLER_78_629 ();
 sg13g2_fill_1 FILLER_78_631 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_fill_1 FILLER_78_677 ();
 sg13g2_fill_1 FILLER_78_709 ();
 sg13g2_fill_2 FILLER_78_719 ();
 sg13g2_fill_2 FILLER_78_753 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_decap_4 FILLER_78_862 ();
 sg13g2_fill_1 FILLER_78_866 ();
 sg13g2_fill_2 FILLER_78_875 ();
 sg13g2_fill_1 FILLER_78_877 ();
 sg13g2_fill_1 FILLER_78_907 ();
 sg13g2_fill_1 FILLER_78_943 ();
 sg13g2_fill_2 FILLER_78_984 ();
 sg13g2_decap_8 FILLER_78_1022 ();
 sg13g2_decap_8 FILLER_78_1029 ();
 sg13g2_decap_8 FILLER_78_1036 ();
 sg13g2_decap_8 FILLER_78_1043 ();
 sg13g2_decap_8 FILLER_78_1050 ();
 sg13g2_decap_8 FILLER_78_1057 ();
 sg13g2_decap_8 FILLER_78_1064 ();
 sg13g2_decap_8 FILLER_78_1071 ();
 sg13g2_decap_8 FILLER_78_1078 ();
 sg13g2_decap_8 FILLER_78_1085 ();
 sg13g2_decap_8 FILLER_78_1092 ();
 sg13g2_decap_8 FILLER_78_1099 ();
 sg13g2_decap_8 FILLER_78_1106 ();
 sg13g2_decap_8 FILLER_78_1113 ();
 sg13g2_decap_8 FILLER_78_1120 ();
 sg13g2_decap_8 FILLER_78_1127 ();
 sg13g2_decap_8 FILLER_78_1134 ();
 sg13g2_decap_8 FILLER_78_1141 ();
 sg13g2_decap_8 FILLER_78_1148 ();
 sg13g2_decap_8 FILLER_78_1155 ();
 sg13g2_decap_8 FILLER_78_1162 ();
 sg13g2_decap_8 FILLER_78_1169 ();
 sg13g2_decap_8 FILLER_78_1176 ();
 sg13g2_decap_8 FILLER_78_1183 ();
 sg13g2_decap_8 FILLER_78_1190 ();
 sg13g2_decap_8 FILLER_78_1197 ();
 sg13g2_decap_8 FILLER_78_1204 ();
 sg13g2_decap_8 FILLER_78_1211 ();
 sg13g2_decap_8 FILLER_78_1218 ();
 sg13g2_decap_8 FILLER_78_1225 ();
 sg13g2_decap_8 FILLER_78_1232 ();
 sg13g2_decap_8 FILLER_78_1239 ();
 sg13g2_decap_8 FILLER_78_1246 ();
 sg13g2_decap_8 FILLER_78_1253 ();
 sg13g2_decap_8 FILLER_78_1260 ();
 sg13g2_decap_8 FILLER_78_1267 ();
 sg13g2_decap_8 FILLER_78_1274 ();
 sg13g2_decap_8 FILLER_78_1281 ();
 sg13g2_decap_8 FILLER_78_1288 ();
 sg13g2_decap_8 FILLER_78_1295 ();
 sg13g2_decap_8 FILLER_78_1302 ();
 sg13g2_decap_4 FILLER_78_1309 ();
 sg13g2_fill_2 FILLER_78_1313 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_fill_2 FILLER_79_35 ();
 sg13g2_fill_1 FILLER_79_92 ();
 sg13g2_fill_1 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_155 ();
 sg13g2_decap_8 FILLER_79_162 ();
 sg13g2_decap_8 FILLER_79_169 ();
 sg13g2_decap_8 FILLER_79_176 ();
 sg13g2_fill_2 FILLER_79_187 ();
 sg13g2_fill_1 FILLER_79_220 ();
 sg13g2_decap_8 FILLER_79_236 ();
 sg13g2_decap_4 FILLER_79_243 ();
 sg13g2_fill_2 FILLER_79_247 ();
 sg13g2_decap_8 FILLER_79_253 ();
 sg13g2_decap_8 FILLER_79_260 ();
 sg13g2_decap_8 FILLER_79_267 ();
 sg13g2_decap_8 FILLER_79_274 ();
 sg13g2_fill_2 FILLER_79_281 ();
 sg13g2_fill_2 FILLER_79_288 ();
 sg13g2_fill_1 FILLER_79_290 ();
 sg13g2_decap_8 FILLER_79_295 ();
 sg13g2_decap_8 FILLER_79_302 ();
 sg13g2_decap_8 FILLER_79_309 ();
 sg13g2_decap_8 FILLER_79_316 ();
 sg13g2_fill_2 FILLER_79_323 ();
 sg13g2_fill_2 FILLER_79_329 ();
 sg13g2_fill_1 FILLER_79_335 ();
 sg13g2_decap_8 FILLER_79_340 ();
 sg13g2_fill_1 FILLER_79_351 ();
 sg13g2_decap_8 FILLER_79_369 ();
 sg13g2_decap_4 FILLER_79_376 ();
 sg13g2_fill_2 FILLER_79_380 ();
 sg13g2_fill_2 FILLER_79_450 ();
 sg13g2_fill_1 FILLER_79_452 ();
 sg13g2_decap_4 FILLER_79_478 ();
 sg13g2_fill_2 FILLER_79_495 ();
 sg13g2_decap_8 FILLER_79_505 ();
 sg13g2_fill_2 FILLER_79_512 ();
 sg13g2_fill_1 FILLER_79_514 ();
 sg13g2_fill_1 FILLER_79_572 ();
 sg13g2_fill_2 FILLER_79_607 ();
 sg13g2_decap_8 FILLER_79_652 ();
 sg13g2_decap_4 FILLER_79_659 ();
 sg13g2_fill_2 FILLER_79_667 ();
 sg13g2_fill_2 FILLER_79_826 ();
 sg13g2_fill_2 FILLER_79_842 ();
 sg13g2_fill_2 FILLER_79_875 ();
 sg13g2_fill_1 FILLER_79_877 ();
 sg13g2_fill_2 FILLER_79_944 ();
 sg13g2_fill_2 FILLER_79_977 ();
 sg13g2_decap_8 FILLER_79_1014 ();
 sg13g2_decap_8 FILLER_79_1021 ();
 sg13g2_decap_8 FILLER_79_1028 ();
 sg13g2_decap_8 FILLER_79_1035 ();
 sg13g2_decap_8 FILLER_79_1042 ();
 sg13g2_decap_8 FILLER_79_1049 ();
 sg13g2_decap_8 FILLER_79_1056 ();
 sg13g2_decap_8 FILLER_79_1063 ();
 sg13g2_decap_8 FILLER_79_1070 ();
 sg13g2_decap_8 FILLER_79_1077 ();
 sg13g2_decap_8 FILLER_79_1084 ();
 sg13g2_decap_8 FILLER_79_1091 ();
 sg13g2_decap_8 FILLER_79_1098 ();
 sg13g2_decap_8 FILLER_79_1105 ();
 sg13g2_decap_8 FILLER_79_1112 ();
 sg13g2_decap_8 FILLER_79_1119 ();
 sg13g2_decap_8 FILLER_79_1126 ();
 sg13g2_decap_8 FILLER_79_1133 ();
 sg13g2_decap_8 FILLER_79_1140 ();
 sg13g2_decap_8 FILLER_79_1147 ();
 sg13g2_decap_8 FILLER_79_1154 ();
 sg13g2_decap_8 FILLER_79_1161 ();
 sg13g2_decap_8 FILLER_79_1168 ();
 sg13g2_decap_8 FILLER_79_1175 ();
 sg13g2_decap_8 FILLER_79_1182 ();
 sg13g2_decap_8 FILLER_79_1189 ();
 sg13g2_decap_8 FILLER_79_1196 ();
 sg13g2_decap_8 FILLER_79_1203 ();
 sg13g2_decap_8 FILLER_79_1210 ();
 sg13g2_decap_8 FILLER_79_1217 ();
 sg13g2_decap_8 FILLER_79_1224 ();
 sg13g2_decap_8 FILLER_79_1231 ();
 sg13g2_decap_8 FILLER_79_1238 ();
 sg13g2_decap_8 FILLER_79_1245 ();
 sg13g2_decap_8 FILLER_79_1252 ();
 sg13g2_decap_8 FILLER_79_1259 ();
 sg13g2_decap_8 FILLER_79_1266 ();
 sg13g2_decap_8 FILLER_79_1273 ();
 sg13g2_decap_8 FILLER_79_1280 ();
 sg13g2_decap_8 FILLER_79_1287 ();
 sg13g2_decap_8 FILLER_79_1294 ();
 sg13g2_decap_8 FILLER_79_1301 ();
 sg13g2_decap_8 FILLER_79_1308 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_fill_1 FILLER_80_98 ();
 sg13g2_fill_2 FILLER_80_111 ();
 sg13g2_fill_1 FILLER_80_135 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_4 FILLER_80_194 ();
 sg13g2_decap_4 FILLER_80_214 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_decap_8 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_decap_8 FILLER_80_249 ();
 sg13g2_decap_8 FILLER_80_256 ();
 sg13g2_decap_8 FILLER_80_263 ();
 sg13g2_decap_8 FILLER_80_270 ();
 sg13g2_decap_8 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_284 ();
 sg13g2_decap_8 FILLER_80_291 ();
 sg13g2_decap_8 FILLER_80_298 ();
 sg13g2_decap_8 FILLER_80_305 ();
 sg13g2_decap_8 FILLER_80_312 ();
 sg13g2_decap_8 FILLER_80_319 ();
 sg13g2_decap_8 FILLER_80_326 ();
 sg13g2_decap_8 FILLER_80_333 ();
 sg13g2_decap_8 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_347 ();
 sg13g2_decap_4 FILLER_80_354 ();
 sg13g2_fill_2 FILLER_80_358 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_fill_1 FILLER_80_379 ();
 sg13g2_fill_1 FILLER_80_423 ();
 sg13g2_fill_2 FILLER_80_485 ();
 sg13g2_decap_8 FILLER_80_513 ();
 sg13g2_decap_8 FILLER_80_520 ();
 sg13g2_decap_8 FILLER_80_527 ();
 sg13g2_fill_1 FILLER_80_534 ();
 sg13g2_decap_8 FILLER_80_539 ();
 sg13g2_decap_8 FILLER_80_546 ();
 sg13g2_decap_8 FILLER_80_553 ();
 sg13g2_decap_8 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_567 ();
 sg13g2_decap_8 FILLER_80_574 ();
 sg13g2_fill_2 FILLER_80_581 ();
 sg13g2_fill_2 FILLER_80_587 ();
 sg13g2_fill_1 FILLER_80_589 ();
 sg13g2_fill_1 FILLER_80_608 ();
 sg13g2_decap_8 FILLER_80_613 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_631 ();
 sg13g2_decap_8 FILLER_80_678 ();
 sg13g2_decap_8 FILLER_80_689 ();
 sg13g2_fill_2 FILLER_80_731 ();
 sg13g2_fill_2 FILLER_80_751 ();
 sg13g2_fill_1 FILLER_80_784 ();
 sg13g2_fill_2 FILLER_80_799 ();
 sg13g2_fill_1 FILLER_80_801 ();
 sg13g2_decap_8 FILLER_80_836 ();
 sg13g2_decap_8 FILLER_80_843 ();
 sg13g2_decap_4 FILLER_80_850 ();
 sg13g2_fill_1 FILLER_80_854 ();
 sg13g2_decap_8 FILLER_80_859 ();
 sg13g2_decap_8 FILLER_80_866 ();
 sg13g2_fill_1 FILLER_80_873 ();
 sg13g2_fill_2 FILLER_80_976 ();
 sg13g2_fill_1 FILLER_80_978 ();
 sg13g2_decap_8 FILLER_80_1023 ();
 sg13g2_decap_8 FILLER_80_1030 ();
 sg13g2_decap_8 FILLER_80_1037 ();
 sg13g2_decap_8 FILLER_80_1044 ();
 sg13g2_decap_8 FILLER_80_1051 ();
 sg13g2_decap_8 FILLER_80_1058 ();
 sg13g2_decap_8 FILLER_80_1065 ();
 sg13g2_decap_8 FILLER_80_1072 ();
 sg13g2_decap_8 FILLER_80_1079 ();
 sg13g2_decap_8 FILLER_80_1086 ();
 sg13g2_decap_8 FILLER_80_1093 ();
 sg13g2_decap_8 FILLER_80_1100 ();
 sg13g2_decap_8 FILLER_80_1107 ();
 sg13g2_decap_8 FILLER_80_1114 ();
 sg13g2_decap_8 FILLER_80_1121 ();
 sg13g2_decap_8 FILLER_80_1128 ();
 sg13g2_decap_8 FILLER_80_1135 ();
 sg13g2_decap_8 FILLER_80_1142 ();
 sg13g2_decap_8 FILLER_80_1149 ();
 sg13g2_decap_8 FILLER_80_1156 ();
 sg13g2_decap_8 FILLER_80_1163 ();
 sg13g2_decap_8 FILLER_80_1170 ();
 sg13g2_decap_8 FILLER_80_1177 ();
 sg13g2_decap_8 FILLER_80_1184 ();
 sg13g2_decap_8 FILLER_80_1191 ();
 sg13g2_decap_8 FILLER_80_1198 ();
 sg13g2_decap_8 FILLER_80_1205 ();
 sg13g2_decap_8 FILLER_80_1212 ();
 sg13g2_decap_8 FILLER_80_1219 ();
 sg13g2_decap_8 FILLER_80_1226 ();
 sg13g2_decap_8 FILLER_80_1233 ();
 sg13g2_decap_8 FILLER_80_1240 ();
 sg13g2_decap_8 FILLER_80_1247 ();
 sg13g2_decap_8 FILLER_80_1254 ();
 sg13g2_decap_8 FILLER_80_1261 ();
 sg13g2_decap_8 FILLER_80_1268 ();
 sg13g2_decap_8 FILLER_80_1275 ();
 sg13g2_decap_8 FILLER_80_1282 ();
 sg13g2_decap_8 FILLER_80_1289 ();
 sg13g2_decap_8 FILLER_80_1296 ();
 sg13g2_decap_8 FILLER_80_1303 ();
 sg13g2_decap_4 FILLER_80_1310 ();
 sg13g2_fill_1 FILLER_80_1314 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule

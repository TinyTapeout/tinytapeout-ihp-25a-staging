module tt_um_wokwi_group_6 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire \proj_10.net10 ;
 wire \proj_10.net11 ;
 wire \proj_10.net17 ;
 wire \proj_10.net18 ;
 wire \proj_10.net19 ;
 wire \proj_10.net20 ;
 wire \proj_10.net21 ;
 wire \proj_10.net22 ;
 wire \proj_10.net23 ;
 wire \proj_10.net24 ;
 wire \proj_10.net25 ;
 wire \proj_10.net26 ;
 wire \proj_10.net27 ;
 wire \proj_10.net8 ;
 wire \proj_10.net9 ;
 wire \proj_11.net15 ;
 wire \proj_11.net16 ;
 wire \proj_11.net17 ;
 wire \proj_11.net18 ;
 wire \proj_11.net19 ;
 wire \proj_11.net20 ;
 wire \proj_11.net6 ;
 wire \proj_11.net7 ;
 wire \proj_11.net8 ;
 wire \proj_11.net9 ;
 wire \proj_12.net15 ;
 wire \proj_12.net16 ;
 wire \proj_12.net17 ;
 wire \proj_12.net18 ;
 wire \proj_12.net19 ;
 wire \proj_12.net20 ;
 wire \proj_12.net21 ;
 wire \proj_12.net22 ;
 wire \proj_12.net23 ;
 wire \proj_12.net24 ;
 wire \proj_12.net25 ;
 wire \proj_12.net26 ;
 wire \proj_12.net27 ;
 wire \proj_12.net28 ;
 wire \proj_12.net29 ;
 wire \proj_12.net30 ;
 wire \proj_12.net31 ;
 wire \proj_12.net32 ;
 wire \proj_12.net33 ;
 wire \proj_12.net6 ;
 wire \proj_12.net7 ;
 wire \proj_12.net8 ;
 wire \proj_12.net9 ;
 wire \proj_13.net10 ;
 wire \proj_13.net100 ;
 wire \proj_13.net101 ;
 wire \proj_13.net102 ;
 wire \proj_13.net103 ;
 wire \proj_13.net104 ;
 wire \proj_13.net105 ;
 wire \proj_13.net106 ;
 wire \proj_13.net107 ;
 wire \proj_13.net108 ;
 wire \proj_13.net109 ;
 wire \proj_13.net110 ;
 wire \proj_13.net111 ;
 wire \proj_13.net112 ;
 wire \proj_13.net113 ;
 wire \proj_13.net114 ;
 wire \proj_13.net115 ;
 wire \proj_13.net116 ;
 wire \proj_13.net117 ;
 wire \proj_13.net118 ;
 wire \proj_13.net119 ;
 wire \proj_13.net120 ;
 wire \proj_13.net121 ;
 wire \proj_13.net122 ;
 wire \proj_13.net123 ;
 wire \proj_13.net124 ;
 wire \proj_13.net125 ;
 wire \proj_13.net126 ;
 wire \proj_13.net127 ;
 wire \proj_13.net128 ;
 wire \proj_13.net129 ;
 wire \proj_13.net130 ;
 wire \proj_13.net131 ;
 wire \proj_13.net132 ;
 wire \proj_13.net133 ;
 wire \proj_13.net134 ;
 wire \proj_13.net135 ;
 wire \proj_13.net136 ;
 wire \proj_13.net137 ;
 wire \proj_13.net138 ;
 wire \proj_13.net139 ;
 wire \proj_13.net140 ;
 wire \proj_13.net141 ;
 wire \proj_13.net142 ;
 wire \proj_13.net143 ;
 wire \proj_13.net144 ;
 wire \proj_13.net145 ;
 wire \proj_13.net146 ;
 wire \proj_13.net147 ;
 wire \proj_13.net148 ;
 wire \proj_13.net149 ;
 wire \proj_13.net150 ;
 wire \proj_13.net151 ;
 wire \proj_13.net152 ;
 wire \proj_13.net153 ;
 wire \proj_13.net154 ;
 wire \proj_13.net155 ;
 wire \proj_13.net156 ;
 wire \proj_13.net157 ;
 wire \proj_13.net158 ;
 wire \proj_13.net159 ;
 wire \proj_13.net16 ;
 wire \proj_13.net160 ;
 wire \proj_13.net161 ;
 wire \proj_13.net162 ;
 wire \proj_13.net163 ;
 wire \proj_13.net164 ;
 wire \proj_13.net165 ;
 wire \proj_13.net166 ;
 wire \proj_13.net167 ;
 wire \proj_13.net168 ;
 wire \proj_13.net169 ;
 wire \proj_13.net17 ;
 wire \proj_13.net170 ;
 wire \proj_13.net171 ;
 wire \proj_13.net172 ;
 wire \proj_13.net173 ;
 wire \proj_13.net174 ;
 wire \proj_13.net175 ;
 wire \proj_13.net176 ;
 wire \proj_13.net177 ;
 wire \proj_13.net178 ;
 wire \proj_13.net179 ;
 wire \proj_13.net18 ;
 wire \proj_13.net180 ;
 wire \proj_13.net181 ;
 wire \proj_13.net182 ;
 wire \proj_13.net183 ;
 wire \proj_13.net184 ;
 wire \proj_13.net185 ;
 wire \proj_13.net186 ;
 wire \proj_13.net187 ;
 wire \proj_13.net188 ;
 wire \proj_13.net189 ;
 wire \proj_13.net19 ;
 wire \proj_13.net190 ;
 wire \proj_13.net191 ;
 wire \proj_13.net192 ;
 wire \proj_13.net193 ;
 wire \proj_13.net194 ;
 wire \proj_13.net195 ;
 wire \proj_13.net196 ;
 wire \proj_13.net197 ;
 wire \proj_13.net198 ;
 wire \proj_13.net199 ;
 wire \proj_13.net20 ;
 wire \proj_13.net200 ;
 wire \proj_13.net201 ;
 wire \proj_13.net202 ;
 wire \proj_13.net203 ;
 wire \proj_13.net204 ;
 wire \proj_13.net205 ;
 wire \proj_13.net206 ;
 wire \proj_13.net207 ;
 wire \proj_13.net208 ;
 wire \proj_13.net209 ;
 wire \proj_13.net21 ;
 wire \proj_13.net210 ;
 wire \proj_13.net211 ;
 wire \proj_13.net212 ;
 wire \proj_13.net213 ;
 wire \proj_13.net214 ;
 wire \proj_13.net215 ;
 wire \proj_13.net216 ;
 wire \proj_13.net217 ;
 wire \proj_13.net218 ;
 wire \proj_13.net22 ;
 wire \proj_13.net23 ;
 wire \proj_13.net24 ;
 wire \proj_13.net25 ;
 wire \proj_13.net26 ;
 wire \proj_13.net27 ;
 wire \proj_13.net28 ;
 wire \proj_13.net29 ;
 wire \proj_13.net3 ;
 wire \proj_13.net30 ;
 wire \proj_13.net31 ;
 wire \proj_13.net32 ;
 wire \proj_13.net33 ;
 wire \proj_13.net34 ;
 wire \proj_13.net35 ;
 wire \proj_13.net36 ;
 wire \proj_13.net37 ;
 wire \proj_13.net38 ;
 wire \proj_13.net39 ;
 wire \proj_13.net4 ;
 wire \proj_13.net40 ;
 wire \proj_13.net41 ;
 wire \proj_13.net42 ;
 wire \proj_13.net43 ;
 wire \proj_13.net44 ;
 wire \proj_13.net45 ;
 wire \proj_13.net46 ;
 wire \proj_13.net47 ;
 wire \proj_13.net48 ;
 wire \proj_13.net49 ;
 wire \proj_13.net5 ;
 wire \proj_13.net50 ;
 wire \proj_13.net51 ;
 wire \proj_13.net52 ;
 wire \proj_13.net53 ;
 wire \proj_13.net54 ;
 wire \proj_13.net55 ;
 wire \proj_13.net56 ;
 wire \proj_13.net57 ;
 wire \proj_13.net58 ;
 wire \proj_13.net59 ;
 wire \proj_13.net6 ;
 wire \proj_13.net60 ;
 wire \proj_13.net61 ;
 wire \proj_13.net62 ;
 wire \proj_13.net63 ;
 wire \proj_13.net64 ;
 wire \proj_13.net65 ;
 wire \proj_13.net66 ;
 wire \proj_13.net67 ;
 wire \proj_13.net68 ;
 wire \proj_13.net69 ;
 wire \proj_13.net7 ;
 wire \proj_13.net70 ;
 wire \proj_13.net71 ;
 wire \proj_13.net72 ;
 wire \proj_13.net73 ;
 wire \proj_13.net74 ;
 wire \proj_13.net75 ;
 wire \proj_13.net76 ;
 wire \proj_13.net77 ;
 wire \proj_13.net78 ;
 wire \proj_13.net79 ;
 wire \proj_13.net8 ;
 wire \proj_13.net80 ;
 wire \proj_13.net81 ;
 wire \proj_13.net82 ;
 wire \proj_13.net83 ;
 wire \proj_13.net84 ;
 wire \proj_13.net85 ;
 wire \proj_13.net86 ;
 wire \proj_13.net87 ;
 wire \proj_13.net88 ;
 wire \proj_13.net89 ;
 wire \proj_13.net9 ;
 wire \proj_13.net90 ;
 wire \proj_13.net91 ;
 wire \proj_13.net92 ;
 wire \proj_13.net93 ;
 wire \proj_13.net94 ;
 wire \proj_13.net95 ;
 wire \proj_13.net96 ;
 wire \proj_13.net97 ;
 wire \proj_13.net98 ;
 wire \proj_13.net99 ;
 wire \proj_14.net10 ;
 wire \proj_14.net11 ;
 wire \proj_14.net12 ;
 wire \proj_14.net4 ;
 wire \proj_14.net5 ;
 wire \proj__0.net15 ;
 wire \proj__0.net16 ;
 wire \proj__0.net17 ;
 wire \proj__0.net18 ;
 wire \proj__0.net19 ;
 wire \proj__0.net20 ;
 wire \proj__0.net9 ;
 wire \proj__1.net10 ;
 wire \proj__1.net11 ;
 wire \proj__1.net12 ;
 wire \proj__1.net9 ;
 wire \proj__2.net4 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net14 ;
 wire \proj__4.net10 ;
 wire \proj__4.net9 ;
 wire \proj__5.net10 ;
 wire \proj__5.net11 ;
 wire \proj__5.net9 ;
 wire \proj__6.net11 ;
 wire \proj__6.net12 ;
 wire \proj__6.net13 ;
 wire \proj__6.net14 ;
 wire \proj__6.net16 ;
 wire \proj__6.net17 ;
 wire \proj__6.net18 ;
 wire \proj__6.net9 ;
 wire \proj__7.net10 ;
 wire \proj__7.net11 ;
 wire \proj__7.net12 ;
 wire \proj__7.net13 ;
 wire \proj__7.net14 ;
 wire \proj__8.net3 ;
 wire \proj__8.net4 ;
 wire \proj__8.net5 ;
 wire \proj__8.net6 ;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire \proj_12.flop1/q ;
 wire net29;
 wire \proj_12.flop10/q ;
 wire net30;
 wire \proj_12.flop11/q ;
 wire net31;
 wire \proj_12.flop12/q ;
 wire net32;
 wire \proj_12.flop13/q ;
 wire net33;
 wire \proj_12.flop14/q ;
 wire net34;
 wire \proj_12.flop15/q ;
 wire net35;
 wire \proj_12.flop16/q ;
 wire net36;
 wire \proj_12.flop2/q ;
 wire net49;
 wire \proj_12.flop3/q ;
 wire net50;
 wire \proj_12.flop4/q ;
 wire net51;
 wire \proj_12.flop5/q ;
 wire net52;
 wire \proj_12.flop6/q ;
 wire net53;
 wire \proj_12.flop7/q ;
 wire net54;
 wire \proj_12.flop8/q ;
 wire net55;
 wire \proj_12.flop9/q ;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire \proj__8.flop1/notq ;
 wire net155;
 wire \proj__8.flop2/notq ;
 wire net156;
 wire \proj__8.flop3/notq ;
 wire clk_regs;
 wire \proj__8.flop4/notq ;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_1_0__leaf_clk_regs;
 wire clknet_1_1__leaf_clk_regs;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;

 sg13g2_and2_2 _062_ (.A(_034_),
    .B(_036_),
    .X(_037_));
 sg13g2_nand2_2 _063_ (.Y(_038_),
    .A(net8),
    .B(net7));
 sg13g2_nand2b_2 _064_ (.Y(_039_),
    .B(net10),
    .A_N(net9));
 sg13g2_nor2_2 _065_ (.A(_038_),
    .B(_039_),
    .Y(_040_));
 sg13g2_nand2b_2 _066_ (.Y(_041_),
    .B(net7),
    .A_N(net8));
 sg13g2_nor2_1 _067_ (.A(_039_),
    .B(_041_),
    .Y(_042_));
 sg13g2_a22oi_1 _068_ (.Y(_043_),
    .B1(_042_),
    .B2(net38),
    .A2(_040_),
    .A1(\proj_11.net6 ));
 sg13g2_nor2b_1 _069_ (.A(net10),
    .B_N(net9),
    .Y(_044_));
 sg13g2_nand2b_2 _070_ (.Y(_045_),
    .B(net9),
    .A_N(net10));
 sg13g2_nand2_1 _071_ (.Y(_046_),
    .A(\proj__6.net9 ),
    .B(_044_));
 sg13g2_nand2_2 _072_ (.Y(_047_),
    .A(net9),
    .B(net10));
 sg13g2_o21ai_1 _073_ (.B1(_046_),
    .Y(_048_),
    .A1(_031_),
    .A2(_047_));
 sg13g2_nor2_2 _074_ (.A(_041_),
    .B(_045_),
    .Y(_049_));
 sg13g2_nor3_2 _075_ (.A(net9),
    .B(net10),
    .C(_038_),
    .Y(_050_));
 sg13g2_nor3_2 _076_ (.A(_030_),
    .B(net7),
    .C(_039_),
    .Y(_051_));
 sg13g2_a22oi_1 _077_ (.Y(_052_),
    .B1(_051_),
    .B2(\proj_10.net8 ),
    .A2(_050_),
    .A1(\proj__3.net11 ));
 sg13g2_nor3_2 _078_ (.A(net9),
    .B(net10),
    .C(_041_),
    .Y(_053_));
 sg13g2_nor2_2 _079_ (.A(_041_),
    .B(_047_),
    .Y(_054_));
 sg13g2_a22oi_1 _080_ (.Y(_055_),
    .B1(_054_),
    .B2(\proj_13.net3 ),
    .A2(_053_),
    .A1(\proj__1.net9 ));
 sg13g2_nor3_2 _081_ (.A(net8),
    .B(net7),
    .C(_039_),
    .Y(_056_));
 sg13g2_nor2_2 _082_ (.A(_038_),
    .B(_045_),
    .Y(_057_));
 sg13g2_a22oi_1 _083_ (.Y(_058_),
    .B1(_057_),
    .B2(net47),
    .A2(_048_),
    .A1(_033_));
 sg13g2_a22oi_1 _084_ (.Y(_059_),
    .B1(_056_),
    .B2(\proj__8.net3 ),
    .A2(_049_),
    .A1(\proj__5.net9 ));
 sg13g2_and3_1 _085_ (.X(_060_),
    .A(_052_),
    .B(_055_),
    .C(_059_));
 sg13g2_nand4_1 _086_ (.B(_043_),
    .C(_058_),
    .A(_037_),
    .Y(uo_out[0]),
    .D(_060_));
 sg13g2_a22oi_1 _087_ (.Y(_061_),
    .B1(_054_),
    .B2(\proj_13.net4 ),
    .A2(_040_),
    .A1(\proj_11.net7 ));
 sg13g2_a22oi_1 _088_ (.Y(_000_),
    .B1(_057_),
    .B2(net40),
    .A2(_053_),
    .A1(\proj__1.net10 ));
 sg13g2_a22oi_1 _089_ (.Y(_001_),
    .B1(_050_),
    .B2(\proj__3.net12 ),
    .A2(_049_),
    .A1(\proj__5.net9 ));
 sg13g2_a22oi_1 _090_ (.Y(_002_),
    .B1(_056_),
    .B2(\proj__8.net4 ),
    .A2(_051_),
    .A1(\proj_10.net9 ));
 sg13g2_a22oi_1 _091_ (.Y(_003_),
    .B1(_035_),
    .B2(\proj_12.net6 ),
    .A2(_033_),
    .A1(\proj_14.net5 ));
 sg13g2_or2_1 _092_ (.X(_004_),
    .B(_003_),
    .A(_047_));
 sg13g2_and4_1 _093_ (.A(_037_),
    .B(_001_),
    .C(_002_),
    .D(_004_),
    .X(_005_));
 sg13g2_nor3_2 _094_ (.A(net8),
    .B(net7),
    .C(_047_),
    .Y(_006_));
 sg13g2_nand3_1 _095_ (.B(_000_),
    .C(_005_),
    .A(_061_),
    .Y(uo_out[1]));
 sg13g2_nand3_1 _096_ (.B(_035_),
    .C(_044_),
    .A(\proj__4.net9 ),
    .Y(_007_));
 sg13g2_a22oi_1 _097_ (.Y(_008_),
    .B1(_054_),
    .B2(\proj_13.net5 ),
    .A2(_049_),
    .A1(\proj__5.net10 ));
 sg13g2_a22oi_1 _098_ (.Y(_009_),
    .B1(_057_),
    .B2(\proj__7.net10 ),
    .A2(_050_),
    .A1(\proj__3.net13 ));
 sg13g2_a22oi_1 _099_ (.Y(_010_),
    .B1(_056_),
    .B2(\proj__8.net5 ),
    .A2(_040_),
    .A1(\proj_11.net8 ));
 sg13g2_a22oi_1 _100_ (.Y(_011_),
    .B1(_053_),
    .B2(\proj__1.net11 ),
    .A2(_051_),
    .A1(\proj_10.net10 ));
 sg13g2_and4_1 _101_ (.A(_037_),
    .B(_008_),
    .C(_009_),
    .D(_011_),
    .X(_012_));
 sg13g2_nand3_1 _102_ (.B(_010_),
    .C(_012_),
    .A(_007_),
    .Y(uo_out[2]));
 sg13g2_nand3_1 _103_ (.B(_035_),
    .C(_044_),
    .A(\proj__4.net10 ),
    .Y(_013_));
 sg13g2_a22oi_1 _104_ (.Y(_014_),
    .B1(_049_),
    .B2(\proj__5.net11 ),
    .A2(_040_),
    .A1(\proj_11.net9 ));
 sg13g2_a22oi_1 _105_ (.Y(_015_),
    .B1(_054_),
    .B2(\proj_13.net6 ),
    .A2(_053_),
    .A1(\proj__1.net12 ));
 sg13g2_a22oi_1 _106_ (.Y(_016_),
    .B1(_051_),
    .B2(\proj_10.net11 ),
    .A2(_050_),
    .A1(\proj__3.net14 ));
 sg13g2_a22oi_1 _107_ (.Y(_017_),
    .B1(_057_),
    .B2(\proj__7.net11 ),
    .A2(_056_),
    .A1(\proj__8.net6 ));
 sg13g2_and4_1 _108_ (.A(_037_),
    .B(_015_),
    .C(_016_),
    .D(_017_),
    .X(_018_));
 sg13g2_nand3_1 _109_ (.B(_014_),
    .C(_018_),
    .A(_013_),
    .Y(uo_out[3]));
 sg13g2_nand2_1 _110_ (.Y(_019_),
    .A(net7),
    .B(_032_));
 sg13g2_o21ai_1 _111_ (.B1(_019_),
    .Y(_020_),
    .A1(net8),
    .A2(_045_));
 sg13g2_a22oi_1 _112_ (.Y(_021_),
    .B1(_020_),
    .B2(net37),
    .A2(_057_),
    .A1(net4));
 sg13g2_a22oi_1 _113_ (.Y(_022_),
    .B1(_006_),
    .B2(\proj_12.net7 ),
    .A2(_054_),
    .A1(\proj_13.net7 ));
 sg13g2_nand3_1 _114_ (.B(_021_),
    .C(_022_),
    .A(_037_),
    .Y(uo_out[4]));
 sg13g2_a22oi_1 _115_ (.Y(_023_),
    .B1(_020_),
    .B2(net4),
    .A2(_006_),
    .A1(\proj_12.net8 ));
 sg13g2_a22oi_1 _116_ (.Y(_024_),
    .B1(_057_),
    .B2(\proj__7.net12 ),
    .A2(_054_),
    .A1(\proj_13.net8 ));
 sg13g2_nand3_1 _117_ (.B(_023_),
    .C(_024_),
    .A(_037_),
    .Y(uo_out[5]));
 sg13g2_nand2_1 _118_ (.Y(_025_),
    .A(\proj__7.net13 ),
    .B(_057_));
 sg13g2_a22oi_1 _119_ (.Y(_026_),
    .B1(_020_),
    .B2(net5),
    .A2(_054_),
    .A1(\proj_13.net9 ));
 sg13g2_nand3_1 _120_ (.B(_025_),
    .C(_026_),
    .A(_037_),
    .Y(uo_out[6]));
 sg13g2_nand2_1 _121_ (.Y(_027_),
    .A(net6),
    .B(_020_));
 sg13g2_nand2_1 _122_ (.Y(_028_),
    .A(\proj_13.net10 ),
    .B(_054_));
 sg13g2_a22oi_1 _123_ (.Y(_029_),
    .B1(_006_),
    .B2(\proj_12.net9 ),
    .A2(_057_),
    .A1(\proj__7.net14 ));
 sg13g2_nand4_1 _124_ (.B(_027_),
    .C(_028_),
    .A(_034_),
    .Y(uo_out[7]),
    .D(_029_));
 sg13g2_inv_1 _125_ (.Y(_030_),
    .A(net8));
 sg13g2_inv_1 _126_ (.Y(_031_),
    .A(\proj_14.net4 ));
 sg13g2_nor2_1 _127_ (.A(net9),
    .B(net10),
    .Y(_032_));
 sg13g2_nor2b_1 _128_ (.A(net7),
    .B_N(net8),
    .Y(_033_));
 sg13g2_nand3_1 _129_ (.B(_032_),
    .C(_033_),
    .A(\proj__2.net4 ),
    .Y(_034_));
 sg13g2_nor2_2 _130_ (.A(net8),
    .B(net7),
    .Y(_035_));
 sg13g2_nand3_1 _131_ (.B(_032_),
    .C(_035_),
    .A(\proj__0.net9 ),
    .Y(_036_));
 sg13g2_tielo tt_um_wokwi_group_6_12 (.L_LO(net12));
 sg13g2_tielo tt_um_wokwi_group_6_13 (.L_LO(net13));
 sg13g2_tielo tt_um_wokwi_group_6_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wokwi_group_6_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_group_6_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_group_6_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_group_6_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_group_6_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_group_6_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_group_6_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_group_6_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_group_6_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_group_6_24 (.L_LO(net24));
 sg13g2_tielo tt_um_wokwi_group_6_25 (.L_LO(net25));
 sg13g2_tielo tt_um_wokwi_group_6_26 (.L_LO(net26));
 sg13g2_tiehi \proj_12.flop1/_1__27  (.L_HI(net27));
 sg13g2_and2_1 \proj_10.and1/_0_  (.A(net47),
    .B(net38),
    .X(\proj_10.net18 ));
 sg13g2_and2_1 \proj_10.and2/_0_  (.A(net5),
    .B(\proj_10.net17 ),
    .X(\proj_10.net19 ));
 sg13g2_and2_1 \proj_10.and3/_0_  (.A(net43),
    .B(net37),
    .X(\proj_10.net22 ));
 sg13g2_and2_1 \proj_10.and4/_0_  (.A(\proj_10.net20 ),
    .B(\proj_10.net21 ),
    .X(\proj_10.net23 ));
 sg13g2_and2_1 \proj_10.and5/_0_  (.A(net40),
    .B(net4),
    .X(\proj_10.net26 ));
 sg13g2_and2_1 \proj_10.and6/_0_  (.A(\proj_10.net24 ),
    .B(\proj_10.net25 ),
    .X(\proj_10.net27 ));
 sg13g2_or2_1 \proj_10.or1/_0_  (.X(\proj_10.net20 ),
    .B(\proj_10.net19 ),
    .A(\proj_10.net18 ));
 sg13g2_or2_1 \proj_10.or2/_0_  (.X(\proj_10.net24 ),
    .B(\proj_10.net22 ),
    .A(\proj_10.net23 ));
 sg13g2_or2_1 \proj_10.or3/_0_  (.X(\proj_10.net11 ),
    .B(\proj_10.net26 ),
    .A(\proj_10.net27 ));
 sg13g2_xor2_1 \proj_10.xor1/_0_  (.B(net47),
    .A(net39),
    .X(\proj_10.net17 ));
 sg13g2_xor2_1 \proj_10.xor2/_0_  (.B(\proj_10.net17 ),
    .A(net5),
    .X(\proj_10.net8 ));
 sg13g2_xor2_1 \proj_10.xor3/_0_  (.B(net42),
    .A(net37),
    .X(\proj_10.net21 ));
 sg13g2_xor2_1 \proj_10.xor4/_0_  (.B(\proj_10.net21 ),
    .A(\proj_10.net20 ),
    .X(\proj_10.net9 ));
 sg13g2_xor2_1 \proj_10.xor5/_0_  (.B(net40),
    .A(net4),
    .X(\proj_10.net25 ));
 sg13g2_xor2_1 \proj_10.xor6/_0_  (.B(\proj_10.net25 ),
    .A(\proj_10.net24 ),
    .X(\proj_10.net10 ));
 sg13g2_and2_1 \proj_11.and1/_0_  (.A(net39),
    .B(net43),
    .X(\proj_11.net16 ));
 sg13g2_and2_1 \proj_11.and2/_0_  (.A(net37),
    .B(net40),
    .X(\proj_11.net18 ));
 sg13g2_and2_1 \proj_11.and3/_0_  (.A(net47),
    .B(\proj_11.net15 ),
    .X(\proj_11.net19 ));
 sg13g2_and2_1 \proj_11.and4/_0_  (.A(\proj_11.net7 ),
    .B(\proj_11.net17 ),
    .X(\proj_11.net20 ));
 sg13g2_or2_1 \proj_11.or1/_0_  (.X(\proj_11.net8 ),
    .B(\proj_11.net20 ),
    .A(\proj_11.net18 ));
 sg13g2_or2_1 \proj_11.or2/_0_  (.X(\proj_11.net7 ),
    .B(\proj_11.net19 ),
    .A(\proj_11.net16 ));
 sg13g2_xor2_1 \proj_11.xor1/_0_  (.B(net42),
    .A(net39),
    .X(\proj_11.net15 ));
 sg13g2_xor2_1 \proj_11.xor2/_0_  (.B(net40),
    .A(net37),
    .X(\proj_11.net17 ));
 sg13g2_xor2_1 \proj_11.xor3/_0_  (.B(\proj_11.net15 ),
    .A(net48),
    .X(\proj_11.net6 ));
 sg13g2_xor2_1 \proj_11.xor4/_0_  (.B(\proj_11.net17 ),
    .A(\proj_11.net7 ),
    .X(\proj_11.net9 ));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net39),
    .B(net43),
    .X(\proj_12.net15 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(net41),
    .B(net47),
    .X(\proj_12.net17 ));
 sg13g2_and2_1 \proj_12.and3/_0_  (.A(\proj_12.net16 ),
    .B(\proj_12.net15 ),
    .X(\proj_12.net18 ));
 sg13g2_dfrbp_1 \proj_12.flop1/_1_  (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net27),
    .D(net158),
    .Q_N(\proj_12.net19 ),
    .Q(\proj_12.flop1/q ));
 sg13g2_tiehi \proj_12.flop10/_1__28  (.L_HI(net28));
 sg13g2_dfrbp_1 \proj_12.flop10/_1_  (.CLK(\proj_12.net27 ),
    .RESET_B(net28),
    .D(\proj_12.net28 ),
    .Q_N(\proj_12.net28 ),
    .Q(\proj_12.flop10/q ));
 sg13g2_tiehi \proj_12.flop11/_1__29  (.L_HI(net29));
 sg13g2_dfrbp_1 \proj_12.flop11/_1_  (.CLK(\proj_12.net28 ),
    .RESET_B(net29),
    .D(\proj_12.net29 ),
    .Q_N(\proj_12.net29 ),
    .Q(\proj_12.flop11/q ));
 sg13g2_tiehi \proj_12.flop12/_1__30  (.L_HI(net30));
 sg13g2_dfrbp_1 \proj_12.flop12/_1_  (.CLK(\proj_12.net29 ),
    .RESET_B(net30),
    .D(\proj_12.net30 ),
    .Q_N(\proj_12.net30 ),
    .Q(\proj_12.flop12/q ));
 sg13g2_tiehi \proj_12.flop13/_1__31  (.L_HI(net31));
 sg13g2_dfrbp_1 \proj_12.flop13/_1_  (.CLK(\proj_12.net30 ),
    .RESET_B(net31),
    .D(\proj_12.net31 ),
    .Q_N(\proj_12.net31 ),
    .Q(\proj_12.flop13/q ));
 sg13g2_tiehi \proj_12.flop14/_1__32  (.L_HI(net32));
 sg13g2_dfrbp_1 \proj_12.flop14/_1_  (.CLK(\proj_12.net31 ),
    .RESET_B(net32),
    .D(\proj_12.net32 ),
    .Q_N(\proj_12.net32 ),
    .Q(\proj_12.flop14/q ));
 sg13g2_tiehi \proj_12.flop15/_1__33  (.L_HI(net33));
 sg13g2_dfrbp_1 \proj_12.flop15/_1_  (.CLK(\proj_12.net32 ),
    .RESET_B(net33),
    .D(\proj_12.net33 ),
    .Q_N(\proj_12.net33 ),
    .Q(\proj_12.flop15/q ));
 sg13g2_tiehi \proj_12.flop16/_1__34  (.L_HI(net34));
 sg13g2_dfrbp_1 \proj_12.flop16/_1_  (.CLK(\proj_12.net33 ),
    .RESET_B(net34),
    .D(\proj_12.net9 ),
    .Q_N(\proj_12.net9 ),
    .Q(\proj_12.flop16/q ));
 sg13g2_tiehi \proj_12.flop2/_1__35  (.L_HI(net35));
 sg13g2_dfrbp_1 \proj_12.flop2/_1_  (.CLK(\proj_12.net19 ),
    .RESET_B(net35),
    .D(\proj_12.net20 ),
    .Q_N(\proj_12.net20 ),
    .Q(\proj_12.flop2/q ));
 sg13g2_tiehi \proj_12.flop3/_1__36  (.L_HI(net36));
 sg13g2_dfrbp_1 \proj_12.flop3/_1_  (.CLK(\proj_12.net20 ),
    .RESET_B(net36),
    .D(\proj_12.net21 ),
    .Q_N(\proj_12.net21 ),
    .Q(\proj_12.flop3/q ));
 sg13g2_tiehi \proj_12.flop4/_1__37  (.L_HI(net49));
 sg13g2_dfrbp_1 \proj_12.flop4/_1_  (.CLK(\proj_12.net21 ),
    .RESET_B(net49),
    .D(\proj_12.net22 ),
    .Q_N(\proj_12.net22 ),
    .Q(\proj_12.flop4/q ));
 sg13g2_tiehi \proj_12.flop5/_1__38  (.L_HI(net50));
 sg13g2_dfrbp_1 \proj_12.flop5/_1_  (.CLK(\proj_12.net22 ),
    .RESET_B(net50),
    .D(\proj_12.net23 ),
    .Q_N(\proj_12.net23 ),
    .Q(\proj_12.flop5/q ));
 sg13g2_tiehi \proj_12.flop6/_1__39  (.L_HI(net51));
 sg13g2_dfrbp_1 \proj_12.flop6/_1_  (.CLK(\proj_12.net23 ),
    .RESET_B(net51),
    .D(\proj_12.net24 ),
    .Q_N(\proj_12.net24 ),
    .Q(\proj_12.flop6/q ));
 sg13g2_tiehi \proj_12.flop7/_1__40  (.L_HI(net52));
 sg13g2_dfrbp_1 \proj_12.flop7/_1_  (.CLK(\proj_12.net24 ),
    .RESET_B(net52),
    .D(\proj_12.net25 ),
    .Q_N(\proj_12.net25 ),
    .Q(\proj_12.flop7/q ));
 sg13g2_tiehi \proj_12.flop8/_1__41  (.L_HI(net53));
 sg13g2_dfrbp_1 \proj_12.flop8/_1_  (.CLK(\proj_12.net25 ),
    .RESET_B(net53),
    .D(\proj_12.net26 ),
    .Q_N(\proj_12.net26 ),
    .Q(\proj_12.flop8/q ));
 sg13g2_tiehi \proj_12.flop9/_1__42  (.L_HI(net54));
 sg13g2_dfrbp_1 \proj_12.flop9/_1_  (.CLK(\proj_12.net26 ),
    .RESET_B(net54),
    .D(\proj_12.net27 ),
    .Q_N(\proj_12.net27 ),
    .Q(\proj_12.flop9/q ));
 sg13g2_tiehi \proj_13.flop1/_1__43  (.L_HI(net55));
 sg13g2_or2_1 \proj_12.or1/_0_  (.X(\proj_12.net8 ),
    .B(\proj_12.net18 ),
    .A(\proj_12.net17 ));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net42),
    .A(net38),
    .X(\proj_12.net7 ));
 sg13g2_xor2_1 \proj_12.xor2/_0_  (.B(net48),
    .A(net41),
    .X(\proj_12.net16 ));
 sg13g2_xor2_1 \proj_12.xor3/_0_  (.B(\proj_12.net15 ),
    .A(\proj_12.net16 ),
    .X(\proj_12.net6 ));
 sg13g2_dfrbp_1 \proj_13.flop1/_1_  (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net55),
    .D(net157),
    .Q_N(\proj_13.net16 ),
    .Q(\proj_13.net17 ));
 sg13g2_tiehi \proj_13.flop10/_1__44  (.L_HI(net56));
 sg13g2_dfrbp_1 \proj_13.flop10/_1_  (.CLK(\proj_13.net29 ),
    .RESET_B(net56),
    .D(\proj_13.net30 ),
    .Q_N(\proj_13.net30 ),
    .Q(\proj_13.net31 ));
 sg13g2_tiehi \proj_13.flop11/_1__45  (.L_HI(net57));
 sg13g2_dfrbp_1 \proj_13.flop11/_1_  (.CLK(\proj_13.net31 ),
    .RESET_B(net57),
    .D(\proj_13.net32 ),
    .Q_N(\proj_13.net32 ),
    .Q(\proj_13.net33 ));
 sg13g2_tiehi \proj_13.flop12/_1__46  (.L_HI(net58));
 sg13g2_dfrbp_1 \proj_13.flop12/_1_  (.CLK(\proj_13.net33 ),
    .RESET_B(net58),
    .D(\proj_13.net34 ),
    .Q_N(\proj_13.net34 ),
    .Q(\proj_13.net35 ));
 sg13g2_tiehi \proj_13.flop13/_1__47  (.L_HI(net59));
 sg13g2_dfrbp_1 \proj_13.flop13/_1_  (.CLK(\proj_13.net35 ),
    .RESET_B(net59),
    .D(\proj_13.net36 ),
    .Q_N(\proj_13.net36 ),
    .Q(\proj_13.net37 ));
 sg13g2_tiehi \proj_13.flop14/_1__48  (.L_HI(net60));
 sg13g2_dfrbp_1 \proj_13.flop14/_1_  (.CLK(\proj_13.net37 ),
    .RESET_B(net60),
    .D(\proj_13.net38 ),
    .Q_N(\proj_13.net38 ),
    .Q(\proj_13.net39 ));
 sg13g2_tiehi \proj_13.flop15/_1__49  (.L_HI(net61));
 sg13g2_dfrbp_1 \proj_13.flop15/_1_  (.CLK(\proj_13.net39 ),
    .RESET_B(net61),
    .D(\proj_13.net40 ),
    .Q_N(\proj_13.net40 ),
    .Q(\proj_13.net41 ));
 sg13g2_tiehi \proj_13.flop16/_1__50  (.L_HI(net62));
 sg13g2_dfrbp_1 \proj_13.flop16/_1_  (.CLK(\proj_13.net41 ),
    .RESET_B(net62),
    .D(\proj_13.net42 ),
    .Q_N(\proj_13.net42 ),
    .Q(\proj_13.net43 ));
 sg13g2_tiehi \proj_13.flop17/_1__51  (.L_HI(net63));
 sg13g2_dfrbp_1 \proj_13.flop17/_1_  (.CLK(\proj_13.net54 ),
    .RESET_B(net63),
    .D(\proj_13.net55 ),
    .Q_N(\proj_13.net55 ),
    .Q(\proj_13.net56 ));
 sg13g2_tiehi \proj_13.flop18/_1__52  (.L_HI(net64));
 sg13g2_dfrbp_1 \proj_13.flop18/_1_  (.CLK(\proj_13.net56 ),
    .RESET_B(net64),
    .D(\proj_13.net57 ),
    .Q_N(\proj_13.net57 ),
    .Q(\proj_13.net58 ));
 sg13g2_tiehi \proj_13.flop19/_1__53  (.L_HI(net65));
 sg13g2_dfrbp_1 \proj_13.flop19/_1_  (.CLK(\proj_13.net58 ),
    .RESET_B(net65),
    .D(\proj_13.net59 ),
    .Q_N(\proj_13.net59 ),
    .Q(\proj_13.net60 ));
 sg13g2_tiehi \proj_13.flop2/_1__54  (.L_HI(net66));
 sg13g2_dfrbp_1 \proj_13.flop2/_1_  (.CLK(\proj_13.net43 ),
    .RESET_B(net66),
    .D(\proj_13.net51 ),
    .Q_N(\proj_13.net51 ),
    .Q(\proj_13.net52 ));
 sg13g2_tiehi \proj_13.flop20/_1__55  (.L_HI(net67));
 sg13g2_dfrbp_1 \proj_13.flop20/_1_  (.CLK(\proj_13.net60 ),
    .RESET_B(net67),
    .D(\proj_13.net61 ),
    .Q_N(\proj_13.net61 ),
    .Q(\proj_13.net62 ));
 sg13g2_tiehi \proj_13.flop21/_1__56  (.L_HI(net68));
 sg13g2_dfrbp_1 \proj_13.flop21/_1_  (.CLK(\proj_13.net62 ),
    .RESET_B(net68),
    .D(\proj_13.net63 ),
    .Q_N(\proj_13.net63 ),
    .Q(\proj_13.net64 ));
 sg13g2_tiehi \proj_13.flop22/_1__57  (.L_HI(net69));
 sg13g2_dfrbp_1 \proj_13.flop22/_1_  (.CLK(\proj_13.net64 ),
    .RESET_B(net69),
    .D(\proj_13.net65 ),
    .Q_N(\proj_13.net65 ),
    .Q(\proj_13.net66 ));
 sg13g2_tiehi \proj_13.flop23/_1__58  (.L_HI(net70));
 sg13g2_dfrbp_1 \proj_13.flop23/_1_  (.CLK(\proj_13.net66 ),
    .RESET_B(net70),
    .D(\proj_13.net67 ),
    .Q_N(\proj_13.net67 ),
    .Q(\proj_13.net68 ));
 sg13g2_tiehi \proj_13.flop24/_1__59  (.L_HI(net71));
 sg13g2_dfrbp_1 \proj_13.flop24/_1_  (.CLK(\proj_13.net68 ),
    .RESET_B(net71),
    .D(\proj_13.net69 ),
    .Q_N(\proj_13.net69 ),
    .Q(\proj_13.net70 ));
 sg13g2_tiehi \proj_13.flop25/_1__60  (.L_HI(net72));
 sg13g2_dfrbp_1 \proj_13.flop25/_1_  (.CLK(\proj_13.net70 ),
    .RESET_B(net72),
    .D(\proj_13.net71 ),
    .Q_N(\proj_13.net71 ),
    .Q(\proj_13.net72 ));
 sg13g2_tiehi \proj_13.flop26/_1__61  (.L_HI(net73));
 sg13g2_dfrbp_1 \proj_13.flop26/_1_  (.CLK(\proj_13.net72 ),
    .RESET_B(net73),
    .D(\proj_13.net73 ),
    .Q_N(\proj_13.net73 ),
    .Q(\proj_13.net74 ));
 sg13g2_tiehi \proj_13.flop27/_1__62  (.L_HI(net74));
 sg13g2_dfrbp_1 \proj_13.flop27/_1_  (.CLK(\proj_13.net74 ),
    .RESET_B(net74),
    .D(\proj_13.net75 ),
    .Q_N(\proj_13.net75 ),
    .Q(\proj_13.net76 ));
 sg13g2_tiehi \proj_13.flop28/_1__63  (.L_HI(net75));
 sg13g2_dfrbp_1 \proj_13.flop28/_1_  (.CLK(\proj_13.net76 ),
    .RESET_B(net75),
    .D(\proj_13.net77 ),
    .Q_N(\proj_13.net77 ),
    .Q(\proj_13.net78 ));
 sg13g2_tiehi \proj_13.flop29/_1__64  (.L_HI(net76));
 sg13g2_dfrbp_1 \proj_13.flop29/_1_  (.CLK(\proj_13.net78 ),
    .RESET_B(net76),
    .D(\proj_13.net79 ),
    .Q_N(\proj_13.net79 ),
    .Q(\proj_13.net80 ));
 sg13g2_tiehi \proj_13.flop3/_1__65  (.L_HI(net77));
 sg13g2_dfrbp_1 \proj_13.flop3/_1_  (.CLK(\proj_13.net52 ),
    .RESET_B(net77),
    .D(\proj_13.net53 ),
    .Q_N(\proj_13.net53 ),
    .Q(\proj_13.net54 ));
 sg13g2_tiehi \proj_13.flop30/_1__66  (.L_HI(net78));
 sg13g2_dfrbp_1 \proj_13.flop30/_1_  (.CLK(\proj_13.net80 ),
    .RESET_B(net78),
    .D(\proj_13.net81 ),
    .Q_N(\proj_13.net81 ),
    .Q(\proj_13.net82 ));
 sg13g2_tiehi \proj_13.flop31/_1__67  (.L_HI(net79));
 sg13g2_dfrbp_1 \proj_13.flop31/_1_  (.CLK(\proj_13.net82 ),
    .RESET_B(net79),
    .D(\proj_13.net83 ),
    .Q_N(\proj_13.net83 ),
    .Q(\proj_13.net84 ));
 sg13g2_tiehi \proj_13.flop32/_1__68  (.L_HI(net80));
 sg13g2_dfrbp_1 \proj_13.flop32/_1_  (.CLK(\proj_13.net84 ),
    .RESET_B(net80),
    .D(\proj_13.net85 ),
    .Q_N(\proj_13.net85 ),
    .Q(\proj_13.net86 ));
 sg13g2_tiehi \proj_13.flop33/_1__69  (.L_HI(net81));
 sg13g2_dfrbp_1 \proj_13.flop33/_1_  (.CLK(\proj_13.net86 ),
    .RESET_B(net81),
    .D(\proj_13.net87 ),
    .Q_N(\proj_13.net87 ),
    .Q(\proj_13.net88 ));
 sg13g2_tiehi \proj_13.flop34/_1__70  (.L_HI(net82));
 sg13g2_dfrbp_1 \proj_13.flop34/_1_  (.CLK(\proj_13.net88 ),
    .RESET_B(net82),
    .D(\proj_13.net89 ),
    .Q_N(\proj_13.net89 ),
    .Q(\proj_13.net90 ));
 sg13g2_tiehi \proj_13.flop35/_1__71  (.L_HI(net83));
 sg13g2_dfrbp_1 \proj_13.flop35/_1_  (.CLK(\proj_13.net90 ),
    .RESET_B(net83),
    .D(\proj_13.net91 ),
    .Q_N(\proj_13.net91 ),
    .Q(\proj_13.net92 ));
 sg13g2_tiehi \proj_13.flop36/_1__72  (.L_HI(net84));
 sg13g2_dfrbp_1 \proj_13.flop36/_1_  (.CLK(\proj_13.net92 ),
    .RESET_B(net84),
    .D(\proj_13.net93 ),
    .Q_N(\proj_13.net93 ),
    .Q(\proj_13.net94 ));
 sg13g2_tiehi \proj_13.flop37/_1__73  (.L_HI(net85));
 sg13g2_dfrbp_1 \proj_13.flop37/_1_  (.CLK(\proj_13.net94 ),
    .RESET_B(net85),
    .D(\proj_13.net95 ),
    .Q_N(\proj_13.net95 ),
    .Q(\proj_13.net96 ));
 sg13g2_tiehi \proj_13.flop38/_1__74  (.L_HI(net86));
 sg13g2_dfrbp_1 \proj_13.flop38/_1_  (.CLK(\proj_13.net96 ),
    .RESET_B(net86),
    .D(\proj_13.net97 ),
    .Q_N(\proj_13.net97 ),
    .Q(\proj_13.net98 ));
 sg13g2_tiehi \proj_13.flop39/_1__75  (.L_HI(net87));
 sg13g2_dfrbp_1 \proj_13.flop39/_1_  (.CLK(\proj_13.net98 ),
    .RESET_B(net87),
    .D(\proj_13.net99 ),
    .Q_N(\proj_13.net99 ),
    .Q(\proj_13.net100 ));
 sg13g2_tiehi \proj_13.flop4/_1__76  (.L_HI(net88));
 sg13g2_dfrbp_1 \proj_13.flop4/_1_  (.CLK(\proj_13.net17 ),
    .RESET_B(net88),
    .D(\proj_13.net18 ),
    .Q_N(\proj_13.net18 ),
    .Q(\proj_13.net19 ));
 sg13g2_tiehi \proj_13.flop40/_1__77  (.L_HI(net89));
 sg13g2_dfrbp_1 \proj_13.flop40/_1_  (.CLK(\proj_13.net100 ),
    .RESET_B(net89),
    .D(\proj_13.net101 ),
    .Q_N(\proj_13.net101 ),
    .Q(\proj_13.net102 ));
 sg13g2_tiehi \proj_13.flop41/_1__78  (.L_HI(net90));
 sg13g2_dfrbp_1 \proj_13.flop41/_1_  (.CLK(\proj_13.net102 ),
    .RESET_B(net90),
    .D(\proj_13.net103 ),
    .Q_N(\proj_13.net103 ),
    .Q(\proj_13.net104 ));
 sg13g2_tiehi \proj_13.flop42/_1__79  (.L_HI(net91));
 sg13g2_dfrbp_1 \proj_13.flop42/_1_  (.CLK(\proj_13.net104 ),
    .RESET_B(net91),
    .D(\proj_13.net105 ),
    .Q_N(\proj_13.net105 ),
    .Q(\proj_13.net106 ));
 sg13g2_tiehi \proj_13.flop43/_1__80  (.L_HI(net92));
 sg13g2_dfrbp_1 \proj_13.flop43/_1_  (.CLK(\proj_13.net106 ),
    .RESET_B(net92),
    .D(\proj_13.net107 ),
    .Q_N(\proj_13.net107 ),
    .Q(\proj_13.net108 ));
 sg13g2_tiehi \proj_13.flop44/_1__81  (.L_HI(net93));
 sg13g2_dfrbp_1 \proj_13.flop44/_1_  (.CLK(\proj_13.net108 ),
    .RESET_B(net93),
    .D(\proj_13.net109 ),
    .Q_N(\proj_13.net109 ),
    .Q(\proj_13.net110 ));
 sg13g2_tiehi \proj_13.flop45/_1__82  (.L_HI(net94));
 sg13g2_dfrbp_1 \proj_13.flop45/_1_  (.CLK(\proj_13.net110 ),
    .RESET_B(net94),
    .D(\proj_13.net111 ),
    .Q_N(\proj_13.net111 ),
    .Q(\proj_13.net112 ));
 sg13g2_tiehi \proj_13.flop46/_1__83  (.L_HI(net95));
 sg13g2_dfrbp_1 \proj_13.flop46/_1_  (.CLK(\proj_13.net112 ),
    .RESET_B(net95),
    .D(\proj_13.net113 ),
    .Q_N(\proj_13.net113 ),
    .Q(\proj_13.net114 ));
 sg13g2_tiehi \proj_13.flop47/_1__84  (.L_HI(net96));
 sg13g2_dfrbp_1 \proj_13.flop47/_1_  (.CLK(\proj_13.net114 ),
    .RESET_B(net96),
    .D(\proj_13.net115 ),
    .Q_N(\proj_13.net115 ),
    .Q(\proj_13.net116 ));
 sg13g2_tiehi \proj_13.flop48/_1__85  (.L_HI(net97));
 sg13g2_dfrbp_1 \proj_13.flop48/_1_  (.CLK(\proj_13.net116 ),
    .RESET_B(net97),
    .D(\proj_13.net117 ),
    .Q_N(\proj_13.net117 ),
    .Q(\proj_13.net118 ));
 sg13g2_tiehi \proj_13.flop49/_1__86  (.L_HI(net98));
 sg13g2_dfrbp_1 \proj_13.flop49/_1_  (.CLK(\proj_13.net118 ),
    .RESET_B(net98),
    .D(\proj_13.net119 ),
    .Q_N(\proj_13.net119 ),
    .Q(\proj_13.net120 ));
 sg13g2_tiehi \proj_13.flop5/_1__87  (.L_HI(net99));
 sg13g2_dfrbp_1 \proj_13.flop5/_1_  (.CLK(\proj_13.net23 ),
    .RESET_B(net99),
    .D(\proj_13.net24 ),
    .Q_N(\proj_13.net24 ),
    .Q(\proj_13.net25 ));
 sg13g2_tiehi \proj_13.flop50/_1__88  (.L_HI(net100));
 sg13g2_dfrbp_1 \proj_13.flop50/_1_  (.CLK(\proj_13.net120 ),
    .RESET_B(net100),
    .D(\proj_13.net121 ),
    .Q_N(\proj_13.net121 ),
    .Q(\proj_13.net122 ));
 sg13g2_tiehi \proj_13.flop51/_1__89  (.L_HI(net101));
 sg13g2_dfrbp_1 \proj_13.flop51/_1_  (.CLK(\proj_13.net122 ),
    .RESET_B(net101),
    .D(\proj_13.net123 ),
    .Q_N(\proj_13.net123 ),
    .Q(\proj_13.net124 ));
 sg13g2_tiehi \proj_13.flop52/_1__90  (.L_HI(net102));
 sg13g2_dfrbp_1 \proj_13.flop52/_1_  (.CLK(\proj_13.net124 ),
    .RESET_B(net102),
    .D(\proj_13.net125 ),
    .Q_N(\proj_13.net125 ),
    .Q(\proj_13.net126 ));
 sg13g2_tiehi \proj_13.flop53/_1__91  (.L_HI(net103));
 sg13g2_dfrbp_1 \proj_13.flop53/_1_  (.CLK(\proj_13.net126 ),
    .RESET_B(net103),
    .D(\proj_13.net127 ),
    .Q_N(\proj_13.net127 ),
    .Q(\proj_13.net128 ));
 sg13g2_tiehi \proj_13.flop54/_1__92  (.L_HI(net104));
 sg13g2_dfrbp_1 \proj_13.flop54/_1_  (.CLK(\proj_13.net128 ),
    .RESET_B(net104),
    .D(\proj_13.net129 ),
    .Q_N(\proj_13.net129 ),
    .Q(\proj_13.net130 ));
 sg13g2_tiehi \proj_13.flop55/_1__93  (.L_HI(net105));
 sg13g2_dfrbp_1 \proj_13.flop55/_1_  (.CLK(\proj_13.net130 ),
    .RESET_B(net105),
    .D(\proj_13.net131 ),
    .Q_N(\proj_13.net131 ),
    .Q(\proj_13.net132 ));
 sg13g2_tiehi \proj_13.flop56/_1__94  (.L_HI(net106));
 sg13g2_dfrbp_1 \proj_13.flop56/_1_  (.CLK(\proj_13.net132 ),
    .RESET_B(net106),
    .D(\proj_13.net133 ),
    .Q_N(\proj_13.net133 ),
    .Q(\proj_13.net134 ));
 sg13g2_tiehi \proj_13.flop57/_1__95  (.L_HI(net107));
 sg13g2_dfrbp_1 \proj_13.flop57/_1_  (.CLK(\proj_13.net136 ),
    .RESET_B(net107),
    .D(\proj_13.net135 ),
    .Q_N(\proj_13.net135 ),
    .Q(\proj_13.net137 ));
 sg13g2_tiehi \proj_13.flop58/_1__96  (.L_HI(net108));
 sg13g2_dfrbp_1 \proj_13.flop58/_1_  (.CLK(\proj_13.net137 ),
    .RESET_B(net108),
    .D(\proj_13.net138 ),
    .Q_N(\proj_13.net138 ),
    .Q(\proj_13.net139 ));
 sg13g2_tiehi \proj_13.flop59/_1__97  (.L_HI(net109));
 sg13g2_dfrbp_1 \proj_13.flop59/_1_  (.CLK(\proj_13.net139 ),
    .RESET_B(net109),
    .D(\proj_13.net140 ),
    .Q_N(\proj_13.net140 ),
    .Q(\proj_13.net141 ));
 sg13g2_tiehi \proj_13.flop6/_1__98  (.L_HI(net110));
 sg13g2_dfrbp_1 \proj_13.flop6/_1_  (.CLK(\proj_13.net19 ),
    .RESET_B(net110),
    .D(\proj_13.net20 ),
    .Q_N(\proj_13.net20 ),
    .Q(\proj_13.net21 ));
 sg13g2_tiehi \proj_13.flop60/_1__99  (.L_HI(net111));
 sg13g2_dfrbp_1 \proj_13.flop60/_1_  (.CLK(\proj_13.net141 ),
    .RESET_B(net111),
    .D(\proj_13.net142 ),
    .Q_N(\proj_13.net142 ),
    .Q(\proj_13.net143 ));
 sg13g2_tiehi \proj_13.flop61/_1__100  (.L_HI(net112));
 sg13g2_dfrbp_1 \proj_13.flop61/_1_  (.CLK(\proj_13.net143 ),
    .RESET_B(net112),
    .D(\proj_13.net144 ),
    .Q_N(\proj_13.net144 ),
    .Q(\proj_13.net145 ));
 sg13g2_tiehi \proj_13.flop62/_1__101  (.L_HI(net113));
 sg13g2_dfrbp_1 \proj_13.flop62/_1_  (.CLK(\proj_13.net145 ),
    .RESET_B(net113),
    .D(\proj_13.net146 ),
    .Q_N(\proj_13.net146 ),
    .Q(\proj_13.net147 ));
 sg13g2_tiehi \proj_13.flop63/_1__102  (.L_HI(net114));
 sg13g2_dfrbp_1 \proj_13.flop63/_1_  (.CLK(\proj_13.net147 ),
    .RESET_B(net114),
    .D(\proj_13.net148 ),
    .Q_N(\proj_13.net148 ),
    .Q(\proj_13.net149 ));
 sg13g2_tiehi \proj_13.flop64/_1__103  (.L_HI(net115));
 sg13g2_dfrbp_1 \proj_13.flop64/_1_  (.CLK(\proj_13.net149 ),
    .RESET_B(net115),
    .D(\proj_13.net150 ),
    .Q_N(\proj_13.net150 ),
    .Q(\proj_13.net151 ));
 sg13g2_tiehi \proj_13.flop65/_1__104  (.L_HI(net116));
 sg13g2_dfrbp_1 \proj_13.flop65/_1_  (.CLK(\proj_13.net151 ),
    .RESET_B(net116),
    .D(\proj_13.net152 ),
    .Q_N(\proj_13.net152 ),
    .Q(\proj_13.net153 ));
 sg13g2_tiehi \proj_13.flop66/_1__105  (.L_HI(net117));
 sg13g2_dfrbp_1 \proj_13.flop66/_1_  (.CLK(\proj_13.net153 ),
    .RESET_B(net117),
    .D(\proj_13.net154 ),
    .Q_N(\proj_13.net154 ),
    .Q(\proj_13.net155 ));
 sg13g2_tiehi \proj_13.flop67/_1__106  (.L_HI(net118));
 sg13g2_dfrbp_1 \proj_13.flop67/_1_  (.CLK(\proj_13.net155 ),
    .RESET_B(net118),
    .D(\proj_13.net156 ),
    .Q_N(\proj_13.net156 ),
    .Q(\proj_13.net157 ));
 sg13g2_tiehi \proj_13.flop68/_1__107  (.L_HI(net119));
 sg13g2_dfrbp_1 \proj_13.flop68/_1_  (.CLK(\proj_13.net157 ),
    .RESET_B(net119),
    .D(\proj_13.net158 ),
    .Q_N(\proj_13.net158 ),
    .Q(\proj_13.net159 ));
 sg13g2_tiehi \proj_13.flop69/_1__108  (.L_HI(net120));
 sg13g2_dfrbp_1 \proj_13.flop69/_1_  (.CLK(\proj_13.net159 ),
    .RESET_B(net120),
    .D(\proj_13.net160 ),
    .Q_N(\proj_13.net160 ),
    .Q(\proj_13.net161 ));
 sg13g2_tiehi \proj_13.flop7/_1__109  (.L_HI(net121));
 sg13g2_dfrbp_1 \proj_13.flop7/_1_  (.CLK(\proj_13.net21 ),
    .RESET_B(net121),
    .D(\proj_13.net22 ),
    .Q_N(\proj_13.net22 ),
    .Q(\proj_13.net23 ));
 sg13g2_tiehi \proj_13.flop70/_1__110  (.L_HI(net122));
 sg13g2_dfrbp_1 \proj_13.flop70/_1_  (.CLK(\proj_13.net161 ),
    .RESET_B(net122),
    .D(\proj_13.net162 ),
    .Q_N(\proj_13.net162 ),
    .Q(\proj_13.net163 ));
 sg13g2_tiehi \proj_13.flop71/_1__111  (.L_HI(net123));
 sg13g2_dfrbp_1 \proj_13.flop71/_1_  (.CLK(\proj_13.net165 ),
    .RESET_B(net123),
    .D(\proj_13.net164 ),
    .Q_N(\proj_13.net164 ),
    .Q(\proj_13.net166 ));
 sg13g2_tiehi \proj_13.flop72/_1__112  (.L_HI(net124));
 sg13g2_dfrbp_1 \proj_13.flop72/_1_  (.CLK(\proj_13.net166 ),
    .RESET_B(net124),
    .D(\proj_13.net167 ),
    .Q_N(\proj_13.net167 ),
    .Q(\proj_13.net168 ));
 sg13g2_tiehi \proj_13.flop73/_1__113  (.L_HI(net125));
 sg13g2_dfrbp_1 \proj_13.flop73/_1_  (.CLK(\proj_13.net168 ),
    .RESET_B(net125),
    .D(\proj_13.net169 ),
    .Q_N(\proj_13.net169 ),
    .Q(\proj_13.net170 ));
 sg13g2_tiehi \proj_13.flop74/_1__114  (.L_HI(net126));
 sg13g2_dfrbp_1 \proj_13.flop74/_1_  (.CLK(\proj_13.net170 ),
    .RESET_B(net126),
    .D(\proj_13.net171 ),
    .Q_N(\proj_13.net171 ),
    .Q(\proj_13.net172 ));
 sg13g2_tiehi \proj_13.flop75/_1__115  (.L_HI(net127));
 sg13g2_dfrbp_1 \proj_13.flop75/_1_  (.CLK(\proj_13.net172 ),
    .RESET_B(net127),
    .D(\proj_13.net173 ),
    .Q_N(\proj_13.net173 ),
    .Q(\proj_13.net174 ));
 sg13g2_tiehi \proj_13.flop76/_1__116  (.L_HI(net128));
 sg13g2_dfrbp_1 \proj_13.flop76/_1_  (.CLK(\proj_13.net174 ),
    .RESET_B(net128),
    .D(\proj_13.net175 ),
    .Q_N(\proj_13.net175 ),
    .Q(\proj_13.net176 ));
 sg13g2_tiehi \proj_13.flop77/_1__117  (.L_HI(net129));
 sg13g2_dfrbp_1 \proj_13.flop77/_1_  (.CLK(\proj_13.net176 ),
    .RESET_B(net129),
    .D(\proj_13.net177 ),
    .Q_N(\proj_13.net177 ),
    .Q(\proj_13.net178 ));
 sg13g2_tiehi \proj_13.flop78/_1__118  (.L_HI(net130));
 sg13g2_dfrbp_1 \proj_13.flop78/_1_  (.CLK(\proj_13.net178 ),
    .RESET_B(net130),
    .D(\proj_13.net179 ),
    .Q_N(\proj_13.net179 ),
    .Q(\proj_13.net180 ));
 sg13g2_tiehi \proj_13.flop79/_1__119  (.L_HI(net131));
 sg13g2_dfrbp_1 \proj_13.flop79/_1_  (.CLK(\proj_13.net180 ),
    .RESET_B(net131),
    .D(\proj_13.net181 ),
    .Q_N(\proj_13.net181 ),
    .Q(\proj_13.net182 ));
 sg13g2_tiehi \proj_13.flop8/_1__120  (.L_HI(net132));
 sg13g2_dfrbp_1 \proj_13.flop8/_1_  (.CLK(\proj_13.net25 ),
    .RESET_B(net132),
    .D(\proj_13.net26 ),
    .Q_N(\proj_13.net26 ),
    .Q(\proj_13.net27 ));
 sg13g2_tiehi \proj_13.flop80/_1__121  (.L_HI(net133));
 sg13g2_dfrbp_1 \proj_13.flop80/_1_  (.CLK(\proj_13.net182 ),
    .RESET_B(net133),
    .D(\proj_13.net183 ),
    .Q_N(\proj_13.net183 ),
    .Q(\proj_13.net184 ));
 sg13g2_tiehi \proj_13.flop81/_1__122  (.L_HI(net134));
 sg13g2_dfrbp_1 \proj_13.flop81/_1_  (.CLK(\proj_13.net184 ),
    .RESET_B(net134),
    .D(\proj_13.net185 ),
    .Q_N(\proj_13.net185 ),
    .Q(\proj_13.net186 ));
 sg13g2_tiehi \proj_13.flop82/_1__123  (.L_HI(net135));
 sg13g2_dfrbp_1 \proj_13.flop82/_1_  (.CLK(\proj_13.net186 ),
    .RESET_B(net135),
    .D(\proj_13.net187 ),
    .Q_N(\proj_13.net187 ),
    .Q(\proj_13.net188 ));
 sg13g2_tiehi \proj_13.flop83/_1__124  (.L_HI(net136));
 sg13g2_dfrbp_1 \proj_13.flop83/_1_  (.CLK(\proj_13.net188 ),
    .RESET_B(net136),
    .D(\proj_13.net189 ),
    .Q_N(\proj_13.net189 ),
    .Q(\proj_13.net190 ));
 sg13g2_tiehi \proj_13.flop84/_1__125  (.L_HI(net137));
 sg13g2_dfrbp_1 \proj_13.flop84/_1_  (.CLK(\proj_13.net190 ),
    .RESET_B(net137),
    .D(\proj_13.net191 ),
    .Q_N(\proj_13.net191 ),
    .Q(\proj_13.net136 ));
 sg13g2_tiehi \proj_13.flop85/_1__126  (.L_HI(net138));
 sg13g2_dfrbp_1 \proj_13.flop85/_1_  (.CLK(\proj_13.net134 ),
    .RESET_B(net138),
    .D(\proj_13.net192 ),
    .Q_N(\proj_13.net192 ),
    .Q(\proj_13.net193 ));
 sg13g2_tiehi \proj_13.flop86/_1__127  (.L_HI(net139));
 sg13g2_dfrbp_1 \proj_13.flop86/_1_  (.CLK(\proj_13.net193 ),
    .RESET_B(net139),
    .D(\proj_13.net194 ),
    .Q_N(\proj_13.net194 ),
    .Q(\proj_13.net195 ));
 sg13g2_tiehi \proj_13.flop87/_1__128  (.L_HI(net140));
 sg13g2_dfrbp_1 \proj_13.flop87/_1_  (.CLK(\proj_13.net195 ),
    .RESET_B(net140),
    .D(\proj_13.net196 ),
    .Q_N(\proj_13.net196 ),
    .Q(\proj_13.net197 ));
 sg13g2_tiehi \proj_13.flop88/_1__129  (.L_HI(net141));
 sg13g2_dfrbp_1 \proj_13.flop88/_1_  (.CLK(\proj_13.net197 ),
    .RESET_B(net141),
    .D(\proj_13.net198 ),
    .Q_N(\proj_13.net198 ),
    .Q(\proj_13.net199 ));
 sg13g2_tiehi \proj_13.flop89/_1__130  (.L_HI(net142));
 sg13g2_dfrbp_1 \proj_13.flop89/_1_  (.CLK(\proj_13.net199 ),
    .RESET_B(net142),
    .D(\proj_13.net200 ),
    .Q_N(\proj_13.net200 ),
    .Q(\proj_13.net201 ));
 sg13g2_tiehi \proj_13.flop9/_1__131  (.L_HI(net143));
 sg13g2_dfrbp_1 \proj_13.flop9/_1_  (.CLK(\proj_13.net27 ),
    .RESET_B(net143),
    .D(\proj_13.net28 ),
    .Q_N(\proj_13.net28 ),
    .Q(\proj_13.net29 ));
 sg13g2_tiehi \proj_13.flop90/_1__132  (.L_HI(net144));
 sg13g2_dfrbp_1 \proj_13.flop90/_1_  (.CLK(\proj_13.net201 ),
    .RESET_B(net144),
    .D(\proj_13.net202 ),
    .Q_N(\proj_13.net202 ),
    .Q(\proj_13.net203 ));
 sg13g2_tiehi \proj_13.flop91/_1__133  (.L_HI(net145));
 sg13g2_dfrbp_1 \proj_13.flop91/_1_  (.CLK(\proj_13.net203 ),
    .RESET_B(net145),
    .D(\proj_13.net204 ),
    .Q_N(\proj_13.net204 ),
    .Q(\proj_13.net205 ));
 sg13g2_tiehi \proj_13.flop92/_1__134  (.L_HI(net146));
 sg13g2_dfrbp_1 \proj_13.flop92/_1_  (.CLK(\proj_13.net205 ),
    .RESET_B(net146),
    .D(\proj_13.net206 ),
    .Q_N(\proj_13.net206 ),
    .Q(\proj_13.net207 ));
 sg13g2_tiehi \proj_13.flop93/_1__135  (.L_HI(net147));
 sg13g2_dfrbp_1 \proj_13.flop93/_1_  (.CLK(\proj_13.net207 ),
    .RESET_B(net147),
    .D(\proj_13.net208 ),
    .Q_N(\proj_13.net208 ),
    .Q(\proj_13.net209 ));
 sg13g2_tiehi \proj_13.flop94/_1__136  (.L_HI(net148));
 sg13g2_dfrbp_1 \proj_13.flop94/_1_  (.CLK(\proj_13.net209 ),
    .RESET_B(net148),
    .D(\proj_13.net210 ),
    .Q_N(\proj_13.net210 ),
    .Q(\proj_13.net211 ));
 sg13g2_tiehi \proj_13.flop95/_1__137  (.L_HI(net149));
 sg13g2_dfrbp_1 \proj_13.flop95/_1_  (.CLK(\proj_13.net211 ),
    .RESET_B(net149),
    .D(\proj_13.net212 ),
    .Q_N(\proj_13.net212 ),
    .Q(\proj_13.net213 ));
 sg13g2_tiehi \proj_13.flop96/_1__138  (.L_HI(net150));
 sg13g2_dfrbp_1 \proj_13.flop96/_1_  (.CLK(\proj_13.net213 ),
    .RESET_B(net150),
    .D(\proj_13.net214 ),
    .Q_N(\proj_13.net214 ),
    .Q(\proj_13.net215 ));
 sg13g2_tiehi \proj_13.flop97/_1__139  (.L_HI(net151));
 sg13g2_dfrbp_1 \proj_13.flop97/_1_  (.CLK(\proj_13.net215 ),
    .RESET_B(net151),
    .D(\proj_13.net216 ),
    .Q_N(\proj_13.net216 ),
    .Q(\proj_13.net217 ));
 sg13g2_tiehi \proj_13.flop98/_1__140  (.L_HI(net152));
 sg13g2_dfrbp_1 \proj_13.flop98/_1_  (.CLK(\proj_13.net217 ),
    .RESET_B(net152),
    .D(\proj_13.net218 ),
    .Q_N(\proj_13.net218 ),
    .Q(\proj_13.net165 ));
 sg13g2_tiehi \proj__8.flop1/_1__141  (.L_HI(net153));
 sg13g2_mux2_1 \proj_13.mux1/_0_  (.A0(net45),
    .A1(net45),
    .S(\proj_13.net43 ),
    .X(\proj_13.net3 ));
 sg13g2_mux2_1 \proj_13.mux2/_0_  (.A0(net44),
    .A1(\proj_13.net44 ),
    .S(\proj_13.net43 ),
    .X(\proj_13.net4 ));
 sg13g2_mux2_1 \proj_13.mux3/_0_  (.A0(net45),
    .A1(\proj_13.net45 ),
    .S(\proj_13.net43 ),
    .X(\proj_13.net5 ));
 sg13g2_mux2_1 \proj_13.mux4/_0_  (.A0(net45),
    .A1(net45),
    .S(\proj_13.net43 ),
    .X(\proj_13.net6 ));
 sg13g2_mux2_1 \proj_13.mux5/_0_  (.A0(\proj_13.net46 ),
    .A1(\proj_13.net47 ),
    .S(\proj_13.net43 ),
    .X(\proj_13.net7 ));
 sg13g2_mux2_1 \proj_13.mux6/_0_  (.A0(net46),
    .A1(\proj_13.net48 ),
    .S(\proj_13.net43 ),
    .X(\proj_13.net8 ));
 sg13g2_mux2_1 \proj_13.mux7/_0_  (.A0(\proj_13.net49 ),
    .A1(\proj_13.net50 ),
    .S(\proj_13.net43 ),
    .X(\proj_13.net9 ));
 sg13g2_inv_1 \proj_13.not1/_0_  (.Y(\proj_13.net44 ),
    .A(net44));
 sg13g2_inv_1 \proj_13.not2/_0_  (.Y(\proj_13.net45 ),
    .A(net44));
 sg13g2_inv_1 \proj_13.not3/_0_  (.Y(\proj_13.net47 ),
    .A(net44));
 sg13g2_inv_1 \proj_13.not4/_0_  (.Y(\proj_13.net46 ),
    .A(net44));
 sg13g2_inv_1 \proj_13.not5/_0_  (.Y(\proj_13.net48 ),
    .A(net44));
 sg13g2_inv_1 \proj_13.not6/_0_  (.Y(\proj_13.net50 ),
    .A(net44));
 sg13g2_inv_1 \proj_13.not7/_0_  (.Y(\proj_13.net49 ),
    .A(net44));
 sg13g2_inv_1 \proj_13.not8/_0_  (.Y(\proj_13.net10 ),
    .A(\proj_13.net163 ));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(net41),
    .B(\proj_14.net10 ),
    .X(\proj_14.net11 ));
 sg13g2_and2_1 \proj_14.and2/_0_  (.A(net43),
    .B(net48),
    .X(\proj_14.net12 ));
 sg13g2_or2_1 \proj_14.or1/_0_  (.X(\proj_14.net5 ),
    .B(\proj_14.net11 ),
    .A(\proj_14.net12 ));
 sg13g2_xor2_1 \proj_14.xor1/_0_  (.B(net48),
    .A(net43),
    .X(\proj_14.net10 ));
 sg13g2_xor2_1 \proj_14.xor2/_0_  (.B(\proj_14.net10 ),
    .A(net41),
    .X(\proj_14.net4 ));
 sg13g2_and2_1 \proj__0.and1/_0_  (.A(net43),
    .B(net48),
    .X(\proj__0.net15 ));
 sg13g2_and2_1 \proj__0.and2/_0_  (.A(net41),
    .B(\proj__0.net15 ),
    .X(\proj__0.net16 ));
 sg13g2_and2_1 \proj__0.and3/_0_  (.A(net39),
    .B(\proj__0.net16 ),
    .X(\proj__0.net17 ));
 sg13g2_and2_1 \proj__0.and4/_0_  (.A(net3),
    .B(\proj__0.net17 ),
    .X(\proj__0.net18 ));
 sg13g2_and2_1 \proj__0.and5/_0_  (.A(net4),
    .B(\proj__0.net18 ),
    .X(\proj__0.net19 ));
 sg13g2_and2_1 \proj__0.and6/_0_  (.A(net5),
    .B(\proj__0.net19 ),
    .X(\proj__0.net20 ));
 sg13g2_and2_1 \proj__0.and7/_0_  (.A(net6),
    .B(\proj__0.net20 ),
    .X(\proj__0.net9 ));
 sg13g2_inv_1 \proj__1.not1/_0_  (.Y(\proj__1.net9 ),
    .A(net46));
 sg13g2_inv_1 \proj__1.not2/_0_  (.Y(\proj__1.net10 ),
    .A(net42));
 sg13g2_inv_1 \proj__1.not3/_0_  (.Y(\proj__1.net11 ),
    .A(net40));
 sg13g2_inv_1 \proj__1.not4/_0_  (.Y(\proj__1.net12 ),
    .A(net38));
 sg13g2_mux2_1 \proj__2.mux1/_0_  (.A0(net37),
    .A1(net5),
    .S(net6),
    .X(\proj__2.net4 ));
 sg13g2_nand2_1 \proj__3.nand1/_0_  (.Y(\proj__3.net11 ),
    .A(net1),
    .B(clknet_1_0__leaf_clk));
 sg13g2_nand2_1 \proj__3.nand2/_0_  (.Y(\proj__3.net12 ),
    .A(net42),
    .B(net47));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net13 ),
    .A(net40));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net14 ),
    .A(net38));
 sg13g2_and2_1 \proj__4.and1/_0_  (.A(net38),
    .B(net41),
    .X(\proj__4.net10 ));
 sg13g2_or2_1 \proj__4.or1/_0_  (.X(\proj__4.net9 ),
    .B(net47),
    .A(net42));
 sg13g2_nand2_1 \proj__5.nand1/_0_  (.Y(\proj__5.net9 ),
    .A(net42),
    .B(net47));
 sg13g2_inv_1 \proj__5.not3/_0_  (.Y(\proj__5.net10 ),
    .A(net40));
 sg13g2_inv_1 \proj__5.not4/_0_  (.Y(\proj__5.net11 ),
    .A(net38));
 sg13g2_and2_1 \proj__6.gate1/_0_  (.A(net39),
    .B(net48),
    .X(\proj__6.net11 ));
 sg13g2_and2_1 \proj__6.gate10/_0_  (.A(\proj__6.net16 ),
    .B(\proj__6.net11 ),
    .X(\proj__6.net12 ));
 sg13g2_and2_1 \proj__6.gate11/_0_  (.A(\proj__6.net17 ),
    .B(\proj__6.net18 ),
    .X(\proj__6.net13 ));
 sg13g2_and2_1 \proj__6.gate12/_0_  (.A(net6),
    .B(\proj__6.net14 ),
    .X(\proj__6.net9 ));
 sg13g2_xor2_1 \proj__6.gate3/_0_  (.B(\proj__6.net12 ),
    .A(\proj__6.net13 ),
    .X(\proj__6.net14 ));
 sg13g2_or2_1 \proj__6.gate7/_0_  (.X(\proj__6.net16 ),
    .B(net37),
    .A(net5));
 sg13g2_or2_1 \proj__6.gate8/_0_  (.X(\proj__6.net17 ),
    .B(net4),
    .A(net5));
 sg13g2_and2_1 \proj__6.gate9/_0_  (.A(net41),
    .B(net43),
    .X(\proj__6.net18 ));
 sg13g2_and2_1 \proj__7.and1/_0_  (.A(net5),
    .B(net38),
    .X(\proj__7.net13 ));
 sg13g2_nand2_1 \proj__7.nand1/_0_  (.Y(\proj__7.net10 ),
    .A(\proj__7.net14 ),
    .B(\proj__7.net11 ));
 sg13g2_inv_1 \proj__7.not1/_0_  (.Y(\proj__7.net11 ),
    .A(net6));
 sg13g2_or2_1 \proj__7.or1/_0_  (.X(\proj__7.net12 ),
    .B(net1),
    .A(\proj__7.net13 ));
 sg13g2_xor2_1 \proj__7.xor1/_0_  (.B(net42),
    .A(net37),
    .X(\proj__7.net14 ));
 sg13g2_dfrbp_1 \proj__8.flop1/_1_  (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net153),
    .D(net2),
    .Q_N(\proj__8.flop1/notq ),
    .Q(\proj__8.net3 ));
 sg13g2_tiehi \proj__8.flop2/_1__142  (.L_HI(net154));
 sg13g2_dfrbp_1 \proj__8.flop2/_1_  (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net154),
    .D(net160),
    .Q_N(\proj__8.flop2/notq ),
    .Q(\proj__8.net5 ));
 sg13g2_tiehi \proj__8.flop3/_1__143  (.L_HI(net155));
 sg13g2_dfrbp_1 \proj__8.flop3/_1_  (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net155),
    .D(net161),
    .Q_N(\proj__8.flop3/notq ),
    .Q(\proj__8.net4 ));
 sg13g2_tiehi \proj__8.flop4/_1__144  (.L_HI(net156));
 sg13g2_dfrbp_1 \proj__8.flop4/_1_  (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net156),
    .D(net159),
    .Q_N(\proj__8.flop4/notq ),
    .Q(\proj__8.net6 ));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_buf_4 fanout37 (.X(net37),
    .A(net3));
 sg13g2_buf_2 fanout38 (.A(net39),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(ui_in[3]),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(net41),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(ui_in[2]),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(net43),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(ui_in[1]),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(net46),
    .X(net44));
 sg13g2_buf_1 fanout45 (.A(net46),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net2),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(net2),
    .X(net48));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_4 input7 (.X(net7),
    .A(uio_in[0]));
 sg13g2_buf_4 input8 (.X(net8),
    .A(uio_in[1]));
 sg13g2_buf_4 input9 (.X(net9),
    .A(uio_in[2]));
 sg13g2_buf_4 input10 (.X(net10),
    .A(uio_in[3]));
 sg13g2_tielo tt_um_wokwi_group_6_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_1_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_1_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_1__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\proj_13.net16 ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold2 (.A(\proj_12.net19 ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold3 (.A(\proj__8.net5 ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold4 (.A(\proj__8.net4 ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold5 (.A(\proj__8.net3 ),
    .X(net161));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_fill_1 FILLER_14_168 ();
 sg13g2_fill_2 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_227 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_decap_8 FILLER_14_262 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_8 FILLER_14_276 ();
 sg13g2_decap_8 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_decap_8 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_8 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_262 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_decap_8 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_283 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_decap_4 FILLER_16_111 ();
 sg13g2_fill_2 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_4 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_fill_2 FILLER_17_146 ();
 sg13g2_fill_1 FILLER_17_148 ();
 sg13g2_decap_4 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_167 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_decap_8 FILLER_17_174 ();
 sg13g2_decap_8 FILLER_17_181 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_260 ();
 sg13g2_decap_8 FILLER_17_267 ();
 sg13g2_decap_8 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_decap_8 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_302 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_316 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_344 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_155 ();
 sg13g2_decap_8 FILLER_18_162 ();
 sg13g2_decap_8 FILLER_18_169 ();
 sg13g2_decap_8 FILLER_18_176 ();
 sg13g2_decap_8 FILLER_18_183 ();
 sg13g2_decap_4 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_decap_8 FILLER_18_267 ();
 sg13g2_decap_8 FILLER_18_274 ();
 sg13g2_decap_8 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_288 ();
 sg13g2_decap_8 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_decap_8 FILLER_18_316 ();
 sg13g2_decap_8 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_18_337 ();
 sg13g2_decap_8 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_4 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_114 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_4 FILLER_19_133 ();
 sg13g2_fill_2 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_4 FILLER_20_144 ();
 sg13g2_fill_2 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_154 ();
 sg13g2_fill_1 FILLER_20_156 ();
 sg13g2_fill_2 FILLER_20_209 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_147 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_decap_4 FILLER_21_188 ();
 sg13g2_fill_2 FILLER_21_192 ();
 sg13g2_decap_8 FILLER_21_198 ();
 sg13g2_decap_8 FILLER_21_205 ();
 sg13g2_decap_8 FILLER_21_212 ();
 sg13g2_decap_8 FILLER_21_219 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_decap_4 FILLER_21_244 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_decap_4 FILLER_21_284 ();
 sg13g2_fill_2 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_4 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_269 ();
 sg13g2_decap_8 FILLER_22_276 ();
 sg13g2_decap_8 FILLER_22_283 ();
 sg13g2_decap_8 FILLER_22_290 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_334 ();
 sg13g2_fill_1 FILLER_22_336 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_4 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_decap_4 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_205 ();
 sg13g2_decap_8 FILLER_23_236 ();
 sg13g2_decap_8 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_250 ();
 sg13g2_decap_8 FILLER_23_257 ();
 sg13g2_decap_4 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_275 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_4 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_157 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_227 ();
 sg13g2_fill_1 FILLER_25_301 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_4 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_4 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_146 ();
 sg13g2_decap_8 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_decap_4 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_decap_4 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_4 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_219 ();
 sg13g2_decap_8 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_240 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_264 ();
 sg13g2_fill_2 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_fill_1 FILLER_26_376 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_decap_8 FILLER_27_149 ();
 sg13g2_fill_2 FILLER_27_156 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_decap_8 FILLER_27_244 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_4 FILLER_27_372 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_190 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_254 ();
 sg13g2_fill_2 FILLER_28_291 ();
 sg13g2_fill_2 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_fill_2 FILLER_28_375 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_366 ();
 sg13g2_decap_4 FILLER_29_373 ();
 sg13g2_fill_1 FILLER_29_377 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_69 ();
 sg13g2_decap_8 FILLER_30_76 ();
 sg13g2_fill_2 FILLER_30_83 ();
 sg13g2_decap_8 FILLER_30_89 ();
 sg13g2_decap_4 FILLER_30_96 ();
 sg13g2_fill_2 FILLER_30_100 ();
 sg13g2_decap_4 FILLER_30_188 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_229 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_fill_2 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_369 ();
 sg13g2_decap_8 FILLER_30_376 ();
 sg13g2_decap_4 FILLER_30_383 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_40 ();
 sg13g2_decap_4 FILLER_31_47 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_152 ();
 sg13g2_decap_8 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_4 FILLER_31_252 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_4 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_208 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_4 FILLER_32_249 ();
 sg13g2_decap_4 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_374 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_68 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_fill_1 FILLER_33_106 ();
 sg13g2_decap_4 FILLER_33_111 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_180 ();
 sg13g2_decap_4 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_197 ();
 sg13g2_decap_8 FILLER_33_241 ();
 sg13g2_decap_8 FILLER_33_248 ();
 sg13g2_decap_4 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_decap_4 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_344 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_39 ();
 sg13g2_decap_8 FILLER_34_46 ();
 sg13g2_decap_8 FILLER_34_53 ();
 sg13g2_decap_8 FILLER_34_60 ();
 sg13g2_decap_4 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_71 ();
 sg13g2_decap_8 FILLER_34_99 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_decap_4 FILLER_34_135 ();
 sg13g2_fill_1 FILLER_34_139 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_184 ();
 sg13g2_decap_8 FILLER_34_191 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_decap_4 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_253 ();
 sg13g2_decap_8 FILLER_34_260 ();
 sg13g2_decap_4 FILLER_34_267 ();
 sg13g2_decap_4 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_decap_8 FILLER_34_334 ();
 sg13g2_decap_8 FILLER_34_341 ();
 sg13g2_fill_2 FILLER_34_348 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_34 ();
 sg13g2_fill_2 FILLER_35_38 ();
 sg13g2_decap_8 FILLER_35_66 ();
 sg13g2_decap_4 FILLER_35_73 ();
 sg13g2_fill_1 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_104 ();
 sg13g2_decap_8 FILLER_35_111 ();
 sg13g2_fill_2 FILLER_35_118 ();
 sg13g2_decap_8 FILLER_35_124 ();
 sg13g2_decap_8 FILLER_35_131 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_decap_4 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_decap_8 FILLER_35_162 ();
 sg13g2_decap_8 FILLER_35_169 ();
 sg13g2_decap_8 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_183 ();
 sg13g2_decap_8 FILLER_35_190 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_decap_8 FILLER_35_204 ();
 sg13g2_decap_8 FILLER_35_211 ();
 sg13g2_decap_8 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_225 ();
 sg13g2_decap_4 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_262 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_fill_2 FILLER_35_276 ();
 sg13g2_fill_1 FILLER_35_278 ();
 sg13g2_decap_8 FILLER_35_299 ();
 sg13g2_decap_8 FILLER_35_306 ();
 sg13g2_fill_1 FILLER_35_313 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_18 ();
 sg13g2_decap_8 FILLER_36_23 ();
 sg13g2_decap_8 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_37 ();
 sg13g2_decap_8 FILLER_36_44 ();
 sg13g2_decap_8 FILLER_36_55 ();
 sg13g2_decap_8 FILLER_36_62 ();
 sg13g2_decap_8 FILLER_36_69 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_decap_8 FILLER_36_104 ();
 sg13g2_decap_8 FILLER_36_111 ();
 sg13g2_decap_8 FILLER_36_118 ();
 sg13g2_decap_8 FILLER_36_125 ();
 sg13g2_decap_8 FILLER_36_132 ();
 sg13g2_decap_8 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_decap_8 FILLER_36_160 ();
 sg13g2_decap_8 FILLER_36_167 ();
 sg13g2_decap_8 FILLER_36_174 ();
 sg13g2_decap_8 FILLER_36_181 ();
 sg13g2_decap_8 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_195 ();
 sg13g2_decap_8 FILLER_36_202 ();
 sg13g2_decap_8 FILLER_36_209 ();
 sg13g2_decap_8 FILLER_36_216 ();
 sg13g2_decap_8 FILLER_36_223 ();
 sg13g2_decap_8 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_fill_2 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_251 ();
 sg13g2_fill_2 FILLER_36_279 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_286 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_fill_2 FILLER_36_297 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_fill_1 FILLER_37_88 ();
 sg13g2_decap_8 FILLER_37_97 ();
 sg13g2_decap_8 FILLER_37_104 ();
 sg13g2_decap_8 FILLER_37_111 ();
 sg13g2_decap_8 FILLER_37_118 ();
 sg13g2_decap_8 FILLER_37_125 ();
 sg13g2_decap_8 FILLER_37_132 ();
 sg13g2_decap_8 FILLER_37_139 ();
 sg13g2_decap_8 FILLER_37_146 ();
 sg13g2_decap_8 FILLER_37_153 ();
 sg13g2_decap_8 FILLER_37_160 ();
 sg13g2_decap_8 FILLER_37_167 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_decap_8 FILLER_37_181 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_decap_8 FILLER_37_195 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_decap_8 FILLER_37_216 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_decap_8 FILLER_37_230 ();
 sg13g2_decap_8 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_251 ();
 sg13g2_decap_4 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_fill_1 FILLER_37_270 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net11;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_oe[7] = net18;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
 assign uio_out[6] = net25;
 assign uio_out[7] = net26;
endmodule

module tt_um_alphaonesoc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire clk_regs;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire \addr[0] ;
 wire \addr[10] ;
 wire \addr[11] ;
 wire \addr[12] ;
 wire \addr[13] ;
 wire \addr[14] ;
 wire \addr[15] ;
 wire \addr[16] ;
 wire \addr[17] ;
 wire \addr[18] ;
 wire \addr[19] ;
 wire \addr[1] ;
 wire \addr[20] ;
 wire \addr[21] ;
 wire \addr[22] ;
 wire \addr[23] ;
 wire \addr[24] ;
 wire \addr[25] ;
 wire \addr[26] ;
 wire \addr[27] ;
 wire \addr[2] ;
 wire \addr[3] ;
 wire \addr[4] ;
 wire \addr[5] ;
 wire \addr[6] ;
 wire \addr[7] ;
 wire \addr[8] ;
 wire \addr[9] ;
 wire \data_to_write[0] ;
 wire \data_to_write[10] ;
 wire \data_to_write[11] ;
 wire \data_to_write[12] ;
 wire \data_to_write[13] ;
 wire \data_to_write[14] ;
 wire \data_to_write[15] ;
 wire \data_to_write[16] ;
 wire \data_to_write[17] ;
 wire \data_to_write[18] ;
 wire \data_to_write[19] ;
 wire \data_to_write[1] ;
 wire \data_to_write[20] ;
 wire \data_to_write[21] ;
 wire \data_to_write[22] ;
 wire \data_to_write[23] ;
 wire \data_to_write[24] ;
 wire \data_to_write[25] ;
 wire \data_to_write[26] ;
 wire \data_to_write[27] ;
 wire \data_to_write[28] ;
 wire \data_to_write[29] ;
 wire \data_to_write[2] ;
 wire \data_to_write[30] ;
 wire \data_to_write[31] ;
 wire \data_to_write[3] ;
 wire \data_to_write[4] ;
 wire \data_to_write[5] ;
 wire \data_to_write[6] ;
 wire \data_to_write[7] ;
 wire \data_to_write[8] ;
 wire \data_to_write[9] ;
 wire debug_data_continue;
 wire debug_instr_valid;
 wire \debug_rd[0] ;
 wire \debug_rd[1] ;
 wire \debug_rd[2] ;
 wire \debug_rd[3] ;
 wire \debug_rd_r[0] ;
 wire \debug_rd_r[1] ;
 wire \debug_rd_r[2] ;
 wire \debug_rd_r[3] ;
 wire debug_register_data;
 wire debug_uart_txd;
 wire \gpio_out[0] ;
 wire \gpio_out[1] ;
 wire \gpio_out[2] ;
 wire \gpio_out[3] ;
 wire \gpio_out[4] ;
 wire \gpio_out[5] ;
 wire \gpio_out[6] ;
 wire \gpio_out[7] ;
 wire \gpio_out_sel[0] ;
 wire \gpio_out_sel[1] ;
 wire \gpio_out_sel[2] ;
 wire \gpio_out_sel[3] ;
 wire \gpio_out_sel[4] ;
 wire \gpio_out_sel[5] ;
 wire \gpio_out_sel[6] ;
 wire \gpio_out_sel[7] ;
 wire \i_core.cpu.additional_mem_ops[0] ;
 wire \i_core.cpu.additional_mem_ops[1] ;
 wire \i_core.cpu.additional_mem_ops[2] ;
 wire \i_core.cpu.alu_op[0] ;
 wire \i_core.cpu.alu_op[1] ;
 wire \i_core.cpu.alu_op[2] ;
 wire \i_core.cpu.alu_op[3] ;
 wire \i_core.cpu.counter[2] ;
 wire \i_core.cpu.counter[3] ;
 wire \i_core.cpu.counter[4] ;
 wire \i_core.cpu.data_read_n[0] ;
 wire \i_core.cpu.data_read_n[1] ;
 wire \i_core.cpu.data_ready_core ;
 wire \i_core.cpu.data_ready_latch ;
 wire \i_core.cpu.data_write_n[0] ;
 wire \i_core.cpu.data_write_n[1] ;
 wire \i_core.cpu.i_core.cmp ;
 wire \i_core.cpu.i_core.cmp_out ;
 wire \i_core.cpu.i_core.cy ;
 wire \i_core.cpu.i_core.cy_out ;
 wire \i_core.cpu.i_core.cycle[0] ;
 wire \i_core.cpu.i_core.cycle[1] ;
 wire \i_core.cpu.i_core.cycle_count[0] ;
 wire \i_core.cpu.i_core.cycle_count[1] ;
 wire \i_core.cpu.i_core.cycle_count[2] ;
 wire \i_core.cpu.i_core.cycle_count[3] ;
 wire \i_core.cpu.i_core.i_cycles.cy ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_cycles.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_cycles.rstn ;
 wire \i_core.cpu.i_core.i_instrret.add ;
 wire \i_core.cpu.i_core.i_instrret.cy ;
 wire \i_core.cpu.i_core.i_instrret.data[0] ;
 wire \i_core.cpu.i_core.i_instrret.data[1] ;
 wire \i_core.cpu.i_core.i_instrret.data[2] ;
 wire \i_core.cpu.i_core.i_instrret.data[3] ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_instrret.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[10].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[11].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[12].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[13].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[14].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[15].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[16].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[17].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[18].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[19].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[20].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[21].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[22].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[23].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[24].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[25].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[26].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[27].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[28].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[29].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[30].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[31].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[4].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[5].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[6].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[7].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[8].A ;
 wire \i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[9].A ;
 wire \i_core.cpu.i_core.i_registers.rd[0] ;
 wire \i_core.cpu.i_core.i_registers.rd[1] ;
 wire \i_core.cpu.i_core.i_registers.rd[2] ;
 wire \i_core.cpu.i_core.i_registers.rd[3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[10][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[10][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[10][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[10][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[11][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[11][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[11][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[11][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[12][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[12][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[12][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[12][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[13][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[13][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[13][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[13][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[14][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[14][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[14][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[14][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[15][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[15][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[15][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[15][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[1][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[1][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[1][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[1][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[2][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[2][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[2][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[2][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[5][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[5][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[5][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[5][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[6][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[6][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[6][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[6][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[7][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[7][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[7][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[7][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[8][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[8][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[8][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[8][3] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[9][0] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[9][1] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[9][2] ;
 wire \i_core.cpu.i_core.i_registers.reg_access[9][3] ;
 wire \i_core.cpu.i_core.i_registers.rs1[0] ;
 wire \i_core.cpu.i_core.i_registers.rs1[1] ;
 wire \i_core.cpu.i_core.i_registers.rs1[2] ;
 wire \i_core.cpu.i_core.i_registers.rs1[3] ;
 wire \i_core.cpu.i_core.i_registers.rs2[0] ;
 wire \i_core.cpu.i_core.i_registers.rs2[1] ;
 wire \i_core.cpu.i_core.i_registers.rs2[2] ;
 wire \i_core.cpu.i_core.i_registers.rs2[3] ;
 wire \i_core.cpu.i_core.i_shift.a[0] ;
 wire \i_core.cpu.i_core.i_shift.a[10] ;
 wire \i_core.cpu.i_core.i_shift.a[11] ;
 wire \i_core.cpu.i_core.i_shift.a[12] ;
 wire \i_core.cpu.i_core.i_shift.a[13] ;
 wire \i_core.cpu.i_core.i_shift.a[14] ;
 wire \i_core.cpu.i_core.i_shift.a[15] ;
 wire \i_core.cpu.i_core.i_shift.a[16] ;
 wire \i_core.cpu.i_core.i_shift.a[17] ;
 wire \i_core.cpu.i_core.i_shift.a[18] ;
 wire \i_core.cpu.i_core.i_shift.a[19] ;
 wire \i_core.cpu.i_core.i_shift.a[1] ;
 wire \i_core.cpu.i_core.i_shift.a[20] ;
 wire \i_core.cpu.i_core.i_shift.a[21] ;
 wire \i_core.cpu.i_core.i_shift.a[22] ;
 wire \i_core.cpu.i_core.i_shift.a[23] ;
 wire \i_core.cpu.i_core.i_shift.a[24] ;
 wire \i_core.cpu.i_core.i_shift.a[25] ;
 wire \i_core.cpu.i_core.i_shift.a[26] ;
 wire \i_core.cpu.i_core.i_shift.a[27] ;
 wire \i_core.cpu.i_core.i_shift.a[28] ;
 wire \i_core.cpu.i_core.i_shift.a[29] ;
 wire \i_core.cpu.i_core.i_shift.a[2] ;
 wire \i_core.cpu.i_core.i_shift.a[30] ;
 wire \i_core.cpu.i_core.i_shift.a[31] ;
 wire \i_core.cpu.i_core.i_shift.a[3] ;
 wire \i_core.cpu.i_core.i_shift.a[4] ;
 wire \i_core.cpu.i_core.i_shift.a[5] ;
 wire \i_core.cpu.i_core.i_shift.a[6] ;
 wire \i_core.cpu.i_core.i_shift.a[7] ;
 wire \i_core.cpu.i_core.i_shift.a[8] ;
 wire \i_core.cpu.i_core.i_shift.a[9] ;
 wire \i_core.cpu.i_core.i_shift.adjusted_shift_amt[0] ;
 wire \i_core.cpu.i_core.i_shift.adjusted_shift_amt[1] ;
 wire \i_core.cpu.i_core.i_shift.b[2] ;
 wire \i_core.cpu.i_core.i_shift.b[3] ;
 wire \i_core.cpu.i_core.i_shift.b[4] ;
 wire \i_core.cpu.i_core.imm_lo[0] ;
 wire \i_core.cpu.i_core.imm_lo[10] ;
 wire \i_core.cpu.i_core.imm_lo[11] ;
 wire \i_core.cpu.i_core.imm_lo[1] ;
 wire \i_core.cpu.i_core.imm_lo[2] ;
 wire \i_core.cpu.i_core.imm_lo[3] ;
 wire \i_core.cpu.i_core.imm_lo[4] ;
 wire \i_core.cpu.i_core.imm_lo[5] ;
 wire \i_core.cpu.i_core.imm_lo[6] ;
 wire \i_core.cpu.i_core.imm_lo[7] ;
 wire \i_core.cpu.i_core.imm_lo[8] ;
 wire \i_core.cpu.i_core.imm_lo[9] ;
 wire \i_core.cpu.i_core.interrupt_req[0] ;
 wire \i_core.cpu.i_core.interrupt_req[1] ;
 wire \i_core.cpu.i_core.is_double_fault_r ;
 wire \i_core.cpu.i_core.is_interrupt ;
 wire \i_core.cpu.i_core.last_interrupt_req[0] ;
 wire \i_core.cpu.i_core.last_interrupt_req[1] ;
 wire \i_core.cpu.i_core.load_done ;
 wire \i_core.cpu.i_core.load_top_bit ;
 wire \i_core.cpu.i_core.mcause[0] ;
 wire \i_core.cpu.i_core.mcause[1] ;
 wire \i_core.cpu.i_core.mcause[3] ;
 wire \i_core.cpu.i_core.mcause[4] ;
 wire \i_core.cpu.i_core.mem_op[0] ;
 wire \i_core.cpu.i_core.mem_op[1] ;
 wire \i_core.cpu.i_core.mem_op[2] ;
 wire \i_core.cpu.i_core.mepc[0] ;
 wire \i_core.cpu.i_core.mepc[10] ;
 wire \i_core.cpu.i_core.mepc[11] ;
 wire \i_core.cpu.i_core.mepc[12] ;
 wire \i_core.cpu.i_core.mepc[13] ;
 wire \i_core.cpu.i_core.mepc[14] ;
 wire \i_core.cpu.i_core.mepc[15] ;
 wire \i_core.cpu.i_core.mepc[16] ;
 wire \i_core.cpu.i_core.mepc[17] ;
 wire \i_core.cpu.i_core.mepc[18] ;
 wire \i_core.cpu.i_core.mepc[19] ;
 wire \i_core.cpu.i_core.mepc[1] ;
 wire \i_core.cpu.i_core.mepc[20] ;
 wire \i_core.cpu.i_core.mepc[21] ;
 wire \i_core.cpu.i_core.mepc[22] ;
 wire \i_core.cpu.i_core.mepc[23] ;
 wire \i_core.cpu.i_core.mepc[2] ;
 wire \i_core.cpu.i_core.mepc[3] ;
 wire \i_core.cpu.i_core.mepc[4] ;
 wire \i_core.cpu.i_core.mepc[5] ;
 wire \i_core.cpu.i_core.mepc[6] ;
 wire \i_core.cpu.i_core.mepc[7] ;
 wire \i_core.cpu.i_core.mepc[8] ;
 wire \i_core.cpu.i_core.mepc[9] ;
 wire \i_core.cpu.i_core.mie[16] ;
 wire \i_core.cpu.i_core.mie[17] ;
 wire \i_core.cpu.i_core.mie[18] ;
 wire \i_core.cpu.i_core.mie[19] ;
 wire \i_core.cpu.i_core.mip[16] ;
 wire \i_core.cpu.i_core.mip[17] ;
 wire \i_core.cpu.i_core.mstatus_mie ;
 wire \i_core.cpu.i_core.mstatus_mpie ;
 wire \i_core.cpu.i_core.mstatus_mte ;
 wire \i_core.cpu.i_core.multiplier.accum[0] ;
 wire \i_core.cpu.i_core.multiplier.accum[10] ;
 wire \i_core.cpu.i_core.multiplier.accum[11] ;
 wire \i_core.cpu.i_core.multiplier.accum[12] ;
 wire \i_core.cpu.i_core.multiplier.accum[13] ;
 wire \i_core.cpu.i_core.multiplier.accum[14] ;
 wire \i_core.cpu.i_core.multiplier.accum[15] ;
 wire \i_core.cpu.i_core.multiplier.accum[1] ;
 wire \i_core.cpu.i_core.multiplier.accum[2] ;
 wire \i_core.cpu.i_core.multiplier.accum[3] ;
 wire \i_core.cpu.i_core.multiplier.accum[4] ;
 wire \i_core.cpu.i_core.multiplier.accum[5] ;
 wire \i_core.cpu.i_core.multiplier.accum[6] ;
 wire \i_core.cpu.i_core.multiplier.accum[7] ;
 wire \i_core.cpu.i_core.multiplier.accum[8] ;
 wire \i_core.cpu.i_core.multiplier.accum[9] ;
 wire \i_core.cpu.i_core.time_hi[0] ;
 wire \i_core.cpu.i_core.time_hi[1] ;
 wire \i_core.cpu.i_core.time_hi[2] ;
 wire \i_core.cpu.imm[12] ;
 wire \i_core.cpu.imm[13] ;
 wire \i_core.cpu.imm[14] ;
 wire \i_core.cpu.imm[15] ;
 wire \i_core.cpu.imm[16] ;
 wire \i_core.cpu.imm[17] ;
 wire \i_core.cpu.imm[18] ;
 wire \i_core.cpu.imm[19] ;
 wire \i_core.cpu.imm[20] ;
 wire \i_core.cpu.imm[21] ;
 wire \i_core.cpu.imm[22] ;
 wire \i_core.cpu.imm[23] ;
 wire \i_core.cpu.imm[24] ;
 wire \i_core.cpu.imm[25] ;
 wire \i_core.cpu.imm[26] ;
 wire \i_core.cpu.imm[27] ;
 wire \i_core.cpu.imm[28] ;
 wire \i_core.cpu.imm[29] ;
 wire \i_core.cpu.imm[30] ;
 wire \i_core.cpu.imm[31] ;
 wire \i_core.cpu.instr_data[0][0] ;
 wire \i_core.cpu.instr_data[0][10] ;
 wire \i_core.cpu.instr_data[0][11] ;
 wire \i_core.cpu.instr_data[0][12] ;
 wire \i_core.cpu.instr_data[0][13] ;
 wire \i_core.cpu.instr_data[0][14] ;
 wire \i_core.cpu.instr_data[0][15] ;
 wire \i_core.cpu.instr_data[0][1] ;
 wire \i_core.cpu.instr_data[0][2] ;
 wire \i_core.cpu.instr_data[0][3] ;
 wire \i_core.cpu.instr_data[0][4] ;
 wire \i_core.cpu.instr_data[0][5] ;
 wire \i_core.cpu.instr_data[0][6] ;
 wire \i_core.cpu.instr_data[0][7] ;
 wire \i_core.cpu.instr_data[0][8] ;
 wire \i_core.cpu.instr_data[0][9] ;
 wire \i_core.cpu.instr_data[1][0] ;
 wire \i_core.cpu.instr_data[1][10] ;
 wire \i_core.cpu.instr_data[1][11] ;
 wire \i_core.cpu.instr_data[1][12] ;
 wire \i_core.cpu.instr_data[1][13] ;
 wire \i_core.cpu.instr_data[1][14] ;
 wire \i_core.cpu.instr_data[1][15] ;
 wire \i_core.cpu.instr_data[1][1] ;
 wire \i_core.cpu.instr_data[1][2] ;
 wire \i_core.cpu.instr_data[1][3] ;
 wire \i_core.cpu.instr_data[1][4] ;
 wire \i_core.cpu.instr_data[1][5] ;
 wire \i_core.cpu.instr_data[1][6] ;
 wire \i_core.cpu.instr_data[1][7] ;
 wire \i_core.cpu.instr_data[1][8] ;
 wire \i_core.cpu.instr_data[1][9] ;
 wire \i_core.cpu.instr_data[2][0] ;
 wire \i_core.cpu.instr_data[2][10] ;
 wire \i_core.cpu.instr_data[2][11] ;
 wire \i_core.cpu.instr_data[2][12] ;
 wire \i_core.cpu.instr_data[2][13] ;
 wire \i_core.cpu.instr_data[2][14] ;
 wire \i_core.cpu.instr_data[2][15] ;
 wire \i_core.cpu.instr_data[2][1] ;
 wire \i_core.cpu.instr_data[2][2] ;
 wire \i_core.cpu.instr_data[2][3] ;
 wire \i_core.cpu.instr_data[2][4] ;
 wire \i_core.cpu.instr_data[2][5] ;
 wire \i_core.cpu.instr_data[2][6] ;
 wire \i_core.cpu.instr_data[2][7] ;
 wire \i_core.cpu.instr_data[2][8] ;
 wire \i_core.cpu.instr_data[2][9] ;
 wire \i_core.cpu.instr_data[3][0] ;
 wire \i_core.cpu.instr_data[3][10] ;
 wire \i_core.cpu.instr_data[3][11] ;
 wire \i_core.cpu.instr_data[3][12] ;
 wire \i_core.cpu.instr_data[3][13] ;
 wire \i_core.cpu.instr_data[3][14] ;
 wire \i_core.cpu.instr_data[3][15] ;
 wire \i_core.cpu.instr_data[3][1] ;
 wire \i_core.cpu.instr_data[3][2] ;
 wire \i_core.cpu.instr_data[3][3] ;
 wire \i_core.cpu.instr_data[3][4] ;
 wire \i_core.cpu.instr_data[3][5] ;
 wire \i_core.cpu.instr_data[3][6] ;
 wire \i_core.cpu.instr_data[3][7] ;
 wire \i_core.cpu.instr_data[3][8] ;
 wire \i_core.cpu.instr_data[3][9] ;
 wire \i_core.cpu.instr_data_in[0] ;
 wire \i_core.cpu.instr_data_in[10] ;
 wire \i_core.cpu.instr_data_in[11] ;
 wire \i_core.cpu.instr_data_in[12] ;
 wire \i_core.cpu.instr_data_in[13] ;
 wire \i_core.cpu.instr_data_in[14] ;
 wire \i_core.cpu.instr_data_in[15] ;
 wire \i_core.cpu.instr_data_in[1] ;
 wire \i_core.cpu.instr_data_in[2] ;
 wire \i_core.cpu.instr_data_in[3] ;
 wire \i_core.cpu.instr_data_in[4] ;
 wire \i_core.cpu.instr_data_in[5] ;
 wire \i_core.cpu.instr_data_in[6] ;
 wire \i_core.cpu.instr_data_in[7] ;
 wire \i_core.cpu.instr_data_in[8] ;
 wire \i_core.cpu.instr_data_in[9] ;
 wire \i_core.cpu.instr_data_start[10] ;
 wire \i_core.cpu.instr_data_start[11] ;
 wire \i_core.cpu.instr_data_start[12] ;
 wire \i_core.cpu.instr_data_start[13] ;
 wire \i_core.cpu.instr_data_start[14] ;
 wire \i_core.cpu.instr_data_start[15] ;
 wire \i_core.cpu.instr_data_start[16] ;
 wire \i_core.cpu.instr_data_start[17] ;
 wire \i_core.cpu.instr_data_start[18] ;
 wire \i_core.cpu.instr_data_start[19] ;
 wire \i_core.cpu.instr_data_start[20] ;
 wire \i_core.cpu.instr_data_start[21] ;
 wire \i_core.cpu.instr_data_start[22] ;
 wire \i_core.cpu.instr_data_start[23] ;
 wire \i_core.cpu.instr_data_start[3] ;
 wire \i_core.cpu.instr_data_start[4] ;
 wire \i_core.cpu.instr_data_start[5] ;
 wire \i_core.cpu.instr_data_start[6] ;
 wire \i_core.cpu.instr_data_start[7] ;
 wire \i_core.cpu.instr_data_start[8] ;
 wire \i_core.cpu.instr_data_start[9] ;
 wire \i_core.cpu.instr_fetch_running ;
 wire \i_core.cpu.instr_fetch_started ;
 wire \i_core.cpu.instr_fetch_stopped ;
 wire \i_core.cpu.instr_len[1] ;
 wire \i_core.cpu.instr_len[2] ;
 wire \i_core.cpu.instr_write_offset[1] ;
 wire \i_core.cpu.instr_write_offset[2] ;
 wire \i_core.cpu.instr_write_offset[3] ;
 wire \i_core.cpu.is_alu_imm ;
 wire \i_core.cpu.is_alu_reg ;
 wire \i_core.cpu.is_auipc ;
 wire \i_core.cpu.is_branch ;
 wire \i_core.cpu.is_jal ;
 wire \i_core.cpu.is_jalr ;
 wire \i_core.cpu.is_load ;
 wire \i_core.cpu.is_lui ;
 wire \i_core.cpu.is_store ;
 wire \i_core.cpu.is_system ;
 wire \i_core.cpu.load_started ;
 wire \i_core.cpu.mem_op_increment_reg ;
 wire \i_core.cpu.no_write_in_progress ;
 wire \i_core.cpu.pc[1] ;
 wire \i_core.cpu.pc[2] ;
 wire \i_core.cpu.was_early_branch ;
 wire \i_core.mem.data_from_read[16] ;
 wire \i_core.mem.data_from_read[17] ;
 wire \i_core.mem.data_from_read[18] ;
 wire \i_core.mem.data_from_read[19] ;
 wire \i_core.mem.data_from_read[20] ;
 wire \i_core.mem.data_from_read[21] ;
 wire \i_core.mem.data_from_read[22] ;
 wire \i_core.mem.data_from_read[23] ;
 wire \i_core.mem.data_stall ;
 wire \i_core.mem.instr_active ;
 wire \i_core.mem.q_ctrl.addr[0] ;
 wire \i_core.mem.q_ctrl.addr[10] ;
 wire \i_core.mem.q_ctrl.addr[11] ;
 wire \i_core.mem.q_ctrl.addr[12] ;
 wire \i_core.mem.q_ctrl.addr[13] ;
 wire \i_core.mem.q_ctrl.addr[14] ;
 wire \i_core.mem.q_ctrl.addr[15] ;
 wire \i_core.mem.q_ctrl.addr[16] ;
 wire \i_core.mem.q_ctrl.addr[17] ;
 wire \i_core.mem.q_ctrl.addr[18] ;
 wire \i_core.mem.q_ctrl.addr[19] ;
 wire \i_core.mem.q_ctrl.addr[1] ;
 wire \i_core.mem.q_ctrl.addr[20] ;
 wire \i_core.mem.q_ctrl.addr[21] ;
 wire \i_core.mem.q_ctrl.addr[22] ;
 wire \i_core.mem.q_ctrl.addr[23] ;
 wire \i_core.mem.q_ctrl.addr[2] ;
 wire \i_core.mem.q_ctrl.addr[3] ;
 wire \i_core.mem.q_ctrl.addr[4] ;
 wire \i_core.mem.q_ctrl.addr[5] ;
 wire \i_core.mem.q_ctrl.addr[6] ;
 wire \i_core.mem.q_ctrl.addr[7] ;
 wire \i_core.mem.q_ctrl.addr[8] ;
 wire \i_core.mem.q_ctrl.addr[9] ;
 wire \i_core.mem.q_ctrl.data_ready ;
 wire \i_core.mem.q_ctrl.data_req ;
 wire \i_core.mem.q_ctrl.delay_cycles_cfg[0] ;
 wire \i_core.mem.q_ctrl.delay_cycles_cfg[1] ;
 wire \i_core.mem.q_ctrl.delay_cycles_cfg[2] ;
 wire \i_core.mem.q_ctrl.fsm_state[0] ;
 wire \i_core.mem.q_ctrl.fsm_state[1] ;
 wire \i_core.mem.q_ctrl.fsm_state[2] ;
 wire \i_core.mem.q_ctrl.is_writing ;
 wire \i_core.mem.q_ctrl.last_ram_a_sel ;
 wire \i_core.mem.q_ctrl.last_ram_b_sel ;
 wire \i_core.mem.q_ctrl.nibbles_remaining[0] ;
 wire \i_core.mem.q_ctrl.nibbles_remaining[1] ;
 wire \i_core.mem.q_ctrl.nibbles_remaining[2] ;
 wire \i_core.mem.q_ctrl.read_cycles_count[0] ;
 wire \i_core.mem.q_ctrl.read_cycles_count[1] ;
 wire \i_core.mem.q_ctrl.read_cycles_count[2] ;
 wire \i_core.mem.q_ctrl.rstn ;
 wire \i_core.mem.q_ctrl.spi_clk_out ;
 wire \i_core.mem.q_ctrl.spi_data_oe[0] ;
 wire \i_core.mem.q_ctrl.spi_flash_select ;
 wire \i_core.mem.q_ctrl.spi_in_buffer[0] ;
 wire \i_core.mem.q_ctrl.spi_in_buffer[1] ;
 wire \i_core.mem.q_ctrl.spi_in_buffer[2] ;
 wire \i_core.mem.q_ctrl.spi_in_buffer[3] ;
 wire \i_core.mem.q_ctrl.spi_in_buffer[4] ;
 wire \i_core.mem.q_ctrl.spi_in_buffer[5] ;
 wire \i_core.mem.q_ctrl.spi_in_buffer[6] ;
 wire \i_core.mem.q_ctrl.spi_in_buffer[7] ;
 wire \i_core.mem.q_ctrl.spi_ram_a_select ;
 wire \i_core.mem.q_ctrl.spi_ram_b_select ;
 wire \i_core.mem.q_ctrl.stop_txn_reg ;
 wire \i_core.mem.qspi_data_buf[10] ;
 wire \i_core.mem.qspi_data_buf[11] ;
 wire \i_core.mem.qspi_data_buf[12] ;
 wire \i_core.mem.qspi_data_buf[13] ;
 wire \i_core.mem.qspi_data_buf[14] ;
 wire \i_core.mem.qspi_data_buf[15] ;
 wire \i_core.mem.qspi_data_buf[24] ;
 wire \i_core.mem.qspi_data_buf[25] ;
 wire \i_core.mem.qspi_data_buf[26] ;
 wire \i_core.mem.qspi_data_buf[27] ;
 wire \i_core.mem.qspi_data_buf[28] ;
 wire \i_core.mem.qspi_data_buf[29] ;
 wire \i_core.mem.qspi_data_buf[30] ;
 wire \i_core.mem.qspi_data_buf[31] ;
 wire \i_core.mem.qspi_data_buf[8] ;
 wire \i_core.mem.qspi_data_buf[9] ;
 wire \i_core.mem.qspi_data_byte_idx[0] ;
 wire \i_core.mem.qspi_data_byte_idx[1] ;
 wire \i_core.mem.qspi_write_done ;
 wire \i_debug_uart_tx.cycle_counter[0] ;
 wire \i_debug_uart_tx.cycle_counter[1] ;
 wire \i_debug_uart_tx.cycle_counter[2] ;
 wire \i_debug_uart_tx.cycle_counter[3] ;
 wire \i_debug_uart_tx.cycle_counter[4] ;
 wire \i_debug_uart_tx.data_to_send[0] ;
 wire \i_debug_uart_tx.data_to_send[1] ;
 wire \i_debug_uart_tx.data_to_send[2] ;
 wire \i_debug_uart_tx.data_to_send[3] ;
 wire \i_debug_uart_tx.data_to_send[4] ;
 wire \i_debug_uart_tx.data_to_send[5] ;
 wire \i_debug_uart_tx.data_to_send[6] ;
 wire \i_debug_uart_tx.data_to_send[7] ;
 wire \i_debug_uart_tx.fsm_state[0] ;
 wire \i_debug_uart_tx.fsm_state[1] ;
 wire \i_debug_uart_tx.fsm_state[2] ;
 wire \i_debug_uart_tx.fsm_state[3] ;
 wire \i_spi.bits_remaining[0] ;
 wire \i_spi.bits_remaining[1] ;
 wire \i_spi.bits_remaining[2] ;
 wire \i_spi.bits_remaining[3] ;
 wire \i_spi.busy ;
 wire \i_spi.clock_count[0] ;
 wire \i_spi.clock_count[1] ;
 wire \i_spi.clock_divider[0] ;
 wire \i_spi.clock_divider[1] ;
 wire \i_spi.data[0] ;
 wire \i_spi.data[1] ;
 wire \i_spi.data[2] ;
 wire \i_spi.data[3] ;
 wire \i_spi.data[4] ;
 wire \i_spi.data[5] ;
 wire \i_spi.data[6] ;
 wire \i_spi.data[7] ;
 wire \i_spi.end_txn_reg ;
 wire \i_spi.read_latency ;
 wire \i_spi.spi_clk_out ;
 wire \i_spi.spi_dc ;
 wire \i_spi.spi_select ;
 wire \i_uart_rx.bit_sample ;
 wire \i_uart_rx.cycle_counter[0] ;
 wire \i_uart_rx.cycle_counter[10] ;
 wire \i_uart_rx.cycle_counter[1] ;
 wire \i_uart_rx.cycle_counter[2] ;
 wire \i_uart_rx.cycle_counter[3] ;
 wire \i_uart_rx.cycle_counter[4] ;
 wire \i_uart_rx.cycle_counter[5] ;
 wire \i_uart_rx.cycle_counter[6] ;
 wire \i_uart_rx.cycle_counter[7] ;
 wire \i_uart_rx.cycle_counter[8] ;
 wire \i_uart_rx.cycle_counter[9] ;
 wire \i_uart_rx.fsm_state[0] ;
 wire \i_uart_rx.fsm_state[1] ;
 wire \i_uart_rx.fsm_state[2] ;
 wire \i_uart_rx.fsm_state[3] ;
 wire \i_uart_rx.recieved_data[0] ;
 wire \i_uart_rx.recieved_data[1] ;
 wire \i_uart_rx.recieved_data[2] ;
 wire \i_uart_rx.recieved_data[3] ;
 wire \i_uart_rx.recieved_data[4] ;
 wire \i_uart_rx.recieved_data[5] ;
 wire \i_uart_rx.recieved_data[6] ;
 wire \i_uart_rx.recieved_data[7] ;
 wire \i_uart_rx.rxd_reg[0] ;
 wire \i_uart_rx.rxd_reg[1] ;
 wire \i_uart_rx.uart_rts ;
 wire \i_uart_tx.cycle_counter[0] ;
 wire \i_uart_tx.cycle_counter[10] ;
 wire \i_uart_tx.cycle_counter[1] ;
 wire \i_uart_tx.cycle_counter[2] ;
 wire \i_uart_tx.cycle_counter[3] ;
 wire \i_uart_tx.cycle_counter[4] ;
 wire \i_uart_tx.cycle_counter[5] ;
 wire \i_uart_tx.cycle_counter[6] ;
 wire \i_uart_tx.cycle_counter[7] ;
 wire \i_uart_tx.cycle_counter[8] ;
 wire \i_uart_tx.cycle_counter[9] ;
 wire \i_uart_tx.data_to_send[0] ;
 wire \i_uart_tx.data_to_send[1] ;
 wire \i_uart_tx.data_to_send[2] ;
 wire \i_uart_tx.data_to_send[3] ;
 wire \i_uart_tx.data_to_send[4] ;
 wire \i_uart_tx.data_to_send[5] ;
 wire \i_uart_tx.data_to_send[6] ;
 wire \i_uart_tx.data_to_send[7] ;
 wire \i_uart_tx.fsm_state[0] ;
 wire \i_uart_tx.fsm_state[1] ;
 wire \i_uart_tx.fsm_state[2] ;
 wire \i_uart_tx.fsm_state[3] ;
 wire \i_uart_tx.txd_reg ;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_57_clk_regs;
 wire clknet_leaf_58_clk_regs;
 wire clknet_leaf_59_clk_regs;
 wire clknet_leaf_60_clk_regs;
 wire clknet_leaf_61_clk_regs;
 wire clknet_leaf_62_clk_regs;
 wire clknet_leaf_63_clk_regs;
 wire clknet_leaf_64_clk_regs;
 wire clknet_leaf_65_clk_regs;
 wire clknet_leaf_66_clk_regs;
 wire clknet_leaf_67_clk_regs;
 wire clknet_leaf_68_clk_regs;
 wire clknet_leaf_69_clk_regs;
 wire clknet_leaf_70_clk_regs;
 wire clknet_leaf_71_clk_regs;
 wire clknet_leaf_72_clk_regs;
 wire clknet_leaf_73_clk_regs;
 wire clknet_leaf_74_clk_regs;
 wire clknet_leaf_75_clk_regs;
 wire clknet_leaf_76_clk_regs;
 wire clknet_leaf_77_clk_regs;
 wire clknet_leaf_78_clk_regs;
 wire clknet_leaf_79_clk_regs;
 wire clknet_leaf_80_clk_regs;
 wire clknet_leaf_81_clk_regs;
 wire clknet_leaf_82_clk_regs;
 wire clknet_leaf_83_clk_regs;
 wire clknet_leaf_84_clk_regs;
 wire clknet_leaf_85_clk_regs;
 wire clknet_leaf_86_clk_regs;
 wire clknet_leaf_87_clk_regs;
 wire clknet_leaf_88_clk_regs;
 wire clknet_leaf_89_clk_regs;
 wire clknet_leaf_90_clk_regs;
 wire clknet_leaf_91_clk_regs;
 wire clknet_leaf_92_clk_regs;
 wire clknet_leaf_93_clk_regs;
 wire clknet_leaf_94_clk_regs;
 wire clknet_leaf_95_clk_regs;
 wire clknet_leaf_96_clk_regs;
 wire clknet_leaf_97_clk_regs;
 wire clknet_leaf_98_clk_regs;
 wire clknet_leaf_99_clk_regs;
 wire clknet_leaf_100_clk_regs;
 wire clknet_leaf_101_clk_regs;
 wire clknet_leaf_102_clk_regs;
 wire clknet_leaf_103_clk_regs;
 wire clknet_leaf_104_clk_regs;
 wire clknet_leaf_105_clk_regs;
 wire clknet_leaf_106_clk_regs;
 wire clknet_leaf_107_clk_regs;
 wire clknet_leaf_108_clk_regs;
 wire clknet_leaf_109_clk_regs;
 wire clknet_leaf_110_clk_regs;
 wire clknet_leaf_111_clk_regs;
 wire clknet_leaf_112_clk_regs;
 wire clknet_leaf_113_clk_regs;
 wire clknet_leaf_114_clk_regs;
 wire clknet_leaf_115_clk_regs;
 wire clknet_leaf_116_clk_regs;
 wire clknet_leaf_117_clk_regs;
 wire clknet_leaf_118_clk_regs;
 wire clknet_leaf_119_clk_regs;
 wire clknet_leaf_120_clk_regs;
 wire clknet_leaf_121_clk_regs;
 wire clknet_leaf_122_clk_regs;
 wire clknet_leaf_123_clk_regs;
 wire clknet_leaf_124_clk_regs;
 wire clknet_leaf_125_clk_regs;
 wire clknet_leaf_126_clk_regs;
 wire clknet_leaf_128_clk_regs;
 wire clknet_leaf_129_clk_regs;
 wire clknet_leaf_130_clk_regs;
 wire clknet_leaf_131_clk_regs;
 wire clknet_leaf_132_clk_regs;
 wire clknet_leaf_133_clk_regs;
 wire clknet_leaf_134_clk_regs;
 wire clknet_leaf_135_clk_regs;
 wire clknet_leaf_136_clk_regs;
 wire clknet_leaf_137_clk_regs;
 wire clknet_leaf_138_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire delaynet_1_clk;
 wire delaynet_2_clk;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;

 sg13g2_inv_4 _05945_ (.A(net1393),
    .Y(_00747_));
 sg13g2_inv_1 _05946_ (.Y(_00748_),
    .A(net2320));
 sg13g2_inv_1 _05947_ (.Y(_00749_),
    .A(\i_core.cpu.additional_mem_ops[0] ));
 sg13g2_inv_1 _05948_ (.Y(_00750_),
    .A(net2262));
 sg13g2_inv_1 _05949_ (.Y(_00751_),
    .A(\i_core.cpu.is_jalr ));
 sg13g2_inv_1 _05950_ (.Y(_00752_),
    .A(net2486));
 sg13g2_inv_1 _05951_ (.Y(_00753_),
    .A(\i_core.cpu.is_auipc ));
 sg13g2_inv_1 _05952_ (.Y(_00754_),
    .A(net1920));
 sg13g2_inv_1 _05953_ (.Y(_00755_),
    .A(net1419));
 sg13g2_inv_1 _05954_ (.Y(_00756_),
    .A(\i_core.cpu.instr_data_start[22] ));
 sg13g2_inv_1 _05955_ (.Y(_00757_),
    .A(net1423));
 sg13g2_inv_1 _05956_ (.Y(_00758_),
    .A(\i_core.cpu.instr_data_start[18] ));
 sg13g2_inv_1 _05957_ (.Y(_00759_),
    .A(net1424));
 sg13g2_inv_1 _05958_ (.Y(_00760_),
    .A(net2621));
 sg13g2_inv_1 _05959_ (.Y(_00761_),
    .A(net2579));
 sg13g2_inv_1 _05960_ (.Y(_00762_),
    .A(net2662));
 sg13g2_inv_2 _05961_ (.Y(_00763_),
    .A(net2477));
 sg13g2_inv_1 _05962_ (.Y(_00764_),
    .A(net2656));
 sg13g2_inv_2 _05963_ (.Y(_00765_),
    .A(net2555));
 sg13g2_inv_1 _05964_ (.Y(_00766_),
    .A(net2063));
 sg13g2_inv_1 _05965_ (.Y(_00767_),
    .A(\i_core.mem.q_ctrl.spi_flash_select ));
 sg13g2_inv_1 _05966_ (.Y(_00768_),
    .A(net1430));
 sg13g2_inv_1 _05967_ (.Y(_00769_),
    .A(\i_core.mem.q_ctrl.nibbles_remaining[2] ));
 sg13g2_inv_1 _05968_ (.Y(_00770_),
    .A(\i_core.mem.instr_active ));
 sg13g2_inv_1 _05969_ (.Y(_00771_),
    .A(\i_core.cpu.i_core.mie[17] ));
 sg13g2_inv_1 _05970_ (.Y(_00772_),
    .A(net2313));
 sg13g2_inv_1 _05971_ (.Y(_00773_),
    .A(net2338));
 sg13g2_inv_1 _05972_ (.Y(_00774_),
    .A(net2420));
 sg13g2_inv_1 _05973_ (.Y(_00775_),
    .A(\data_to_write[0] ));
 sg13g2_inv_1 _05974_ (.Y(_00776_),
    .A(\i_spi.bits_remaining[3] ));
 sg13g2_inv_1 _05975_ (.Y(_00777_),
    .A(\i_spi.bits_remaining[0] ));
 sg13g2_inv_1 _05976_ (.Y(_00778_),
    .A(net1454));
 sg13g2_inv_1 _05977_ (.Y(_00779_),
    .A(net2535));
 sg13g2_inv_1 _05978_ (.Y(_00780_),
    .A(net2569));
 sg13g2_inv_1 _05979_ (.Y(_00781_),
    .A(net2023));
 sg13g2_inv_1 _05980_ (.Y(_00782_),
    .A(\i_uart_tx.cycle_counter[9] ));
 sg13g2_inv_1 _05981_ (.Y(_00783_),
    .A(net1461));
 sg13g2_inv_1 _05982_ (.Y(_00784_),
    .A(\i_core.cpu.i_core.time_hi[0] ));
 sg13g2_inv_2 _05983_ (.Y(_00785_),
    .A(\i_core.cpu.i_core.cycle[0] ));
 sg13g2_inv_1 _05984_ (.Y(_00786_),
    .A(net1405));
 sg13g2_inv_4 _05985_ (.A(net1409),
    .Y(_00787_));
 sg13g2_inv_1 _05986_ (.Y(_00788_),
    .A(net1415));
 sg13g2_inv_1 _05987_ (.Y(_00789_),
    .A(net2189));
 sg13g2_inv_1 _05988_ (.Y(_00790_),
    .A(net1394));
 sg13g2_inv_1 _05989_ (.Y(_00791_),
    .A(net1402));
 sg13g2_inv_2 _05990_ (.Y(_00792_),
    .A(net2675));
 sg13g2_inv_2 _05991_ (.Y(_00793_),
    .A(\i_core.cpu.instr_write_offset[2] ));
 sg13g2_inv_1 _05992_ (.Y(_00794_),
    .A(\i_core.mem.q_ctrl.data_ready ));
 sg13g2_inv_1 _05993_ (.Y(_00795_),
    .A(\i_uart_rx.cycle_counter[0] ));
 sg13g2_inv_1 _05994_ (.Y(_00796_),
    .A(net2482));
 sg13g2_inv_1 _05995_ (.Y(_00797_),
    .A(net2614));
 sg13g2_inv_1 _05996_ (.Y(_00798_),
    .A(net2563));
 sg13g2_inv_1 _05997_ (.Y(_00799_),
    .A(net2028));
 sg13g2_inv_1 _05998_ (.Y(_00800_),
    .A(net1956));
 sg13g2_inv_1 _05999_ (.Y(_00801_),
    .A(net2586));
 sg13g2_inv_1 _06000_ (.Y(_00802_),
    .A(net1973));
 sg13g2_inv_1 _06001_ (.Y(_00803_),
    .A(\i_core.cpu.i_core.imm_lo[0] ));
 sg13g2_inv_1 _06002_ (.Y(_00804_),
    .A(net2065));
 sg13g2_inv_1 _06003_ (.Y(_00805_),
    .A(net1992));
 sg13g2_inv_1 _06004_ (.Y(_00806_),
    .A(\i_core.cpu.i_core.cmp ));
 sg13g2_inv_1 _06005_ (.Y(_00807_),
    .A(_00090_));
 sg13g2_inv_1 _06006_ (.Y(_00808_),
    .A(net2045));
 sg13g2_inv_1 _06007_ (.Y(_00809_),
    .A(net1946));
 sg13g2_inv_1 _06008_ (.Y(_00810_),
    .A(_00102_));
 sg13g2_inv_1 _06009_ (.Y(_00811_),
    .A(_00139_));
 sg13g2_inv_1 _06010_ (.Y(_00812_),
    .A(_00143_));
 sg13g2_inv_1 _06011_ (.Y(_00813_),
    .A(_00089_));
 sg13g2_inv_1 _06012_ (.Y(_00814_),
    .A(\i_uart_rx.cycle_counter[2] ));
 sg13g2_inv_1 _06013_ (.Y(_00815_),
    .A(\i_uart_rx.cycle_counter[8] ));
 sg13g2_inv_1 _06014_ (.Y(_00816_),
    .A(net2051));
 sg13g2_inv_1 _06015_ (.Y(_00817_),
    .A(\addr[6] ));
 sg13g2_inv_1 _06016_ (.Y(_00818_),
    .A(net1321));
 sg13g2_inv_1 _06017_ (.Y(_00819_),
    .A(\i_core.cpu.instr_fetch_stopped ));
 sg13g2_inv_1 _06018_ (.Y(_00820_),
    .A(net2503));
 sg13g2_inv_1 _06019_ (.Y(_00821_),
    .A(net2327));
 sg13g2_inv_1 _06020_ (.Y(_00822_),
    .A(net2237));
 sg13g2_inv_1 _06021_ (.Y(_00823_),
    .A(net2619));
 sg13g2_inv_1 _06022_ (.Y(_00824_),
    .A(\i_core.cpu.i_core.i_instrret.data[0] ));
 sg13g2_inv_1 _06023_ (.Y(_00825_),
    .A(net2547));
 sg13g2_inv_1 _06024_ (.Y(_00826_),
    .A(net2483));
 sg13g2_inv_1 _06025_ (.Y(_00827_),
    .A(net2469));
 sg13g2_inv_1 _06026_ (.Y(_00828_),
    .A(\gpio_out[4] ));
 sg13g2_inv_1 _06027_ (.Y(_00829_),
    .A(net1438));
 sg13g2_inv_1 _06028_ (.Y(_00830_),
    .A(net2639));
 sg13g2_inv_1 _06029_ (.Y(_00831_),
    .A(net2417));
 sg13g2_inv_1 _06030_ (.Y(_00832_),
    .A(net2374));
 sg13g2_inv_2 _06031_ (.Y(_00833_),
    .A(net2290));
 sg13g2_inv_1 _06032_ (.Y(_00834_),
    .A(net6));
 sg13g2_inv_1 _06033_ (.Y(_00835_),
    .A(net2659));
 sg13g2_inv_1 _06034_ (.Y(_00836_),
    .A(net2422));
 sg13g2_inv_2 _06035_ (.Y(_00837_),
    .A(net1470));
 sg13g2_inv_1 _06036_ (.Y(_00838_),
    .A(net2462));
 sg13g2_inv_1 _06037_ (.Y(_00839_),
    .A(\gpio_out[7] ));
 sg13g2_inv_1 _06038_ (.Y(_00840_),
    .A(\i_core.cpu.i_core.multiplier.accum[3] ));
 sg13g2_inv_1 _06039_ (.Y(_00841_),
    .A(net2147));
 sg13g2_inv_1 _06040_ (.Y(_00842_),
    .A(net2297));
 sg13g2_inv_1 _06041_ (.Y(_00843_),
    .A(net2410));
 sg13g2_inv_2 _06042_ (.Y(_00844_),
    .A(_00202_));
 sg13g2_inv_1 _06043_ (.Y(_00845_),
    .A(_00205_));
 sg13g2_inv_1 _06044_ (.Y(_00846_),
    .A(net2354));
 sg13g2_inv_1 _06045_ (.Y(_00847_),
    .A(net2305));
 sg13g2_inv_1 _06046_ (.Y(_00848_),
    .A(_00207_));
 sg13g2_inv_1 _06047_ (.Y(_00849_),
    .A(net2179));
 sg13g2_inv_1 _06048_ (.Y(_00850_),
    .A(_00213_));
 sg13g2_inv_1 _06049_ (.Y(_00851_),
    .A(net2157));
 sg13g2_inv_1 _06050_ (.Y(_00852_),
    .A(net2033));
 sg13g2_inv_2 _06051_ (.Y(_00853_),
    .A(net9));
 sg13g2_inv_1 _06052_ (.Y(_00854_),
    .A(net10));
 sg13g2_inv_1 _06053_ (.Y(_00855_),
    .A(\i_core.mem.q_ctrl.spi_in_buffer[6] ));
 sg13g2_inv_1 _06054_ (.Y(_00856_),
    .A(net12));
 sg13g2_inv_1 _06055_ (.Y(_00857_),
    .A(net1790));
 sg13g2_inv_1 _06056_ (.Y(_00858_),
    .A(net1814));
 sg13g2_inv_1 _06057_ (.Y(_00859_),
    .A(net1755));
 sg13g2_inv_1 _06058_ (.Y(_00860_),
    .A(net1758));
 sg13g2_inv_1 _06059_ (.Y(_00861_),
    .A(\i_core.cpu.i_core.multiplier.accum[4] ));
 sg13g2_inv_1 _06060_ (.Y(_00862_),
    .A(\i_core.cpu.i_core.multiplier.accum[5] ));
 sg13g2_inv_1 _06061_ (.Y(_00863_),
    .A(\i_core.cpu.i_core.multiplier.accum[6] ));
 sg13g2_inv_1 _06062_ (.Y(_00864_),
    .A(\i_core.cpu.i_core.multiplier.accum[7] ));
 sg13g2_inv_1 _06063_ (.Y(_00865_),
    .A(\i_core.cpu.i_core.multiplier.accum[8] ));
 sg13g2_inv_1 _06064_ (.Y(_00866_),
    .A(\i_core.cpu.i_core.multiplier.accum[9] ));
 sg13g2_inv_1 _06065_ (.Y(_00867_),
    .A(\i_core.cpu.i_core.multiplier.accum[10] ));
 sg13g2_inv_1 _06066_ (.Y(_00868_),
    .A(\i_core.cpu.i_core.multiplier.accum[11] ));
 sg13g2_inv_1 _06067_ (.Y(_00869_),
    .A(\i_core.cpu.i_core.multiplier.accum[12] ));
 sg13g2_inv_1 _06068_ (.Y(_00870_),
    .A(\i_core.cpu.i_core.multiplier.accum[13] ));
 sg13g2_inv_1 _06069_ (.Y(_00871_),
    .A(\i_core.cpu.i_core.multiplier.accum[14] ));
 sg13g2_inv_1 _06070_ (.Y(_00872_),
    .A(\i_core.cpu.i_core.multiplier.accum[15] ));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_o21ai_1 _06072_ (.B1(net1390),
    .Y(_00873_),
    .A1(\i_core.cpu.is_jal ),
    .A2(\i_core.cpu.is_auipc ));
 sg13g2_nor2_1 _06073_ (.A(net1408),
    .B(net1414),
    .Y(_00874_));
 sg13g2_nand2_2 _06074_ (.Y(_00875_),
    .A(_00787_),
    .B(net1377));
 sg13g2_and2_1 _06075_ (.A(net1409),
    .B(net1412),
    .X(_00876_));
 sg13g2_nand2_2 _06076_ (.Y(_00877_),
    .A(net1410),
    .B(net1416));
 sg13g2_a22oi_1 _06077_ (.Y(_00878_),
    .B1(net1364),
    .B2(net1425),
    .A2(net1367),
    .A1(net1428));
 sg13g2_nor2b_1 _06078_ (.A(net1408),
    .B_N(net1414),
    .Y(_00879_));
 sg13g2_nand2_2 _06079_ (.Y(_00880_),
    .A(_00787_),
    .B(net1412));
 sg13g2_nor2b_1 _06080_ (.A(net1414),
    .B_N(net1408),
    .Y(_00881_));
 sg13g2_nand2_2 _06081_ (.Y(_00882_),
    .A(net1409),
    .B(net1377));
 sg13g2_a22oi_1 _06082_ (.Y(_00883_),
    .B1(net1358),
    .B2(\i_core.cpu.instr_data_start[11] ),
    .A2(net1362),
    .A1(net1427));
 sg13g2_a21oi_1 _06083_ (.A1(_00878_),
    .A2(_00883_),
    .Y(_00884_),
    .B1(net1406));
 sg13g2_nor2_2 _06084_ (.A(net1381),
    .B(net1410),
    .Y(_00885_));
 sg13g2_nand2_2 _06085_ (.Y(_00886_),
    .A(net1405),
    .B(_00787_));
 sg13g2_mux2_1 _06086_ (.A0(\i_core.cpu.instr_data_start[19] ),
    .A1(\i_core.cpu.instr_data_start[23] ),
    .S(net1415),
    .X(_00887_));
 sg13g2_a21oi_2 _06087_ (.B1(_00884_),
    .Y(_00888_),
    .A2(_00887_),
    .A1(_00885_));
 sg13g2_nor2_1 _06088_ (.A(_00873_),
    .B(_00888_),
    .Y(_00889_));
 sg13g2_nor2b_2 _06089_ (.A(\i_core.cpu.i_core.i_registers.rs1[3] ),
    .B_N(\i_core.cpu.i_core.i_registers.rs1[2] ),
    .Y(_00890_));
 sg13g2_nor2b_2 _06090_ (.A(\i_core.cpu.i_core.i_registers.rs1[0] ),
    .B_N(\i_core.cpu.i_core.i_registers.rs1[1] ),
    .Y(_00891_));
 sg13g2_and2_2 _06091_ (.A(_00890_),
    .B(_00891_),
    .X(_00892_));
 sg13g2_nor2b_1 _06092_ (.A(\i_core.cpu.i_core.i_registers.rs1[2] ),
    .B_N(\i_core.cpu.i_core.i_registers.rs1[3] ),
    .Y(_00893_));
 sg13g2_and2_1 _06093_ (.A(net1356),
    .B(net1355),
    .X(_00894_));
 sg13g2_nand3_1 _06094_ (.B(net1356),
    .C(net1355),
    .A(\i_core.cpu.i_core.i_registers.reg_access[10][3] ),
    .Y(_00895_));
 sg13g2_nor2b_2 _06095_ (.A(\i_core.cpu.i_core.i_registers.rs1[1] ),
    .B_N(\i_core.cpu.i_core.i_registers.rs1[0] ),
    .Y(_00896_));
 sg13g2_and2_1 _06096_ (.A(_00890_),
    .B(_00896_),
    .X(_00897_));
 sg13g2_nor2_2 _06097_ (.A(\i_core.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_core.cpu.i_core.i_registers.rs1[1] ),
    .Y(_00898_));
 sg13g2_and2_2 _06098_ (.A(_00893_),
    .B(_00898_),
    .X(_00899_));
 sg13g2_and2_2 _06099_ (.A(\i_core.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_core.cpu.i_core.i_registers.rs1[2] ),
    .X(_00900_));
 sg13g2_nand3_1 _06100_ (.B(net1356),
    .C(_00900_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[14][3] ),
    .Y(_00901_));
 sg13g2_and2_1 _06101_ (.A(_00893_),
    .B(_00896_),
    .X(_00902_));
 sg13g2_nand3_1 _06102_ (.B(net1355),
    .C(_00896_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[9][3] ),
    .Y(_00903_));
 sg13g2_and2_1 _06103_ (.A(_00898_),
    .B(_00900_),
    .X(_00904_));
 sg13g2_and2_2 _06104_ (.A(_00896_),
    .B(_00900_),
    .X(_00905_));
 sg13g2_a22oi_1 _06105_ (.Y(_00906_),
    .B1(_00905_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[13][3] ),
    .A2(_00904_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[12][3] ));
 sg13g2_and2_2 _06106_ (.A(net1404),
    .B(net1408),
    .X(_00907_));
 sg13g2_nand2_1 _06107_ (.Y(_00908_),
    .A(net1407),
    .B(net1410));
 sg13g2_nand4_1 _06108_ (.B(_00890_),
    .C(_00898_),
    .A(net1379),
    .Y(_00909_),
    .D(_00907_));
 sg13g2_and2_2 _06109_ (.A(\i_core.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_core.cpu.i_core.i_registers.rs1[1] ),
    .X(_00910_));
 sg13g2_and2_1 _06110_ (.A(net1355),
    .B(_00910_),
    .X(_00911_));
 sg13g2_nand3_1 _06111_ (.B(net1355),
    .C(_00910_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[11][3] ),
    .Y(_00912_));
 sg13g2_and2_1 _06112_ (.A(_00890_),
    .B(_00910_),
    .X(_00913_));
 sg13g2_nand4_1 _06113_ (.B(\i_core.cpu.i_core.i_registers.rs1[1] ),
    .C(\i_core.cpu.i_core.i_registers.rs1[3] ),
    .A(\i_core.cpu.i_core.i_registers.rs1[0] ),
    .Y(_00914_),
    .D(\i_core.cpu.i_core.i_registers.rs1[2] ));
 sg13g2_nor2_1 _06114_ (.A(_00091_),
    .B(_00914_),
    .Y(_00915_));
 sg13g2_a21oi_1 _06115_ (.A1(\i_core.cpu.i_core.i_registers.reg_access[7][3] ),
    .A2(_00913_),
    .Y(_00916_),
    .B1(_00915_));
 sg13g2_nor2_2 _06116_ (.A(\i_core.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_core.cpu.i_core.i_registers.rs1[2] ),
    .Y(_00917_));
 sg13g2_and2_1 _06117_ (.A(_00896_),
    .B(_00917_),
    .X(_00918_));
 sg13g2_and3_1 _06118_ (.X(_00919_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[1][3] ),
    .B(_00896_),
    .C(_00917_));
 sg13g2_nand3_1 _06119_ (.B(_00891_),
    .C(_00917_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[2][3] ),
    .Y(_00920_));
 sg13g2_nand2_1 _06120_ (.Y(_00921_),
    .A(_00901_),
    .B(_00909_));
 sg13g2_a21oi_2 _06121_ (.B1(_00921_),
    .Y(_00922_),
    .A2(_00892_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[6][3] ));
 sg13g2_and4_1 _06122_ (.A(_00895_),
    .B(_00903_),
    .C(_00912_),
    .D(_00920_),
    .X(_00923_));
 sg13g2_a221oi_1 _06123_ (.B2(\i_core.cpu.i_core.i_registers.reg_access[8][3] ),
    .C1(_00919_),
    .B1(_00899_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[5][3] ),
    .Y(_00924_),
    .A2(_00897_));
 sg13g2_and4_1 _06124_ (.A(_00906_),
    .B(_00916_),
    .C(_00923_),
    .D(_00924_),
    .X(_00925_));
 sg13g2_nand2_2 _06125_ (.Y(_00926_),
    .A(_00922_),
    .B(_00925_));
 sg13g2_inv_1 _06126_ (.Y(_00927_),
    .A(_00926_));
 sg13g2_a21oi_2 _06127_ (.B1(_00889_),
    .Y(_00928_),
    .A2(_00926_),
    .A1(_00873_));
 sg13g2_nor2_2 _06128_ (.A(net1402),
    .B(\i_core.cpu.alu_op[3] ),
    .Y(_00929_));
 sg13g2_and2_1 _06129_ (.A(net1390),
    .B(\i_core.cpu.is_branch ),
    .X(_00930_));
 sg13g2_nand2_1 _06130_ (.Y(_00931_),
    .A(net1392),
    .B(\i_core.cpu.is_branch ));
 sg13g2_o21ai_1 _06131_ (.B1(net1391),
    .Y(_00932_),
    .A1(\i_core.cpu.is_branch ),
    .A2(\i_core.cpu.is_alu_reg ));
 sg13g2_inv_1 _06132_ (.Y(_00933_),
    .A(_00932_));
 sg13g2_nor2b_1 _06133_ (.A(\i_core.cpu.i_core.i_registers.rs2[1] ),
    .B_N(\i_core.cpu.i_core.i_registers.rs2[0] ),
    .Y(_00934_));
 sg13g2_nor2b_1 _06134_ (.A(\i_core.cpu.i_core.i_registers.rs2[2] ),
    .B_N(\i_core.cpu.i_core.i_registers.rs2[3] ),
    .Y(_00935_));
 sg13g2_and2_1 _06135_ (.A(net1341),
    .B(_00935_),
    .X(_00936_));
 sg13g2_nand2_1 _06136_ (.Y(_00937_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[9][3] ),
    .B(_00936_));
 sg13g2_and2_1 _06137_ (.A(\i_core.cpu.i_core.i_registers.rs2[3] ),
    .B(\i_core.cpu.i_core.i_registers.rs2[2] ),
    .X(_00938_));
 sg13g2_nor2b_2 _06138_ (.A(\i_core.cpu.i_core.i_registers.rs2[0] ),
    .B_N(\i_core.cpu.i_core.i_registers.rs2[1] ),
    .Y(_00939_));
 sg13g2_nand3_1 _06139_ (.B(net1339),
    .C(net1338),
    .A(\i_core.cpu.i_core.i_registers.reg_access[14][3] ),
    .Y(_00940_));
 sg13g2_nor2_2 _06140_ (.A(\i_core.cpu.i_core.i_registers.rs2[3] ),
    .B(\i_core.cpu.i_core.i_registers.rs2[2] ),
    .Y(_00941_));
 sg13g2_and2_1 _06141_ (.A(net1338),
    .B(_00941_),
    .X(_00942_));
 sg13g2_and2_1 _06142_ (.A(_00935_),
    .B(_00939_),
    .X(_00943_));
 sg13g2_a22oi_1 _06143_ (.Y(_00944_),
    .B1(_00943_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[10][3] ),
    .A2(_00942_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[2][3] ));
 sg13g2_and2_1 _06144_ (.A(net1341),
    .B(_00941_),
    .X(_00945_));
 sg13g2_nand3_1 _06145_ (.B(net1341),
    .C(_00941_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[1][3] ),
    .Y(_00946_));
 sg13g2_nor2_2 _06146_ (.A(\i_core.cpu.i_core.i_registers.rs2[1] ),
    .B(\i_core.cpu.i_core.i_registers.rs2[0] ),
    .Y(_00947_));
 sg13g2_nand3_1 _06147_ (.B(_00935_),
    .C(_00947_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[8][3] ),
    .Y(_00948_));
 sg13g2_and2_1 _06148_ (.A(\i_core.cpu.i_core.i_registers.rs2[1] ),
    .B(\i_core.cpu.i_core.i_registers.rs2[0] ),
    .X(_00949_));
 sg13g2_and2_1 _06149_ (.A(net1340),
    .B(net1337),
    .X(_00950_));
 sg13g2_nand3_1 _06150_ (.B(net1340),
    .C(_00949_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[11][3] ),
    .Y(_00951_));
 sg13g2_nor2b_2 _06151_ (.A(\i_core.cpu.i_core.i_registers.rs2[3] ),
    .B_N(\i_core.cpu.i_core.i_registers.rs2[2] ),
    .Y(_00952_));
 sg13g2_nand3_1 _06152_ (.B(net1338),
    .C(_00952_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[6][3] ),
    .Y(_00953_));
 sg13g2_and4_1 _06153_ (.A(_00946_),
    .B(_00948_),
    .C(_00951_),
    .D(_00953_),
    .X(_00954_));
 sg13g2_and4_1 _06154_ (.A(_00937_),
    .B(_00940_),
    .C(_00944_),
    .D(_00954_),
    .X(_00955_));
 sg13g2_nand3_1 _06155_ (.B(_00907_),
    .C(_00947_),
    .A(net1379),
    .Y(_00956_));
 sg13g2_a22oi_1 _06156_ (.Y(_00957_),
    .B1(_00949_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[7][3] ),
    .A2(net1341),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[5][3] ));
 sg13g2_nand2_1 _06157_ (.Y(_00958_),
    .A(_00956_),
    .B(_00957_));
 sg13g2_nand2_1 _06158_ (.Y(_00959_),
    .A(_00952_),
    .B(_00958_));
 sg13g2_nand3_1 _06159_ (.B(net1342),
    .C(_00938_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[13][3] ),
    .Y(_00960_));
 sg13g2_nand2_1 _06160_ (.Y(_00961_),
    .A(net1339),
    .B(net1337));
 sg13g2_nor2_1 _06161_ (.A(_00091_),
    .B(_00961_),
    .Y(_00962_));
 sg13g2_and2_1 _06162_ (.A(net1339),
    .B(_00947_),
    .X(_00963_));
 sg13g2_a21oi_1 _06163_ (.A1(\i_core.cpu.i_core.i_registers.reg_access[12][3] ),
    .A2(_00963_),
    .Y(_00964_),
    .B1(_00962_));
 sg13g2_nand4_1 _06164_ (.B(_00959_),
    .C(_00960_),
    .A(_00955_),
    .Y(_00965_),
    .D(_00964_));
 sg13g2_a21oi_1 _06165_ (.A1(\i_core.cpu.imm[15] ),
    .A2(net1363),
    .Y(_00966_),
    .B1(net1406));
 sg13g2_nand2_1 _06166_ (.Y(_00967_),
    .A(\i_core.cpu.i_core.imm_lo[7] ),
    .B(net1361));
 sg13g2_a22oi_1 _06167_ (.Y(_00968_),
    .B1(net1358),
    .B2(\i_core.cpu.i_core.imm_lo[11] ),
    .A2(net1366),
    .A1(\i_core.cpu.i_core.imm_lo[3] ));
 sg13g2_nand3_1 _06168_ (.B(_00967_),
    .C(_00968_),
    .A(_00966_),
    .Y(_00969_));
 sg13g2_nand2_1 _06169_ (.Y(_00970_),
    .A(\i_core.cpu.imm[23] ),
    .B(_00879_));
 sg13g2_a22oi_1 _06170_ (.Y(_00971_),
    .B1(net1357),
    .B2(\i_core.cpu.imm[27] ),
    .A2(net1363),
    .A1(\i_core.cpu.imm[31] ));
 sg13g2_a21oi_1 _06171_ (.A1(\i_core.cpu.imm[19] ),
    .A2(net1368),
    .Y(_00972_),
    .B1(net1380));
 sg13g2_nand3_1 _06172_ (.B(_00971_),
    .C(_00972_),
    .A(_00970_),
    .Y(_00973_));
 sg13g2_nand2_2 _06173_ (.Y(_00974_),
    .A(_00969_),
    .B(_00973_));
 sg13g2_nand2_1 _06174_ (.Y(_00975_),
    .A(_00932_),
    .B(_00974_));
 sg13g2_o21ai_1 _06175_ (.B1(_00975_),
    .Y(_00976_),
    .A1(_00932_),
    .A2(_00965_));
 sg13g2_xor2_1 _06176_ (.B(_00976_),
    .A(_00929_),
    .X(_00977_));
 sg13g2_inv_1 _06177_ (.Y(_00978_),
    .A(_00977_));
 sg13g2_nand2_1 _06178_ (.Y(_00979_),
    .A(_00928_),
    .B(_00978_));
 sg13g2_nor2_1 _06179_ (.A(_00928_),
    .B(_00978_),
    .Y(_00980_));
 sg13g2_nor2_1 _06180_ (.A(\i_core.cpu.instr_data_start[18] ),
    .B(net1413),
    .Y(_00981_));
 sg13g2_a21oi_1 _06181_ (.A1(_00756_),
    .A2(net1413),
    .Y(_00982_),
    .B1(_00981_));
 sg13g2_a22oi_1 _06182_ (.Y(_00983_),
    .B1(net1364),
    .B2(net1426),
    .A2(net1366),
    .A1(\i_core.cpu.pc[2] ));
 sg13g2_a22oi_1 _06183_ (.Y(_00984_),
    .B1(net1358),
    .B2(\i_core.cpu.instr_data_start[10] ),
    .A2(net1362),
    .A1(\i_core.cpu.instr_data_start[6] ));
 sg13g2_nand2_1 _06184_ (.Y(_00985_),
    .A(_00983_),
    .B(_00984_));
 sg13g2_a22oi_1 _06185_ (.Y(_00986_),
    .B1(_00985_),
    .B2(net1381),
    .A2(_00982_),
    .A1(_00885_));
 sg13g2_nor2_1 _06186_ (.A(_00873_),
    .B(_00986_),
    .Y(_00987_));
 sg13g2_or2_1 _06187_ (.X(_00988_),
    .B(_00914_),
    .A(_00093_));
 sg13g2_nand3_1 _06188_ (.B(net1356),
    .C(_00917_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[2][2] ),
    .Y(_00989_));
 sg13g2_nand3_1 _06189_ (.B(_00898_),
    .C(_00900_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[12][2] ),
    .Y(_00990_));
 sg13g2_nand2_1 _06190_ (.Y(_00991_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[7][2] ),
    .B(_00913_));
 sg13g2_nand2_1 _06191_ (.Y(_00992_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[13][2] ),
    .B(_00905_));
 sg13g2_nand3_1 _06192_ (.B(net1356),
    .C(_00900_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[14][2] ),
    .Y(_00993_));
 sg13g2_nand2_1 _06193_ (.Y(_00994_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[8][2] ),
    .B(_00899_));
 sg13g2_nor2_2 _06194_ (.A(net1406),
    .B(_00882_),
    .Y(_00995_));
 sg13g2_nand4_1 _06195_ (.B(net1359),
    .C(_00910_),
    .A(net1382),
    .Y(_00996_),
    .D(_00917_));
 sg13g2_a22oi_1 _06196_ (.Y(_00997_),
    .B1(_00897_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[5][2] ),
    .A2(_00892_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[6][2] ));
 sg13g2_a22oi_1 _06197_ (.Y(_00998_),
    .B1(_00902_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[9][2] ),
    .A2(_00894_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[10][2] ));
 sg13g2_a22oi_1 _06198_ (.Y(_00999_),
    .B1(_00918_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[1][2] ),
    .A2(_00911_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[11][2] ));
 sg13g2_and4_1 _06199_ (.A(_00988_),
    .B(_00989_),
    .C(_00990_),
    .D(_00993_),
    .X(_01000_));
 sg13g2_and4_1 _06200_ (.A(_00992_),
    .B(_00994_),
    .C(_00997_),
    .D(_01000_),
    .X(_01001_));
 sg13g2_and4_1 _06201_ (.A(_00991_),
    .B(_00996_),
    .C(_00998_),
    .D(_00999_),
    .X(_01002_));
 sg13g2_nand2_2 _06202_ (.Y(_01003_),
    .A(_01001_),
    .B(_01002_));
 sg13g2_a21oi_2 _06203_ (.B1(_00987_),
    .Y(_01004_),
    .A2(_01003_),
    .A1(_00873_));
 sg13g2_a21oi_1 _06204_ (.A1(\i_core.cpu.imm[14] ),
    .A2(net1363),
    .Y(_01005_),
    .B1(net1406));
 sg13g2_nand2_1 _06205_ (.Y(_01006_),
    .A(\i_core.cpu.i_core.imm_lo[6] ),
    .B(net1361));
 sg13g2_a22oi_1 _06206_ (.Y(_01007_),
    .B1(net1358),
    .B2(\i_core.cpu.i_core.imm_lo[10] ),
    .A2(net1366),
    .A1(\i_core.cpu.i_core.imm_lo[2] ));
 sg13g2_nand3_1 _06207_ (.B(_01006_),
    .C(_01007_),
    .A(_01005_),
    .Y(_01008_));
 sg13g2_a21oi_1 _06208_ (.A1(\i_core.cpu.imm[22] ),
    .A2(net1360),
    .Y(_01009_),
    .B1(net1380));
 sg13g2_nand2_1 _06209_ (.Y(_01010_),
    .A(\i_core.cpu.imm[26] ),
    .B(net1359));
 sg13g2_a22oi_1 _06210_ (.Y(_01011_),
    .B1(net1365),
    .B2(\i_core.cpu.imm[30] ),
    .A2(net1368),
    .A1(\i_core.cpu.imm[18] ));
 sg13g2_nand3_1 _06211_ (.B(_01010_),
    .C(_01011_),
    .A(_01009_),
    .Y(_01012_));
 sg13g2_nand2_2 _06212_ (.Y(_01013_),
    .A(_01008_),
    .B(_01012_));
 sg13g2_nand3_1 _06213_ (.B(net1341),
    .C(net1340),
    .A(\i_core.cpu.i_core.i_registers.reg_access[9][2] ),
    .Y(_01014_));
 sg13g2_nand3_1 _06214_ (.B(net1340),
    .C(_00947_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[8][2] ),
    .Y(_01015_));
 sg13g2_nand2_1 _06215_ (.Y(_01016_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[1][2] ),
    .B(_00945_));
 sg13g2_nand3_1 _06216_ (.B(net1342),
    .C(net1339),
    .A(\i_core.cpu.i_core.i_registers.reg_access[13][2] ),
    .Y(_01017_));
 sg13g2_nand3_1 _06217_ (.B(_00939_),
    .C(_00952_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[6][2] ),
    .Y(_01018_));
 sg13g2_nand3_1 _06218_ (.B(_00949_),
    .C(_00995_),
    .A(_00941_),
    .Y(_01019_));
 sg13g2_nand3_1 _06219_ (.B(net1339),
    .C(net1338),
    .A(\i_core.cpu.i_core.i_registers.reg_access[14][2] ),
    .Y(_01020_));
 sg13g2_and2_1 _06220_ (.A(net1341),
    .B(_00952_),
    .X(_01021_));
 sg13g2_and2_1 _06221_ (.A(net1337),
    .B(_00952_),
    .X(_01022_));
 sg13g2_a22oi_1 _06222_ (.Y(_01023_),
    .B1(_01022_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[7][2] ),
    .A2(_00963_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[12][2] ));
 sg13g2_and2_1 _06223_ (.A(_01017_),
    .B(_01020_),
    .X(_01024_));
 sg13g2_o21ai_1 _06224_ (.B1(_01014_),
    .Y(_01025_),
    .A1(_00093_),
    .A2(_00961_));
 sg13g2_a221oi_1 _06225_ (.B2(\i_core.cpu.i_core.i_registers.reg_access[11][2] ),
    .C1(_01025_),
    .B1(_00950_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[2][2] ),
    .Y(_01026_),
    .A2(_00942_));
 sg13g2_nand4_1 _06226_ (.B(_01018_),
    .C(_01024_),
    .A(_01015_),
    .Y(_01027_),
    .D(_01026_));
 sg13g2_a22oi_1 _06227_ (.Y(_01028_),
    .B1(_01021_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[5][2] ),
    .A2(_00943_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[10][2] ));
 sg13g2_nand4_1 _06228_ (.B(_01019_),
    .C(_01023_),
    .A(_01016_),
    .Y(_01029_),
    .D(_01028_));
 sg13g2_nor2_2 _06229_ (.A(_01027_),
    .B(_01029_),
    .Y(_01030_));
 sg13g2_mux2_2 _06230_ (.A0(_01013_),
    .A1(_01030_),
    .S(_00933_),
    .X(_01031_));
 sg13g2_xnor2_1 _06231_ (.Y(_01032_),
    .A(_00929_),
    .B(_01031_));
 sg13g2_or2_1 _06232_ (.X(_01033_),
    .B(_01032_),
    .A(_01004_));
 sg13g2_a22oi_1 _06233_ (.Y(_01034_),
    .B1(net1364),
    .B2(\i_core.cpu.instr_data_start[13] ),
    .A2(net1366),
    .A1(\i_core.cpu.pc[1] ));
 sg13g2_a22oi_1 _06234_ (.Y(_01035_),
    .B1(net1358),
    .B2(\i_core.cpu.instr_data_start[9] ),
    .A2(net1362),
    .A1(\i_core.cpu.instr_data_start[5] ));
 sg13g2_nand2_1 _06235_ (.Y(_01036_),
    .A(_01034_),
    .B(_01035_));
 sg13g2_mux2_1 _06236_ (.A0(\i_core.cpu.instr_data_start[17] ),
    .A1(\i_core.cpu.instr_data_start[21] ),
    .S(net1413),
    .X(_01037_));
 sg13g2_a22oi_1 _06237_ (.Y(_01038_),
    .B1(_01037_),
    .B2(_00885_),
    .A2(_01036_),
    .A1(net1381));
 sg13g2_nor2_1 _06238_ (.A(_00873_),
    .B(_01038_),
    .Y(_01039_));
 sg13g2_a22oi_1 _06239_ (.Y(_01040_),
    .B1(_00918_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[1][1] ),
    .A2(_00892_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[6][1] ));
 sg13g2_nand3_1 _06240_ (.B(net1355),
    .C(_00910_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[11][1] ),
    .Y(_01041_));
 sg13g2_nand2_1 _06241_ (.Y(_01042_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[13][1] ),
    .B(_00905_));
 sg13g2_nand3_1 _06242_ (.B(net1356),
    .C(_00900_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[14][1] ),
    .Y(_01043_));
 sg13g2_nand3_1 _06243_ (.B(_00891_),
    .C(_00917_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[2][1] ),
    .Y(_01044_));
 sg13g2_nor2_1 _06244_ (.A(_00094_),
    .B(_00914_),
    .Y(_01045_));
 sg13g2_a22oi_1 _06245_ (.Y(_01046_),
    .B1(_00902_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[9][1] ),
    .A2(_00899_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[8][1] ));
 sg13g2_a22oi_1 _06246_ (.Y(_01047_),
    .B1(_00904_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[12][1] ),
    .A2(_00894_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[10][1] ));
 sg13g2_nand4_1 _06247_ (.B(_01044_),
    .C(_01046_),
    .A(_01043_),
    .Y(_01048_),
    .D(_01047_));
 sg13g2_a221oi_1 _06248_ (.B2(\i_core.cpu.i_core.i_registers.reg_access[7][1] ),
    .C1(_01045_),
    .B1(_00913_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[5][1] ),
    .Y(_01049_),
    .A2(_00897_));
 sg13g2_nand4_1 _06249_ (.B(_01041_),
    .C(_01042_),
    .A(_01040_),
    .Y(_01050_),
    .D(_01049_));
 sg13g2_or2_2 _06250_ (.X(_01051_),
    .B(_01050_),
    .A(_01048_));
 sg13g2_a21oi_2 _06251_ (.B1(_01039_),
    .Y(_01052_),
    .A2(_01051_),
    .A1(_00873_));
 sg13g2_a22oi_1 _06252_ (.Y(_01053_),
    .B1(_01022_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[7][1] ),
    .A2(_00936_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[9][1] ));
 sg13g2_a22oi_1 _06253_ (.Y(_01054_),
    .B1(_01021_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[5][1] ),
    .A2(_00945_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[1][1] ));
 sg13g2_a22oi_1 _06254_ (.Y(_01055_),
    .B1(_00950_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[11][1] ),
    .A2(_00943_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[10][1] ));
 sg13g2_nand3_1 _06255_ (.B(_01054_),
    .C(_01055_),
    .A(_01053_),
    .Y(_01056_));
 sg13g2_and2_1 _06256_ (.A(\i_core.cpu.i_core.i_registers.reg_access[12][1] ),
    .B(_00963_),
    .X(_01057_));
 sg13g2_nand3_1 _06257_ (.B(net1338),
    .C(_00952_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[6][1] ),
    .Y(_01058_));
 sg13g2_o21ai_1 _06258_ (.B1(_01058_),
    .Y(_01059_),
    .A1(_00094_),
    .A2(_00961_));
 sg13g2_nand2_1 _06259_ (.Y(_01060_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[2][1] ),
    .B(_00942_));
 sg13g2_nand3_1 _06260_ (.B(net1342),
    .C(_00938_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[13][1] ),
    .Y(_01061_));
 sg13g2_nand3_1 _06261_ (.B(net1340),
    .C(_00947_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[8][1] ),
    .Y(_01062_));
 sg13g2_nand3_1 _06262_ (.B(net1339),
    .C(net1338),
    .A(\i_core.cpu.i_core.i_registers.reg_access[14][1] ),
    .Y(_01063_));
 sg13g2_nand4_1 _06263_ (.B(_01061_),
    .C(_01062_),
    .A(_01060_),
    .Y(_01064_),
    .D(_01063_));
 sg13g2_nor4_2 _06264_ (.A(_01056_),
    .B(_01057_),
    .C(_01059_),
    .Y(_01065_),
    .D(_01064_));
 sg13g2_a22oi_1 _06265_ (.Y(_01066_),
    .B1(net1361),
    .B2(\i_core.cpu.i_core.imm_lo[5] ),
    .A2(net1363),
    .A1(\i_core.cpu.imm[13] ));
 sg13g2_a221oi_1 _06266_ (.B2(\i_core.cpu.i_core.imm_lo[9] ),
    .C1(net1406),
    .B1(net1358),
    .A1(\i_core.cpu.i_core.imm_lo[1] ),
    .Y(_01067_),
    .A2(net1366));
 sg13g2_and2_1 _06267_ (.A(\i_core.cpu.imm[29] ),
    .B(net1363),
    .X(_01068_));
 sg13g2_a21oi_1 _06268_ (.A1(\i_core.cpu.imm[21] ),
    .A2(net1361),
    .Y(_01069_),
    .B1(net1381));
 sg13g2_a221oi_1 _06269_ (.B2(\i_core.cpu.imm[25] ),
    .C1(_01068_),
    .B1(net1359),
    .A1(\i_core.cpu.imm[17] ),
    .Y(_01070_),
    .A2(net1367));
 sg13g2_a22oi_1 _06270_ (.Y(_01071_),
    .B1(_01069_),
    .B2(_01070_),
    .A2(_01067_),
    .A1(_01066_));
 sg13g2_nand2_1 _06271_ (.Y(_01072_),
    .A(_00932_),
    .B(_01071_));
 sg13g2_o21ai_1 _06272_ (.B1(_01072_),
    .Y(_01073_),
    .A1(_00932_),
    .A2(_01065_));
 sg13g2_inv_1 _06273_ (.Y(_01074_),
    .A(_01073_));
 sg13g2_xnor2_1 _06274_ (.Y(_01075_),
    .A(_00929_),
    .B(_01073_));
 sg13g2_nor2b_1 _06275_ (.A(_01052_),
    .B_N(_01075_),
    .Y(_01076_));
 sg13g2_nand3_1 _06276_ (.B(net1356),
    .C(_00900_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[14][0] ),
    .Y(_01077_));
 sg13g2_nand3_1 _06277_ (.B(net1355),
    .C(_00910_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[11][0] ),
    .Y(_01078_));
 sg13g2_nand3_1 _06278_ (.B(net1356),
    .C(_00917_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[2][0] ),
    .Y(_01079_));
 sg13g2_nand4_1 _06279_ (.B(_00907_),
    .C(_00910_),
    .A(net1379),
    .Y(_01080_),
    .D(_00917_));
 sg13g2_nand3_1 _06280_ (.B(net1355),
    .C(_00896_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[9][0] ),
    .Y(_01081_));
 sg13g2_nand3_1 _06281_ (.B(_00900_),
    .C(_00910_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[15][0] ),
    .Y(_01082_));
 sg13g2_a22oi_1 _06282_ (.Y(_01083_),
    .B1(_00904_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[12][0] ),
    .A2(_00899_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[8][0] ));
 sg13g2_a22oi_1 _06283_ (.Y(_01084_),
    .B1(_00918_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[1][0] ),
    .A2(_00897_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[5][0] ));
 sg13g2_and2_1 _06284_ (.A(_01078_),
    .B(_01079_),
    .X(_01085_));
 sg13g2_a22oi_1 _06285_ (.Y(_01086_),
    .B1(_00905_),
    .B2(\i_core.cpu.i_core.i_registers.reg_access[13][0] ),
    .A2(_00892_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[6][0] ));
 sg13g2_and4_1 _06286_ (.A(_01083_),
    .B(_01084_),
    .C(_01085_),
    .D(_01086_),
    .X(_01087_));
 sg13g2_nand4_1 _06287_ (.B(_01080_),
    .C(_01081_),
    .A(_01077_),
    .Y(_01088_),
    .D(_01082_));
 sg13g2_a221oi_1 _06288_ (.B2(\i_core.cpu.i_core.i_registers.reg_access[7][0] ),
    .C1(_01088_),
    .B1(_00913_),
    .A1(\i_core.cpu.i_core.i_registers.reg_access[10][0] ),
    .Y(_01089_),
    .A2(_00894_));
 sg13g2_nand2_2 _06289_ (.Y(_01090_),
    .A(_01087_),
    .B(_01089_));
 sg13g2_a21oi_1 _06290_ (.A1(_00757_),
    .A2(net1413),
    .Y(_01091_),
    .B1(_00886_));
 sg13g2_o21ai_1 _06291_ (.B1(_01091_),
    .Y(_01092_),
    .A1(net1424),
    .A2(net1413));
 sg13g2_nor2_1 _06292_ (.A(_00761_),
    .B(_00877_),
    .Y(_01093_));
 sg13g2_a221oi_1 _06293_ (.B2(\i_core.cpu.instr_data_start[8] ),
    .C1(_01093_),
    .B1(net1358),
    .A1(\i_core.cpu.instr_data_start[4] ),
    .Y(_01094_),
    .A2(net1361));
 sg13g2_o21ai_1 _06294_ (.B1(_01092_),
    .Y(_01095_),
    .A1(net1406),
    .A2(_01094_));
 sg13g2_mux2_2 _06295_ (.A0(_01095_),
    .A1(_01090_),
    .S(_00873_),
    .X(_01096_));
 sg13g2_and2_1 _06296_ (.A(\i_core.cpu.i_core.imm_lo[8] ),
    .B(net1358),
    .X(_01097_));
 sg13g2_a221oi_1 _06297_ (.B2(\i_core.cpu.i_core.imm_lo[4] ),
    .C1(_01097_),
    .B1(net1361),
    .A1(\i_core.cpu.i_core.imm_lo[0] ),
    .Y(_01098_),
    .A2(net1366));
 sg13g2_a21oi_1 _06298_ (.A1(\i_core.cpu.imm[12] ),
    .A2(net1363),
    .Y(_01099_),
    .B1(net1406));
 sg13g2_a22oi_1 _06299_ (.Y(_01100_),
    .B1(net1363),
    .B2(\i_core.cpu.imm[28] ),
    .A2(net1367),
    .A1(\i_core.cpu.imm[16] ));
 sg13g2_a221oi_1 _06300_ (.B2(\i_core.cpu.imm[24] ),
    .C1(net1381),
    .B1(net1359),
    .A1(\i_core.cpu.imm[20] ),
    .Y(_01101_),
    .A2(net1361));
 sg13g2_a22oi_1 _06301_ (.Y(_01102_),
    .B1(_01100_),
    .B2(_01101_),
    .A2(_01099_),
    .A1(_01098_));
 sg13g2_nand3_1 _06302_ (.B(net1342),
    .C(_00938_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[13][0] ),
    .Y(_01103_));
 sg13g2_nand3_1 _06303_ (.B(net1340),
    .C(net1337),
    .A(\i_core.cpu.i_core.i_registers.reg_access[11][0] ),
    .Y(_01104_));
 sg13g2_nand3_1 _06304_ (.B(net1341),
    .C(net1340),
    .A(\i_core.cpu.i_core.i_registers.reg_access[9][0] ),
    .Y(_01105_));
 sg13g2_nand3_1 _06305_ (.B(net1338),
    .C(_00952_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[6][0] ),
    .Y(_01106_));
 sg13g2_nand3_1 _06306_ (.B(net1339),
    .C(net1337),
    .A(\i_core.cpu.i_core.i_registers.reg_access[15][0] ),
    .Y(_01107_));
 sg13g2_nand2_1 _06307_ (.Y(_01108_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[7][0] ),
    .B(_01022_));
 sg13g2_nand4_1 _06308_ (.B(net1354),
    .C(_00941_),
    .A(net1379),
    .Y(_01109_),
    .D(net1337));
 sg13g2_nand3_1 _06309_ (.B(net1339),
    .C(net1338),
    .A(\i_core.cpu.i_core.i_registers.reg_access[14][0] ),
    .Y(_01110_));
 sg13g2_nand2_1 _06310_ (.Y(_01111_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[12][0] ),
    .B(_00963_));
 sg13g2_nand2_1 _06311_ (.Y(_01112_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[10][0] ),
    .B(_00943_));
 sg13g2_nand3_1 _06312_ (.B(net1340),
    .C(_00947_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[8][0] ),
    .Y(_01113_));
 sg13g2_nand3_1 _06313_ (.B(_00939_),
    .C(_00941_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[2][0] ),
    .Y(_01114_));
 sg13g2_nand2_1 _06314_ (.Y(_01115_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[5][0] ),
    .B(_01021_));
 sg13g2_nand3_1 _06315_ (.B(net1341),
    .C(_00941_),
    .A(\i_core.cpu.i_core.i_registers.reg_access[1][0] ),
    .Y(_01116_));
 sg13g2_nand4_1 _06316_ (.B(_01111_),
    .C(_01112_),
    .A(_01108_),
    .Y(_01117_),
    .D(_01115_));
 sg13g2_nand4_1 _06317_ (.B(_01106_),
    .C(_01110_),
    .A(_01103_),
    .Y(_01118_),
    .D(_01114_));
 sg13g2_nand3_1 _06318_ (.B(_01109_),
    .C(_01113_),
    .A(_01104_),
    .Y(_01119_));
 sg13g2_nand3_1 _06319_ (.B(_01107_),
    .C(_01116_),
    .A(_01105_),
    .Y(_01120_));
 sg13g2_nor3_2 _06320_ (.A(_01118_),
    .B(_01119_),
    .C(_01120_),
    .Y(_01121_));
 sg13g2_nand2b_2 _06321_ (.Y(_01122_),
    .B(_01121_),
    .A_N(_01117_));
 sg13g2_nand3b_1 _06322_ (.B(_01121_),
    .C(_00933_),
    .Y(_01123_),
    .A_N(_01117_));
 sg13g2_nand2b_1 _06323_ (.Y(_01124_),
    .B(_00932_),
    .A_N(_01102_));
 sg13g2_and2_1 _06324_ (.A(_01123_),
    .B(_01124_),
    .X(_01125_));
 sg13g2_and3_1 _06325_ (.X(_01126_),
    .A(_00929_),
    .B(_01123_),
    .C(_01124_));
 sg13g2_a21oi_1 _06326_ (.A1(_01123_),
    .A2(_01124_),
    .Y(_01127_),
    .B1(_00929_));
 sg13g2_nor2_1 _06327_ (.A(_01126_),
    .B(_01127_),
    .Y(_01128_));
 sg13g2_o21ai_1 _06328_ (.B1(_01096_),
    .Y(_01129_),
    .A1(_01126_),
    .A2(_01127_));
 sg13g2_nor3_1 _06329_ (.A(_01096_),
    .B(_01126_),
    .C(_01127_),
    .Y(_01130_));
 sg13g2_xnor2_1 _06330_ (.Y(_01131_),
    .A(_01096_),
    .B(_01128_));
 sg13g2_nor2_1 _06331_ (.A(net1404),
    .B(_00875_),
    .Y(_01132_));
 sg13g2_nand2_1 _06332_ (.Y(_01133_),
    .A(net1380),
    .B(net1368));
 sg13g2_nor3_1 _06333_ (.A(net1403),
    .B(\i_core.cpu.alu_op[3] ),
    .C(net1312),
    .Y(_01134_));
 sg13g2_a21oi_1 _06334_ (.A1(_00095_),
    .A2(net1312),
    .Y(_01135_),
    .B1(_01134_));
 sg13g2_inv_1 _06335_ (.Y(_01136_),
    .A(_01135_));
 sg13g2_o21ai_1 _06336_ (.B1(_01129_),
    .Y(_01137_),
    .A1(_01130_),
    .A2(_01136_));
 sg13g2_xnor2_1 _06337_ (.Y(_01138_),
    .A(_01052_),
    .B(_01075_));
 sg13g2_a21oi_2 _06338_ (.B1(_01076_),
    .Y(_01139_),
    .A2(_01138_),
    .A1(_01137_));
 sg13g2_xnor2_1 _06339_ (.Y(_01140_),
    .A(_01004_),
    .B(_01032_));
 sg13g2_o21ai_1 _06340_ (.B1(_01033_),
    .Y(_01141_),
    .A1(_01139_),
    .A2(_01140_));
 sg13g2_a21o_1 _06341_ (.A2(_01141_),
    .A1(_00979_),
    .B1(_00980_),
    .X(\i_core.cpu.i_core.cy_out ));
 sg13g2_nor2_1 _06342_ (.A(_00928_),
    .B(_00976_),
    .Y(_01142_));
 sg13g2_xnor2_1 _06343_ (.Y(_01143_),
    .A(_00928_),
    .B(_00976_));
 sg13g2_nand2_1 _06344_ (.Y(_01144_),
    .A(net1403),
    .B(_01143_));
 sg13g2_a221oi_1 _06345_ (.B2(_00792_),
    .C1(_00980_),
    .B1(_01144_),
    .A1(_00979_),
    .Y(_01145_),
    .A2(_01141_));
 sg13g2_o21ai_1 _06346_ (.B1(_01143_),
    .Y(_01146_),
    .A1(\i_core.cpu.i_core.cmp ),
    .A2(net1279));
 sg13g2_nor2_1 _06347_ (.A(_01052_),
    .B(_01074_),
    .Y(_01147_));
 sg13g2_xor2_1 _06348_ (.B(_01073_),
    .A(_01052_),
    .X(_01148_));
 sg13g2_nor2_1 _06349_ (.A(_01004_),
    .B(_01031_),
    .Y(_01149_));
 sg13g2_xnor2_1 _06350_ (.Y(_01150_),
    .A(_01004_),
    .B(_01031_));
 sg13g2_xnor2_1 _06351_ (.Y(_01151_),
    .A(_01096_),
    .B(_01125_));
 sg13g2_nand3_1 _06352_ (.B(_01150_),
    .C(_01151_),
    .A(_01148_),
    .Y(_01152_));
 sg13g2_or2_1 _06353_ (.X(_01153_),
    .B(_01152_),
    .A(_01146_));
 sg13g2_o21ai_1 _06354_ (.B1(_00792_),
    .Y(_01154_),
    .A1(_00791_),
    .A2(_00980_));
 sg13g2_a21oi_1 _06355_ (.A1(_00791_),
    .A2(_01153_),
    .Y(_01155_),
    .B1(_01154_));
 sg13g2_or2_1 _06356_ (.X(\i_core.cpu.i_core.cmp_out ),
    .B(_01155_),
    .A(_01145_));
 sg13g2_nor2_1 _06357_ (.A(_00747_),
    .B(_00083_),
    .Y(_01156_));
 sg13g2_nor3_1 _06358_ (.A(_00747_),
    .B(\i_core.cpu.is_store ),
    .C(\i_core.cpu.is_load ),
    .Y(_01157_));
 sg13g2_or2_1 _06359_ (.X(_01158_),
    .B(_01157_),
    .A(_01156_));
 sg13g2_nor2_2 _06360_ (.A(_00084_),
    .B(_00877_),
    .Y(_01159_));
 sg13g2_nand2b_1 _06361_ (.Y(_01160_),
    .B(net1365),
    .A_N(_00084_));
 sg13g2_nor3_1 _06362_ (.A(net1394),
    .B(net1374),
    .C(\i_core.cpu.alu_op[3] ),
    .Y(_01161_));
 sg13g2_nor2_2 _06363_ (.A(net1402),
    .B(\i_core.cpu.alu_op[0] ),
    .Y(_01162_));
 sg13g2_and2_2 _06364_ (.A(net1403),
    .B(\i_core.cpu.alu_op[3] ),
    .X(_01163_));
 sg13g2_nand2_2 _06365_ (.Y(_01164_),
    .A(net1402),
    .B(\i_core.cpu.alu_op[3] ));
 sg13g2_nor2_1 _06366_ (.A(net1402),
    .B(_00792_),
    .Y(_01165_));
 sg13g2_nand2_2 _06367_ (.Y(_01166_),
    .A(net1374),
    .B(\i_core.cpu.alu_op[0] ));
 sg13g2_nor2_1 _06368_ (.A(_01163_),
    .B(net1306),
    .Y(_01167_));
 sg13g2_nor3_1 _06369_ (.A(_01161_),
    .B(_01163_),
    .C(net1307),
    .Y(_01168_));
 sg13g2_xor2_1 _06370_ (.B(_01168_),
    .A(_00085_),
    .X(_01169_));
 sg13g2_nand2_2 _06371_ (.Y(_01170_),
    .A(net1390),
    .B(\i_core.cpu.is_alu_imm ));
 sg13g2_o21ai_1 _06372_ (.B1(net1390),
    .Y(_01171_),
    .A1(\i_core.cpu.is_alu_reg ),
    .A2(\i_core.cpu.is_alu_imm ));
 sg13g2_nor3_1 _06373_ (.A(\i_core.cpu.i_core.cycle[1] ),
    .B(_01169_),
    .C(_01171_),
    .Y(_01172_));
 sg13g2_and2_1 _06374_ (.A(\i_core.cpu.is_store ),
    .B(\i_core.cpu.no_write_in_progress ),
    .X(_01173_));
 sg13g2_nand2_2 _06375_ (.Y(_01174_),
    .A(\i_core.cpu.is_store ),
    .B(net2392));
 sg13g2_o21ai_1 _06376_ (.B1(net1390),
    .Y(_01175_),
    .A1(\i_core.cpu.is_branch ),
    .A2(_01173_));
 sg13g2_nand2_2 _06377_ (.Y(_01176_),
    .A(net1390),
    .B(\i_core.cpu.is_lui ));
 sg13g2_and2_2 _06378_ (.A(net1391),
    .B(\i_core.cpu.is_system ),
    .X(_01177_));
 sg13g2_nand2_1 _06379_ (.Y(_01178_),
    .A(net1391),
    .B(\i_core.cpu.is_system ));
 sg13g2_o21ai_1 _06380_ (.B1(net1390),
    .Y(_01179_),
    .A1(\i_core.cpu.is_system ),
    .A2(\i_core.cpu.is_jalr ));
 sg13g2_nand3_1 _06381_ (.B(\i_core.cpu.i_core.load_done ),
    .C(_01171_),
    .A(\i_core.cpu.is_load ),
    .Y(_01180_));
 sg13g2_and4_1 _06382_ (.A(_01158_),
    .B(_01176_),
    .C(_01179_),
    .D(_01180_),
    .X(_01181_));
 sg13g2_nand4_1 _06383_ (.B(_00873_),
    .C(_01175_),
    .A(_00086_),
    .Y(_01182_),
    .D(_01181_));
 sg13g2_o21ai_1 _06384_ (.B1(_01159_),
    .Y(_01183_),
    .A1(_01172_),
    .A2(_01182_));
 sg13g2_nand2b_2 _06385_ (.Y(_01184_),
    .B(_01158_),
    .A_N(_01183_));
 sg13g2_o21ai_1 _06386_ (.B1(_01184_),
    .Y(_00029_),
    .A1(net2424),
    .A2(_01183_));
 sg13g2_nor3_2 _06387_ (.A(\addr[27] ),
    .B(\addr[26] ),
    .C(\addr[25] ),
    .Y(_01185_));
 sg13g2_or3_2 _06388_ (.A(\addr[27] ),
    .B(\addr[26] ),
    .C(\addr[25] ),
    .X(_01186_));
 sg13g2_a21oi_2 _06389_ (.B1(_01186_),
    .Y(_01187_),
    .A2(\i_core.cpu.data_write_n[1] ),
    .A1(\i_core.cpu.data_read_n[1] ));
 sg13g2_xnor2_1 _06390_ (.Y(_01188_),
    .A(\i_core.mem.qspi_data_byte_idx[1] ),
    .B(_01187_));
 sg13g2_nand2_1 _06391_ (.Y(_01189_),
    .A(\i_core.cpu.data_read_n[0] ),
    .B(\i_core.cpu.data_write_n[0] ));
 sg13g2_nand2_2 _06392_ (.Y(_01190_),
    .A(_01187_),
    .B(_01189_));
 sg13g2_xnor2_1 _06393_ (.Y(_01191_),
    .A(_00157_),
    .B(_01190_));
 sg13g2_nor2_1 _06394_ (.A(_01188_),
    .B(_01191_),
    .Y(_01192_));
 sg13g2_and2_1 _06395_ (.A(net2505),
    .B(_01192_),
    .X(_00082_));
 sg13g2_mux2_2 _06396_ (.A0(\i_uart_tx.txd_reg ),
    .A1(\gpio_out[0] ),
    .S(\gpio_out_sel[0] ),
    .X(uo_out[0]));
 sg13g2_nand2b_1 _06397_ (.Y(_01193_),
    .B(\i_spi.spi_select ),
    .A_N(debug_register_data));
 sg13g2_a21oi_1 _06398_ (.A1(\debug_rd_r[2] ),
    .A2(debug_register_data),
    .Y(_01194_),
    .B1(\gpio_out_sel[4] ));
 sg13g2_a22oi_1 _06399_ (.Y(uo_out[4]),
    .B1(_01193_),
    .B2(_01194_),
    .A2(_00828_),
    .A1(\gpio_out_sel[4] ));
 sg13g2_o21ai_1 _06400_ (.B1(_01171_),
    .Y(_01195_),
    .A1(_00747_),
    .A2(_00753_));
 sg13g2_nand3_1 _06401_ (.B(\i_core.cpu.data_ready_core ),
    .C(_01156_),
    .A(\i_core.cpu.is_load ),
    .Y(_01196_));
 sg13g2_nor2b_1 _06402_ (.A(_01195_),
    .B_N(_01196_),
    .Y(_01197_));
 sg13g2_o21ai_1 _06403_ (.B1(net1392),
    .Y(_01198_),
    .A1(\i_core.cpu.is_jal ),
    .A2(\i_core.cpu.is_jalr ));
 sg13g2_a21oi_2 _06404_ (.B1(_00747_),
    .Y(_01199_),
    .A2(_00751_),
    .A1(_00750_));
 sg13g2_nand2_1 _06405_ (.Y(_01200_),
    .A(\i_core.cpu.instr_len[2] ),
    .B(\i_core.cpu.pc[2] ));
 sg13g2_nor2_1 _06406_ (.A(\i_core.cpu.instr_len[2] ),
    .B(\i_core.cpu.pc[2] ),
    .Y(_01201_));
 sg13g2_xor2_1 _06407_ (.B(\i_core.cpu.pc[2] ),
    .A(\i_core.cpu.instr_len[2] ),
    .X(_01202_));
 sg13g2_nand2_1 _06408_ (.Y(_01203_),
    .A(\i_core.cpu.instr_len[1] ),
    .B(\i_core.cpu.pc[1] ));
 sg13g2_o21ai_1 _06409_ (.B1(_01200_),
    .Y(_01204_),
    .A1(_01201_),
    .A2(_01203_));
 sg13g2_nand2_2 _06410_ (.Y(_01205_),
    .A(\i_core.cpu.instr_data_start[3] ),
    .B(_01204_));
 sg13g2_nor2_1 _06411_ (.A(_00163_),
    .B(_01205_),
    .Y(_01206_));
 sg13g2_nor4_2 _06412_ (.A(_00764_),
    .B(_00765_),
    .C(_00163_),
    .Y(_01207_),
    .D(_01205_));
 sg13g2_nand3_1 _06413_ (.B(net1427),
    .C(_01207_),
    .A(\i_core.cpu.instr_data_start[8] ),
    .Y(_01208_));
 sg13g2_nor2_1 _06414_ (.A(_00763_),
    .B(_01208_),
    .Y(_01209_));
 sg13g2_nor3_2 _06415_ (.A(_00762_),
    .B(_00763_),
    .C(_01208_),
    .Y(_01210_));
 sg13g2_nand3_1 _06416_ (.B(\i_core.cpu.instr_data_start[11] ),
    .C(_01210_),
    .A(\i_core.cpu.instr_data_start[12] ),
    .Y(_01211_));
 sg13g2_a21o_1 _06417_ (.A2(_01210_),
    .A1(\i_core.cpu.instr_data_start[11] ),
    .B1(\i_core.cpu.instr_data_start[12] ),
    .X(_01212_));
 sg13g2_nand2_1 _06418_ (.Y(_01213_),
    .A(_01211_),
    .B(_01212_));
 sg13g2_inv_1 _06419_ (.Y(_01214_),
    .A(_01213_));
 sg13g2_a21o_1 _06420_ (.A2(_01207_),
    .A1(net1427),
    .B1(\i_core.cpu.instr_data_start[8] ),
    .X(_01215_));
 sg13g2_nand2_1 _06421_ (.Y(_01216_),
    .A(_01208_),
    .B(_01215_));
 sg13g2_xor2_1 _06422_ (.B(_01205_),
    .A(_00163_),
    .X(_01217_));
 sg13g2_a22oi_1 _06423_ (.Y(_01218_),
    .B1(_01217_),
    .B2(net1361),
    .A2(_01214_),
    .A1(net1364));
 sg13g2_o21ai_1 _06424_ (.B1(_01218_),
    .Y(_01219_),
    .A1(_00882_),
    .A2(_01216_));
 sg13g2_nor2_1 _06425_ (.A(_00760_),
    .B(_01211_),
    .Y(_01220_));
 sg13g2_and3_1 _06426_ (.X(_01221_),
    .A(\i_core.cpu.instr_data_start[15] ),
    .B(\i_core.cpu.instr_data_start[14] ),
    .C(_01220_));
 sg13g2_nand3_1 _06427_ (.B(\i_core.cpu.instr_data_start[16] ),
    .C(_01221_),
    .A(\i_core.cpu.instr_data_start[17] ),
    .Y(_01222_));
 sg13g2_nor2_1 _06428_ (.A(_00758_),
    .B(_01222_),
    .Y(_01223_));
 sg13g2_nor3_1 _06429_ (.A(_00758_),
    .B(_00165_),
    .C(_01222_),
    .Y(_01224_));
 sg13g2_xnor2_1 _06430_ (.Y(_01225_),
    .A(\i_core.cpu.instr_data_start[20] ),
    .B(_01224_));
 sg13g2_nand2_1 _06431_ (.Y(_01226_),
    .A(net1413),
    .B(_01225_));
 sg13g2_nand2_2 _06432_ (.Y(_01227_),
    .A(net1405),
    .B(_00092_));
 sg13g2_xnor2_1 _06433_ (.Y(_01228_),
    .A(\i_core.cpu.instr_data_start[16] ),
    .B(_01221_));
 sg13g2_a21oi_1 _06434_ (.A1(net1378),
    .A2(_01228_),
    .Y(_01229_),
    .B1(_01227_));
 sg13g2_a22oi_1 _06435_ (.Y(_01230_),
    .B1(_01226_),
    .B2(_01229_),
    .A2(_01219_),
    .A1(net1381));
 sg13g2_nor2_1 _06436_ (.A(_01162_),
    .B(_01178_),
    .Y(_01231_));
 sg13g2_nand2b_2 _06437_ (.Y(_01232_),
    .B(_01177_),
    .A_N(_01162_));
 sg13g2_nor2_2 _06438_ (.A(_01199_),
    .B(_01232_),
    .Y(_01233_));
 sg13g2_nor2_2 _06439_ (.A(_00084_),
    .B(_00875_),
    .Y(_01234_));
 sg13g2_nand2b_2 _06440_ (.Y(_01235_),
    .B(net1366),
    .A_N(_00084_));
 sg13g2_nand2_1 _06441_ (.Y(_01236_),
    .A(\i_core.cpu.i_core.imm_lo[8] ),
    .B(\i_core.cpu.i_core.imm_lo[9] ));
 sg13g2_nor3_2 _06442_ (.A(\i_core.cpu.i_core.imm_lo[11] ),
    .B(\i_core.cpu.i_core.imm_lo[10] ),
    .C(_01236_),
    .Y(_01237_));
 sg13g2_nor3_2 _06443_ (.A(\i_core.cpu.i_core.imm_lo[7] ),
    .B(\i_core.cpu.i_core.imm_lo[5] ),
    .C(\i_core.cpu.i_core.imm_lo[4] ),
    .Y(_01238_));
 sg13g2_nand3_1 _06444_ (.B(_01237_),
    .C(_01238_),
    .A(\i_core.cpu.i_core.imm_lo[6] ),
    .Y(_01239_));
 sg13g2_nor2_1 _06445_ (.A(\i_core.cpu.i_core.imm_lo[1] ),
    .B(\i_core.cpu.i_core.imm_lo[0] ),
    .Y(_01240_));
 sg13g2_nand3_1 _06446_ (.B(\i_core.cpu.i_core.imm_lo[2] ),
    .C(_01240_),
    .A(_00797_),
    .Y(_01241_));
 sg13g2_inv_1 _06447_ (.Y(_01242_),
    .A(_01241_));
 sg13g2_nor3_2 _06448_ (.A(_01235_),
    .B(_01239_),
    .C(_01241_),
    .Y(_01243_));
 sg13g2_nor2_1 _06449_ (.A(\i_core.cpu.i_core.imm_lo[3] ),
    .B(\i_core.cpu.i_core.imm_lo[2] ),
    .Y(_01244_));
 sg13g2_nand3_1 _06450_ (.B(_00803_),
    .C(_01244_),
    .A(\i_core.cpu.i_core.imm_lo[1] ),
    .Y(_01245_));
 sg13g2_nor2_1 _06451_ (.A(_01239_),
    .B(_01245_),
    .Y(_01246_));
 sg13g2_nor3_2 _06452_ (.A(net1311),
    .B(_01239_),
    .C(_01245_),
    .Y(_01247_));
 sg13g2_a22oi_1 _06453_ (.Y(_01248_),
    .B1(_01247_),
    .B2(\i_core.cpu.i_core.mcause[0] ),
    .A2(_01243_),
    .A1(\i_core.cpu.i_core.mip[16] ));
 sg13g2_and2_1 _06454_ (.A(_00801_),
    .B(_01238_),
    .X(_01249_));
 sg13g2_and2_1 _06455_ (.A(_01237_),
    .B(_01249_),
    .X(_01250_));
 sg13g2_and3_2 _06456_ (.X(_01251_),
    .A(_01234_),
    .B(_01242_),
    .C(_01250_));
 sg13g2_nor3_1 _06457_ (.A(\i_core.cpu.i_core.imm_lo[3] ),
    .B(\i_core.cpu.i_core.imm_lo[2] ),
    .C(\i_core.cpu.i_core.imm_lo[1] ),
    .Y(_01252_));
 sg13g2_inv_1 _06458_ (.Y(_01253_),
    .A(_01252_));
 sg13g2_nor2_1 _06459_ (.A(_00803_),
    .B(_01253_),
    .Y(_01254_));
 sg13g2_nand2b_1 _06460_ (.Y(_01255_),
    .B(_01254_),
    .A_N(_01239_));
 sg13g2_nor2_2 _06461_ (.A(net1354),
    .B(_01255_),
    .Y(_01256_));
 sg13g2_a22oi_1 _06462_ (.Y(_01257_),
    .B1(_01256_),
    .B2(\i_core.cpu.i_core.mepc[0] ),
    .A2(_01251_),
    .A1(\i_core.cpu.i_core.mie[16] ));
 sg13g2_nor2_1 _06463_ (.A(\i_core.cpu.i_core.imm_lo[8] ),
    .B(\i_core.cpu.i_core.imm_lo[9] ),
    .Y(_01258_));
 sg13g2_nand4_1 _06464_ (.B(\i_core.cpu.i_core.imm_lo[10] ),
    .C(_01249_),
    .A(\i_core.cpu.i_core.imm_lo[11] ),
    .Y(_01259_),
    .D(_01258_));
 sg13g2_nor3_2 _06465_ (.A(_00803_),
    .B(_01253_),
    .C(_01259_),
    .Y(_01260_));
 sg13g2_nor3_2 _06466_ (.A(\i_core.cpu.i_core.imm_lo[0] ),
    .B(_01253_),
    .C(_01259_),
    .Y(_01261_));
 sg13g2_nor2_1 _06467_ (.A(_01245_),
    .B(_01259_),
    .Y(_01262_));
 sg13g2_nor3_1 _06468_ (.A(_00164_),
    .B(_01245_),
    .C(_01259_),
    .Y(_01263_));
 sg13g2_a221oi_1 _06469_ (.B2(\i_core.cpu.i_core.cycle_count[0] ),
    .C1(_01263_),
    .B1(_01261_),
    .A1(\i_core.cpu.i_core.cycle_count[3] ),
    .Y(_01264_),
    .A2(_01260_));
 sg13g2_nand2_1 _06470_ (.Y(_01265_),
    .A(_00084_),
    .B(net1362));
 sg13g2_nand2_1 _06471_ (.Y(_01266_),
    .A(_01250_),
    .B(_01254_));
 sg13g2_and3_1 _06472_ (.X(_01267_),
    .A(\i_core.cpu.i_core.mcause[4] ),
    .B(net1311),
    .C(_01246_));
 sg13g2_nand3_1 _06473_ (.B(net1311),
    .C(_01246_),
    .A(\i_core.cpu.i_core.mcause[4] ),
    .Y(_01268_));
 sg13g2_a21o_1 _06474_ (.A2(_01268_),
    .A1(_01266_),
    .B1(_01265_),
    .X(_01269_));
 sg13g2_nand4_1 _06475_ (.B(_01257_),
    .C(_01264_),
    .A(_01248_),
    .Y(_01270_),
    .D(_01269_));
 sg13g2_a22oi_1 _06476_ (.Y(_01271_),
    .B1(_01233_),
    .B2(_01270_),
    .A2(\i_core.cpu.is_lui ),
    .A1(net1391));
 sg13g2_o21ai_1 _06477_ (.B1(_01271_),
    .Y(_01272_),
    .A1(_01198_),
    .A2(_01230_));
 sg13g2_o21ai_1 _06478_ (.B1(_01272_),
    .Y(_01273_),
    .A1(_01102_),
    .A2(_01176_));
 sg13g2_nor3_2 _06479_ (.A(net1394),
    .B(net1402),
    .C(\i_core.cpu.alu_op[0] ),
    .Y(_01274_));
 sg13g2_nand2_2 _06480_ (.Y(_01275_),
    .A(net1375),
    .B(_01162_));
 sg13g2_a21oi_1 _06481_ (.A1(_01131_),
    .A2(_01135_),
    .Y(_01276_),
    .B1(_01275_));
 sg13g2_o21ai_1 _06482_ (.B1(_01276_),
    .Y(_01277_),
    .A1(_01131_),
    .A2(_01135_));
 sg13g2_nand3_1 _06483_ (.B(_01096_),
    .C(_01125_),
    .A(net1374),
    .Y(_01278_));
 sg13g2_nand2_2 _06484_ (.Y(_01279_),
    .A(net1394),
    .B(_00792_));
 sg13g2_o21ai_1 _06485_ (.B1(_01278_),
    .Y(_01280_),
    .A1(_01096_),
    .A2(_01125_));
 sg13g2_nor3_2 _06486_ (.A(net1375),
    .B(net1374),
    .C(_00792_),
    .Y(_01281_));
 sg13g2_nand3_1 _06487_ (.B(_01125_),
    .C(_01281_),
    .A(_01096_),
    .Y(_01282_));
 sg13g2_o21ai_1 _06488_ (.B1(_01282_),
    .Y(_01283_),
    .A1(_01279_),
    .A2(_01280_));
 sg13g2_nor2b_1 _06489_ (.A(_01283_),
    .B_N(_01277_),
    .Y(_01284_));
 sg13g2_a21o_1 _06490_ (.A2(_00166_),
    .A1(net1403),
    .B1(net1307),
    .X(_01285_));
 sg13g2_or2_1 _06491_ (.X(_01286_),
    .B(_01285_),
    .A(_01284_));
 sg13g2_nand2_1 _06492_ (.Y(_01287_),
    .A(\i_core.cpu.alu_op[3] ),
    .B(\i_core.cpu.i_core.i_shift.a[31] ));
 sg13g2_xnor2_1 _06493_ (.Y(_01288_),
    .A(net1407),
    .B(net1394));
 sg13g2_xnor2_1 _06494_ (.Y(_01289_),
    .A(net1410),
    .B(net1394));
 sg13g2_nand2_1 _06495_ (.Y(_01290_),
    .A(\i_core.cpu.i_core.i_shift.b[3] ),
    .B(_01289_));
 sg13g2_xor2_1 _06496_ (.B(_01289_),
    .A(\i_core.cpu.i_core.i_shift.b[3] ),
    .X(_01291_));
 sg13g2_xnor2_1 _06497_ (.Y(_01292_),
    .A(net1416),
    .B(net1401));
 sg13g2_nand2_1 _06498_ (.Y(_01293_),
    .A(\i_core.cpu.i_core.i_shift.b[2] ),
    .B(_01292_));
 sg13g2_nand3_1 _06499_ (.B(_01291_),
    .C(_01292_),
    .A(\i_core.cpu.i_core.i_shift.b[2] ),
    .Y(_01294_));
 sg13g2_nand2_1 _06500_ (.Y(_01295_),
    .A(_01290_),
    .B(_01294_));
 sg13g2_a21o_1 _06501_ (.A2(_01288_),
    .A1(\i_core.cpu.i_core.i_shift.b[4] ),
    .B1(_01295_),
    .X(_01296_));
 sg13g2_o21ai_1 _06502_ (.B1(_01296_),
    .Y(_01297_),
    .A1(\i_core.cpu.i_core.i_shift.b[4] ),
    .A2(_01288_));
 sg13g2_nand2b_2 _06503_ (.Y(_01298_),
    .B(_01287_),
    .A_N(_01297_));
 sg13g2_and2_1 _06504_ (.A(net1399),
    .B(_00186_),
    .X(_01299_));
 sg13g2_a21oi_1 _06505_ (.A1(net1376),
    .A2(_00185_),
    .Y(_01300_),
    .B1(_01299_));
 sg13g2_mux2_1 _06506_ (.A0(_00183_),
    .A1(_00184_),
    .S(net1398),
    .X(_01301_));
 sg13g2_nand2_1 _06507_ (.Y(_01302_),
    .A(net1448),
    .B(_01301_));
 sg13g2_o21ai_1 _06508_ (.B1(_01302_),
    .Y(_01303_),
    .A1(net1448),
    .A2(_01300_));
 sg13g2_xor2_1 _06509_ (.B(_01292_),
    .A(\i_core.cpu.i_core.i_shift.b[2] ),
    .X(_01304_));
 sg13g2_xnor2_1 _06510_ (.Y(_01305_),
    .A(\i_core.cpu.i_core.i_shift.b[2] ),
    .B(_01292_));
 sg13g2_mux4_1 _06511_ (.S0(net1399),
    .A0(_00181_),
    .A1(_00182_),
    .A2(_00179_),
    .A3(_00180_),
    .S1(net1448),
    .X(_01306_));
 sg13g2_nand2_1 _06512_ (.Y(_01307_),
    .A(net1440),
    .B(_01306_));
 sg13g2_a21oi_1 _06513_ (.A1(net1372),
    .A2(_01303_),
    .Y(_01308_),
    .B1(net1305));
 sg13g2_xnor2_1 _06514_ (.Y(_01309_),
    .A(\i_core.cpu.i_core.i_shift.b[4] ),
    .B(_01288_));
 sg13g2_nor2b_2 _06515_ (.A(_01295_),
    .B_N(_01309_),
    .Y(_01310_));
 sg13g2_nand3_1 _06516_ (.B(_01294_),
    .C(_01309_),
    .A(_01290_),
    .Y(_01311_));
 sg13g2_mux4_1 _06517_ (.S0(net1398),
    .A0(_00173_),
    .A1(_00174_),
    .A2(_00171_),
    .A3(_00172_),
    .S1(net1449),
    .X(_01312_));
 sg13g2_mux4_1 _06518_ (.S0(net1396),
    .A0(_00177_),
    .A1(_00178_),
    .A2(_00175_),
    .A3(_00176_),
    .S1(net1447),
    .X(_01313_));
 sg13g2_nand2_1 _06519_ (.Y(_01314_),
    .A(net1371),
    .B(_01313_));
 sg13g2_a21oi_1 _06520_ (.A1(net1441),
    .A2(_01312_),
    .Y(_01315_),
    .B1(net1302));
 sg13g2_a221oi_1 _06521_ (.B2(_01315_),
    .C1(_01310_),
    .B1(_01314_),
    .A1(_01307_),
    .Y(_01316_),
    .A2(_01308_));
 sg13g2_mux4_1 _06522_ (.S0(net1398),
    .A0(_00172_),
    .A1(_00171_),
    .A2(_00174_),
    .A3(_00173_),
    .S1(net1449),
    .X(_01317_));
 sg13g2_inv_1 _06523_ (.Y(_01318_),
    .A(_01317_));
 sg13g2_nor2_1 _06524_ (.A(net1373),
    .B(_01318_),
    .Y(_01319_));
 sg13g2_mux4_1 _06525_ (.S0(net1395),
    .A0(_00167_),
    .A1(_00168_),
    .A2(_00170_),
    .A3(_00169_),
    .S1(net1443),
    .X(_01320_));
 sg13g2_a21oi_1 _06526_ (.A1(net1373),
    .A2(_01320_),
    .Y(_01321_),
    .B1(_01319_));
 sg13g2_mux4_1 _06527_ (.S0(net1396),
    .A0(_00176_),
    .A1(_00175_),
    .A2(_00178_),
    .A3(_00177_),
    .S1(net1447),
    .X(_01322_));
 sg13g2_nand2_1 _06528_ (.Y(_01323_),
    .A(net1373),
    .B(_01322_));
 sg13g2_mux4_1 _06529_ (.S0(net1398),
    .A0(_00180_),
    .A1(_00179_),
    .A2(_00182_),
    .A3(_00181_),
    .S1(net1448),
    .X(_01324_));
 sg13g2_a21oi_1 _06530_ (.A1(net1440),
    .A2(_01324_),
    .Y(_01325_),
    .B1(net1301));
 sg13g2_a221oi_1 _06531_ (.B2(_01325_),
    .C1(_01311_),
    .B1(_01323_),
    .A1(net1302),
    .Y(_01326_),
    .A2(_01321_));
 sg13g2_xnor2_1 _06532_ (.Y(_01327_),
    .A(_01291_),
    .B(_01293_));
 sg13g2_nor3_1 _06533_ (.A(_01316_),
    .B(_01326_),
    .C(_01327_),
    .Y(_01328_));
 sg13g2_mux2_1 _06534_ (.A0(_00194_),
    .A1(_00193_),
    .S(net1401),
    .X(_01329_));
 sg13g2_nor2_1 _06535_ (.A(net1442),
    .B(_01329_),
    .Y(_01330_));
 sg13g2_and2_1 _06536_ (.A(net1395),
    .B(_00195_),
    .X(_01331_));
 sg13g2_a21oi_1 _06537_ (.A1(net1376),
    .A2(_00196_),
    .Y(_01332_),
    .B1(_01331_));
 sg13g2_a21oi_1 _06538_ (.A1(net1442),
    .A2(_01332_),
    .Y(_01333_),
    .B1(_01330_));
 sg13g2_nand2_1 _06539_ (.Y(_01334_),
    .A(net1438),
    .B(_01333_));
 sg13g2_mux2_1 _06540_ (.A0(_00169_),
    .A1(_00170_),
    .S(net1395),
    .X(_01335_));
 sg13g2_nor2_1 _06541_ (.A(net1443),
    .B(_01335_),
    .Y(_01336_));
 sg13g2_and2_1 _06542_ (.A(net1395),
    .B(_00167_),
    .X(_01337_));
 sg13g2_a21oi_1 _06543_ (.A1(net1376),
    .A2(_00168_),
    .Y(_01338_),
    .B1(_01337_));
 sg13g2_a21oi_1 _06544_ (.A1(net1443),
    .A2(_01338_),
    .Y(_01339_),
    .B1(_01336_));
 sg13g2_a21oi_1 _06545_ (.A1(net1369),
    .A2(_01339_),
    .Y(_01340_),
    .B1(net1304));
 sg13g2_a21oi_1 _06546_ (.A1(net1438),
    .A2(_01287_),
    .Y(_01341_),
    .B1(net1303));
 sg13g2_mux2_1 _06547_ (.A0(_00198_),
    .A1(_00197_),
    .S(net1395),
    .X(_01342_));
 sg13g2_nand3_1 _06548_ (.B(\i_core.cpu.i_core.i_shift.a[31] ),
    .C(net1444),
    .A(\i_core.cpu.alu_op[3] ),
    .Y(_01343_));
 sg13g2_o21ai_1 _06549_ (.B1(_01343_),
    .Y(_01344_),
    .A1(net1442),
    .A2(_01342_));
 sg13g2_nand2b_1 _06550_ (.Y(_01345_),
    .B(net1369),
    .A_N(_01344_));
 sg13g2_a221oi_1 _06551_ (.B2(_01345_),
    .C1(_01310_),
    .B1(_01341_),
    .A1(_01334_),
    .Y(_01346_),
    .A2(_01340_));
 sg13g2_mux2_1 _06552_ (.A0(_00184_),
    .A1(_00183_),
    .S(net1399),
    .X(_01347_));
 sg13g2_nor2_1 _06553_ (.A(net1448),
    .B(_01347_),
    .Y(_01348_));
 sg13g2_and2_1 _06554_ (.A(net1399),
    .B(_00185_),
    .X(_01349_));
 sg13g2_a21oi_1 _06555_ (.A1(net1376),
    .A2(_00186_),
    .Y(_01350_),
    .B1(_01349_));
 sg13g2_a21oi_1 _06556_ (.A1(net1448),
    .A2(_01350_),
    .Y(_01351_),
    .B1(_01348_));
 sg13g2_mux2_1 _06557_ (.A0(_00188_),
    .A1(_00187_),
    .S(net1397),
    .X(_01352_));
 sg13g2_mux2_1 _06558_ (.A0(_00190_),
    .A1(_00189_),
    .S(net1397),
    .X(_01353_));
 sg13g2_mux2_1 _06559_ (.A0(_01352_),
    .A1(_01353_),
    .S(net1445),
    .X(_01354_));
 sg13g2_a21o_1 _06560_ (.A2(_01354_),
    .A1(net1440),
    .B1(net1305),
    .X(_01355_));
 sg13g2_a21oi_1 _06561_ (.A1(net1371),
    .A2(_01351_),
    .Y(_01356_),
    .B1(_01355_));
 sg13g2_mux2_1 _06562_ (.A0(_00192_),
    .A1(_00191_),
    .S(net1397),
    .X(_01357_));
 sg13g2_nor2_1 _06563_ (.A(net1445),
    .B(_01357_),
    .Y(_01358_));
 sg13g2_and2_1 _06564_ (.A(net1397),
    .B(_00192_),
    .X(_01359_));
 sg13g2_a21oi_1 _06565_ (.A1(net1376),
    .A2(_00191_),
    .Y(_01360_),
    .B1(_01359_));
 sg13g2_a21oi_1 _06566_ (.A1(net1446),
    .A2(_01360_),
    .Y(_01361_),
    .B1(_01358_));
 sg13g2_mux2_1 _06567_ (.A0(_00189_),
    .A1(_00190_),
    .S(net1396),
    .X(_01362_));
 sg13g2_mux2_1 _06568_ (.A0(_00187_),
    .A1(_00188_),
    .S(net1396),
    .X(_01363_));
 sg13g2_mux2_1 _06569_ (.A0(_01362_),
    .A1(_01363_),
    .S(net1445),
    .X(_01364_));
 sg13g2_mux2_1 _06570_ (.A0(_01361_),
    .A1(_01364_),
    .S(net1440),
    .X(_01365_));
 sg13g2_o21ai_1 _06571_ (.B1(_01310_),
    .Y(_01366_),
    .A1(net1301),
    .A2(_01365_));
 sg13g2_o21ai_1 _06572_ (.B1(net1277),
    .Y(_01367_),
    .A1(_01356_),
    .A2(_01366_));
 sg13g2_o21ai_1 _06573_ (.B1(_01297_),
    .Y(_01368_),
    .A1(_01346_),
    .A2(_01367_));
 sg13g2_o21ai_1 _06574_ (.B1(_01298_),
    .Y(_01369_),
    .A1(_01328_),
    .A2(_01368_));
 sg13g2_nor2_2 _06575_ (.A(\i_core.cpu.i_core.cycle[1] ),
    .B(_00785_),
    .Y(_01370_));
 sg13g2_and2_1 _06576_ (.A(net1306),
    .B(_01370_),
    .X(_01371_));
 sg13g2_nand2_1 _06577_ (.Y(_01372_),
    .A(net1306),
    .B(_01370_));
 sg13g2_nand2_1 _06578_ (.Y(_01373_),
    .A(net1445),
    .B(_01362_));
 sg13g2_o21ai_1 _06579_ (.B1(_01373_),
    .Y(_01374_),
    .A1(net1445),
    .A2(_01360_));
 sg13g2_nor2_1 _06580_ (.A(net1445),
    .B(_01363_),
    .Y(_01375_));
 sg13g2_a21oi_2 _06581_ (.B1(_01375_),
    .Y(_01376_),
    .A2(_01300_),
    .A1(net1448));
 sg13g2_nand2_1 _06582_ (.Y(_01377_),
    .A(net1439),
    .B(_01376_));
 sg13g2_a21oi_1 _06583_ (.A1(net1372),
    .A2(_01374_),
    .Y(_01378_),
    .B1(net1305));
 sg13g2_mux4_1 _06584_ (.S0(net1396),
    .A0(_00179_),
    .A1(_00180_),
    .A2(_00177_),
    .A3(_00178_),
    .S1(net1446),
    .X(_01379_));
 sg13g2_nand2_1 _06585_ (.Y(_01380_),
    .A(net1439),
    .B(_01379_));
 sg13g2_mux4_1 _06586_ (.S0(net1398),
    .A0(_00183_),
    .A1(_00184_),
    .A2(_00181_),
    .A3(_00182_),
    .S1(net1449),
    .X(_01381_));
 sg13g2_a21oi_1 _06587_ (.A1(net1371),
    .A2(_01381_),
    .Y(_01382_),
    .B1(net1301));
 sg13g2_a221oi_1 _06588_ (.B2(_01382_),
    .C1(net1277),
    .B1(_01380_),
    .A1(_01377_),
    .Y(_01383_),
    .A2(_01378_));
 sg13g2_nand2_1 _06589_ (.Y(_01384_),
    .A(net1442),
    .B(_01342_));
 sg13g2_o21ai_1 _06590_ (.B1(_01384_),
    .Y(_01385_),
    .A1(net1442),
    .A2(_01332_));
 sg13g2_nand2_1 _06591_ (.Y(_01386_),
    .A(net1438),
    .B(_01385_));
 sg13g2_nand2_1 _06592_ (.Y(_01387_),
    .A(net1443),
    .B(_01329_));
 sg13g2_o21ai_1 _06593_ (.B1(_01387_),
    .Y(_01388_),
    .A1(net1443),
    .A2(_01338_));
 sg13g2_a21oi_1 _06594_ (.A1(net1369),
    .A2(_01388_),
    .Y(_01389_),
    .B1(net1303));
 sg13g2_mux4_1 _06595_ (.S0(net1396),
    .A0(_00175_),
    .A1(_00176_),
    .A2(_00173_),
    .A3(_00174_),
    .S1(net1447),
    .X(_01390_));
 sg13g2_mux4_1 _06596_ (.S0(net1398),
    .A0(_00171_),
    .A1(_00172_),
    .A2(_00169_),
    .A3(_00170_),
    .S1(net1449),
    .X(_01391_));
 sg13g2_mux2_1 _06597_ (.A0(_01390_),
    .A1(_01391_),
    .S(net1438),
    .X(_01392_));
 sg13g2_o21ai_1 _06598_ (.B1(net1277),
    .Y(_01393_),
    .A1(net1304),
    .A2(_01392_));
 sg13g2_a21oi_1 _06599_ (.A1(_01386_),
    .A2(_01389_),
    .Y(_01394_),
    .B1(_01393_));
 sg13g2_or3_1 _06600_ (.A(_01310_),
    .B(_01383_),
    .C(_01394_),
    .X(_01395_));
 sg13g2_mux4_1 _06601_ (.S0(net1395),
    .A0(_00193_),
    .A1(_00194_),
    .A2(_00167_),
    .A3(_00168_),
    .S1(net1442),
    .X(_01396_));
 sg13g2_mux4_1 _06602_ (.S0(net1395),
    .A0(_00197_),
    .A1(_00198_),
    .A2(_00195_),
    .A3(_00196_),
    .S1(net1442),
    .X(_01397_));
 sg13g2_mux4_1 _06603_ (.S0(net1396),
    .A0(_00174_),
    .A1(_00173_),
    .A2(_00176_),
    .A3(_00175_),
    .S1(net1447),
    .X(_01398_));
 sg13g2_mux4_1 _06604_ (.S0(net1398),
    .A0(_00170_),
    .A1(_00169_),
    .A2(_00172_),
    .A3(_00171_),
    .S1(net1449),
    .X(_01399_));
 sg13g2_mux4_1 _06605_ (.S0(net1369),
    .A0(_01396_),
    .A1(_01397_),
    .A2(_01398_),
    .A3(_01399_),
    .S1(net1304),
    .X(_01400_));
 sg13g2_nand2b_1 _06606_ (.Y(_01401_),
    .B(_01400_),
    .A_N(net1277));
 sg13g2_nand2_1 _06607_ (.Y(_01402_),
    .A(net1445),
    .B(_01352_));
 sg13g2_o21ai_1 _06608_ (.B1(_01402_),
    .Y(_01403_),
    .A1(net1448),
    .A2(_01350_));
 sg13g2_inv_1 _06609_ (.Y(_01404_),
    .A(_01403_));
 sg13g2_mux2_1 _06610_ (.A0(_01353_),
    .A1(_01357_),
    .S(net1445),
    .X(_01405_));
 sg13g2_a21oi_1 _06611_ (.A1(net1439),
    .A2(_01405_),
    .Y(_01406_),
    .B1(net1301));
 sg13g2_o21ai_1 _06612_ (.B1(_01406_),
    .Y(_01407_),
    .A1(net1439),
    .A2(_01404_));
 sg13g2_mux4_1 _06613_ (.S0(net1398),
    .A0(_00182_),
    .A1(_00181_),
    .A2(_00184_),
    .A3(_00183_),
    .S1(net1449),
    .X(_01408_));
 sg13g2_mux4_1 _06614_ (.S0(net1396),
    .A0(_00178_),
    .A1(_00177_),
    .A2(_00180_),
    .A3(_00179_),
    .S1(net1446),
    .X(_01409_));
 sg13g2_inv_1 _06615_ (.Y(_01410_),
    .A(_01409_));
 sg13g2_a21oi_1 _06616_ (.A1(net1440),
    .A2(_01408_),
    .Y(_01411_),
    .B1(net1305));
 sg13g2_o21ai_1 _06617_ (.B1(_01411_),
    .Y(_01412_),
    .A1(net1439),
    .A2(_01410_));
 sg13g2_nand3_1 _06618_ (.B(_01407_),
    .C(_01412_),
    .A(net1277),
    .Y(_01413_));
 sg13g2_nand3_1 _06619_ (.B(_01401_),
    .C(_01413_),
    .A(_01310_),
    .Y(_01414_));
 sg13g2_nand3_1 _06620_ (.B(_01395_),
    .C(_01414_),
    .A(_01297_),
    .Y(_01415_));
 sg13g2_and2_1 _06621_ (.A(_01298_),
    .B(_01415_),
    .X(_01416_));
 sg13g2_o21ai_1 _06622_ (.B1(_01371_),
    .Y(_01417_),
    .A1(net1375),
    .A2(_01416_));
 sg13g2_a21oi_1 _06623_ (.A1(net1375),
    .A2(_01369_),
    .Y(_01418_),
    .B1(_01417_));
 sg13g2_a21oi_2 _06624_ (.B1(_00085_),
    .Y(_01419_),
    .A2(_01089_),
    .A1(_01087_));
 sg13g2_a21oi_1 _06625_ (.A1(\i_core.cpu.i_core.i_shift.a[0] ),
    .A2(net1238),
    .Y(_01420_),
    .B1(\i_core.cpu.i_core.multiplier.accum[0] ));
 sg13g2_nand3_1 _06626_ (.B(\i_core.cpu.i_core.multiplier.accum[0] ),
    .C(net1238),
    .A(\i_core.cpu.i_core.i_shift.a[0] ),
    .Y(_01421_));
 sg13g2_nor2_1 _06627_ (.A(_01164_),
    .B(_01420_),
    .Y(_01422_));
 sg13g2_a21oi_1 _06628_ (.A1(_01421_),
    .A2(_01422_),
    .Y(_01423_),
    .B1(_01418_));
 sg13g2_o21ai_1 _06629_ (.B1(_01423_),
    .Y(_01424_),
    .A1(_01163_),
    .A2(_01286_));
 sg13g2_nand3_1 _06630_ (.B(_01161_),
    .C(_01370_),
    .A(net1279),
    .Y(_01425_));
 sg13g2_o21ai_1 _06631_ (.B1(_01195_),
    .Y(_01426_),
    .A1(_00806_),
    .A2(_01425_));
 sg13g2_nor2_1 _06632_ (.A(_01424_),
    .B(_01426_),
    .Y(_01427_));
 sg13g2_nand2_1 _06633_ (.Y(_01428_),
    .A(\i_core.mem.q_ctrl.data_ready ),
    .B(_01192_));
 sg13g2_a21oi_1 _06634_ (.A1(_00151_),
    .A2(_01428_),
    .Y(_01429_),
    .B1(_00813_));
 sg13g2_a21o_2 _06635_ (.A2(_01428_),
    .A1(_00151_),
    .B1(_00813_),
    .X(_01430_));
 sg13g2_nor2_2 _06636_ (.A(_01190_),
    .B(_01430_),
    .Y(_01431_));
 sg13g2_and4_1 _06637_ (.A(\i_core.cpu.data_read_n[0] ),
    .B(\i_core.cpu.data_write_n[0] ),
    .C(_01187_),
    .D(_01429_),
    .X(_01432_));
 sg13g2_nand4_1 _06638_ (.B(\i_core.cpu.data_write_n[0] ),
    .C(_01187_),
    .A(\i_core.cpu.data_read_n[0] ),
    .Y(_01433_),
    .D(net1202));
 sg13g2_nand2_2 _06639_ (.Y(_01434_),
    .A(net1408),
    .B(net1335));
 sg13g2_mux4_1 _06640_ (.S0(net1411),
    .A0(\i_core.cpu.instr_data_in[8] ),
    .A1(\i_core.cpu.instr_data_in[12] ),
    .A2(\i_core.mem.qspi_data_buf[8] ),
    .A3(\i_core.mem.qspi_data_buf[12] ),
    .S1(net1190),
    .X(_01435_));
 sg13g2_nand2_1 _06641_ (.Y(_01436_),
    .A(net1408),
    .B(_01435_));
 sg13g2_mux4_1 _06642_ (.S0(_01431_),
    .A0(\i_core.cpu.instr_data_in[0] ),
    .A1(\i_core.cpu.instr_data_in[8] ),
    .A2(\i_core.cpu.instr_data_in[4] ),
    .A3(\i_core.cpu.instr_data_in[12] ),
    .S1(net1411),
    .X(_01437_));
 sg13g2_a21oi_1 _06643_ (.A1(_00787_),
    .A2(_01437_),
    .Y(_01438_),
    .B1(_01186_));
 sg13g2_nor4_1 _06644_ (.A(\addr[24] ),
    .B(\addr[1] ),
    .C(\addr[7] ),
    .D(\addr[6] ),
    .Y(_01439_));
 sg13g2_nor3_1 _06645_ (.A(\addr[0] ),
    .B(\addr[26] ),
    .C(\addr[25] ),
    .Y(_01440_));
 sg13g2_nand3_1 _06646_ (.B(_01439_),
    .C(_01440_),
    .A(\addr[27] ),
    .Y(_01441_));
 sg13g2_nor4_1 _06647_ (.A(\addr[13] ),
    .B(\addr[12] ),
    .C(\addr[15] ),
    .D(\addr[14] ),
    .Y(_01442_));
 sg13g2_nor4_1 _06648_ (.A(\addr[9] ),
    .B(\addr[8] ),
    .C(\addr[11] ),
    .D(\addr[10] ),
    .Y(_01443_));
 sg13g2_nor4_1 _06649_ (.A(\addr[17] ),
    .B(\addr[16] ),
    .C(\addr[19] ),
    .D(\addr[18] ),
    .Y(_01444_));
 sg13g2_nor4_2 _06650_ (.A(\addr[21] ),
    .B(\addr[20] ),
    .C(\addr[23] ),
    .Y(_01445_),
    .D(\addr[22] ));
 sg13g2_nand4_1 _06651_ (.B(_01443_),
    .C(_01444_),
    .A(_01442_),
    .Y(_01446_),
    .D(_01445_));
 sg13g2_nor3_2 _06652_ (.A(\addr[3] ),
    .B(_01441_),
    .C(_01446_),
    .Y(_01447_));
 sg13g2_inv_2 _06653_ (.Y(_01448_),
    .A(_01447_));
 sg13g2_nand2_2 _06654_ (.Y(_01449_),
    .A(net1451),
    .B(_01447_));
 sg13g2_nor3_2 _06655_ (.A(\addr[5] ),
    .B(_01441_),
    .C(_01446_),
    .Y(_01450_));
 sg13g2_nor2_1 _06656_ (.A(\addr[9] ),
    .B(\addr[10] ),
    .Y(_01451_));
 sg13g2_nor2_1 _06657_ (.A(\addr[17] ),
    .B(\addr[18] ),
    .Y(_01452_));
 sg13g2_nand4_1 _06658_ (.B(_01445_),
    .C(_01451_),
    .A(_01442_),
    .Y(_01453_),
    .D(_01452_));
 sg13g2_or4_1 _06659_ (.A(\addr[8] ),
    .B(\addr[11] ),
    .C(\addr[16] ),
    .D(\addr[19] ),
    .X(_01454_));
 sg13g2_nor3_1 _06660_ (.A(_01441_),
    .B(_01453_),
    .C(_01454_),
    .Y(_01455_));
 sg13g2_nand2b_1 _06661_ (.Y(_01456_),
    .B(_01455_),
    .A_N(\addr[5] ));
 sg13g2_nor4_1 _06662_ (.A(net1450),
    .B(_00156_),
    .C(_01449_),
    .D(_01450_),
    .Y(_01457_));
 sg13g2_nor4_2 _06663_ (.A(net1451),
    .B(net1450),
    .C(_01448_),
    .Y(_01458_),
    .D(_01450_));
 sg13g2_and2_1 _06664_ (.A(\i_spi.data[0] ),
    .B(_01458_),
    .X(_01459_));
 sg13g2_or3_2 _06665_ (.A(\i_uart_tx.fsm_state[3] ),
    .B(\i_uart_tx.fsm_state[2] ),
    .C(\i_uart_tx.fsm_state[1] ),
    .X(_01460_));
 sg13g2_nor2_2 _06666_ (.A(\i_uart_tx.fsm_state[0] ),
    .B(_01460_),
    .Y(_01461_));
 sg13g2_or2_1 _06667_ (.X(_01462_),
    .B(_01460_),
    .A(\i_uart_tx.fsm_state[0] ));
 sg13g2_nand2_2 _06668_ (.Y(_01463_),
    .A(net1450),
    .B(_01450_));
 sg13g2_nor2_1 _06669_ (.A(_01449_),
    .B(_01463_),
    .Y(_01464_));
 sg13g2_nor3_1 _06670_ (.A(_01449_),
    .B(_01461_),
    .C(_01463_),
    .Y(_01465_));
 sg13g2_nor2b_1 _06671_ (.A(\addr[3] ),
    .B_N(_01455_),
    .Y(_01466_));
 sg13g2_nand2_1 _06672_ (.Y(_01467_),
    .A(net1451),
    .B(_01448_));
 sg13g2_or3_2 _06673_ (.A(\i_debug_uart_tx.fsm_state[3] ),
    .B(\i_debug_uart_tx.fsm_state[2] ),
    .C(\i_debug_uart_tx.fsm_state[1] ),
    .X(_01468_));
 sg13g2_nor2_2 _06674_ (.A(\i_debug_uart_tx.fsm_state[0] ),
    .B(_01468_),
    .Y(_01469_));
 sg13g2_or2_2 _06675_ (.X(_01470_),
    .B(_01468_),
    .A(\i_debug_uart_tx.fsm_state[0] ));
 sg13g2_nor3_1 _06676_ (.A(_01463_),
    .B(_01467_),
    .C(_01469_),
    .Y(_01471_));
 sg13g2_nor4_1 _06677_ (.A(_01457_),
    .B(_01459_),
    .C(_01465_),
    .D(_01471_),
    .Y(_01472_));
 sg13g2_nor2_1 _06678_ (.A(net1451),
    .B(_01463_),
    .Y(_01473_));
 sg13g2_nor3_2 _06679_ (.A(net1451),
    .B(_01448_),
    .C(_01463_),
    .Y(_01474_));
 sg13g2_nand2_1 _06680_ (.Y(_01475_),
    .A(\i_uart_rx.recieved_data[0] ),
    .B(net1235));
 sg13g2_nand2b_2 _06681_ (.Y(_01476_),
    .B(_01450_),
    .A_N(net1450));
 sg13g2_nor3_2 _06682_ (.A(net1451),
    .B(_01448_),
    .C(_01476_),
    .Y(_01477_));
 sg13g2_a21oi_1 _06683_ (.A1(uo_out[0]),
    .A2(_01477_),
    .Y(_01478_),
    .B1(net1416));
 sg13g2_nor2_2 _06684_ (.A(_01449_),
    .B(_01476_),
    .Y(_01479_));
 sg13g2_nor2_2 _06685_ (.A(_01467_),
    .B(_01476_),
    .Y(_01480_));
 sg13g2_a22oi_1 _06686_ (.Y(_01481_),
    .B1(_01480_),
    .B2(\gpio_out_sel[0] ),
    .A2(_01479_),
    .A1(net2));
 sg13g2_nor2b_1 _06687_ (.A(net1451),
    .B_N(_01466_),
    .Y(_01482_));
 sg13g2_nor2_1 _06688_ (.A(net1450),
    .B(_01456_),
    .Y(_01483_));
 sg13g2_nand4_1 _06689_ (.B(_01475_),
    .C(_01478_),
    .A(_01472_),
    .Y(_01484_),
    .D(_01481_));
 sg13g2_nand2_1 _06690_ (.Y(_01485_),
    .A(uo_out[4]),
    .B(_01477_));
 sg13g2_a22oi_1 _06691_ (.Y(_01486_),
    .B1(_01480_),
    .B2(\gpio_out_sel[4] ),
    .A2(net1236),
    .A1(\i_spi.data[4] ));
 sg13g2_a22oi_1 _06692_ (.Y(_01487_),
    .B1(_01479_),
    .B2(net5),
    .A2(net1235),
    .A1(\i_uart_rx.recieved_data[4] ));
 sg13g2_nand4_1 _06693_ (.B(_01485_),
    .C(_01486_),
    .A(net1416),
    .Y(_01488_),
    .D(_01487_));
 sg13g2_nand3_1 _06694_ (.B(_01484_),
    .C(_01488_),
    .A(_00787_),
    .Y(_01489_));
 sg13g2_nor2b_1 _06695_ (.A(_01450_),
    .B_N(net1450),
    .Y(_01490_));
 sg13g2_inv_1 _06696_ (.Y(_01491_),
    .A(_01490_));
 sg13g2_a21oi_1 _06697_ (.A1(net1452),
    .A2(_01450_),
    .Y(_01492_),
    .B1(_01447_));
 sg13g2_nor2_2 _06698_ (.A(_01490_),
    .B(_01492_),
    .Y(_01493_));
 sg13g2_a22oi_1 _06699_ (.Y(_01494_),
    .B1(_01491_),
    .B2(_01447_),
    .A2(_01450_),
    .A1(net1451));
 sg13g2_a22oi_1 _06700_ (.Y(_01495_),
    .B1(_01489_),
    .B2(net1234),
    .A2(_01438_),
    .A1(_01436_));
 sg13g2_nand2b_1 _06701_ (.Y(_01496_),
    .B(net1409),
    .A_N(\i_core.cpu.i_core.mem_op[0] ));
 sg13g2_a21oi_2 _06702_ (.B1(\i_core.cpu.i_core.mem_op[1] ),
    .Y(_01497_),
    .A2(_01496_),
    .A1(net1380));
 sg13g2_mux4_1 _06703_ (.S0(net1411),
    .A0(\i_core.cpu.instr_data_in[8] ),
    .A1(\i_core.cpu.instr_data_in[12] ),
    .A2(\i_core.mem.qspi_data_buf[24] ),
    .A3(\i_core.mem.qspi_data_buf[28] ),
    .S1(_01430_),
    .X(_01498_));
 sg13g2_nor2b_1 _06704_ (.A(_01434_),
    .B_N(_01498_),
    .Y(_01499_));
 sg13g2_a22oi_1 _06705_ (.Y(_01500_),
    .B1(net1360),
    .B2(\i_core.mem.data_from_read[20] ),
    .A2(net1368),
    .A1(\i_core.mem.data_from_read[16] ));
 sg13g2_a21oi_1 _06706_ (.A1(net1335),
    .A2(_01500_),
    .Y(_01501_),
    .B1(net1234));
 sg13g2_nor3_1 _06707_ (.A(net1380),
    .B(_01499_),
    .C(_01501_),
    .Y(_01502_));
 sg13g2_nor2_1 _06708_ (.A(_01497_),
    .B(_01502_),
    .Y(_01503_));
 sg13g2_o21ai_1 _06709_ (.B1(_01503_),
    .Y(_01504_),
    .A1(net1404),
    .A2(_01495_));
 sg13g2_a21oi_2 _06710_ (.B1(_01196_),
    .Y(_01505_),
    .A2(_01497_),
    .A1(\i_core.cpu.i_core.load_top_bit ));
 sg13g2_nor2b_1 _06711_ (.A(_01195_),
    .B_N(_01505_),
    .Y(_01506_));
 sg13g2_a221oi_1 _06712_ (.B2(_01506_),
    .C1(_01427_),
    .B1(_01504_),
    .A1(_01197_),
    .Y(\debug_rd[0] ),
    .A2(_01273_));
 sg13g2_nand2_2 _06713_ (.Y(_01507_),
    .A(\i_core.cpu.i_core.i_registers.rd[1] ),
    .B(\i_core.cpu.i_core.i_registers.rd[0] ));
 sg13g2_nand4_1 _06714_ (.B(_01197_),
    .C(_01198_),
    .A(_01176_),
    .Y(_01508_),
    .D(_01232_));
 sg13g2_nand3_1 _06715_ (.B(_01163_),
    .C(_01195_),
    .A(_00085_),
    .Y(_01509_));
 sg13g2_nand2_2 _06716_ (.Y(_01510_),
    .A(_01508_),
    .B(_01509_));
 sg13g2_inv_1 _06717_ (.Y(_01511_),
    .A(_01510_));
 sg13g2_nand3_1 _06718_ (.B(\i_core.cpu.i_core.i_registers.rd[3] ),
    .C(_01511_),
    .A(\i_core.cpu.i_core.i_registers.rd[2] ),
    .Y(_01512_));
 sg13g2_nor2_2 _06719_ (.A(_01507_),
    .B(_01512_),
    .Y(_01513_));
 sg13g2_mux2_1 _06720_ (.A0(net2453),
    .A1(net1165),
    .S(_01513_),
    .X(_00050_));
 sg13g2_mux2_2 _06721_ (.A0(\i_uart_rx.uart_rts ),
    .A1(\gpio_out[1] ),
    .S(\gpio_out_sel[1] ),
    .X(uo_out[1]));
 sg13g2_mux2_1 _06722_ (.A0(\i_spi.spi_clk_out ),
    .A1(\debug_rd_r[3] ),
    .S(debug_register_data),
    .X(_01514_));
 sg13g2_mux2_2 _06723_ (.A0(_01514_),
    .A1(\gpio_out[5] ),
    .S(\gpio_out_sel[5] ),
    .X(uo_out[5]));
 sg13g2_nand3_1 _06724_ (.B(\i_core.cpu.instr_data_start[19] ),
    .C(_01223_),
    .A(\i_core.cpu.instr_data_start[20] ),
    .Y(_01515_));
 sg13g2_nand4_1 _06725_ (.B(net1423),
    .C(\i_core.cpu.instr_data_start[19] ),
    .A(\i_core.cpu.instr_data_start[21] ),
    .Y(_01516_),
    .D(_01223_));
 sg13g2_xor2_1 _06726_ (.B(_01515_),
    .A(\i_core.cpu.instr_data_start[21] ),
    .X(_01517_));
 sg13g2_a21o_1 _06727_ (.A2(_01221_),
    .A1(net1424),
    .B1(\i_core.cpu.instr_data_start[17] ),
    .X(_01518_));
 sg13g2_and2_1 _06728_ (.A(_01222_),
    .B(_01518_),
    .X(_01519_));
 sg13g2_or2_1 _06729_ (.X(_01520_),
    .B(_01519_),
    .A(net1416));
 sg13g2_a21oi_1 _06730_ (.A1(net1414),
    .A2(_01517_),
    .Y(_01521_),
    .B1(_01227_));
 sg13g2_xnor2_1 _06731_ (.Y(_01522_),
    .A(_00760_),
    .B(_01211_));
 sg13g2_nand2_1 _06732_ (.Y(_01523_),
    .A(net1364),
    .B(_01522_));
 sg13g2_xnor2_1 _06733_ (.Y(_01524_),
    .A(_00765_),
    .B(_01206_));
 sg13g2_nor2_1 _06734_ (.A(_00880_),
    .B(_01524_),
    .Y(_01525_));
 sg13g2_xor2_1 _06735_ (.B(\i_core.cpu.pc[1] ),
    .A(\i_core.cpu.instr_len[1] ),
    .X(_01526_));
 sg13g2_o21ai_1 _06736_ (.B1(net1381),
    .Y(_01527_),
    .A1(_00875_),
    .A2(_01526_));
 sg13g2_xnor2_1 _06737_ (.Y(_01528_),
    .A(\i_core.cpu.instr_data_start[9] ),
    .B(_01208_));
 sg13g2_nor2_1 _06738_ (.A(_00882_),
    .B(_01528_),
    .Y(_01529_));
 sg13g2_nor3_1 _06739_ (.A(_01525_),
    .B(_01527_),
    .C(_01529_),
    .Y(_01530_));
 sg13g2_a22oi_1 _06740_ (.Y(_01531_),
    .B1(_01523_),
    .B2(_01530_),
    .A2(_01521_),
    .A1(_01520_));
 sg13g2_nand2_1 _06741_ (.Y(_01532_),
    .A(\i_core.cpu.i_core.i_cycles.i_regbuf[4].A ),
    .B(net1308));
 sg13g2_o21ai_1 _06742_ (.B1(_01532_),
    .Y(_01533_),
    .A1(_00784_),
    .A2(net1308));
 sg13g2_nor3_1 _06743_ (.A(_00199_),
    .B(_01245_),
    .C(_01259_),
    .Y(_01534_));
 sg13g2_a221oi_1 _06744_ (.B2(_01260_),
    .C1(_01534_),
    .B1(_01533_),
    .A1(\i_core.cpu.i_core.cycle_count[1] ),
    .Y(_01535_),
    .A2(_01261_));
 sg13g2_a22oi_1 _06745_ (.Y(_01536_),
    .B1(_01256_),
    .B2(\i_core.cpu.i_core.mepc[1] ),
    .A2(_01243_),
    .A1(\i_core.cpu.i_core.mip[17] ));
 sg13g2_a22oi_1 _06746_ (.Y(_01537_),
    .B1(_01251_),
    .B2(\i_core.cpu.i_core.mie[17] ),
    .A2(_01247_),
    .A1(\i_core.cpu.i_core.mcause[1] ));
 sg13g2_nand3_1 _06747_ (.B(_01536_),
    .C(_01537_),
    .A(_01535_),
    .Y(_01538_));
 sg13g2_a22oi_1 _06748_ (.Y(_01539_),
    .B1(_01233_),
    .B2(_01538_),
    .A2(\i_core.cpu.is_lui ),
    .A1(net1390));
 sg13g2_o21ai_1 _06749_ (.B1(_01539_),
    .Y(_01540_),
    .A1(_01198_),
    .A2(_01531_));
 sg13g2_o21ai_1 _06750_ (.B1(_01540_),
    .Y(_01541_),
    .A1(_01071_),
    .A2(_01176_));
 sg13g2_o21ai_1 _06751_ (.B1(net1365),
    .Y(_01542_),
    .A1(_00833_),
    .A2(net1190));
 sg13g2_a21oi_1 _06752_ (.A1(\i_core.mem.qspi_data_buf[13] ),
    .A2(net1190),
    .Y(_01543_),
    .B1(_01542_));
 sg13g2_mux2_1 _06753_ (.A0(_00832_),
    .A1(_00833_),
    .S(net1411),
    .X(_01544_));
 sg13g2_mux4_1 _06754_ (.S0(_01431_),
    .A0(\i_core.cpu.instr_data_in[1] ),
    .A1(\i_core.cpu.instr_data_in[9] ),
    .A2(\i_core.cpu.instr_data_in[5] ),
    .A3(\i_core.cpu.instr_data_in[13] ),
    .S1(net1411),
    .X(_01545_));
 sg13g2_nor2_1 _06755_ (.A(net1408),
    .B(_01545_),
    .Y(_01546_));
 sg13g2_o21ai_1 _06756_ (.B1(net1357),
    .Y(_01547_),
    .A1(_00832_),
    .A2(net1190));
 sg13g2_a21oi_1 _06757_ (.A1(\i_core.mem.qspi_data_buf[9] ),
    .A2(net1190),
    .Y(_01548_),
    .B1(_01547_));
 sg13g2_or3_1 _06758_ (.A(_01543_),
    .B(_01546_),
    .C(_01548_),
    .X(_01549_));
 sg13g2_nand2_1 _06759_ (.Y(_01550_),
    .A(\i_spi.data[5] ),
    .B(net1236));
 sg13g2_a22oi_1 _06760_ (.Y(_01551_),
    .B1(_01480_),
    .B2(\gpio_out_sel[5] ),
    .A2(_01479_),
    .A1(net6));
 sg13g2_a22oi_1 _06761_ (.Y(_01552_),
    .B1(_01477_),
    .B2(uo_out[5]),
    .A2(net1235),
    .A1(\i_uart_rx.recieved_data[5] ));
 sg13g2_nand4_1 _06762_ (.B(_01550_),
    .C(_01551_),
    .A(net1415),
    .Y(_01553_),
    .D(_01552_));
 sg13g2_nor2_2 _06763_ (.A(_00780_),
    .B(\i_uart_rx.fsm_state[2] ),
    .Y(_01554_));
 sg13g2_and2_2 _06764_ (.A(\i_uart_rx.fsm_state[1] ),
    .B(\i_uart_rx.fsm_state[0] ),
    .X(_01555_));
 sg13g2_nand2_1 _06765_ (.Y(_01556_),
    .A(\i_uart_rx.fsm_state[1] ),
    .B(_01554_));
 sg13g2_and2_2 _06766_ (.A(_01554_),
    .B(_01555_),
    .X(_01557_));
 sg13g2_nand2_2 _06767_ (.Y(_01558_),
    .A(_01554_),
    .B(_01555_));
 sg13g2_a22oi_1 _06768_ (.Y(_01559_),
    .B1(_01557_),
    .B2(_01464_),
    .A2(uo_out[1]),
    .A1(_01477_));
 sg13g2_a22oi_1 _06769_ (.Y(_01560_),
    .B1(_01479_),
    .B2(net3),
    .A2(net1236),
    .A1(\i_spi.data[1] ));
 sg13g2_a22oi_1 _06770_ (.Y(_01561_),
    .B1(_01480_),
    .B2(\gpio_out_sel[1] ),
    .A2(net1235),
    .A1(\i_uart_rx.recieved_data[1] ));
 sg13g2_nand4_1 _06771_ (.B(_01559_),
    .C(_01560_),
    .A(net1378),
    .Y(_01562_),
    .D(_01561_));
 sg13g2_nand3_1 _06772_ (.B(_01553_),
    .C(_01562_),
    .A(_00787_),
    .Y(_01563_));
 sg13g2_a22oi_1 _06773_ (.Y(_01564_),
    .B1(_01563_),
    .B2(net1234),
    .A2(_01549_),
    .A1(net1335));
 sg13g2_nand2_1 _06774_ (.Y(_01565_),
    .A(net1377),
    .B(\i_core.mem.qspi_data_buf[25] ));
 sg13g2_a21oi_1 _06775_ (.A1(net1411),
    .A2(\i_core.mem.qspi_data_buf[29] ),
    .Y(_01566_),
    .B1(net1202));
 sg13g2_a221oi_1 _06776_ (.B2(_01566_),
    .C1(_01434_),
    .B1(_01565_),
    .A1(net1202),
    .Y(_01567_),
    .A2(_01544_));
 sg13g2_a22oi_1 _06777_ (.Y(_01568_),
    .B1(net1360),
    .B2(\i_core.mem.data_from_read[21] ),
    .A2(net1368),
    .A1(\i_core.mem.data_from_read[17] ));
 sg13g2_a21oi_1 _06778_ (.A1(net1335),
    .A2(_01568_),
    .Y(_01569_),
    .B1(net1234));
 sg13g2_nor3_1 _06779_ (.A(net1380),
    .B(_01567_),
    .C(_01569_),
    .Y(_01570_));
 sg13g2_nor2_1 _06780_ (.A(_01497_),
    .B(_01570_),
    .Y(_01571_));
 sg13g2_o21ai_1 _06781_ (.B1(_01571_),
    .Y(_01572_),
    .A1(net1404),
    .A2(_01564_));
 sg13g2_a221oi_1 _06782_ (.B2(_01505_),
    .C1(_01195_),
    .B1(_01572_),
    .A1(_01196_),
    .Y(_01573_),
    .A2(_01541_));
 sg13g2_xnor2_1 _06783_ (.Y(_01574_),
    .A(_01137_),
    .B(_01138_));
 sg13g2_nand2_1 _06784_ (.Y(_01575_),
    .A(net1374),
    .B(_01147_));
 sg13g2_a21oi_1 _06785_ (.A1(_01052_),
    .A2(_01074_),
    .Y(_01576_),
    .B1(_01279_));
 sg13g2_nand2_1 _06786_ (.Y(_01577_),
    .A(_01575_),
    .B(_01576_));
 sg13g2_o21ai_1 _06787_ (.B1(_01577_),
    .Y(_01578_),
    .A1(_01275_),
    .A2(_01574_));
 sg13g2_a21oi_1 _06788_ (.A1(_01147_),
    .A2(_01281_),
    .Y(_01579_),
    .B1(_01578_));
 sg13g2_nor2_1 _06789_ (.A(_01285_),
    .B(_01579_),
    .Y(_01580_));
 sg13g2_nor2b_2 _06790_ (.A(_00085_),
    .B_N(_01051_),
    .Y(_01581_));
 sg13g2_nand2_1 _06791_ (.Y(_01582_),
    .A(\i_core.cpu.i_core.i_shift.a[0] ),
    .B(net1217));
 sg13g2_nand2_1 _06792_ (.Y(_01583_),
    .A(\i_core.cpu.i_core.i_shift.a[1] ),
    .B(net1238));
 sg13g2_or2_1 _06793_ (.X(_01584_),
    .B(_01583_),
    .A(_00200_));
 sg13g2_xor2_1 _06794_ (.B(_01583_),
    .A(_00200_),
    .X(_01585_));
 sg13g2_nand2b_1 _06795_ (.Y(_01586_),
    .B(_01585_),
    .A_N(_01421_));
 sg13g2_xor2_1 _06796_ (.B(_01585_),
    .A(_01421_),
    .X(_01587_));
 sg13g2_or2_1 _06797_ (.X(_01588_),
    .B(_01587_),
    .A(_01582_));
 sg13g2_a21oi_1 _06798_ (.A1(_01582_),
    .A2(_01587_),
    .Y(_01589_),
    .B1(_01164_));
 sg13g2_a22oi_1 _06799_ (.Y(_01590_),
    .B1(_01588_),
    .B2(_01589_),
    .A2(_01580_),
    .A1(_01164_));
 sg13g2_nand2_1 _06800_ (.Y(_01591_),
    .A(net1439),
    .B(_01381_));
 sg13g2_a21oi_1 _06801_ (.A1(net1371),
    .A2(_01376_),
    .Y(_01592_),
    .B1(net1304));
 sg13g2_nand2_1 _06802_ (.Y(_01593_),
    .A(net1441),
    .B(_01390_));
 sg13g2_a21oi_1 _06803_ (.A1(_00829_),
    .A2(_01379_),
    .Y(_01594_),
    .B1(net1301));
 sg13g2_a221oi_1 _06804_ (.B2(_01594_),
    .C1(_01310_),
    .B1(_01593_),
    .A1(_01591_),
    .Y(_01595_),
    .A2(_01592_));
 sg13g2_nand2_1 _06805_ (.Y(_01596_),
    .A(net1373),
    .B(_01398_));
 sg13g2_a21oi_1 _06806_ (.A1(net1441),
    .A2(_01409_),
    .Y(_01597_),
    .B1(net1302));
 sg13g2_nand2_1 _06807_ (.Y(_01598_),
    .A(\i_core.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .B(_01399_));
 sg13g2_a21oi_1 _06808_ (.A1(net1369),
    .A2(_01396_),
    .Y(_01599_),
    .B1(net1304));
 sg13g2_a221oi_1 _06809_ (.B2(_01599_),
    .C1(_01311_),
    .B1(_01598_),
    .A1(_01596_),
    .Y(_01600_),
    .A2(_01597_));
 sg13g2_or3_1 _06810_ (.A(net1277),
    .B(_01595_),
    .C(_01600_),
    .X(_01601_));
 sg13g2_nand2_1 _06811_ (.Y(_01602_),
    .A(net1438),
    .B(_01388_));
 sg13g2_a21oi_1 _06812_ (.A1(net1369),
    .A2(_01391_),
    .Y(_01603_),
    .B1(net1304));
 sg13g2_nand2_1 _06813_ (.Y(_01604_),
    .A(net1369),
    .B(_01385_));
 sg13g2_a221oi_1 _06814_ (.B2(_01341_),
    .C1(_01310_),
    .B1(_01604_),
    .A1(_01602_),
    .Y(_01605_),
    .A2(_01603_));
 sg13g2_nor2_1 _06815_ (.A(net1371),
    .B(_01404_),
    .Y(_01606_));
 sg13g2_a21oi_1 _06816_ (.A1(net1372),
    .A2(_01408_),
    .Y(_01607_),
    .B1(_01606_));
 sg13g2_nand2_1 _06817_ (.Y(_01608_),
    .A(net1439),
    .B(_01374_));
 sg13g2_a21oi_1 _06818_ (.A1(net1371),
    .A2(_01405_),
    .Y(_01609_),
    .B1(net1301));
 sg13g2_a221oi_1 _06819_ (.B2(_01609_),
    .C1(_01311_),
    .B1(_01608_),
    .A1(net1302),
    .Y(_01610_),
    .A2(_01607_));
 sg13g2_nor2b_1 _06820_ (.A(_01610_),
    .B_N(_01327_),
    .Y(_01611_));
 sg13g2_nand2b_1 _06821_ (.Y(_01612_),
    .B(_01611_),
    .A_N(_01605_));
 sg13g2_nand3_1 _06822_ (.B(_01601_),
    .C(_01612_),
    .A(_01297_),
    .Y(_01613_));
 sg13g2_nand3_1 _06823_ (.B(_01298_),
    .C(_01613_),
    .A(net1375),
    .Y(_01614_));
 sg13g2_a21oi_1 _06824_ (.A1(net1441),
    .A2(_01322_),
    .Y(_01615_),
    .B1(net1302));
 sg13g2_o21ai_1 _06825_ (.B1(_01615_),
    .Y(_01616_),
    .A1(net1441),
    .A2(_01318_));
 sg13g2_mux4_1 _06826_ (.S0(net1395),
    .A0(_00195_),
    .A1(_00196_),
    .A2(_00193_),
    .A3(_00194_),
    .S1(net1442),
    .X(_01617_));
 sg13g2_and2_1 _06827_ (.A(net1370),
    .B(_01617_),
    .X(_01618_));
 sg13g2_a21oi_1 _06828_ (.A1(net1438),
    .A2(_01320_),
    .Y(_01619_),
    .B1(_01618_));
 sg13g2_and2_1 _06829_ (.A(net1371),
    .B(_01324_),
    .X(_01620_));
 sg13g2_a21oi_1 _06830_ (.A1(net1439),
    .A2(_01351_),
    .Y(_01621_),
    .B1(_01620_));
 sg13g2_nand2_1 _06831_ (.Y(_01622_),
    .A(net1371),
    .B(_01354_));
 sg13g2_a21oi_1 _06832_ (.A1(net1440),
    .A2(_01361_),
    .Y(_01623_),
    .B1(net1301));
 sg13g2_a21o_1 _06833_ (.A2(_01312_),
    .A1(net1373),
    .B1(net1304),
    .X(_01624_));
 sg13g2_a21oi_1 _06834_ (.A1(net1438),
    .A2(_01339_),
    .Y(_01625_),
    .B1(_01624_));
 sg13g2_o21ai_1 _06835_ (.B1(net1304),
    .Y(_01626_),
    .A1(net1370),
    .A2(_01344_));
 sg13g2_a21oi_1 _06836_ (.A1(net1369),
    .A2(_01333_),
    .Y(_01627_),
    .B1(_01626_));
 sg13g2_mux4_1 _06837_ (.S0(net1305),
    .A0(_01303_),
    .A1(_01313_),
    .A2(_01364_),
    .A3(_01306_),
    .S1(net1372),
    .X(_01628_));
 sg13g2_a21oi_1 _06838_ (.A1(net1303),
    .A2(_01619_),
    .Y(_01629_),
    .B1(_01311_));
 sg13g2_a221oi_1 _06839_ (.B2(_01616_),
    .C1(net1277),
    .B1(_01629_),
    .A1(_01311_),
    .Y(_01630_),
    .A2(_01628_));
 sg13g2_a221oi_1 _06840_ (.B2(_01623_),
    .C1(_01311_),
    .B1(_01622_),
    .A1(net1301),
    .Y(_01631_),
    .A2(_01621_));
 sg13g2_nor3_1 _06841_ (.A(_01310_),
    .B(_01625_),
    .C(_01627_),
    .Y(_01632_));
 sg13g2_nand2b_1 _06842_ (.Y(_01633_),
    .B(net1277),
    .A_N(_01632_));
 sg13g2_o21ai_1 _06843_ (.B1(_01297_),
    .Y(_01634_),
    .A1(_01631_),
    .A2(_01633_));
 sg13g2_o21ai_1 _06844_ (.B1(_01298_),
    .Y(_01635_),
    .A1(_01630_),
    .A2(_01634_));
 sg13g2_inv_1 _06845_ (.Y(_01636_),
    .A(_01635_));
 sg13g2_a21oi_1 _06846_ (.A1(\i_core.cpu.alu_op[2] ),
    .A2(_01636_),
    .Y(_01637_),
    .B1(_01372_));
 sg13g2_nand2_1 _06847_ (.Y(_01638_),
    .A(_01195_),
    .B(_01425_));
 sg13g2_a221oi_1 _06848_ (.B2(_01637_),
    .C1(_01638_),
    .B1(_01614_),
    .A1(_01372_),
    .Y(_01639_),
    .A2(_01590_));
 sg13g2_or2_1 _06849_ (.X(\debug_rd[1] ),
    .B(_01639_),
    .A(_01573_));
 sg13g2_mux2_1 _06850_ (.A0(net2197),
    .A1(net1131),
    .S(_01513_),
    .X(_00051_));
 sg13g2_mux2_1 _06851_ (.A0(\i_spi.spi_dc ),
    .A1(\debug_rd_r[0] ),
    .S(debug_register_data),
    .X(_01640_));
 sg13g2_mux2_2 _06852_ (.A0(_01640_),
    .A1(\gpio_out[2] ),
    .S(\gpio_out_sel[2] ),
    .X(uo_out[2]));
 sg13g2_mux2_2 _06853_ (.A0(debug_uart_txd),
    .A1(\gpio_out[6] ),
    .S(\gpio_out_sel[6] ),
    .X(uo_out[6]));
 sg13g2_o21ai_1 _06854_ (.B1(_01274_),
    .Y(_01641_),
    .A1(_01139_),
    .A2(_01140_));
 sg13g2_a21oi_1 _06855_ (.A1(_01139_),
    .A2(_01140_),
    .Y(_01642_),
    .B1(_01641_));
 sg13g2_nand2_1 _06856_ (.Y(_01643_),
    .A(net1374),
    .B(_01149_));
 sg13g2_a21oi_1 _06857_ (.A1(_01004_),
    .A2(_01031_),
    .Y(_01644_),
    .B1(_01279_));
 sg13g2_a221oi_1 _06858_ (.B2(_01644_),
    .C1(_01642_),
    .B1(_01643_),
    .A1(_01149_),
    .Y(_01645_),
    .A2(_01281_));
 sg13g2_nor2_1 _06859_ (.A(_01285_),
    .B(_01645_),
    .Y(_01646_));
 sg13g2_nand2_1 _06860_ (.Y(_01647_),
    .A(_01586_),
    .B(_01588_));
 sg13g2_nand2_1 _06861_ (.Y(_01648_),
    .A(\i_core.cpu.i_core.i_shift.a[1] ),
    .B(net1217));
 sg13g2_a21oi_2 _06862_ (.B1(_00785_),
    .Y(_01649_),
    .A2(_01002_),
    .A1(_01001_));
 sg13g2_nand2_2 _06863_ (.Y(_01650_),
    .A(\i_core.cpu.i_core.i_shift.a[2] ),
    .B(net1233));
 sg13g2_and4_1 _06864_ (.A(\i_core.cpu.i_core.i_shift.a[0] ),
    .B(\i_core.cpu.i_core.i_shift.a[2] ),
    .C(net1238),
    .D(net1233),
    .X(_01651_));
 sg13g2_a22oi_1 _06865_ (.Y(_01652_),
    .B1(net1233),
    .B2(\i_core.cpu.i_core.i_shift.a[0] ),
    .A2(net1238),
    .A1(\i_core.cpu.i_core.i_shift.a[2] ));
 sg13g2_nor2_1 _06866_ (.A(_01651_),
    .B(_01652_),
    .Y(_01653_));
 sg13g2_and2_1 _06867_ (.A(\i_core.cpu.i_core.multiplier.accum[2] ),
    .B(_01653_),
    .X(_01654_));
 sg13g2_nand2_1 _06868_ (.Y(_01655_),
    .A(\i_core.cpu.i_core.multiplier.accum[2] ),
    .B(_01653_));
 sg13g2_xnor2_1 _06869_ (.Y(_01656_),
    .A(\i_core.cpu.i_core.multiplier.accum[2] ),
    .B(_01653_));
 sg13g2_xor2_1 _06870_ (.B(_01656_),
    .A(_01584_),
    .X(_01657_));
 sg13g2_nand2b_1 _06871_ (.Y(_01658_),
    .B(_01657_),
    .A_N(_01648_));
 sg13g2_xnor2_1 _06872_ (.Y(_01659_),
    .A(_01648_),
    .B(_01657_));
 sg13g2_and2_1 _06873_ (.A(_01647_),
    .B(_01659_),
    .X(_01660_));
 sg13g2_nand2_1 _06874_ (.Y(_01661_),
    .A(_01647_),
    .B(_01659_));
 sg13g2_o21ai_1 _06875_ (.B1(_01163_),
    .Y(_01662_),
    .A1(_01647_),
    .A2(_01659_));
 sg13g2_o21ai_1 _06876_ (.B1(_01372_),
    .Y(_01663_),
    .A1(_01660_),
    .A2(_01662_));
 sg13g2_a21oi_1 _06877_ (.A1(_01164_),
    .A2(_01646_),
    .Y(_01664_),
    .B1(_01663_));
 sg13g2_nand3_1 _06878_ (.B(_01298_),
    .C(_01613_),
    .A(net1394),
    .Y(_01665_));
 sg13g2_nand2_1 _06879_ (.Y(_01666_),
    .A(_01371_),
    .B(_01665_));
 sg13g2_a21oi_1 _06880_ (.A1(net1375),
    .A2(_01636_),
    .Y(_01667_),
    .B1(_01666_));
 sg13g2_nor3_1 _06881_ (.A(_01638_),
    .B(_01664_),
    .C(_01667_),
    .Y(_01668_));
 sg13g2_xnor2_1 _06882_ (.Y(_01669_),
    .A(net1426),
    .B(_01220_));
 sg13g2_inv_1 _06883_ (.Y(_01670_),
    .A(_01669_));
 sg13g2_xnor2_1 _06884_ (.Y(_01671_),
    .A(\i_core.cpu.instr_data_start[10] ),
    .B(_01209_));
 sg13g2_a21oi_1 _06885_ (.A1(\i_core.cpu.instr_data_start[5] ),
    .A2(_01206_),
    .Y(_01672_),
    .B1(\i_core.cpu.instr_data_start[6] ));
 sg13g2_or2_1 _06886_ (.X(_01673_),
    .B(_01672_),
    .A(_01207_));
 sg13g2_nor2_1 _06887_ (.A(_00880_),
    .B(_01673_),
    .Y(_01674_));
 sg13g2_xnor2_1 _06888_ (.Y(_01675_),
    .A(_01202_),
    .B(_01203_));
 sg13g2_a21oi_1 _06889_ (.A1(net1366),
    .A2(_01675_),
    .Y(_01676_),
    .B1(_01674_));
 sg13g2_o21ai_1 _06890_ (.B1(_01676_),
    .Y(_01677_),
    .A1(_00882_),
    .A2(_01671_));
 sg13g2_a21oi_1 _06891_ (.A1(net1363),
    .A2(_01670_),
    .Y(_01678_),
    .B1(_01677_));
 sg13g2_nor2_1 _06892_ (.A(_00756_),
    .B(_01516_),
    .Y(_01679_));
 sg13g2_xnor2_1 _06893_ (.Y(_01680_),
    .A(_00756_),
    .B(_01516_));
 sg13g2_xnor2_1 _06894_ (.Y(_01681_),
    .A(_00758_),
    .B(_01222_));
 sg13g2_inv_1 _06895_ (.Y(_01682_),
    .A(_01681_));
 sg13g2_a21oi_1 _06896_ (.A1(net1415),
    .A2(_01680_),
    .Y(_01683_),
    .B1(_01227_));
 sg13g2_o21ai_1 _06897_ (.B1(_01683_),
    .Y(_01684_),
    .A1(net1415),
    .A2(_01682_));
 sg13g2_o21ai_1 _06898_ (.B1(_01684_),
    .Y(_01685_),
    .A1(net1406),
    .A2(_01678_));
 sg13g2_nand3_1 _06899_ (.B(_01244_),
    .C(_01250_),
    .A(_01240_),
    .Y(_01686_));
 sg13g2_inv_1 _06900_ (.Y(_01687_),
    .A(_01686_));
 sg13g2_and2_2 _06901_ (.A(net2440),
    .B(net1278),
    .X(_01688_));
 sg13g2_a21oi_1 _06902_ (.A1(net1416),
    .A2(net1354),
    .Y(_01689_),
    .B1(net1278));
 sg13g2_nor2_1 _06903_ (.A(_01266_),
    .B(_01689_),
    .Y(_01690_));
 sg13g2_a221oi_1 _06904_ (.B2(_01688_),
    .C1(_01690_),
    .B1(_01687_),
    .A1(\i_core.cpu.i_core.i_instrret.data[2] ),
    .Y(_01691_),
    .A2(_01262_));
 sg13g2_a22oi_1 _06905_ (.Y(_01692_),
    .B1(_01256_),
    .B2(\i_core.cpu.i_core.mepc[2] ),
    .A2(_01251_),
    .A1(\i_core.cpu.i_core.mie[18] ));
 sg13g2_mux2_1 _06906_ (.A0(\i_core.cpu.i_core.time_hi[1] ),
    .A1(\i_core.cpu.i_core.i_cycles.i_regbuf[5].A ),
    .S(net1308),
    .X(_01693_));
 sg13g2_nand2_1 _06907_ (.Y(_01694_),
    .A(_01260_),
    .B(_01693_));
 sg13g2_a22oi_1 _06908_ (.Y(_01695_),
    .B1(_01557_),
    .B2(_01243_),
    .A2(_01261_),
    .A1(\i_core.cpu.i_core.cycle_count[2] ));
 sg13g2_nand4_1 _06909_ (.B(_01692_),
    .C(_01694_),
    .A(_01691_),
    .Y(_01696_),
    .D(_01695_));
 sg13g2_a22oi_1 _06910_ (.Y(_01697_),
    .B1(_01696_),
    .B2(_01233_),
    .A2(_01685_),
    .A1(_01199_));
 sg13g2_mux2_1 _06911_ (.A0(_01013_),
    .A1(_01697_),
    .S(_01176_),
    .X(_01698_));
 sg13g2_a21o_1 _06912_ (.A2(_01432_),
    .A1(\i_core.cpu.instr_data_in[10] ),
    .B1(_00882_),
    .X(_01699_));
 sg13g2_a21oi_1 _06913_ (.A1(\i_core.mem.qspi_data_buf[10] ),
    .A2(_01433_),
    .Y(_01700_),
    .B1(_01699_));
 sg13g2_o21ai_1 _06914_ (.B1(net1365),
    .Y(_01701_),
    .A1(_00835_),
    .A2(net1190));
 sg13g2_a21oi_1 _06915_ (.A1(\i_core.mem.qspi_data_buf[14] ),
    .A2(net1190),
    .Y(_01702_),
    .B1(_01701_));
 sg13g2_or2_1 _06916_ (.X(_01703_),
    .B(\i_core.cpu.instr_data_in[10] ),
    .A(net1412));
 sg13g2_o21ai_1 _06917_ (.B1(_01703_),
    .Y(_01704_),
    .A1(net1377),
    .A2(\i_core.cpu.instr_data_in[14] ));
 sg13g2_mux4_1 _06918_ (.S0(_01431_),
    .A0(\i_core.cpu.instr_data_in[2] ),
    .A1(\i_core.cpu.instr_data_in[10] ),
    .A2(\i_core.cpu.instr_data_in[6] ),
    .A3(\i_core.cpu.instr_data_in[14] ),
    .S1(net1411),
    .X(_01705_));
 sg13g2_nor2_1 _06919_ (.A(net1408),
    .B(_01705_),
    .Y(_01706_));
 sg13g2_or3_1 _06920_ (.A(_01700_),
    .B(_01702_),
    .C(_01706_),
    .X(_01707_));
 sg13g2_nand2_1 _06921_ (.Y(_01708_),
    .A(\i_spi.data[2] ),
    .B(_01458_));
 sg13g2_a22oi_1 _06922_ (.Y(_01709_),
    .B1(uo_out[2]),
    .B2(_01477_),
    .A2(_01479_),
    .A1(net4));
 sg13g2_a22oi_1 _06923_ (.Y(_01710_),
    .B1(_01480_),
    .B2(\gpio_out_sel[2] ),
    .A2(net1235),
    .A1(\i_uart_rx.recieved_data[2] ));
 sg13g2_nand4_1 _06924_ (.B(_01708_),
    .C(_01709_),
    .A(net1378),
    .Y(_01711_),
    .D(_01710_));
 sg13g2_nand2_1 _06925_ (.Y(_01712_),
    .A(_01477_),
    .B(uo_out[6]));
 sg13g2_a22oi_1 _06926_ (.Y(_01713_),
    .B1(_01480_),
    .B2(\gpio_out_sel[6] ),
    .A2(_01479_),
    .A1(net7));
 sg13g2_a22oi_1 _06927_ (.Y(_01714_),
    .B1(net1235),
    .B2(\i_uart_rx.recieved_data[6] ),
    .A2(net1236),
    .A1(\i_spi.data[6] ));
 sg13g2_nand4_1 _06928_ (.B(_01712_),
    .C(_01713_),
    .A(net1415),
    .Y(_01715_),
    .D(_01714_));
 sg13g2_nand3_1 _06929_ (.B(_01711_),
    .C(_01715_),
    .A(_00787_),
    .Y(_01716_));
 sg13g2_a22oi_1 _06930_ (.Y(_01717_),
    .B1(_01716_),
    .B2(net1234),
    .A2(_01707_),
    .A1(net1335));
 sg13g2_nand2_1 _06931_ (.Y(_01718_),
    .A(net1377),
    .B(\i_core.mem.qspi_data_buf[26] ));
 sg13g2_a21oi_1 _06932_ (.A1(net1411),
    .A2(\i_core.mem.qspi_data_buf[30] ),
    .Y(_01719_),
    .B1(net1202));
 sg13g2_a221oi_1 _06933_ (.B2(_01719_),
    .C1(_01434_),
    .B1(_01718_),
    .A1(net1202),
    .Y(_01720_),
    .A2(_01704_));
 sg13g2_a22oi_1 _06934_ (.Y(_01721_),
    .B1(net1360),
    .B2(\i_core.mem.data_from_read[22] ),
    .A2(net1368),
    .A1(\i_core.mem.data_from_read[18] ));
 sg13g2_a21oi_1 _06935_ (.A1(net1335),
    .A2(_01721_),
    .Y(_01722_),
    .B1(net1234));
 sg13g2_nor3_1 _06936_ (.A(net1380),
    .B(_01720_),
    .C(_01722_),
    .Y(_01723_));
 sg13g2_nor2_1 _06937_ (.A(_01497_),
    .B(_01723_),
    .Y(_01724_));
 sg13g2_o21ai_1 _06938_ (.B1(_01724_),
    .Y(_01725_),
    .A1(net1404),
    .A2(_01717_));
 sg13g2_a221oi_1 _06939_ (.B2(_01505_),
    .C1(_01195_),
    .B1(_01725_),
    .A1(_01196_),
    .Y(_01726_),
    .A2(_01698_));
 sg13g2_or2_1 _06940_ (.X(\debug_rd[2] ),
    .B(_01726_),
    .A(_01668_));
 sg13g2_mux2_1 _06941_ (.A0(net2041),
    .A1(net1126),
    .S(_01513_),
    .X(_00052_));
 sg13g2_mux2_1 _06942_ (.A0(\i_spi.data[7] ),
    .A1(\debug_rd_r[1] ),
    .S(debug_register_data),
    .X(_01727_));
 sg13g2_mux2_2 _06943_ (.A0(_01727_),
    .A1(\gpio_out[3] ),
    .S(\gpio_out_sel[3] ),
    .X(uo_out[3]));
 sg13g2_nand2_1 _06944_ (.Y(_01728_),
    .A(\gpio_out_sel[7] ),
    .B(_00839_));
 sg13g2_or3_1 _06945_ (.A(\i_core.cpu.i_core.mem_op[0] ),
    .B(_01145_),
    .C(_01155_),
    .X(_01729_));
 sg13g2_o21ai_1 _06946_ (.B1(\i_core.cpu.i_core.mem_op[0] ),
    .Y(_01730_),
    .A1(_01145_),
    .A2(_01155_));
 sg13g2_nand3_1 _06947_ (.B(_01729_),
    .C(_01730_),
    .A(net1348),
    .Y(_01731_));
 sg13g2_nor3_1 _06948_ (.A(_01178_),
    .B(_01236_),
    .C(_01275_),
    .Y(_01732_));
 sg13g2_nand4_1 _06949_ (.B(\i_core.cpu.i_core.imm_lo[9] ),
    .C(_01177_),
    .A(\i_core.cpu.i_core.imm_lo[8] ),
    .Y(_01733_),
    .D(_01274_));
 sg13g2_nand3_1 _06950_ (.B(_01258_),
    .C(_01274_),
    .A(_01177_),
    .Y(_01734_));
 sg13g2_and2_2 _06951_ (.A(net2424),
    .B(_01734_),
    .X(_01735_));
 sg13g2_nand2_2 _06952_ (.Y(_01736_),
    .A(_00086_),
    .B(_01734_));
 sg13g2_nor3_1 _06953_ (.A(_01199_),
    .B(net1276),
    .C(_01736_),
    .Y(_01737_));
 sg13g2_a21oi_1 _06954_ (.A1(_01731_),
    .A2(_01737_),
    .Y(_01738_),
    .B1(net1309));
 sg13g2_a21o_1 _06955_ (.A2(_01737_),
    .A1(_01731_),
    .B1(net1309),
    .X(_01739_));
 sg13g2_nor2_1 _06956_ (.A(net1393),
    .B(_00098_),
    .Y(_01740_));
 sg13g2_a21oi_2 _06957_ (.B1(_01740_),
    .Y(_01741_),
    .A2(_01675_),
    .A1(net1393));
 sg13g2_a21o_1 _06958_ (.A2(_01675_),
    .A1(net1393),
    .B1(_01740_),
    .X(_01742_));
 sg13g2_nor2_1 _06959_ (.A(net1393),
    .B(_00097_),
    .Y(_01743_));
 sg13g2_a21o_2 _06960_ (.A2(_01526_),
    .A1(net1393),
    .B1(_01743_),
    .X(_01744_));
 sg13g2_a21oi_1 _06961_ (.A1(net1393),
    .A2(_01526_),
    .Y(_01745_),
    .B1(_01743_));
 sg13g2_mux4_1 _06962_ (.S0(net1289),
    .A0(\i_core.cpu.instr_data[1][0] ),
    .A1(\i_core.cpu.instr_data[0][0] ),
    .A2(\i_core.cpu.instr_data[3][0] ),
    .A3(\i_core.cpu.instr_data[2][0] ),
    .S1(net1270),
    .X(_01746_));
 sg13g2_a21o_1 _06963_ (.A2(net1272),
    .A1(_00101_),
    .B1(net1294),
    .X(_01747_));
 sg13g2_a21oi_1 _06964_ (.A1(_00099_),
    .A2(_01741_),
    .Y(_01748_),
    .B1(_01747_));
 sg13g2_a21oi_1 _06965_ (.A1(_00100_),
    .A2(_01741_),
    .Y(_01749_),
    .B1(net1290));
 sg13g2_o21ai_1 _06966_ (.B1(_01749_),
    .Y(_01750_),
    .A1(_00810_),
    .A2(_01741_));
 sg13g2_nand2b_1 _06967_ (.Y(_01751_),
    .B(_01750_),
    .A_N(_01748_));
 sg13g2_nor2b_2 _06968_ (.A(_01748_),
    .B_N(_01750_),
    .Y(_01752_));
 sg13g2_and2_1 _06969_ (.A(_01746_),
    .B(net1215),
    .X(_01753_));
 sg13g2_nand2_1 _06970_ (.Y(_01754_),
    .A(_01746_),
    .B(net1215));
 sg13g2_xnor2_1 _06971_ (.Y(_01755_),
    .A(\i_core.cpu.instr_write_offset[1] ),
    .B(net1291));
 sg13g2_and2_1 _06972_ (.A(_00087_),
    .B(_01744_),
    .X(_01756_));
 sg13g2_nor2b_1 _06973_ (.A(_00096_),
    .B_N(_01204_),
    .Y(_01757_));
 sg13g2_xnor2_1 _06974_ (.Y(_01758_),
    .A(\i_core.cpu.instr_write_offset[3] ),
    .B(_01757_));
 sg13g2_a22oi_1 _06975_ (.Y(_01759_),
    .B1(_01756_),
    .B2(_01758_),
    .A2(net1273),
    .A1(_00793_));
 sg13g2_o21ai_1 _06976_ (.B1(_01758_),
    .Y(_01760_),
    .A1(_00793_),
    .A2(net1273));
 sg13g2_a21oi_1 _06977_ (.A1(_01756_),
    .A2(_01760_),
    .Y(_01761_),
    .B1(_01759_));
 sg13g2_a221oi_1 _06978_ (.B2(_01760_),
    .C1(_01761_),
    .B1(_01759_),
    .A1(net1199),
    .Y(_01762_),
    .A2(_01755_));
 sg13g2_nand2_1 _06979_ (.Y(_01763_),
    .A(\i_core.cpu.i_core.mie[16] ),
    .B(\i_core.cpu.i_core.mip[16] ));
 sg13g2_o21ai_1 _06980_ (.B1(_01763_),
    .Y(_01764_),
    .A1(_00771_),
    .A2(_00774_));
 sg13g2_nand2_1 _06981_ (.Y(_01765_),
    .A(net2168),
    .B(_01461_));
 sg13g2_o21ai_1 _06982_ (.B1(_01765_),
    .Y(_01766_),
    .A1(_00772_),
    .A2(_01558_));
 sg13g2_o21ai_1 _06983_ (.B1(\i_core.cpu.i_core.mstatus_mie ),
    .Y(_01767_),
    .A1(_01764_),
    .A2(_01766_));
 sg13g2_inv_1 _06984_ (.Y(_01768_),
    .A(_01767_));
 sg13g2_nor2_2 _06985_ (.A(_01183_),
    .B(_01767_),
    .Y(_01769_));
 sg13g2_inv_1 _06986_ (.Y(_01770_),
    .A(_01769_));
 sg13g2_nor3_2 _06987_ (.A(_00807_),
    .B(_01762_),
    .C(_01769_),
    .Y(_01771_));
 sg13g2_nor3_2 _06988_ (.A(net2200),
    .B(net2320),
    .C(\i_core.cpu.additional_mem_ops[0] ),
    .Y(_01772_));
 sg13g2_nand2b_2 _06989_ (.Y(_01773_),
    .B(_01772_),
    .A_N(_01184_));
 sg13g2_o21ai_1 _06990_ (.B1(net1189),
    .Y(_01774_),
    .A1(net1392),
    .A2(net1309));
 sg13g2_nor2_1 _06991_ (.A(_01184_),
    .B(_01772_),
    .Y(_01775_));
 sg13g2_or2_1 _06992_ (.X(_01776_),
    .B(_01772_),
    .A(_01184_));
 sg13g2_and4_1 _06993_ (.A(net1465),
    .B(_01771_),
    .C(_01774_),
    .D(_01776_),
    .X(_01777_));
 sg13g2_and2_2 _06994_ (.A(_01746_),
    .B(_01752_),
    .X(_01778_));
 sg13g2_mux4_1 _06995_ (.S0(net1290),
    .A0(_00116_),
    .A1(_00115_),
    .A2(_00118_),
    .A3(_00117_),
    .S1(net1271),
    .X(_01779_));
 sg13g2_inv_4 _06996_ (.A(_01779_),
    .Y(_01780_));
 sg13g2_mux4_1 _06997_ (.S0(net1291),
    .A0(_00120_),
    .A1(_00119_),
    .A2(_00122_),
    .A3(_00121_),
    .S1(net1273),
    .X(_01781_));
 sg13g2_inv_4 _06998_ (.A(net1257),
    .Y(_01782_));
 sg13g2_nor2_2 _06999_ (.A(_01779_),
    .B(_01782_),
    .Y(_01783_));
 sg13g2_nand2_1 _07000_ (.Y(_01784_),
    .A(_01778_),
    .B(net1257));
 sg13g2_nor2_2 _07001_ (.A(_01779_),
    .B(_01784_),
    .Y(_01785_));
 sg13g2_nand2_2 _07002_ (.Y(_01786_),
    .A(_01778_),
    .B(_01783_));
 sg13g2_mux4_1 _07003_ (.S0(net1291),
    .A0(_00108_),
    .A1(_00107_),
    .A2(_00110_),
    .A3(_00109_),
    .S1(net1273),
    .X(_01787_));
 sg13g2_mux4_1 _07004_ (.S0(net1289),
    .A0(_00112_),
    .A1(_00111_),
    .A2(_00114_),
    .A3(_00113_),
    .S1(net1268),
    .X(_01788_));
 sg13g2_nor2_1 _07005_ (.A(net1255),
    .B(net1253),
    .Y(_01789_));
 sg13g2_mux4_1 _07006_ (.S0(net1290),
    .A0(_00104_),
    .A1(_00103_),
    .A2(_00106_),
    .A3(_00105_),
    .S1(net1272),
    .X(_01790_));
 sg13g2_inv_2 _07007_ (.Y(_01791_),
    .A(_01790_));
 sg13g2_mux4_1 _07008_ (.S0(net1290),
    .A0(\i_core.cpu.instr_data[1][2] ),
    .A1(\i_core.cpu.instr_data[0][2] ),
    .A2(\i_core.cpu.instr_data[3][2] ),
    .A3(\i_core.cpu.instr_data[2][2] ),
    .S1(net1271),
    .X(_01792_));
 sg13g2_inv_1 _07009_ (.Y(_01793_),
    .A(net1252));
 sg13g2_nand3_1 _07010_ (.B(_01790_),
    .C(net1252),
    .A(_01789_),
    .Y(_01794_));
 sg13g2_mux4_1 _07011_ (.S0(net1289),
    .A0(\i_core.cpu.instr_data[1][3] ),
    .A1(\i_core.cpu.instr_data[0][3] ),
    .A2(\i_core.cpu.instr_data[3][3] ),
    .A3(\i_core.cpu.instr_data[2][3] ),
    .S1(net1269),
    .X(_01795_));
 sg13g2_nor2b_2 _07012_ (.A(_01794_),
    .B_N(net1250),
    .Y(_01796_));
 sg13g2_nand2b_2 _07013_ (.Y(_01797_),
    .B(net1250),
    .A_N(_01794_));
 sg13g2_o21ai_1 _07014_ (.B1(_01786_),
    .Y(_01798_),
    .A1(net1197),
    .A2(_01797_));
 sg13g2_nand3_1 _07015_ (.B(_01777_),
    .C(_01798_),
    .A(net1176),
    .Y(_01799_));
 sg13g2_nor2_1 _07016_ (.A(_01780_),
    .B(_01782_),
    .Y(_01800_));
 sg13g2_nand2_2 _07017_ (.Y(_01801_),
    .A(_01779_),
    .B(net1257));
 sg13g2_mux4_1 _07018_ (.S0(net1289),
    .A0(_00124_),
    .A1(_00123_),
    .A2(_00126_),
    .A3(_00125_),
    .S1(net1269),
    .X(_01802_));
 sg13g2_or2_2 _07019_ (.X(_01803_),
    .B(_01802_),
    .A(_01746_));
 sg13g2_nor2_2 _07020_ (.A(_01752_),
    .B(_01803_),
    .Y(_01804_));
 sg13g2_nor3_2 _07021_ (.A(_01752_),
    .B(_01801_),
    .C(_01803_),
    .Y(_01805_));
 sg13g2_nand2_1 _07022_ (.Y(_01806_),
    .A(_01800_),
    .B(_01804_));
 sg13g2_or3_2 _07023_ (.A(_01791_),
    .B(net1252),
    .C(net1250),
    .X(_01807_));
 sg13g2_inv_1 _07024_ (.Y(_01808_),
    .A(_01807_));
 sg13g2_nand2_1 _07025_ (.Y(_01809_),
    .A(net1256),
    .B(net1253));
 sg13g2_nor2_2 _07026_ (.A(_01807_),
    .B(_01809_),
    .Y(_01810_));
 sg13g2_and2_1 _07027_ (.A(_01805_),
    .B(_01810_),
    .X(_01811_));
 sg13g2_nand2_2 _07028_ (.Y(_01812_),
    .A(_01805_),
    .B(_01810_));
 sg13g2_a21o_1 _07029_ (.A2(net1271),
    .A1(_00142_),
    .B1(net1290),
    .X(_01813_));
 sg13g2_a21oi_1 _07030_ (.A1(_00140_),
    .A2(_01741_),
    .Y(_01814_),
    .B1(_01813_));
 sg13g2_a21oi_1 _07031_ (.A1(_00141_),
    .A2(net1271),
    .Y(_01815_),
    .B1(net1294));
 sg13g2_o21ai_1 _07032_ (.B1(_01815_),
    .Y(_01816_),
    .A1(_00811_),
    .A2(net1271));
 sg13g2_nor2b_2 _07033_ (.A(_01814_),
    .B_N(_01816_),
    .Y(_01817_));
 sg13g2_nand2b_2 _07034_ (.Y(_01818_),
    .B(_01816_),
    .A_N(_01814_));
 sg13g2_mux4_1 _07035_ (.S0(net1289),
    .A0(_00136_),
    .A1(_00135_),
    .A2(_00138_),
    .A3(_00137_),
    .S1(net1268),
    .X(_01819_));
 sg13g2_nand2_1 _07036_ (.Y(_01820_),
    .A(_01817_),
    .B(_01819_));
 sg13g2_mux4_1 _07037_ (.S0(net1289),
    .A0(_00132_),
    .A1(_00131_),
    .A2(_00134_),
    .A3(_00133_),
    .S1(net1268),
    .X(_01821_));
 sg13g2_inv_1 _07038_ (.Y(_01822_),
    .A(_01821_));
 sg13g2_a21o_1 _07039_ (.A2(net1272),
    .A1(_00146_),
    .B1(net1290),
    .X(_01823_));
 sg13g2_a21oi_1 _07040_ (.A1(_00144_),
    .A2(_01741_),
    .Y(_01824_),
    .B1(_01823_));
 sg13g2_a21oi_1 _07041_ (.A1(_00145_),
    .A2(net1272),
    .Y(_01825_),
    .B1(net1294));
 sg13g2_o21ai_1 _07042_ (.B1(_01825_),
    .Y(_01826_),
    .A1(_00812_),
    .A2(net1272));
 sg13g2_nor2b_1 _07043_ (.A(_01824_),
    .B_N(_01826_),
    .Y(_01827_));
 sg13g2_nand2b_2 _07044_ (.Y(_01828_),
    .B(_01826_),
    .A_N(_01824_));
 sg13g2_mux4_1 _07045_ (.S0(net1289),
    .A0(_00128_),
    .A1(_00127_),
    .A2(_00130_),
    .A3(_00129_),
    .S1(net1270),
    .X(_01829_));
 sg13g2_nand2_1 _07046_ (.Y(_01830_),
    .A(net1249),
    .B(net1213));
 sg13g2_nor4_2 _07047_ (.A(_01812_),
    .B(_01820_),
    .C(_01829_),
    .Y(_01831_),
    .D(_01830_));
 sg13g2_and3_1 _07048_ (.X(_01832_),
    .A(net1176),
    .B(_01777_),
    .C(_01831_));
 sg13g2_nand3_1 _07049_ (.B(_01777_),
    .C(_01831_),
    .A(net1176),
    .Y(_01833_));
 sg13g2_nand2_1 _07050_ (.Y(_01834_),
    .A(_00090_),
    .B(net1179));
 sg13g2_and4_1 _07051_ (.A(_00088_),
    .B(_01799_),
    .C(net1171),
    .D(_01834_),
    .X(_01835_));
 sg13g2_nand2b_1 _07052_ (.Y(_01836_),
    .B(_01204_),
    .A_N(net1189));
 sg13g2_nor2b_1 _07053_ (.A(\i_core.mem.qspi_data_byte_idx[1] ),
    .B_N(\i_core.mem.qspi_data_byte_idx[0] ),
    .Y(_01837_));
 sg13g2_nand2_1 _07054_ (.Y(_01838_),
    .A(\i_core.mem.q_ctrl.data_ready ),
    .B(_01837_));
 sg13g2_inv_1 _07055_ (.Y(_01839_),
    .A(net1288));
 sg13g2_nor3_2 _07056_ (.A(_00770_),
    .B(_00088_),
    .C(net1288),
    .Y(_01840_));
 sg13g2_nor2b_1 _07057_ (.A(_00087_),
    .B_N(_01840_),
    .Y(_01841_));
 sg13g2_nand2_1 _07058_ (.Y(_01842_),
    .A(\i_core.cpu.instr_write_offset[2] ),
    .B(_01841_));
 sg13g2_xor2_1 _07059_ (.B(_01842_),
    .A(\i_core.cpu.instr_write_offset[3] ),
    .X(_01843_));
 sg13g2_xnor2_1 _07060_ (.Y(_01844_),
    .A(_01836_),
    .B(_01843_));
 sg13g2_xnor2_1 _07061_ (.Y(_01845_),
    .A(\i_core.cpu.instr_write_offset[2] ),
    .B(_01841_));
 sg13g2_xnor2_1 _07062_ (.Y(_01846_),
    .A(net2642),
    .B(_01840_));
 sg13g2_xnor2_1 _07063_ (.Y(_01847_),
    .A(_00097_),
    .B(_01846_));
 sg13g2_xor2_1 _07064_ (.B(_01845_),
    .A(_00098_),
    .X(_01848_));
 sg13g2_nor3_2 _07065_ (.A(_01844_),
    .B(_01847_),
    .C(_01848_),
    .Y(_01849_));
 sg13g2_nand4_1 _07066_ (.B(_00794_),
    .C(_01837_),
    .A(\i_core.mem.instr_active ),
    .Y(_01850_),
    .D(_01849_));
 sg13g2_nand2_1 _07067_ (.Y(_01851_),
    .A(\i_core.cpu.instr_fetch_started ),
    .B(_01850_));
 sg13g2_nand2_1 _07068_ (.Y(_01852_),
    .A(_01835_),
    .B(_01851_));
 sg13g2_a21o_1 _07069_ (.A2(\i_core.cpu.data_read_n[0] ),
    .A1(\i_core.cpu.data_read_n[1] ),
    .B1(_01186_),
    .X(_01853_));
 sg13g2_nand2_2 _07070_ (.Y(_01854_),
    .A(\i_core.cpu.data_write_n[1] ),
    .B(\i_core.cpu.data_write_n[0] ));
 sg13g2_nand2_2 _07071_ (.Y(_01855_),
    .A(_01185_),
    .B(_01854_));
 sg13g2_nand2_1 _07072_ (.Y(_01856_),
    .A(_01853_),
    .B(_01855_));
 sg13g2_o21ai_1 _07073_ (.B1(_01856_),
    .Y(_01857_),
    .A1(_01839_),
    .A2(_01849_));
 sg13g2_and2_1 _07074_ (.A(\i_core.mem.instr_active ),
    .B(_01857_),
    .X(_01858_));
 sg13g2_nor2_2 _07075_ (.A(net1431),
    .B(\i_core.mem.q_ctrl.fsm_state[0] ),
    .Y(_01859_));
 sg13g2_and2_2 _07076_ (.A(net1429),
    .B(_01859_),
    .X(_01860_));
 sg13g2_nand2_2 _07077_ (.Y(_01861_),
    .A(net1429),
    .B(_01859_));
 sg13g2_nor2_2 _07078_ (.A(\i_core.mem.q_ctrl.data_ready ),
    .B(\i_core.mem.q_ctrl.data_req ),
    .Y(_01862_));
 sg13g2_nor2_1 _07079_ (.A(debug_data_continue),
    .B(_01862_),
    .Y(_01863_));
 sg13g2_a21oi_1 _07080_ (.A1(_01192_),
    .A2(_01863_),
    .Y(_01864_),
    .B1(net2677));
 sg13g2_a221oi_1 _07081_ (.B2(net2501),
    .C1(_01864_),
    .B1(_01860_),
    .A1(_01852_),
    .Y(_01865_),
    .A2(_01858_));
 sg13g2_a21oi_1 _07082_ (.A1(net1469),
    .A2(_01850_),
    .Y(_01866_),
    .B1(net1468));
 sg13g2_o21ai_1 _07083_ (.B1(_01866_),
    .Y(_01867_),
    .A1(net1469),
    .A2(_01865_));
 sg13g2_o21ai_1 _07084_ (.B1(net1468),
    .Y(_01868_),
    .A1(debug_data_continue),
    .A2(net1470));
 sg13g2_a21oi_1 _07085_ (.A1(net1469),
    .A2(net1312),
    .Y(_01869_),
    .B1(_01868_));
 sg13g2_nor2_1 _07086_ (.A(net6),
    .B(_01869_),
    .Y(_01870_));
 sg13g2_o21ai_1 _07087_ (.B1(net1468),
    .Y(_01871_),
    .A1(_00837_),
    .A2(net1179));
 sg13g2_a21oi_1 _07088_ (.A1(_00837_),
    .A2(_01799_),
    .Y(_01872_),
    .B1(_01871_));
 sg13g2_a21oi_1 _07089_ (.A1(_00837_),
    .A2(_01510_),
    .Y(_01873_),
    .B1(net1468));
 sg13g2_o21ai_1 _07090_ (.B1(_01873_),
    .Y(_01874_),
    .A1(_00837_),
    .A2(net1173));
 sg13g2_nor2_1 _07091_ (.A(_00834_),
    .B(_01872_),
    .Y(_01875_));
 sg13g2_a221oi_1 _07092_ (.B2(_01875_),
    .C1(net7),
    .B1(_01874_),
    .A1(_01867_),
    .Y(_01876_),
    .A2(_01870_));
 sg13g2_a21oi_1 _07093_ (.A1(_00747_),
    .A2(net1469),
    .Y(_01877_),
    .B1(net1468));
 sg13g2_o21ai_1 _07094_ (.B1(_01877_),
    .Y(_01878_),
    .A1(net1469),
    .A2(_01835_));
 sg13g2_a21oi_1 _07095_ (.A1(\i_core.mem.instr_active ),
    .A2(_01839_),
    .Y(_01879_),
    .B1(net1469));
 sg13g2_a21oi_1 _07096_ (.A1(net1469),
    .A2(net1188),
    .Y(_01880_),
    .B1(_01879_));
 sg13g2_a21oi_1 _07097_ (.A1(net1468),
    .A2(_01880_),
    .Y(_01881_),
    .B1(_00834_));
 sg13g2_nand2_2 _07098_ (.Y(_01882_),
    .A(_01185_),
    .B(_01430_));
 sg13g2_and2_2 _07099_ (.A(_01186_),
    .B(_01854_),
    .X(_01883_));
 sg13g2_nand2_1 _07100_ (.Y(_01884_),
    .A(_01186_),
    .B(_01854_));
 sg13g2_a21oi_2 _07101_ (.B1(net1335),
    .Y(_01885_),
    .A2(\i_core.cpu.data_read_n[0] ),
    .A1(\i_core.cpu.data_read_n[1] ));
 sg13g2_mux4_1 _07102_ (.S0(net1469),
    .A0(_01768_),
    .A1(_01882_),
    .A2(_01883_),
    .A3(_01885_),
    .S1(net1468),
    .X(_01886_));
 sg13g2_o21ai_1 _07103_ (.B1(net7),
    .Y(_01887_),
    .A1(net6),
    .A2(_01886_));
 sg13g2_a21oi_1 _07104_ (.A1(_01878_),
    .A2(_01881_),
    .Y(_01888_),
    .B1(_01887_));
 sg13g2_nor3_1 _07105_ (.A(\gpio_out_sel[7] ),
    .B(_01876_),
    .C(_01888_),
    .Y(_01889_));
 sg13g2_a21oi_2 _07106_ (.B1(_01889_),
    .Y(uo_out[7]),
    .A2(_00839_),
    .A1(\gpio_out_sel[7] ));
 sg13g2_nand2_1 _07107_ (.Y(_01890_),
    .A(\i_core.cpu.i_core.i_shift.a[2] ),
    .B(net1217));
 sg13g2_inv_1 _07108_ (.Y(_01891_),
    .A(_01890_));
 sg13g2_nand2_1 _07109_ (.Y(_01892_),
    .A(\i_core.cpu.i_core.i_shift.a[3] ),
    .B(net1238));
 sg13g2_a21oi_2 _07110_ (.B1(_00085_),
    .Y(_01893_),
    .A2(_00925_),
    .A1(_00922_));
 sg13g2_nand2_1 _07111_ (.Y(_01894_),
    .A(\i_core.cpu.i_core.i_shift.a[1] ),
    .B(net1231));
 sg13g2_and4_1 _07112_ (.A(\i_core.cpu.i_core.i_shift.a[0] ),
    .B(\i_core.cpu.i_core.i_shift.a[1] ),
    .C(net1233),
    .D(net1231),
    .X(_01895_));
 sg13g2_a22oi_1 _07113_ (.Y(_01896_),
    .B1(net1231),
    .B2(\i_core.cpu.i_core.i_shift.a[0] ),
    .A2(net1233),
    .A1(\i_core.cpu.i_core.i_shift.a[1] ));
 sg13g2_or3_2 _07114_ (.A(_01892_),
    .B(_01895_),
    .C(_01896_),
    .X(_01897_));
 sg13g2_o21ai_1 _07115_ (.B1(_01892_),
    .Y(_01898_),
    .A1(_01895_),
    .A2(_01896_));
 sg13g2_and3_1 _07116_ (.X(_01899_),
    .A(_01651_),
    .B(_01897_),
    .C(_01898_));
 sg13g2_nand3_1 _07117_ (.B(_01897_),
    .C(_01898_),
    .A(_01651_),
    .Y(_01900_));
 sg13g2_a21oi_1 _07118_ (.A1(_01897_),
    .A2(_01898_),
    .Y(_01901_),
    .B1(_01651_));
 sg13g2_a21o_1 _07119_ (.A2(_01898_),
    .A1(_01897_),
    .B1(_01651_),
    .X(_01902_));
 sg13g2_nor3_1 _07120_ (.A(_00840_),
    .B(_01899_),
    .C(_01901_),
    .Y(_01903_));
 sg13g2_nand3_1 _07121_ (.B(_01900_),
    .C(_01902_),
    .A(\i_core.cpu.i_core.multiplier.accum[3] ),
    .Y(_01904_));
 sg13g2_a21oi_1 _07122_ (.A1(_01900_),
    .A2(_01902_),
    .Y(_01905_),
    .B1(\i_core.cpu.i_core.multiplier.accum[3] ));
 sg13g2_o21ai_1 _07123_ (.B1(_00840_),
    .Y(_01906_),
    .A1(_01899_),
    .A2(_01901_));
 sg13g2_nor3_1 _07124_ (.A(_01655_),
    .B(_01903_),
    .C(_01905_),
    .Y(_01907_));
 sg13g2_nand3_1 _07125_ (.B(_01904_),
    .C(_01906_),
    .A(_01654_),
    .Y(_01908_));
 sg13g2_a21oi_1 _07126_ (.A1(_01904_),
    .A2(_01906_),
    .Y(_01909_),
    .B1(_01654_));
 sg13g2_o21ai_1 _07127_ (.B1(_01655_),
    .Y(_01910_),
    .A1(_01903_),
    .A2(_01905_));
 sg13g2_nor3_1 _07128_ (.A(_01890_),
    .B(_01907_),
    .C(_01909_),
    .Y(_01911_));
 sg13g2_nand3_1 _07129_ (.B(_01908_),
    .C(_01910_),
    .A(_01891_),
    .Y(_01912_));
 sg13g2_a21oi_1 _07130_ (.A1(_01908_),
    .A2(_01910_),
    .Y(_01913_),
    .B1(_01891_));
 sg13g2_o21ai_1 _07131_ (.B1(_01890_),
    .Y(_01914_),
    .A1(_01907_),
    .A2(_01909_));
 sg13g2_o21ai_1 _07132_ (.B1(_01658_),
    .Y(_01915_),
    .A1(_01584_),
    .A2(_01656_));
 sg13g2_nand3_1 _07133_ (.B(_01914_),
    .C(_01915_),
    .A(_01912_),
    .Y(_01916_));
 sg13g2_a21oi_1 _07134_ (.A1(_01912_),
    .A2(_01914_),
    .Y(_01917_),
    .B1(_01915_));
 sg13g2_nor3_1 _07135_ (.A(_01911_),
    .B(_01913_),
    .C(_01915_),
    .Y(_01918_));
 sg13g2_o21ai_1 _07136_ (.B1(_01915_),
    .Y(_01919_),
    .A1(_01911_),
    .A2(_01913_));
 sg13g2_nand2b_1 _07137_ (.Y(_01920_),
    .B(_01919_),
    .A_N(_01918_));
 sg13g2_xnor2_1 _07138_ (.Y(_01921_),
    .A(_01660_),
    .B(_01920_));
 sg13g2_xnor2_1 _07139_ (.Y(_01922_),
    .A(_00928_),
    .B(_00977_));
 sg13g2_a21oi_1 _07140_ (.A1(_01141_),
    .A2(_01922_),
    .Y(_01923_),
    .B1(_01275_));
 sg13g2_o21ai_1 _07141_ (.B1(_01923_),
    .Y(_01924_),
    .A1(_01141_),
    .A2(_01922_));
 sg13g2_nand2_1 _07142_ (.Y(_01925_),
    .A(net1374),
    .B(_01142_));
 sg13g2_a21oi_1 _07143_ (.A1(_00928_),
    .A2(_00976_),
    .Y(_01926_),
    .B1(_01279_));
 sg13g2_a22oi_1 _07144_ (.Y(_01927_),
    .B1(_01925_),
    .B2(_01926_),
    .A2(_01281_),
    .A1(_01142_));
 sg13g2_a21oi_1 _07145_ (.A1(_01924_),
    .A2(_01927_),
    .Y(_01928_),
    .B1(_01285_));
 sg13g2_a21oi_1 _07146_ (.A1(_01164_),
    .A2(_01928_),
    .Y(_01929_),
    .B1(_01371_));
 sg13g2_o21ai_1 _07147_ (.B1(_01929_),
    .Y(_01930_),
    .A1(_01164_),
    .A2(_01921_));
 sg13g2_or2_1 _07148_ (.X(_01931_),
    .B(_01369_),
    .A(net1375));
 sg13g2_a21oi_1 _07149_ (.A1(net1375),
    .A2(_01416_),
    .Y(_01932_),
    .B1(_01372_));
 sg13g2_a21oi_1 _07150_ (.A1(_01931_),
    .A2(_01932_),
    .Y(_01933_),
    .B1(_01638_));
 sg13g2_mux2_1 _07151_ (.A0(\i_core.cpu.instr_data_in[7] ),
    .A1(\i_core.cpu.instr_data_in[15] ),
    .S(_01431_),
    .X(_01934_));
 sg13g2_o21ai_1 _07152_ (.B1(net1360),
    .Y(_01935_),
    .A1(_01186_),
    .A2(_01934_));
 sg13g2_nand3b_1 _07153_ (.B(_01477_),
    .C(_01728_),
    .Y(_01936_),
    .A_N(_01889_));
 sg13g2_a22oi_1 _07154_ (.Y(_01937_),
    .B1(_01480_),
    .B2(\gpio_out_sel[7] ),
    .A2(net1236),
    .A1(\i_spi.data[7] ));
 sg13g2_nand2_1 _07155_ (.Y(_01938_),
    .A(net8),
    .B(_01479_));
 sg13g2_nand3_1 _07156_ (.B(_01937_),
    .C(_01938_),
    .A(_01493_),
    .Y(_01939_));
 sg13g2_a21oi_2 _07157_ (.B1(_01939_),
    .Y(_01940_),
    .A2(net1235),
    .A1(\i_uart_rx.recieved_data[7] ));
 sg13g2_a21o_1 _07158_ (.A2(_01940_),
    .A1(_01936_),
    .B1(_01935_),
    .X(_01941_));
 sg13g2_mux2_1 _07159_ (.A0(\i_core.cpu.instr_data_in[11] ),
    .A1(\i_core.mem.qspi_data_buf[11] ),
    .S(_01433_),
    .X(_01942_));
 sg13g2_nand2b_1 _07160_ (.Y(_01943_),
    .B(net1190),
    .A_N(\i_core.mem.qspi_data_buf[15] ));
 sg13g2_a21oi_1 _07161_ (.A1(_00838_),
    .A2(_01432_),
    .Y(_01944_),
    .B1(net1377));
 sg13g2_a221oi_1 _07162_ (.B2(_01944_),
    .C1(_01186_),
    .B1(_01943_),
    .A1(net1377),
    .Y(_01945_),
    .A2(_01942_));
 sg13g2_nor3_1 _07163_ (.A(_00787_),
    .B(net1234),
    .C(_01945_),
    .Y(_01946_));
 sg13g2_o21ai_1 _07164_ (.B1(\i_core.cpu.instr_data_in[3] ),
    .Y(_01947_),
    .A1(_01190_),
    .A2(_01430_));
 sg13g2_nand2_1 _07165_ (.Y(_01948_),
    .A(\i_core.cpu.instr_data_in[11] ),
    .B(net1202));
 sg13g2_a21oi_1 _07166_ (.A1(\i_core.cpu.instr_data_in[11] ),
    .A2(_01431_),
    .Y(_01949_),
    .B1(_01186_));
 sg13g2_a22oi_1 _07167_ (.Y(_01950_),
    .B1(uo_out[3]),
    .B2(_01477_),
    .A2(_01479_),
    .A1(net1470));
 sg13g2_a22oi_1 _07168_ (.Y(_01951_),
    .B1(_01480_),
    .B2(\gpio_out_sel[3] ),
    .A2(net1236),
    .A1(\i_spi.data[3] ));
 sg13g2_and2_1 _07169_ (.A(_01950_),
    .B(_01951_),
    .X(_01952_));
 sg13g2_a21oi_2 _07170_ (.B1(_01494_),
    .Y(_01953_),
    .A2(_01474_),
    .A1(\i_uart_rx.recieved_data[3] ));
 sg13g2_a221oi_1 _07171_ (.B2(_01953_),
    .C1(_00875_),
    .B1(_01952_),
    .A1(_01947_),
    .Y(_01954_),
    .A2(_01949_));
 sg13g2_nor3_1 _07172_ (.A(net1405),
    .B(_01946_),
    .C(_01954_),
    .Y(_01955_));
 sg13g2_nand2_1 _07173_ (.Y(_01956_),
    .A(\i_core.mem.qspi_data_buf[31] ),
    .B(_01430_));
 sg13g2_a21oi_1 _07174_ (.A1(\i_core.cpu.instr_data_in[15] ),
    .A2(net1202),
    .Y(_01957_),
    .B1(net1377));
 sg13g2_a21oi_1 _07175_ (.A1(\i_core.mem.qspi_data_buf[27] ),
    .A2(_01430_),
    .Y(_01958_),
    .B1(net1412));
 sg13g2_a221oi_1 _07176_ (.B2(_01948_),
    .C1(_01434_),
    .B1(_01958_),
    .A1(_01956_),
    .Y(_01959_),
    .A2(_01957_));
 sg13g2_a22oi_1 _07177_ (.Y(_01960_),
    .B1(net1360),
    .B2(\i_core.mem.data_from_read[23] ),
    .A2(net1368),
    .A1(\i_core.mem.data_from_read[19] ));
 sg13g2_a21oi_1 _07178_ (.A1(net1335),
    .A2(_01960_),
    .Y(_01961_),
    .B1(net1234));
 sg13g2_nor3_1 _07179_ (.A(net1380),
    .B(_01959_),
    .C(_01961_),
    .Y(_01962_));
 sg13g2_a21oi_2 _07180_ (.B1(_01962_),
    .Y(_01963_),
    .A2(_01955_),
    .A1(_01941_));
 sg13g2_nand2b_2 _07181_ (.Y(_01964_),
    .B(_01963_),
    .A_N(_01497_));
 sg13g2_nand2b_1 _07182_ (.Y(_01965_),
    .B(_00974_),
    .A_N(_01176_));
 sg13g2_xnor2_1 _07183_ (.Y(_01966_),
    .A(_00162_),
    .B(_01679_));
 sg13g2_inv_1 _07184_ (.Y(_01967_),
    .A(_01966_));
 sg13g2_xnor2_1 _07185_ (.Y(_01968_),
    .A(_00165_),
    .B(_01223_));
 sg13g2_inv_1 _07186_ (.Y(_01969_),
    .A(_01968_));
 sg13g2_a21oi_1 _07187_ (.A1(net1413),
    .A2(_01967_),
    .Y(_01970_),
    .B1(_01227_));
 sg13g2_o21ai_1 _07188_ (.B1(_01970_),
    .Y(_01971_),
    .A1(net1413),
    .A2(_01968_));
 sg13g2_a21oi_1 _07189_ (.A1(net1426),
    .A2(_01220_),
    .Y(_01972_),
    .B1(net1425));
 sg13g2_or2_1 _07190_ (.X(_01973_),
    .B(_01972_),
    .A(_01221_));
 sg13g2_inv_1 _07191_ (.Y(_01974_),
    .A(_01973_));
 sg13g2_nor2_1 _07192_ (.A(_00877_),
    .B(_01974_),
    .Y(_01975_));
 sg13g2_xnor2_1 _07193_ (.Y(_01976_),
    .A(_00201_),
    .B(_01210_));
 sg13g2_xor2_1 _07194_ (.B(_01207_),
    .A(net1427),
    .X(_01977_));
 sg13g2_nor2_1 _07195_ (.A(_00880_),
    .B(_01977_),
    .Y(_01978_));
 sg13g2_xor2_1 _07196_ (.B(_01204_),
    .A(net1428),
    .X(_01979_));
 sg13g2_nor2_1 _07197_ (.A(_00875_),
    .B(_01979_),
    .Y(_01980_));
 sg13g2_o21ai_1 _07198_ (.B1(net1381),
    .Y(_01981_),
    .A1(_00882_),
    .A2(_01976_));
 sg13g2_or4_1 _07199_ (.A(_01975_),
    .B(_01978_),
    .C(_01980_),
    .D(_01981_),
    .X(_01982_));
 sg13g2_a21oi_1 _07200_ (.A1(_01971_),
    .A2(_01982_),
    .Y(_01983_),
    .B1(_01198_));
 sg13g2_nand2_1 _07201_ (.Y(_01984_),
    .A(_01243_),
    .B(_01461_));
 sg13g2_nor2_1 _07202_ (.A(_01265_),
    .B(_01686_),
    .Y(_01985_));
 sg13g2_a22oi_1 _07203_ (.Y(_01986_),
    .B1(_01985_),
    .B2(\i_core.cpu.i_core.mstatus_mpie ),
    .A2(_01247_),
    .A1(\i_core.cpu.i_core.mcause[3] ));
 sg13g2_nand2_1 _07204_ (.Y(_01987_),
    .A(_01984_),
    .B(_01986_));
 sg13g2_nand2_1 _07205_ (.Y(_01988_),
    .A(\i_core.cpu.i_core.cycle_count[3] ),
    .B(_01261_));
 sg13g2_mux2_1 _07206_ (.A0(\i_core.cpu.i_core.time_hi[2] ),
    .A1(\i_core.cpu.i_core.i_cycles.i_regbuf[6].A ),
    .S(net1308),
    .X(_01989_));
 sg13g2_a22oi_1 _07207_ (.Y(_01990_),
    .B1(_01989_),
    .B2(_01260_),
    .A2(_01262_),
    .A1(\i_core.cpu.i_core.i_instrret.data[3] ));
 sg13g2_a22oi_1 _07208_ (.Y(_01991_),
    .B1(_01267_),
    .B2(_01159_),
    .A2(_01251_),
    .A1(\i_core.cpu.i_core.mie[19] ));
 sg13g2_nor2_1 _07209_ (.A(net1311),
    .B(_01686_),
    .Y(_01992_));
 sg13g2_a22oi_1 _07210_ (.Y(_01993_),
    .B1(_01992_),
    .B2(\i_core.cpu.i_core.mstatus_mie ),
    .A2(_01256_),
    .A1(\i_core.cpu.i_core.mepc[3] ));
 sg13g2_nand4_1 _07211_ (.B(_01990_),
    .C(_01991_),
    .A(_01988_),
    .Y(_01994_),
    .D(_01993_));
 sg13g2_o21ai_1 _07212_ (.B1(_01233_),
    .Y(_01995_),
    .A1(_01987_),
    .A2(_01994_));
 sg13g2_nand2_1 _07213_ (.Y(_01996_),
    .A(_01176_),
    .B(_01995_));
 sg13g2_o21ai_1 _07214_ (.B1(_01965_),
    .Y(_01997_),
    .A1(_01983_),
    .A2(_01996_));
 sg13g2_a221oi_1 _07215_ (.B2(_01196_),
    .C1(_01195_),
    .B1(_01997_),
    .A1(_01505_),
    .Y(_01998_),
    .A2(_01964_));
 sg13g2_a21o_2 _07216_ (.A2(_01933_),
    .A1(_01930_),
    .B1(_01998_),
    .X(\debug_rd[3] ));
 sg13g2_mux2_1 _07217_ (.A0(net2185),
    .A1(net1110),
    .S(_01513_),
    .X(_00053_));
 sg13g2_nand2b_2 _07218_ (.Y(_01999_),
    .B(\i_core.cpu.i_core.i_registers.rd[1] ),
    .A_N(\i_core.cpu.i_core.i_registers.rd[0] ));
 sg13g2_nor2_2 _07219_ (.A(_01512_),
    .B(_01999_),
    .Y(_02000_));
 sg13g2_mux2_1 _07220_ (.A0(net2298),
    .A1(net1165),
    .S(_02000_),
    .X(_00046_));
 sg13g2_mux2_1 _07221_ (.A0(net2296),
    .A1(net1131),
    .S(_02000_),
    .X(_00047_));
 sg13g2_mux2_1 _07222_ (.A0(net2437),
    .A1(net1126),
    .S(_02000_),
    .X(_00048_));
 sg13g2_mux2_1 _07223_ (.A0(net2340),
    .A1(net1110),
    .S(_02000_),
    .X(_00049_));
 sg13g2_nand2_2 _07224_ (.Y(_02001_),
    .A(_00830_),
    .B(\i_core.cpu.i_core.i_registers.rd[0] ));
 sg13g2_nor2_2 _07225_ (.A(_01512_),
    .B(_02001_),
    .Y(_02002_));
 sg13g2_mux2_1 _07226_ (.A0(net2239),
    .A1(net1166),
    .S(_02002_),
    .X(_00042_));
 sg13g2_mux2_1 _07227_ (.A0(net2242),
    .A1(net1132),
    .S(_02002_),
    .X(_00043_));
 sg13g2_mux2_1 _07228_ (.A0(net2530),
    .A1(net1127),
    .S(_02002_),
    .X(_00044_));
 sg13g2_mux2_1 _07229_ (.A0(net2371),
    .A1(net1111),
    .S(_02002_),
    .X(_00045_));
 sg13g2_nor3_2 _07230_ (.A(\i_core.cpu.i_core.i_registers.rd[1] ),
    .B(\i_core.cpu.i_core.i_registers.rd[0] ),
    .C(_01512_),
    .Y(_02003_));
 sg13g2_mux2_1 _07231_ (.A0(net2446),
    .A1(net1165),
    .S(_02003_),
    .X(_00038_));
 sg13g2_mux2_1 _07232_ (.A0(net2380),
    .A1(net1131),
    .S(_02003_),
    .X(_00039_));
 sg13g2_mux2_1 _07233_ (.A0(net2479),
    .A1(net1126),
    .S(_02003_),
    .X(_00040_));
 sg13g2_mux2_1 _07234_ (.A0(net2445),
    .A1(net1110),
    .S(_02003_),
    .X(_00041_));
 sg13g2_nand3b_1 _07235_ (.B(\i_core.cpu.i_core.i_registers.rd[3] ),
    .C(_01511_),
    .Y(_02004_),
    .A_N(\i_core.cpu.i_core.i_registers.rd[2] ));
 sg13g2_nor2_2 _07236_ (.A(_01507_),
    .B(_02004_),
    .Y(_02005_));
 sg13g2_mux2_1 _07237_ (.A0(net2561),
    .A1(net1165),
    .S(_02005_),
    .X(_00034_));
 sg13g2_mux2_1 _07238_ (.A0(net2495),
    .A1(net1131),
    .S(_02005_),
    .X(_00035_));
 sg13g2_mux2_1 _07239_ (.A0(net2548),
    .A1(net1126),
    .S(_02005_),
    .X(_00036_));
 sg13g2_mux2_1 _07240_ (.A0(net2557),
    .A1(net1111),
    .S(_02005_),
    .X(_00037_));
 sg13g2_nor2_2 _07241_ (.A(_01999_),
    .B(_02004_),
    .Y(_02006_));
 sg13g2_mux2_1 _07242_ (.A0(net2084),
    .A1(net1166),
    .S(_02006_),
    .X(_00030_));
 sg13g2_mux2_1 _07243_ (.A0(net2312),
    .A1(net1131),
    .S(_02006_),
    .X(_00031_));
 sg13g2_mux2_1 _07244_ (.A0(net2436),
    .A1(net1127),
    .S(_02006_),
    .X(_00032_));
 sg13g2_mux2_1 _07245_ (.A0(net2360),
    .A1(net1110),
    .S(_02006_),
    .X(_00033_));
 sg13g2_nor2_2 _07246_ (.A(_02001_),
    .B(_02004_),
    .Y(_02007_));
 sg13g2_mux2_1 _07247_ (.A0(net2508),
    .A1(net1165),
    .S(_02007_),
    .X(_00078_));
 sg13g2_mux2_1 _07248_ (.A0(net2390),
    .A1(net1131),
    .S(_02007_),
    .X(_00079_));
 sg13g2_mux2_1 _07249_ (.A0(net2455),
    .A1(net1126),
    .S(_02007_),
    .X(_00080_));
 sg13g2_mux2_1 _07250_ (.A0(net2457),
    .A1(net1110),
    .S(_02007_),
    .X(_00081_));
 sg13g2_nor3_2 _07251_ (.A(\i_core.cpu.i_core.i_registers.rd[1] ),
    .B(\i_core.cpu.i_core.i_registers.rd[0] ),
    .C(_02004_),
    .Y(_02008_));
 sg13g2_mux2_1 _07252_ (.A0(net2322),
    .A1(net1165),
    .S(_02008_),
    .X(_00074_));
 sg13g2_mux2_1 _07253_ (.A0(net2306),
    .A1(net1131),
    .S(_02008_),
    .X(_00075_));
 sg13g2_mux2_1 _07254_ (.A0(net2275),
    .A1(net1127),
    .S(_02008_),
    .X(_00076_));
 sg13g2_mux2_1 _07255_ (.A0(net2454),
    .A1(net1110),
    .S(_02008_),
    .X(_00077_));
 sg13g2_nand2b_1 _07256_ (.Y(_02009_),
    .B(\i_core.cpu.i_core.i_registers.rd[2] ),
    .A_N(\i_core.cpu.i_core.i_registers.rd[3] ));
 sg13g2_nand3_1 _07257_ (.B(\i_core.cpu.i_core.i_registers.rd[0] ),
    .C(\i_core.cpu.i_core.i_registers.rd[2] ),
    .A(\i_core.cpu.i_core.i_registers.rd[1] ),
    .Y(_02010_));
 sg13g2_nor3_2 _07258_ (.A(\i_core.cpu.i_core.i_registers.rd[3] ),
    .B(_01510_),
    .C(_02010_),
    .Y(_02011_));
 sg13g2_mux2_1 _07259_ (.A0(net2029),
    .A1(net1166),
    .S(_02011_),
    .X(_00070_));
 sg13g2_mux2_1 _07260_ (.A0(net2192),
    .A1(net1132),
    .S(_02011_),
    .X(_00071_));
 sg13g2_mux2_1 _07261_ (.A0(net2294),
    .A1(net1126),
    .S(_02011_),
    .X(_00072_));
 sg13g2_mux2_1 _07262_ (.A0(net2245),
    .A1(net1111),
    .S(_02011_),
    .X(_00073_));
 sg13g2_nor3_2 _07263_ (.A(_01510_),
    .B(_01999_),
    .C(_02009_),
    .Y(_02012_));
 sg13g2_mux2_1 _07264_ (.A0(net2507),
    .A1(net1166),
    .S(_02012_),
    .X(_00066_));
 sg13g2_mux2_1 _07265_ (.A0(net2425),
    .A1(net1132),
    .S(_02012_),
    .X(_00067_));
 sg13g2_mux2_1 _07266_ (.A0(net2539),
    .A1(net1127),
    .S(_02012_),
    .X(_00068_));
 sg13g2_mux2_1 _07267_ (.A0(net2385),
    .A1(net1111),
    .S(_02012_),
    .X(_00069_));
 sg13g2_nor3_2 _07268_ (.A(_01510_),
    .B(_02001_),
    .C(_02009_),
    .Y(_02013_));
 sg13g2_mux2_1 _07269_ (.A0(net2574),
    .A1(net1166),
    .S(_02013_),
    .X(_00062_));
 sg13g2_mux2_1 _07270_ (.A0(net2584),
    .A1(net1132),
    .S(_02013_),
    .X(_00063_));
 sg13g2_mux2_1 _07271_ (.A0(net2590),
    .A1(net1126),
    .S(_02013_),
    .X(_00064_));
 sg13g2_mux2_1 _07272_ (.A0(net2567),
    .A1(net1111),
    .S(_02013_),
    .X(_00065_));
 sg13g2_nor4_2 _07273_ (.A(\i_core.cpu.i_core.i_registers.rd[2] ),
    .B(\i_core.cpu.i_core.i_registers.rd[3] ),
    .C(_01510_),
    .Y(_02014_),
    .D(_01999_));
 sg13g2_mux2_1 _07274_ (.A0(net2295),
    .A1(net1165),
    .S(_02014_),
    .X(_00058_));
 sg13g2_mux2_1 _07275_ (.A0(net2207),
    .A1(net1132),
    .S(_02014_),
    .X(_00059_));
 sg13g2_mux2_1 _07276_ (.A0(net2280),
    .A1(net1126),
    .S(_02014_),
    .X(_00060_));
 sg13g2_mux2_1 _07277_ (.A0(net2218),
    .A1(net1110),
    .S(_02014_),
    .X(_00061_));
 sg13g2_nor4_2 _07278_ (.A(\i_core.cpu.i_core.i_registers.rd[2] ),
    .B(\i_core.cpu.i_core.i_registers.rd[3] ),
    .C(_01510_),
    .Y(_02015_),
    .D(_02001_));
 sg13g2_mux2_1 _07279_ (.A0(net2330),
    .A1(net1165),
    .S(_02015_),
    .X(_00054_));
 sg13g2_mux2_1 _07280_ (.A0(net2402),
    .A1(net1131),
    .S(_02015_),
    .X(_00055_));
 sg13g2_mux2_1 _07281_ (.A0(net2257),
    .A1(net1127),
    .S(_02015_),
    .X(_00056_));
 sg13g2_mux2_1 _07282_ (.A0(net2243),
    .A1(net1110),
    .S(_02015_),
    .X(_00057_));
 sg13g2_nor2b_2 _07283_ (.A(\i_core.mem.q_ctrl.fsm_state[0] ),
    .B_N(\i_core.mem.q_ctrl.fsm_state[1] ),
    .Y(_02016_));
 sg13g2_nor2b_2 _07284_ (.A(net1431),
    .B_N(\i_core.mem.q_ctrl.fsm_state[0] ),
    .Y(_02017_));
 sg13g2_or2_1 _07285_ (.X(_02018_),
    .B(net1429),
    .A(net1430));
 sg13g2_a22oi_1 _07286_ (.Y(_02019_),
    .B1(_02017_),
    .B2(_02018_),
    .A2(_02016_),
    .A1(_00768_));
 sg13g2_nand2_1 _07287_ (.Y(_02020_),
    .A(net1429),
    .B(_02017_));
 sg13g2_or2_1 _07288_ (.X(_02021_),
    .B(_02020_),
    .A(\i_core.mem.q_ctrl.nibbles_remaining[0] ));
 sg13g2_nor2_1 _07289_ (.A(net1434),
    .B(_02021_),
    .Y(_02022_));
 sg13g2_and2_1 _07290_ (.A(net1430),
    .B(\i_core.mem.q_ctrl.fsm_state[0] ),
    .X(_02023_));
 sg13g2_nand2_1 _07291_ (.Y(_02024_),
    .A(net1430),
    .B(\i_core.mem.q_ctrl.fsm_state[0] ));
 sg13g2_nor2_2 _07292_ (.A(net1431),
    .B(net1334),
    .Y(_02025_));
 sg13g2_and2_2 _07293_ (.A(_00152_),
    .B(_02016_),
    .X(_02026_));
 sg13g2_a221oi_1 _07294_ (.B2(\i_core.mem.q_ctrl.addr[20] ),
    .C1(_02022_),
    .B1(_02026_),
    .A1(_00845_),
    .Y(_02027_),
    .A2(_02025_));
 sg13g2_nor2_2 _07295_ (.A(_02019_),
    .B(_02027_),
    .Y(uio_out[1]));
 sg13g2_nand2b_1 _07296_ (.Y(_02028_),
    .B(_02025_),
    .A_N(_00206_));
 sg13g2_a21oi_1 _07297_ (.A1(\i_core.mem.q_ctrl.addr[21] ),
    .A2(_02026_),
    .Y(_02029_),
    .B1(_02019_));
 sg13g2_nand3_1 _07298_ (.B(_02028_),
    .C(_02029_),
    .A(_02021_),
    .Y(uio_out[2]));
 sg13g2_a22oi_1 _07299_ (.Y(_02030_),
    .B1(_02026_),
    .B2(\i_core.mem.q_ctrl.addr[22] ),
    .A2(_02025_),
    .A1(\i_core.cpu.instr_data_in[14] ));
 sg13g2_nor2_2 _07300_ (.A(_02019_),
    .B(_02030_),
    .Y(uio_out[4]));
 sg13g2_a221oi_1 _07301_ (.B2(\i_core.mem.q_ctrl.addr[23] ),
    .C1(_02019_),
    .B1(_02026_),
    .A1(_00848_),
    .Y(_02031_),
    .A2(_02025_));
 sg13g2_o21ai_1 _07302_ (.B1(_02031_),
    .Y(uio_out[5]),
    .A1(net1434),
    .A2(_02021_));
 sg13g2_and2_2 _07303_ (.A(\i_core.mem.q_ctrl.spi_data_oe[0] ),
    .B(net1),
    .X(uio_oe[5]));
 sg13g2_nand2_1 _07304_ (.Y(_02032_),
    .A(net1325),
    .B(net2160));
 sg13g2_and3_1 _07305_ (.X(_02033_),
    .A(_01482_),
    .B(_01483_),
    .C(_01883_));
 sg13g2_nand2_1 _07306_ (.Y(_02034_),
    .A(\data_to_write[0] ),
    .B(_02033_));
 sg13g2_o21ai_1 _07307_ (.B1(_02034_),
    .Y(_00000_),
    .A1(_02032_),
    .A2(net1212));
 sg13g2_nand2_1 _07308_ (.Y(_02035_),
    .A(net1326),
    .B(net2004));
 sg13g2_nand2_1 _07309_ (.Y(_02036_),
    .A(\data_to_write[1] ),
    .B(net1212));
 sg13g2_o21ai_1 _07310_ (.B1(_02036_),
    .Y(_00001_),
    .A1(net1212),
    .A2(_02035_));
 sg13g2_nand2_1 _07311_ (.Y(_02037_),
    .A(net1325),
    .B(net2010));
 sg13g2_nand2_1 _07312_ (.Y(_02038_),
    .A(\data_to_write[2] ),
    .B(net1212));
 sg13g2_o21ai_1 _07313_ (.B1(_02038_),
    .Y(_00002_),
    .A1(net1212),
    .A2(_02037_));
 sg13g2_nand2_1 _07314_ (.Y(_02039_),
    .A(net1323),
    .B(net2014));
 sg13g2_nand2_1 _07315_ (.Y(_02040_),
    .A(\data_to_write[3] ),
    .B(net1211));
 sg13g2_o21ai_1 _07316_ (.B1(_02040_),
    .Y(_00003_),
    .A1(net1211),
    .A2(_02039_));
 sg13g2_nand2_1 _07317_ (.Y(_02041_),
    .A(net1322),
    .B(net1986));
 sg13g2_nand2_1 _07318_ (.Y(_02042_),
    .A(\data_to_write[4] ),
    .B(net1211));
 sg13g2_o21ai_1 _07319_ (.B1(_02042_),
    .Y(_00004_),
    .A1(net1211),
    .A2(_02041_));
 sg13g2_nand2_1 _07320_ (.Y(_02043_),
    .A(net1321),
    .B(net2101));
 sg13g2_nand2_1 _07321_ (.Y(_02044_),
    .A(\data_to_write[5] ),
    .B(net1211));
 sg13g2_o21ai_1 _07322_ (.B1(_02044_),
    .Y(_00005_),
    .A1(net1211),
    .A2(_02043_));
 sg13g2_nand2_1 _07323_ (.Y(_02045_),
    .A(net1322),
    .B(net2066));
 sg13g2_nand2_1 _07324_ (.Y(_02046_),
    .A(\data_to_write[6] ),
    .B(net1211));
 sg13g2_o21ai_1 _07325_ (.B1(_02046_),
    .Y(_00006_),
    .A1(net1211),
    .A2(_02045_));
 sg13g2_nand2_1 _07326_ (.Y(_02047_),
    .A(net1323),
    .B(net1988));
 sg13g2_nand2_1 _07327_ (.Y(_02048_),
    .A(\data_to_write[7] ),
    .B(net1212));
 sg13g2_o21ai_1 _07328_ (.B1(_02048_),
    .Y(_00007_),
    .A1(net1212),
    .A2(_02047_));
 sg13g2_nand2_1 _07329_ (.Y(_02049_),
    .A(net1325),
    .B(net2258));
 sg13g2_nor4_1 _07330_ (.A(net1450),
    .B(_01456_),
    .C(_01467_),
    .D(_01884_),
    .Y(_02050_));
 sg13g2_nand2_1 _07331_ (.Y(_02051_),
    .A(\data_to_write[0] ),
    .B(net1210));
 sg13g2_o21ai_1 _07332_ (.B1(_02051_),
    .Y(_00008_),
    .A1(_02049_),
    .A2(net1210));
 sg13g2_nand2_1 _07333_ (.Y(_02052_),
    .A(net1326),
    .B(net2232));
 sg13g2_nand2_1 _07334_ (.Y(_02053_),
    .A(\data_to_write[1] ),
    .B(net1210));
 sg13g2_o21ai_1 _07335_ (.B1(_02053_),
    .Y(_00009_),
    .A1(net1210),
    .A2(_02052_));
 sg13g2_nand2_1 _07336_ (.Y(_02054_),
    .A(net1325),
    .B(net2193));
 sg13g2_nand2_1 _07337_ (.Y(_02055_),
    .A(\data_to_write[2] ),
    .B(net1210));
 sg13g2_o21ai_1 _07338_ (.B1(_02055_),
    .Y(_00010_),
    .A1(net1210),
    .A2(_02054_));
 sg13g2_nand2_1 _07339_ (.Y(_02056_),
    .A(net1323),
    .B(net2195));
 sg13g2_nand2_1 _07340_ (.Y(_02057_),
    .A(\data_to_write[3] ),
    .B(net1209));
 sg13g2_o21ai_1 _07341_ (.B1(_02057_),
    .Y(_00011_),
    .A1(net1209),
    .A2(_02056_));
 sg13g2_nand2_1 _07342_ (.Y(_02058_),
    .A(net1324),
    .B(net2246));
 sg13g2_nand2_1 _07343_ (.Y(_02059_),
    .A(\data_to_write[4] ),
    .B(net1209));
 sg13g2_o21ai_1 _07344_ (.B1(_02059_),
    .Y(_00012_),
    .A1(net1209),
    .A2(_02058_));
 sg13g2_nand2_1 _07345_ (.Y(_02060_),
    .A(net1325),
    .B(net2253));
 sg13g2_nand2_1 _07346_ (.Y(_02061_),
    .A(\data_to_write[5] ),
    .B(net1209));
 sg13g2_o21ai_1 _07347_ (.B1(_02061_),
    .Y(_00013_),
    .A1(net1209),
    .A2(_02060_));
 sg13g2_nand2_1 _07348_ (.Y(_02062_),
    .A(net1323),
    .B(net2310));
 sg13g2_nand2_1 _07349_ (.Y(_02063_),
    .A(\data_to_write[6] ),
    .B(net1209));
 sg13g2_o21ai_1 _07350_ (.B1(_02063_),
    .Y(_00014_),
    .A1(net1209),
    .A2(_02062_));
 sg13g2_nand2_1 _07351_ (.Y(_02064_),
    .A(net1323),
    .B(net2661));
 sg13g2_o21ai_1 _07352_ (.B1(_02064_),
    .Y(_02065_),
    .A1(net1323),
    .A2(net1468));
 sg13g2_mux2_1 _07353_ (.A0(_02065_),
    .A1(net2471),
    .S(net1210),
    .X(_00015_));
 sg13g2_a22oi_1 _07354_ (.Y(_02066_),
    .B1(net1336),
    .B2(net1392),
    .A2(_01156_),
    .A1(\i_core.cpu.is_load ));
 sg13g2_nor2_2 _07355_ (.A(\i_core.cpu.i_core.cycle[1] ),
    .B(\i_core.cpu.i_core.cycle[0] ),
    .Y(_02067_));
 sg13g2_nor4_2 _07356_ (.A(\i_core.cpu.i_core.cycle[1] ),
    .B(\i_core.cpu.i_core.cycle[0] ),
    .C(net1308),
    .Y(_02068_),
    .D(_02066_));
 sg13g2_nand3b_1 _07357_ (.B(_02067_),
    .C(net1310),
    .Y(_02069_),
    .A_N(_02066_));
 sg13g2_nand2_1 _07358_ (.Y(_02070_),
    .A(\i_core.cpu.is_load ),
    .B(net1188));
 sg13g2_nand3_1 _07359_ (.B(net1188),
    .C(_02068_),
    .A(\i_core.cpu.is_load ),
    .Y(_02071_));
 sg13g2_nand2_2 _07360_ (.Y(_02072_),
    .A(\i_core.cpu.is_store ),
    .B(_02068_));
 sg13g2_nand2_1 _07361_ (.Y(_02073_),
    .A(_02071_),
    .B(_02072_));
 sg13g2_nor2_1 _07362_ (.A(net2237),
    .B(_02073_),
    .Y(_02074_));
 sg13g2_a221oi_1 _07363_ (.B2(_01772_),
    .C1(_02074_),
    .B1(_02073_),
    .A1(net1458),
    .Y(_00028_),
    .A2(_02071_));
 sg13g2_o21ai_1 _07364_ (.B1(_01916_),
    .Y(_02075_),
    .A1(_01661_),
    .A2(_01917_));
 sg13g2_nand2_1 _07365_ (.Y(_02076_),
    .A(\i_core.cpu.i_core.i_shift.a[3] ),
    .B(net1217));
 sg13g2_nand2_1 _07366_ (.Y(_02077_),
    .A(_01900_),
    .B(_01904_));
 sg13g2_nand2b_1 _07367_ (.Y(_02078_),
    .B(_01897_),
    .A_N(_01895_));
 sg13g2_nand2_1 _07368_ (.Y(_02079_),
    .A(\i_core.cpu.i_core.i_shift.a[4] ),
    .B(net1238));
 sg13g2_xor2_1 _07369_ (.B(_01894_),
    .A(_01650_),
    .X(_02080_));
 sg13g2_nand2b_1 _07370_ (.Y(_02081_),
    .B(_02080_),
    .A_N(_02079_));
 sg13g2_xnor2_1 _07371_ (.Y(_02082_),
    .A(_02079_),
    .B(_02080_));
 sg13g2_nand2_1 _07372_ (.Y(_02083_),
    .A(_02078_),
    .B(_02082_));
 sg13g2_xnor2_1 _07373_ (.Y(_02084_),
    .A(_02078_),
    .B(_02082_));
 sg13g2_xnor2_1 _07374_ (.Y(_02085_),
    .A(_00861_),
    .B(_02084_));
 sg13g2_nand2b_1 _07375_ (.Y(_02086_),
    .B(_02077_),
    .A_N(_02085_));
 sg13g2_xnor2_1 _07376_ (.Y(_02087_),
    .A(_02077_),
    .B(_02085_));
 sg13g2_nand2b_1 _07377_ (.Y(_02088_),
    .B(_02087_),
    .A_N(_02076_));
 sg13g2_xnor2_1 _07378_ (.Y(_02089_),
    .A(_02076_),
    .B(_02087_));
 sg13g2_nand2_1 _07379_ (.Y(_02090_),
    .A(_01908_),
    .B(_01912_));
 sg13g2_and2_1 _07380_ (.A(_02089_),
    .B(_02090_),
    .X(_02091_));
 sg13g2_xor2_1 _07381_ (.B(_02090_),
    .A(_02089_),
    .X(_02092_));
 sg13g2_xor2_1 _07382_ (.B(_02092_),
    .A(_02075_),
    .X(_00016_));
 sg13g2_a21oi_1 _07383_ (.A1(_02075_),
    .A2(_02092_),
    .Y(_02093_),
    .B1(_02091_));
 sg13g2_nand2_1 _07384_ (.Y(_02094_),
    .A(\i_core.cpu.i_core.i_shift.a[4] ),
    .B(net1217));
 sg13g2_o21ai_1 _07385_ (.B1(_02083_),
    .Y(_02095_),
    .A1(_00861_),
    .A2(_02084_));
 sg13g2_o21ai_1 _07386_ (.B1(_02081_),
    .Y(_02096_),
    .A1(_01650_),
    .A2(_01894_));
 sg13g2_nand2_1 _07387_ (.Y(_02097_),
    .A(\i_core.cpu.i_core.i_shift.a[5] ),
    .B(net1237));
 sg13g2_nand2_2 _07388_ (.Y(_02098_),
    .A(\i_core.cpu.i_core.i_shift.a[3] ),
    .B(net1231));
 sg13g2_nor2_1 _07389_ (.A(_01650_),
    .B(_02098_),
    .Y(_02099_));
 sg13g2_or2_1 _07390_ (.X(_02100_),
    .B(_02098_),
    .A(_01650_));
 sg13g2_a22oi_1 _07391_ (.Y(_02101_),
    .B1(net1231),
    .B2(\i_core.cpu.i_core.i_shift.a[2] ),
    .A2(net1233),
    .A1(\i_core.cpu.i_core.i_shift.a[3] ));
 sg13g2_nor2_1 _07392_ (.A(_02099_),
    .B(_02101_),
    .Y(_02102_));
 sg13g2_xnor2_1 _07393_ (.Y(_02103_),
    .A(_02097_),
    .B(_02102_));
 sg13g2_nand2_1 _07394_ (.Y(_02104_),
    .A(_02096_),
    .B(_02103_));
 sg13g2_xnor2_1 _07395_ (.Y(_02105_),
    .A(_02096_),
    .B(_02103_));
 sg13g2_xnor2_1 _07396_ (.Y(_02106_),
    .A(_00862_),
    .B(_02105_));
 sg13g2_nand2b_1 _07397_ (.Y(_02107_),
    .B(_02095_),
    .A_N(_02106_));
 sg13g2_xor2_1 _07398_ (.B(_02106_),
    .A(_02095_),
    .X(_02108_));
 sg13g2_xor2_1 _07399_ (.B(_02108_),
    .A(_02094_),
    .X(_02109_));
 sg13g2_nand2_1 _07400_ (.Y(_02110_),
    .A(_02086_),
    .B(_02088_));
 sg13g2_nor2_1 _07401_ (.A(_02109_),
    .B(_02110_),
    .Y(_02111_));
 sg13g2_xor2_1 _07402_ (.B(_02110_),
    .A(_02109_),
    .X(_02112_));
 sg13g2_xnor2_1 _07403_ (.Y(_00019_),
    .A(_02093_),
    .B(_02112_));
 sg13g2_nand2_1 _07404_ (.Y(_02113_),
    .A(\i_core.cpu.i_core.i_shift.a[5] ),
    .B(net1217));
 sg13g2_o21ai_1 _07405_ (.B1(_02104_),
    .Y(_02114_),
    .A1(_00862_),
    .A2(_02105_));
 sg13g2_o21ai_1 _07406_ (.B1(_02100_),
    .Y(_02115_),
    .A1(_02097_),
    .A2(_02101_));
 sg13g2_nand2_1 _07407_ (.Y(_02116_),
    .A(\i_core.cpu.i_core.i_shift.a[6] ),
    .B(net1237));
 sg13g2_nand2_1 _07408_ (.Y(_02117_),
    .A(\i_core.cpu.i_core.i_shift.a[4] ),
    .B(net1231));
 sg13g2_nand2_1 _07409_ (.Y(_02118_),
    .A(\i_core.cpu.i_core.i_shift.a[4] ),
    .B(net1233));
 sg13g2_xor2_1 _07410_ (.B(_02118_),
    .A(_02098_),
    .X(_02119_));
 sg13g2_nand2b_1 _07411_ (.Y(_02120_),
    .B(_02119_),
    .A_N(_02116_));
 sg13g2_xnor2_1 _07412_ (.Y(_02121_),
    .A(_02116_),
    .B(_02119_));
 sg13g2_nand2_1 _07413_ (.Y(_02122_),
    .A(_02115_),
    .B(_02121_));
 sg13g2_xnor2_1 _07414_ (.Y(_02123_),
    .A(_02115_),
    .B(_02121_));
 sg13g2_xnor2_1 _07415_ (.Y(_02124_),
    .A(_00863_),
    .B(_02123_));
 sg13g2_nand2b_1 _07416_ (.Y(_02125_),
    .B(_02114_),
    .A_N(_02124_));
 sg13g2_xor2_1 _07417_ (.B(_02124_),
    .A(_02114_),
    .X(_02126_));
 sg13g2_xor2_1 _07418_ (.B(_02126_),
    .A(_02113_),
    .X(_02127_));
 sg13g2_o21ai_1 _07419_ (.B1(_02107_),
    .Y(_02128_),
    .A1(_02094_),
    .A2(_02108_));
 sg13g2_and2_1 _07420_ (.A(_02127_),
    .B(_02128_),
    .X(_02129_));
 sg13g2_inv_1 _07421_ (.Y(_02130_),
    .A(_02129_));
 sg13g2_xnor2_1 _07422_ (.Y(_02131_),
    .A(_02127_),
    .B(_02128_));
 sg13g2_a221oi_1 _07423_ (.B2(_02110_),
    .C1(_02091_),
    .B1(_02109_),
    .A1(_02075_),
    .Y(_02132_),
    .A2(_02092_));
 sg13g2_or3_1 _07424_ (.A(_02111_),
    .B(_02131_),
    .C(_02132_),
    .X(_02133_));
 sg13g2_o21ai_1 _07425_ (.B1(_02131_),
    .Y(_02134_),
    .A1(_02111_),
    .A2(_02132_));
 sg13g2_and2_1 _07426_ (.A(_02133_),
    .B(_02134_),
    .X(_00020_));
 sg13g2_nand2_1 _07427_ (.Y(_02135_),
    .A(\i_core.cpu.i_core.i_shift.a[6] ),
    .B(net1216));
 sg13g2_o21ai_1 _07428_ (.B1(_02122_),
    .Y(_02136_),
    .A1(_00863_),
    .A2(_02123_));
 sg13g2_o21ai_1 _07429_ (.B1(_02120_),
    .Y(_02137_),
    .A1(_02098_),
    .A2(_02118_));
 sg13g2_nand2_1 _07430_ (.Y(_02138_),
    .A(\i_core.cpu.i_core.i_shift.a[7] ),
    .B(net1237));
 sg13g2_nand2_1 _07431_ (.Y(_02139_),
    .A(\i_core.cpu.i_core.i_shift.a[5] ),
    .B(_01893_));
 sg13g2_nand2_1 _07432_ (.Y(_02140_),
    .A(\i_core.cpu.i_core.i_shift.a[5] ),
    .B(_01649_));
 sg13g2_xor2_1 _07433_ (.B(_02140_),
    .A(_02117_),
    .X(_02141_));
 sg13g2_nand2b_1 _07434_ (.Y(_02142_),
    .B(_02141_),
    .A_N(_02138_));
 sg13g2_xnor2_1 _07435_ (.Y(_02143_),
    .A(_02138_),
    .B(_02141_));
 sg13g2_nand2_1 _07436_ (.Y(_02144_),
    .A(_02137_),
    .B(_02143_));
 sg13g2_xnor2_1 _07437_ (.Y(_02145_),
    .A(_02137_),
    .B(_02143_));
 sg13g2_xnor2_1 _07438_ (.Y(_02146_),
    .A(_00864_),
    .B(_02145_));
 sg13g2_nand2b_1 _07439_ (.Y(_02147_),
    .B(_02136_),
    .A_N(_02146_));
 sg13g2_xor2_1 _07440_ (.B(_02146_),
    .A(_02136_),
    .X(_02148_));
 sg13g2_xor2_1 _07441_ (.B(_02148_),
    .A(_02135_),
    .X(_02149_));
 sg13g2_o21ai_1 _07442_ (.B1(_02125_),
    .Y(_02150_),
    .A1(_02113_),
    .A2(_02126_));
 sg13g2_and2_1 _07443_ (.A(_02149_),
    .B(_02150_),
    .X(_02151_));
 sg13g2_xnor2_1 _07444_ (.Y(_02152_),
    .A(_02149_),
    .B(_02150_));
 sg13g2_a21oi_1 _07445_ (.A1(_02130_),
    .A2(_02133_),
    .Y(_02153_),
    .B1(_02152_));
 sg13g2_nand3_1 _07446_ (.B(_02133_),
    .C(_02152_),
    .A(_02130_),
    .Y(_02154_));
 sg13g2_nor2b_1 _07447_ (.A(_02153_),
    .B_N(_02154_),
    .Y(_00021_));
 sg13g2_nor2_1 _07448_ (.A(_02151_),
    .B(_02153_),
    .Y(_02155_));
 sg13g2_nand2_1 _07449_ (.Y(_02156_),
    .A(\i_core.cpu.i_core.i_shift.a[7] ),
    .B(net1216));
 sg13g2_o21ai_1 _07450_ (.B1(_02144_),
    .Y(_02157_),
    .A1(_00864_),
    .A2(_02145_));
 sg13g2_o21ai_1 _07451_ (.B1(_02142_),
    .Y(_02158_),
    .A1(_02117_),
    .A2(_02140_));
 sg13g2_nand2_1 _07452_ (.Y(_02159_),
    .A(\i_core.cpu.i_core.i_shift.a[8] ),
    .B(_01419_));
 sg13g2_nand2_1 _07453_ (.Y(_02160_),
    .A(\i_core.cpu.i_core.i_shift.a[6] ),
    .B(_01893_));
 sg13g2_nand2_1 _07454_ (.Y(_02161_),
    .A(\i_core.cpu.i_core.i_shift.a[6] ),
    .B(_01649_));
 sg13g2_xor2_1 _07455_ (.B(_02161_),
    .A(_02139_),
    .X(_02162_));
 sg13g2_nand2b_1 _07456_ (.Y(_02163_),
    .B(_02162_),
    .A_N(_02159_));
 sg13g2_xnor2_1 _07457_ (.Y(_02164_),
    .A(_02159_),
    .B(_02162_));
 sg13g2_nand2_1 _07458_ (.Y(_02165_),
    .A(_02158_),
    .B(_02164_));
 sg13g2_xnor2_1 _07459_ (.Y(_02166_),
    .A(_02158_),
    .B(_02164_));
 sg13g2_xnor2_1 _07460_ (.Y(_02167_),
    .A(_00865_),
    .B(_02166_));
 sg13g2_nor2b_1 _07461_ (.A(_02167_),
    .B_N(_02157_),
    .Y(_02168_));
 sg13g2_xor2_1 _07462_ (.B(_02167_),
    .A(_02157_),
    .X(_02169_));
 sg13g2_nor2_1 _07463_ (.A(_02156_),
    .B(_02169_),
    .Y(_02170_));
 sg13g2_xor2_1 _07464_ (.B(_02169_),
    .A(_02156_),
    .X(_02171_));
 sg13g2_o21ai_1 _07465_ (.B1(_02147_),
    .Y(_02172_),
    .A1(_02135_),
    .A2(_02148_));
 sg13g2_nand2_1 _07466_ (.Y(_02173_),
    .A(_02171_),
    .B(_02172_));
 sg13g2_xor2_1 _07467_ (.B(_02172_),
    .A(_02171_),
    .X(_02174_));
 sg13g2_o21ai_1 _07468_ (.B1(_02174_),
    .Y(_02175_),
    .A1(_02151_),
    .A2(_02153_));
 sg13g2_xnor2_1 _07469_ (.Y(_00022_),
    .A(_02155_),
    .B(_02174_));
 sg13g2_nand2_1 _07470_ (.Y(_02176_),
    .A(_02173_),
    .B(_02175_));
 sg13g2_nand2_1 _07471_ (.Y(_02177_),
    .A(\i_core.cpu.i_core.i_shift.a[8] ),
    .B(net1216));
 sg13g2_o21ai_1 _07472_ (.B1(_02165_),
    .Y(_02178_),
    .A1(_00865_),
    .A2(_02166_));
 sg13g2_o21ai_1 _07473_ (.B1(_02163_),
    .Y(_02179_),
    .A1(_02139_),
    .A2(_02161_));
 sg13g2_nand2_1 _07474_ (.Y(_02180_),
    .A(\i_core.cpu.i_core.i_shift.a[9] ),
    .B(_01419_));
 sg13g2_nand2_1 _07475_ (.Y(_02181_),
    .A(\i_core.cpu.i_core.i_shift.a[7] ),
    .B(net1231));
 sg13g2_nand2_1 _07476_ (.Y(_02182_),
    .A(\i_core.cpu.i_core.i_shift.a[7] ),
    .B(_01649_));
 sg13g2_xor2_1 _07477_ (.B(_02182_),
    .A(_02160_),
    .X(_02183_));
 sg13g2_nand2b_1 _07478_ (.Y(_02184_),
    .B(_02183_),
    .A_N(_02180_));
 sg13g2_xnor2_1 _07479_ (.Y(_02185_),
    .A(_02180_),
    .B(_02183_));
 sg13g2_nand2_1 _07480_ (.Y(_02186_),
    .A(_02179_),
    .B(_02185_));
 sg13g2_xnor2_1 _07481_ (.Y(_02187_),
    .A(_02179_),
    .B(_02185_));
 sg13g2_xnor2_1 _07482_ (.Y(_02188_),
    .A(_00866_),
    .B(_02187_));
 sg13g2_nand2b_1 _07483_ (.Y(_02189_),
    .B(_02178_),
    .A_N(_02188_));
 sg13g2_xor2_1 _07484_ (.B(_02188_),
    .A(_02178_),
    .X(_02190_));
 sg13g2_xor2_1 _07485_ (.B(_02190_),
    .A(_02177_),
    .X(_02191_));
 sg13g2_nor2_1 _07486_ (.A(_02168_),
    .B(_02170_),
    .Y(_02192_));
 sg13g2_nor3_1 _07487_ (.A(_02168_),
    .B(_02170_),
    .C(_02191_),
    .Y(_02193_));
 sg13g2_nor2b_1 _07488_ (.A(_02192_),
    .B_N(_02191_),
    .Y(_02194_));
 sg13g2_nor2_1 _07489_ (.A(_02193_),
    .B(_02194_),
    .Y(_02195_));
 sg13g2_xor2_1 _07490_ (.B(_02195_),
    .A(_02176_),
    .X(_00023_));
 sg13g2_nand2_1 _07491_ (.Y(_02196_),
    .A(\i_core.cpu.i_core.i_shift.a[9] ),
    .B(net1216));
 sg13g2_o21ai_1 _07492_ (.B1(_02186_),
    .Y(_02197_),
    .A1(_00866_),
    .A2(_02187_));
 sg13g2_o21ai_1 _07493_ (.B1(_02184_),
    .Y(_02198_),
    .A1(_02160_),
    .A2(_02182_));
 sg13g2_nand2_1 _07494_ (.Y(_02199_),
    .A(\i_core.cpu.i_core.i_shift.a[10] ),
    .B(_01419_));
 sg13g2_nand2_1 _07495_ (.Y(_02200_),
    .A(\i_core.cpu.i_core.i_shift.a[8] ),
    .B(net1230));
 sg13g2_nand2_1 _07496_ (.Y(_02201_),
    .A(\i_core.cpu.i_core.i_shift.a[8] ),
    .B(net1232));
 sg13g2_xor2_1 _07497_ (.B(_02201_),
    .A(_02181_),
    .X(_02202_));
 sg13g2_nand2b_1 _07498_ (.Y(_02203_),
    .B(_02202_),
    .A_N(_02199_));
 sg13g2_xnor2_1 _07499_ (.Y(_02204_),
    .A(_02199_),
    .B(_02202_));
 sg13g2_nand2_1 _07500_ (.Y(_02205_),
    .A(_02198_),
    .B(_02204_));
 sg13g2_xnor2_1 _07501_ (.Y(_02206_),
    .A(_02198_),
    .B(_02204_));
 sg13g2_xnor2_1 _07502_ (.Y(_02207_),
    .A(_00867_),
    .B(_02206_));
 sg13g2_nor2b_1 _07503_ (.A(_02207_),
    .B_N(_02197_),
    .Y(_02208_));
 sg13g2_xor2_1 _07504_ (.B(_02207_),
    .A(_02197_),
    .X(_02209_));
 sg13g2_nor2_1 _07505_ (.A(_02196_),
    .B(_02209_),
    .Y(_02210_));
 sg13g2_xor2_1 _07506_ (.B(_02209_),
    .A(_02196_),
    .X(_02211_));
 sg13g2_o21ai_1 _07507_ (.B1(_02189_),
    .Y(_02212_),
    .A1(_02177_),
    .A2(_02190_));
 sg13g2_nand2_1 _07508_ (.Y(_02213_),
    .A(_02211_),
    .B(_02212_));
 sg13g2_xor2_1 _07509_ (.B(_02212_),
    .A(_02211_),
    .X(_02214_));
 sg13g2_a21oi_1 _07510_ (.A1(_02173_),
    .A2(_02175_),
    .Y(_02215_),
    .B1(_02193_));
 sg13g2_o21ai_1 _07511_ (.B1(_02214_),
    .Y(_02216_),
    .A1(_02194_),
    .A2(_02215_));
 sg13g2_or3_1 _07512_ (.A(_02194_),
    .B(_02214_),
    .C(_02215_),
    .X(_02217_));
 sg13g2_and2_1 _07513_ (.A(_02216_),
    .B(_02217_),
    .X(_00024_));
 sg13g2_nand2_1 _07514_ (.Y(_02218_),
    .A(_02213_),
    .B(_02216_));
 sg13g2_nand2_1 _07515_ (.Y(_02219_),
    .A(\i_core.cpu.i_core.i_shift.a[10] ),
    .B(_01581_));
 sg13g2_o21ai_1 _07516_ (.B1(_02205_),
    .Y(_02220_),
    .A1(_00867_),
    .A2(_02206_));
 sg13g2_o21ai_1 _07517_ (.B1(_02203_),
    .Y(_02221_),
    .A1(_02181_),
    .A2(_02201_));
 sg13g2_nand2_1 _07518_ (.Y(_02222_),
    .A(\i_core.cpu.i_core.i_shift.a[11] ),
    .B(net1237));
 sg13g2_nand2_1 _07519_ (.Y(_02223_),
    .A(\i_core.cpu.i_core.i_shift.a[9] ),
    .B(net1230));
 sg13g2_nand2_1 _07520_ (.Y(_02224_),
    .A(\i_core.cpu.i_core.i_shift.a[9] ),
    .B(net1232));
 sg13g2_xor2_1 _07521_ (.B(_02224_),
    .A(_02200_),
    .X(_02225_));
 sg13g2_nand2b_1 _07522_ (.Y(_02226_),
    .B(_02225_),
    .A_N(_02222_));
 sg13g2_xnor2_1 _07523_ (.Y(_02227_),
    .A(_02222_),
    .B(_02225_));
 sg13g2_nand2_1 _07524_ (.Y(_02228_),
    .A(_02221_),
    .B(_02227_));
 sg13g2_xnor2_1 _07525_ (.Y(_02229_),
    .A(_02221_),
    .B(_02227_));
 sg13g2_xnor2_1 _07526_ (.Y(_02230_),
    .A(_00868_),
    .B(_02229_));
 sg13g2_nand2b_1 _07527_ (.Y(_02231_),
    .B(_02220_),
    .A_N(_02230_));
 sg13g2_xor2_1 _07528_ (.B(_02230_),
    .A(_02220_),
    .X(_02232_));
 sg13g2_xor2_1 _07529_ (.B(_02232_),
    .A(_02219_),
    .X(_02233_));
 sg13g2_nor2_1 _07530_ (.A(_02208_),
    .B(_02210_),
    .Y(_02234_));
 sg13g2_nor3_1 _07531_ (.A(_02208_),
    .B(_02210_),
    .C(_02233_),
    .Y(_02235_));
 sg13g2_nor2b_1 _07532_ (.A(_02234_),
    .B_N(_02233_),
    .Y(_02236_));
 sg13g2_nor2_1 _07533_ (.A(_02235_),
    .B(_02236_),
    .Y(_02237_));
 sg13g2_xor2_1 _07534_ (.B(_02237_),
    .A(_02218_),
    .X(_00025_));
 sg13g2_nand2_1 _07535_ (.Y(_02238_),
    .A(\i_core.cpu.i_core.i_shift.a[11] ),
    .B(net1216));
 sg13g2_o21ai_1 _07536_ (.B1(_02228_),
    .Y(_02239_),
    .A1(_00868_),
    .A2(_02229_));
 sg13g2_o21ai_1 _07537_ (.B1(_02226_),
    .Y(_02240_),
    .A1(_02200_),
    .A2(_02224_));
 sg13g2_nand2_1 _07538_ (.Y(_02241_),
    .A(\i_core.cpu.i_core.i_shift.a[12] ),
    .B(net1237));
 sg13g2_nand2_1 _07539_ (.Y(_02242_),
    .A(\i_core.cpu.i_core.i_shift.a[10] ),
    .B(net1230));
 sg13g2_nand2_1 _07540_ (.Y(_02243_),
    .A(\i_core.cpu.i_core.i_shift.a[10] ),
    .B(net1232));
 sg13g2_xor2_1 _07541_ (.B(_02243_),
    .A(_02223_),
    .X(_02244_));
 sg13g2_nand2b_1 _07542_ (.Y(_02245_),
    .B(_02244_),
    .A_N(_02241_));
 sg13g2_xnor2_1 _07543_ (.Y(_02246_),
    .A(_02241_),
    .B(_02244_));
 sg13g2_nand2_1 _07544_ (.Y(_02247_),
    .A(_02240_),
    .B(_02246_));
 sg13g2_xnor2_1 _07545_ (.Y(_02248_),
    .A(_02240_),
    .B(_02246_));
 sg13g2_xnor2_1 _07546_ (.Y(_02249_),
    .A(_00869_),
    .B(_02248_));
 sg13g2_nand2b_1 _07547_ (.Y(_02250_),
    .B(_02239_),
    .A_N(_02249_));
 sg13g2_xor2_1 _07548_ (.B(_02249_),
    .A(_02239_),
    .X(_02251_));
 sg13g2_xor2_1 _07549_ (.B(_02251_),
    .A(_02238_),
    .X(_02252_));
 sg13g2_o21ai_1 _07550_ (.B1(_02231_),
    .Y(_02253_),
    .A1(_02219_),
    .A2(_02232_));
 sg13g2_and2_1 _07551_ (.A(_02252_),
    .B(_02253_),
    .X(_02254_));
 sg13g2_inv_1 _07552_ (.Y(_02255_),
    .A(_02254_));
 sg13g2_xor2_1 _07553_ (.B(_02253_),
    .A(_02252_),
    .X(_02256_));
 sg13g2_a21oi_1 _07554_ (.A1(_02213_),
    .A2(_02216_),
    .Y(_02257_),
    .B1(_02235_));
 sg13g2_o21ai_1 _07555_ (.B1(_02256_),
    .Y(_02258_),
    .A1(_02236_),
    .A2(_02257_));
 sg13g2_or3_1 _07556_ (.A(_02236_),
    .B(_02256_),
    .C(_02257_),
    .X(_02259_));
 sg13g2_and2_1 _07557_ (.A(_02258_),
    .B(_02259_),
    .X(_00026_));
 sg13g2_nand2_1 _07558_ (.Y(_02260_),
    .A(\i_core.cpu.i_core.i_shift.a[12] ),
    .B(net1216));
 sg13g2_o21ai_1 _07559_ (.B1(_02247_),
    .Y(_02261_),
    .A1(_00869_),
    .A2(_02248_));
 sg13g2_o21ai_1 _07560_ (.B1(_02245_),
    .Y(_02262_),
    .A1(_02223_),
    .A2(_02243_));
 sg13g2_nand2_1 _07561_ (.Y(_02263_),
    .A(\i_core.cpu.i_core.i_shift.a[13] ),
    .B(net1237));
 sg13g2_nand2_1 _07562_ (.Y(_02264_),
    .A(\i_core.cpu.i_core.i_shift.a[11] ),
    .B(net1230));
 sg13g2_nand2_1 _07563_ (.Y(_02265_),
    .A(\i_core.cpu.i_core.i_shift.a[11] ),
    .B(net1232));
 sg13g2_xor2_1 _07564_ (.B(_02265_),
    .A(_02242_),
    .X(_02266_));
 sg13g2_nand2b_1 _07565_ (.Y(_02267_),
    .B(_02266_),
    .A_N(_02263_));
 sg13g2_xnor2_1 _07566_ (.Y(_02268_),
    .A(_02263_),
    .B(_02266_));
 sg13g2_nand2_1 _07567_ (.Y(_02269_),
    .A(_02262_),
    .B(_02268_));
 sg13g2_xnor2_1 _07568_ (.Y(_02270_),
    .A(_02262_),
    .B(_02268_));
 sg13g2_xnor2_1 _07569_ (.Y(_02271_),
    .A(_00870_),
    .B(_02270_));
 sg13g2_nand2b_1 _07570_ (.Y(_02272_),
    .B(_02261_),
    .A_N(_02271_));
 sg13g2_xor2_1 _07571_ (.B(_02271_),
    .A(_02261_),
    .X(_02273_));
 sg13g2_xor2_1 _07572_ (.B(_02273_),
    .A(_02260_),
    .X(_02274_));
 sg13g2_o21ai_1 _07573_ (.B1(_02250_),
    .Y(_02275_),
    .A1(_02238_),
    .A2(_02251_));
 sg13g2_and2_1 _07574_ (.A(_02274_),
    .B(_02275_),
    .X(_02276_));
 sg13g2_xor2_1 _07575_ (.B(_02275_),
    .A(_02274_),
    .X(_02277_));
 sg13g2_inv_1 _07576_ (.Y(_02278_),
    .A(_02277_));
 sg13g2_a21oi_2 _07577_ (.B1(_02278_),
    .Y(_02279_),
    .A2(_02258_),
    .A1(_02255_));
 sg13g2_nand3_1 _07578_ (.B(_02258_),
    .C(_02278_),
    .A(_02255_),
    .Y(_02280_));
 sg13g2_nor2b_1 _07579_ (.A(_02279_),
    .B_N(_02280_),
    .Y(_00027_));
 sg13g2_nor2_1 _07580_ (.A(_02276_),
    .B(_02279_),
    .Y(_02281_));
 sg13g2_nand2_1 _07581_ (.Y(_02282_),
    .A(\i_core.cpu.i_core.i_shift.a[13] ),
    .B(net1216));
 sg13g2_o21ai_1 _07582_ (.B1(_02269_),
    .Y(_02283_),
    .A1(_00870_),
    .A2(_02270_));
 sg13g2_o21ai_1 _07583_ (.B1(_02267_),
    .Y(_02284_),
    .A1(_02242_),
    .A2(_02265_));
 sg13g2_nand2_1 _07584_ (.Y(_02285_),
    .A(\i_core.cpu.i_core.i_shift.a[14] ),
    .B(net1237));
 sg13g2_nand2_1 _07585_ (.Y(_02286_),
    .A(\i_core.cpu.i_core.i_shift.a[12] ),
    .B(net1230));
 sg13g2_nand2_1 _07586_ (.Y(_02287_),
    .A(\i_core.cpu.i_core.i_shift.a[12] ),
    .B(net1232));
 sg13g2_xor2_1 _07587_ (.B(_02287_),
    .A(_02264_),
    .X(_02288_));
 sg13g2_nand2b_1 _07588_ (.Y(_02289_),
    .B(_02288_),
    .A_N(_02285_));
 sg13g2_xnor2_1 _07589_ (.Y(_02290_),
    .A(_02285_),
    .B(_02288_));
 sg13g2_nand2_1 _07590_ (.Y(_02291_),
    .A(_02284_),
    .B(_02290_));
 sg13g2_xnor2_1 _07591_ (.Y(_02292_),
    .A(_02284_),
    .B(_02290_));
 sg13g2_xnor2_1 _07592_ (.Y(_02293_),
    .A(_00871_),
    .B(_02292_));
 sg13g2_nor2b_1 _07593_ (.A(_02293_),
    .B_N(_02283_),
    .Y(_02294_));
 sg13g2_xor2_1 _07594_ (.B(_02293_),
    .A(_02283_),
    .X(_02295_));
 sg13g2_nor2_1 _07595_ (.A(_02282_),
    .B(_02295_),
    .Y(_02296_));
 sg13g2_xor2_1 _07596_ (.B(_02295_),
    .A(_02282_),
    .X(_02297_));
 sg13g2_o21ai_1 _07597_ (.B1(_02272_),
    .Y(_02298_),
    .A1(_02260_),
    .A2(_02273_));
 sg13g2_nand2_1 _07598_ (.Y(_02299_),
    .A(_02297_),
    .B(_02298_));
 sg13g2_xor2_1 _07599_ (.B(_02298_),
    .A(_02297_),
    .X(_02300_));
 sg13g2_o21ai_1 _07600_ (.B1(_02300_),
    .Y(_02301_),
    .A1(_02276_),
    .A2(_02279_));
 sg13g2_xnor2_1 _07601_ (.Y(_00017_),
    .A(_02281_),
    .B(_02300_));
 sg13g2_nand2_1 _07602_ (.Y(_02302_),
    .A(\i_core.cpu.i_core.i_shift.a[14] ),
    .B(net1216));
 sg13g2_o21ai_1 _07603_ (.B1(_02291_),
    .Y(_02303_),
    .A1(_00871_),
    .A2(_02292_));
 sg13g2_o21ai_1 _07604_ (.B1(_02289_),
    .Y(_02304_),
    .A1(_02264_),
    .A2(_02287_));
 sg13g2_nand2_1 _07605_ (.Y(_02305_),
    .A(\i_core.cpu.i_core.i_shift.a[15] ),
    .B(net1237));
 sg13g2_nand2_1 _07606_ (.Y(_02306_),
    .A(\i_core.cpu.i_core.i_shift.a[13] ),
    .B(net1230));
 sg13g2_nand2_1 _07607_ (.Y(_02307_),
    .A(\i_core.cpu.i_core.i_shift.a[13] ),
    .B(net1232));
 sg13g2_xor2_1 _07608_ (.B(_02307_),
    .A(_02286_),
    .X(_02308_));
 sg13g2_nand2b_1 _07609_ (.Y(_02309_),
    .B(_02308_),
    .A_N(_02305_));
 sg13g2_xnor2_1 _07610_ (.Y(_02310_),
    .A(_02305_),
    .B(_02308_));
 sg13g2_nand2_1 _07611_ (.Y(_02311_),
    .A(_02304_),
    .B(_02310_));
 sg13g2_xnor2_1 _07612_ (.Y(_02312_),
    .A(_02304_),
    .B(_02310_));
 sg13g2_xnor2_1 _07613_ (.Y(_02313_),
    .A(_00872_),
    .B(_02312_));
 sg13g2_nand2b_1 _07614_ (.Y(_02314_),
    .B(_02303_),
    .A_N(_02313_));
 sg13g2_xor2_1 _07615_ (.B(_02313_),
    .A(_02303_),
    .X(_02315_));
 sg13g2_xor2_1 _07616_ (.B(_02315_),
    .A(_02302_),
    .X(_02316_));
 sg13g2_nor2_1 _07617_ (.A(_02294_),
    .B(_02296_),
    .Y(_02317_));
 sg13g2_nor3_1 _07618_ (.A(_02294_),
    .B(_02296_),
    .C(_02316_),
    .Y(_02318_));
 sg13g2_nor2b_1 _07619_ (.A(_02317_),
    .B_N(_02316_),
    .Y(_02319_));
 sg13g2_nor2_1 _07620_ (.A(_02318_),
    .B(_02319_),
    .Y(_02320_));
 sg13g2_nand2_1 _07621_ (.Y(_02321_),
    .A(_02299_),
    .B(_02301_));
 sg13g2_xor2_1 _07622_ (.B(_02321_),
    .A(_02320_),
    .X(_00018_));
 sg13g2_nand3_1 _07623_ (.B(\i_core.cpu.i_core.cycle[1] ),
    .C(net1278),
    .A(\i_core.cpu.data_ready_core ),
    .Y(_02322_));
 sg13g2_o21ai_1 _07624_ (.B1(_02322_),
    .Y(_00224_),
    .A1(_00789_),
    .A2(net1278));
 sg13g2_nand2_1 _07625_ (.Y(_02323_),
    .A(net1465),
    .B(_01183_));
 sg13g2_nor2_1 _07626_ (.A(net1308),
    .B(_01370_),
    .Y(_02324_));
 sg13g2_a21oi_1 _07627_ (.A1(net2418),
    .A2(net1308),
    .Y(_02325_),
    .B1(_02324_));
 sg13g2_nor2_1 _07628_ (.A(_02323_),
    .B(_02325_),
    .Y(_00225_));
 sg13g2_a21oi_1 _07629_ (.A1(net2418),
    .A2(net1310),
    .Y(_02326_),
    .B1(\i_core.cpu.i_core.cycle[1] ));
 sg13g2_nor2_1 _07630_ (.A(_02323_),
    .B(net2419),
    .Y(_00226_));
 sg13g2_nor2_2 _07631_ (.A(net1312),
    .B(_01735_),
    .Y(_02327_));
 sg13g2_nand2_2 _07632_ (.Y(_02328_),
    .A(net1278),
    .B(_01736_));
 sg13g2_nor2_2 _07633_ (.A(net2139),
    .B(_02328_),
    .Y(_02329_));
 sg13g2_nor2_1 _07634_ (.A(_01071_),
    .B(_01102_),
    .Y(_02330_));
 sg13g2_nand4_1 _07635_ (.B(_01013_),
    .C(_02329_),
    .A(_00974_),
    .Y(_02331_),
    .D(_02330_));
 sg13g2_a21oi_1 _07636_ (.A1(\i_core.cpu.i_core.mie[18] ),
    .A2(_01557_),
    .Y(_02332_),
    .B1(_01765_));
 sg13g2_a21oi_1 _07637_ (.A1(\i_core.cpu.i_core.mie[17] ),
    .A2(\i_core.cpu.i_core.mip[17] ),
    .Y(_02333_),
    .B1(_02332_));
 sg13g2_nand2_1 _07638_ (.Y(_02334_),
    .A(net2139),
    .B(_01763_));
 sg13g2_nor3_1 _07639_ (.A(_02328_),
    .B(_02333_),
    .C(_02334_),
    .Y(_02335_));
 sg13g2_a221oi_1 _07640_ (.B2(_01254_),
    .C1(_02335_),
    .B1(_02329_),
    .A1(net2605),
    .Y(_02336_),
    .A2(_02328_));
 sg13g2_a21oi_1 _07641_ (.A1(_02331_),
    .A2(_02336_),
    .Y(_00227_),
    .B1(net1384));
 sg13g2_nor2_1 _07642_ (.A(_00086_),
    .B(net1311),
    .Y(_02337_));
 sg13g2_nand2b_1 _07643_ (.Y(_02338_),
    .B(_01766_),
    .A_N(_01764_));
 sg13g2_o21ai_1 _07644_ (.B1(net1465),
    .Y(_02339_),
    .A1(net2383),
    .A2(_02327_));
 sg13g2_a21oi_1 _07645_ (.A1(_02337_),
    .A2(_02338_),
    .Y(_00228_),
    .B1(_02339_));
 sg13g2_nand2_1 _07646_ (.Y(_02340_),
    .A(net1966),
    .B(_02328_));
 sg13g2_a21oi_1 _07647_ (.A1(_02331_),
    .A2(_02340_),
    .Y(_00229_),
    .B1(net1384));
 sg13g2_o21ai_1 _07648_ (.B1(net1460),
    .Y(_02341_),
    .A1(net2416),
    .A2(_02327_));
 sg13g2_nor2_1 _07649_ (.A(_02329_),
    .B(_02341_),
    .Y(_00230_));
 sg13g2_nor3_2 _07650_ (.A(net2558),
    .B(net1311),
    .C(_01734_),
    .Y(_02342_));
 sg13g2_a21o_1 _07651_ (.A2(net1311),
    .A1(net2285),
    .B1(_02342_),
    .X(_00231_));
 sg13g2_o21ai_1 _07652_ (.B1(net2523),
    .Y(_02343_),
    .A1(\i_core.cpu.i_core.i_cycles.cy ),
    .A2(net1278));
 sg13g2_nor2_1 _07653_ (.A(_00823_),
    .B(_02343_),
    .Y(_02344_));
 sg13g2_and2_2 _07654_ (.A(net2487),
    .B(_02344_),
    .X(_02345_));
 sg13g2_nand2_2 _07655_ (.Y(_02346_),
    .A(net2413),
    .B(_02345_));
 sg13g2_nand3_1 _07656_ (.B(_01159_),
    .C(_02345_),
    .A(\i_core.cpu.i_core.cycle_count[3] ),
    .Y(_02347_));
 sg13g2_o21ai_1 _07657_ (.B1(net1460),
    .Y(_02348_),
    .A1(net1943),
    .A2(_02347_));
 sg13g2_a21oi_1 _07658_ (.A1(_00784_),
    .A2(_02347_),
    .Y(_00232_),
    .B1(net1944));
 sg13g2_nor3_2 _07659_ (.A(_00784_),
    .B(net1308),
    .C(_02346_),
    .Y(_02349_));
 sg13g2_o21ai_1 _07660_ (.B1(net1460),
    .Y(_02350_),
    .A1(net2128),
    .A2(_02349_));
 sg13g2_a21oi_1 _07661_ (.A1(net2128),
    .A2(_02349_),
    .Y(_00233_),
    .B1(_02350_));
 sg13g2_a21oi_1 _07662_ (.A1(\i_core.cpu.i_core.time_hi[1] ),
    .A2(_02349_),
    .Y(_02351_),
    .B1(net2007));
 sg13g2_and3_1 _07663_ (.X(_02352_),
    .A(net2007),
    .B(\i_core.cpu.i_core.time_hi[1] ),
    .C(_02349_));
 sg13g2_nor3_1 _07664_ (.A(net1384),
    .B(net2008),
    .C(_02352_),
    .Y(_00234_));
 sg13g2_nor3_2 _07665_ (.A(net1458),
    .B(net2285),
    .C(_02342_),
    .Y(_02353_));
 sg13g2_or3_2 _07666_ (.A(net1458),
    .B(net2285),
    .C(_02342_),
    .X(_02354_));
 sg13g2_nor4_2 _07667_ (.A(_00218_),
    .B(_00886_),
    .C(_01234_),
    .Y(_02355_),
    .D(_02354_));
 sg13g2_mux2_1 _07668_ (.A0(net2130),
    .A1(\i_core.cpu.i_core.interrupt_req[0] ),
    .S(_02355_),
    .X(_00235_));
 sg13g2_nand2_1 _07669_ (.Y(_02356_),
    .A(\i_core.cpu.i_core.interrupt_req[1] ),
    .B(_02355_));
 sg13g2_o21ai_1 _07670_ (.B1(_02356_),
    .Y(_00236_),
    .A1(_00841_),
    .A2(_02355_));
 sg13g2_nand2_1 _07671_ (.Y(_02357_),
    .A(net2556),
    .B(net1354));
 sg13g2_nand2_2 _07672_ (.Y(_02358_),
    .A(net1465),
    .B(net1353));
 sg13g2_nor2_1 _07673_ (.A(_01166_),
    .B(_01178_),
    .Y(_02359_));
 sg13g2_nand2_1 _07674_ (.Y(_02360_),
    .A(net1307),
    .B(_01177_));
 sg13g2_nor2_2 _07675_ (.A(_01255_),
    .B(_02360_),
    .Y(_02361_));
 sg13g2_nand2b_1 _07676_ (.Y(_02362_),
    .B(_02361_),
    .A_N(_01090_));
 sg13g2_nor2_1 _07677_ (.A(\i_core.cpu.i_core.mepc[0] ),
    .B(_02361_),
    .Y(_02363_));
 sg13g2_nor2_1 _07678_ (.A(_01736_),
    .B(_02363_),
    .Y(_02364_));
 sg13g2_a22oi_1 _07679_ (.Y(_02365_),
    .B1(_02362_),
    .B2(_02364_),
    .A2(_01736_),
    .A1(_01095_));
 sg13g2_o21ai_1 _07680_ (.B1(_02357_),
    .Y(_00237_),
    .A1(_02358_),
    .A2(_02365_));
 sg13g2_mux2_1 _07681_ (.A0(\i_core.cpu.i_core.mepc[1] ),
    .A1(_01051_),
    .S(_02361_),
    .X(_02366_));
 sg13g2_a21oi_1 _07682_ (.A1(_01038_),
    .A2(_01736_),
    .Y(_02367_),
    .B1(_02358_));
 sg13g2_o21ai_1 _07683_ (.B1(_02367_),
    .Y(_02368_),
    .A1(_01736_),
    .A2(_02366_));
 sg13g2_o21ai_1 _07684_ (.B1(_02368_),
    .Y(_00238_),
    .A1(_00842_),
    .A2(net1352));
 sg13g2_nand2_1 _07685_ (.Y(_02369_),
    .A(net2259),
    .B(net1354));
 sg13g2_nor2_1 _07686_ (.A(_00986_),
    .B(_01735_),
    .Y(_02370_));
 sg13g2_mux2_1 _07687_ (.A0(\i_core.cpu.i_core.mepc[2] ),
    .A1(_01003_),
    .S(_02361_),
    .X(_02371_));
 sg13g2_a21oi_1 _07688_ (.A1(_01735_),
    .A2(_02371_),
    .Y(_02372_),
    .B1(_02370_));
 sg13g2_o21ai_1 _07689_ (.B1(_02369_),
    .Y(_00239_),
    .A1(_02358_),
    .A2(_02372_));
 sg13g2_mux2_1 _07690_ (.A0(\i_core.cpu.i_core.mepc[3] ),
    .A1(_00926_),
    .S(_02361_),
    .X(_02373_));
 sg13g2_a21oi_1 _07691_ (.A1(_00888_),
    .A2(_01736_),
    .Y(_02374_),
    .B1(_02358_));
 sg13g2_o21ai_1 _07692_ (.B1(_02374_),
    .Y(_02375_),
    .A1(_01736_),
    .A2(_02373_));
 sg13g2_o21ai_1 _07693_ (.B1(_02375_),
    .Y(_00240_),
    .A1(_00843_),
    .A2(net1353));
 sg13g2_a21oi_1 _07694_ (.A1(net1402),
    .A2(_00927_),
    .Y(_02376_),
    .B1(_01232_));
 sg13g2_nand3_1 _07695_ (.B(_01985_),
    .C(_02376_),
    .A(net1300),
    .Y(_02377_));
 sg13g2_nand2_1 _07696_ (.Y(_02378_),
    .A(_02328_),
    .B(_02377_));
 sg13g2_and2_1 _07697_ (.A(\i_core.cpu.i_core.mstatus_mie ),
    .B(_02327_),
    .X(_02379_));
 sg13g2_a21oi_2 _07698_ (.B1(_01232_),
    .Y(_02380_),
    .A2(\i_core.cpu.alu_op[0] ),
    .A1(net1402));
 sg13g2_and2_1 _07699_ (.A(_00926_),
    .B(_02380_),
    .X(_02381_));
 sg13g2_a21oi_1 _07700_ (.A1(_02328_),
    .A2(_02381_),
    .Y(_02382_),
    .B1(_02379_));
 sg13g2_o21ai_1 _07701_ (.B1(_02353_),
    .Y(_02383_),
    .A1(net2361),
    .A2(_02378_));
 sg13g2_a21oi_1 _07702_ (.A1(_02378_),
    .A2(_02382_),
    .Y(_00241_),
    .B1(net2362));
 sg13g2_nand2_1 _07703_ (.Y(_02384_),
    .A(\i_core.cpu.i_core.mstatus_mie ),
    .B(net1300));
 sg13g2_a21oi_1 _07704_ (.A1(_01992_),
    .A2(_02376_),
    .Y(_02385_),
    .B1(_02384_));
 sg13g2_a221oi_1 _07705_ (.B2(_02381_),
    .C1(_02385_),
    .B1(_01992_),
    .A1(net2361),
    .Y(_02386_),
    .A2(net1276));
 sg13g2_o21ai_1 _07706_ (.B1(_02353_),
    .Y(_00242_),
    .A1(_02327_),
    .A2(_02386_));
 sg13g2_nor2_1 _07707_ (.A(net2440),
    .B(net1276),
    .Y(_02387_));
 sg13g2_o21ai_1 _07708_ (.B1(_02353_),
    .Y(_00243_),
    .A1(_02327_),
    .A2(_02387_));
 sg13g2_nand2b_1 _07709_ (.Y(_02388_),
    .B(net1176),
    .A_N(_01774_));
 sg13g2_and2_2 _07710_ (.A(_01771_),
    .B(_02388_),
    .X(_02389_));
 sg13g2_nor2_2 _07711_ (.A(net1187),
    .B(_02389_),
    .Y(_02390_));
 sg13g2_nor2_2 _07712_ (.A(net1458),
    .B(_02390_),
    .Y(_02391_));
 sg13g2_nor2_1 _07713_ (.A(\i_core.cpu.i_core.i_registers.rd[0] ),
    .B(net1155),
    .Y(_02392_));
 sg13g2_nand2_1 _07714_ (.Y(_02393_),
    .A(_01753_),
    .B(net1248));
 sg13g2_nand2b_2 _07715_ (.Y(_02394_),
    .B(_01778_),
    .A_N(_01802_));
 sg13g2_nor2_2 _07716_ (.A(_01801_),
    .B(_02394_),
    .Y(_02395_));
 sg13g2_or2_2 _07717_ (.X(_02396_),
    .B(_02394_),
    .A(_01801_));
 sg13g2_nand2_1 _07718_ (.Y(_02397_),
    .A(_01778_),
    .B(_01802_));
 sg13g2_nand3_1 _07719_ (.B(_01779_),
    .C(_01802_),
    .A(_01778_),
    .Y(_02398_));
 sg13g2_nor2b_2 _07720_ (.A(_01746_),
    .B_N(_01802_),
    .Y(_02399_));
 sg13g2_and2_2 _07721_ (.A(_01751_),
    .B(_02399_),
    .X(_02400_));
 sg13g2_nand2_1 _07722_ (.Y(_02401_),
    .A(_01800_),
    .B(_02399_));
 sg13g2_nand2_1 _07723_ (.Y(_02402_),
    .A(_01800_),
    .B(_02400_));
 sg13g2_and2_2 _07724_ (.A(_02398_),
    .B(_02402_),
    .X(_02403_));
 sg13g2_nand2_2 _07725_ (.Y(_02404_),
    .A(_01780_),
    .B(_01782_));
 sg13g2_nor2_2 _07726_ (.A(_02397_),
    .B(_02404_),
    .Y(_02405_));
 sg13g2_or2_2 _07727_ (.X(_02406_),
    .B(_02404_),
    .A(_02397_));
 sg13g2_nand2_1 _07728_ (.Y(_02407_),
    .A(_01783_),
    .B(_01804_));
 sg13g2_and2_2 _07729_ (.A(_01782_),
    .B(_02400_),
    .X(_02408_));
 sg13g2_a21oi_1 _07730_ (.A1(_01783_),
    .A2(_01804_),
    .Y(_02409_),
    .B1(_02408_));
 sg13g2_and3_1 _07731_ (.X(_02410_),
    .A(_02403_),
    .B(_02406_),
    .C(_02409_));
 sg13g2_o21ai_1 _07732_ (.B1(_02410_),
    .Y(_02411_),
    .A1(_01806_),
    .A2(_01810_));
 sg13g2_nor2_1 _07733_ (.A(_02395_),
    .B(_02411_),
    .Y(_02412_));
 sg13g2_nor2_1 _07734_ (.A(net1248),
    .B(_02412_),
    .Y(_02413_));
 sg13g2_nor2_1 _07735_ (.A(_01805_),
    .B(_02400_),
    .Y(_02414_));
 sg13g2_and3_2 _07736_ (.X(_02415_),
    .A(_01784_),
    .B(_02410_),
    .C(_02414_));
 sg13g2_nand2_1 _07737_ (.Y(_02416_),
    .A(_01783_),
    .B(_02400_));
 sg13g2_nand2_1 _07738_ (.Y(_02417_),
    .A(_01805_),
    .B(_01828_));
 sg13g2_a21oi_1 _07739_ (.A1(net1252),
    .A2(_02415_),
    .Y(_02418_),
    .B1(_01753_));
 sg13g2_a22oi_1 _07740_ (.Y(_02419_),
    .B1(_01811_),
    .B2(_01828_),
    .A2(_01802_),
    .A1(_01785_));
 sg13g2_nand3_1 _07741_ (.B(_02418_),
    .C(_02419_),
    .A(_02416_),
    .Y(_02420_));
 sg13g2_a21oi_2 _07742_ (.B1(_02413_),
    .Y(_02421_),
    .A2(_02420_),
    .A1(_02393_));
 sg13g2_nor2_1 _07743_ (.A(net1186),
    .B(_02421_),
    .Y(_02422_));
 sg13g2_a21oi_1 _07744_ (.A1(net1925),
    .A2(net1186),
    .Y(_02423_),
    .B1(_02422_));
 sg13g2_a21oi_1 _07745_ (.A1(net1155),
    .A2(_02423_),
    .Y(_00244_),
    .B1(_02392_));
 sg13g2_nand3_1 _07746_ (.B(_01999_),
    .C(_02001_),
    .A(net1186),
    .Y(_02424_));
 sg13g2_a21o_1 _07747_ (.A2(_02412_),
    .A1(net1198),
    .B1(net1249),
    .X(_02425_));
 sg13g2_nand2_1 _07748_ (.Y(_02426_),
    .A(net1197),
    .B(net1250));
 sg13g2_nand3_1 _07749_ (.B(net1250),
    .C(_02415_),
    .A(net1198),
    .Y(_02427_));
 sg13g2_nand3_1 _07750_ (.B(_02425_),
    .C(_02427_),
    .A(net1185),
    .Y(_02428_));
 sg13g2_nand3_1 _07751_ (.B(_02424_),
    .C(_02428_),
    .A(net1155),
    .Y(_02429_));
 sg13g2_o21ai_1 _07752_ (.B1(_02429_),
    .Y(_00245_),
    .A1(_00830_),
    .A2(net1155));
 sg13g2_xor2_1 _07753_ (.B(_01507_),
    .A(\i_core.cpu.i_core.i_registers.rd[2] ),
    .X(_02430_));
 sg13g2_a21o_1 _07754_ (.A2(_02412_),
    .A1(net1198),
    .B1(_01819_),
    .X(_02431_));
 sg13g2_nor2_1 _07755_ (.A(net1200),
    .B(_01790_),
    .Y(_02432_));
 sg13g2_a21oi_2 _07756_ (.B1(net1187),
    .Y(_02433_),
    .A2(_02432_),
    .A1(_02415_));
 sg13g2_a22oi_1 _07757_ (.Y(_02434_),
    .B1(_02431_),
    .B2(_02433_),
    .A2(_02430_),
    .A1(net1186));
 sg13g2_mux2_1 _07758_ (.A0(net2635),
    .A1(_02434_),
    .S(net1155),
    .X(_00246_));
 sg13g2_xor2_1 _07759_ (.B(_02010_),
    .A(\i_core.cpu.i_core.i_registers.rd[3] ),
    .X(_02435_));
 sg13g2_nand3b_1 _07760_ (.B(net1184),
    .C(net1197),
    .Y(_02436_),
    .A_N(_02411_));
 sg13g2_o21ai_1 _07761_ (.B1(net1197),
    .Y(_02437_),
    .A1(_02395_),
    .A2(_02415_));
 sg13g2_a21oi_2 _07762_ (.B1(net1187),
    .Y(_02438_),
    .A2(_02436_),
    .A1(_01818_));
 sg13g2_a22oi_1 _07763_ (.Y(_02439_),
    .B1(_02437_),
    .B2(_02438_),
    .A2(_02435_),
    .A1(net1186));
 sg13g2_mux2_1 _07764_ (.A0(net2645),
    .A1(_02439_),
    .S(net1155),
    .X(_00247_));
 sg13g2_nor2b_1 _07765_ (.A(net1409),
    .B_N(\i_core.cpu.i_core.mem_op[0] ),
    .Y(_02440_));
 sg13g2_and2_1 _07766_ (.A(net2583),
    .B(net1312),
    .X(_02441_));
 sg13g2_nor4_1 _07767_ (.A(\i_core.cpu.i_core.mem_op[1] ),
    .B(net2287),
    .C(_01196_),
    .D(_02440_),
    .Y(_02442_));
 sg13g2_nand4_1 _07768_ (.B(_00084_),
    .C(_01496_),
    .A(net1414),
    .Y(_02443_),
    .D(_02442_));
 sg13g2_mux2_1 _07769_ (.A0(_01963_),
    .A1(_02441_),
    .S(_02443_),
    .X(_00248_));
 sg13g2_nand3_1 _07770_ (.B(net1235),
    .C(_01883_),
    .A(_01461_),
    .Y(_02444_));
 sg13g2_nor2_1 _07771_ (.A(\data_to_write[0] ),
    .B(net1208),
    .Y(_02445_));
 sg13g2_nand2_1 _07772_ (.Y(_02446_),
    .A(net1968),
    .B(\i_uart_tx.cycle_counter[0] ));
 sg13g2_or2_1 _07773_ (.X(_02447_),
    .B(_02446_),
    .A(\i_uart_tx.cycle_counter[2] ));
 sg13g2_nor2_1 _07774_ (.A(\i_uart_tx.cycle_counter[6] ),
    .B(\i_uart_tx.cycle_counter[4] ),
    .Y(_02448_));
 sg13g2_nor4_1 _07775_ (.A(\i_uart_tx.cycle_counter[10] ),
    .B(_00782_),
    .C(\i_uart_tx.cycle_counter[8] ),
    .D(\i_uart_tx.cycle_counter[7] ),
    .Y(_02449_));
 sg13g2_nand4_1 _07776_ (.B(net2329),
    .C(_02448_),
    .A(net2345),
    .Y(_02450_),
    .D(_02449_));
 sg13g2_nor2_2 _07777_ (.A(_02447_),
    .B(_02450_),
    .Y(_02451_));
 sg13g2_o21ai_1 _07778_ (.B1(\i_uart_tx.fsm_state[3] ),
    .Y(_02452_),
    .A1(net2365),
    .A2(\i_uart_tx.fsm_state[1] ));
 sg13g2_nor2_1 _07779_ (.A(_00782_),
    .B(\i_uart_tx.cycle_counter[7] ),
    .Y(_02453_));
 sg13g2_nand4_1 _07780_ (.B(\i_uart_tx.cycle_counter[3] ),
    .C(_02448_),
    .A(\i_uart_tx.cycle_counter[5] ),
    .Y(_02454_),
    .D(_02453_));
 sg13g2_nor4_1 _07781_ (.A(\i_uart_tx.cycle_counter[10] ),
    .B(\i_uart_tx.cycle_counter[8] ),
    .C(_02447_),
    .D(_02454_),
    .Y(_02455_));
 sg13g2_nand3_1 _07782_ (.B(_02452_),
    .C(_02455_),
    .A(_01460_),
    .Y(_02456_));
 sg13g2_mux2_1 _07783_ (.A0(net2592),
    .A1(net2386),
    .S(_02456_),
    .X(_02457_));
 sg13g2_nor2b_1 _07784_ (.A(_02457_),
    .B_N(net1208),
    .Y(_02458_));
 sg13g2_nor3_1 _07785_ (.A(net1315),
    .B(_02445_),
    .C(_02458_),
    .Y(_00249_));
 sg13g2_nor2_1 _07786_ (.A(\data_to_write[1] ),
    .B(net1208),
    .Y(_02459_));
 sg13g2_mux2_1 _07787_ (.A0(net2581),
    .A1(\i_uart_tx.data_to_send[1] ),
    .S(_02456_),
    .X(_02460_));
 sg13g2_nor2b_1 _07788_ (.A(net2582),
    .B_N(net1208),
    .Y(_02461_));
 sg13g2_nor3_1 _07789_ (.A(net1314),
    .B(_02459_),
    .C(_02461_),
    .Y(_00250_));
 sg13g2_nor2_1 _07790_ (.A(net2684),
    .B(net1207),
    .Y(_02462_));
 sg13g2_mux2_1 _07791_ (.A0(net2634),
    .A1(net2581),
    .S(_02456_),
    .X(_02463_));
 sg13g2_nor2b_1 _07792_ (.A(_02463_),
    .B_N(net1206),
    .Y(_02464_));
 sg13g2_nor3_1 _07793_ (.A(net1315),
    .B(_02462_),
    .C(_02464_),
    .Y(_00251_));
 sg13g2_nor2_1 _07794_ (.A(\data_to_write[3] ),
    .B(net1207),
    .Y(_02465_));
 sg13g2_mux2_1 _07795_ (.A0(net2607),
    .A1(\i_uart_tx.data_to_send[3] ),
    .S(_02456_),
    .X(_02466_));
 sg13g2_nor2b_1 _07796_ (.A(net2608),
    .B_N(net1206),
    .Y(_02467_));
 sg13g2_nor3_1 _07797_ (.A(net1315),
    .B(_02465_),
    .C(_02467_),
    .Y(_00252_));
 sg13g2_nor2_1 _07798_ (.A(net2622),
    .B(net1207),
    .Y(_02468_));
 sg13g2_mux2_1 _07799_ (.A0(net2610),
    .A1(net2607),
    .S(_02456_),
    .X(_02469_));
 sg13g2_nor2b_1 _07800_ (.A(_02469_),
    .B_N(net1207),
    .Y(_02470_));
 sg13g2_nor3_1 _07801_ (.A(net1314),
    .B(_02468_),
    .C(_02470_),
    .Y(_00253_));
 sg13g2_nor2_1 _07802_ (.A(\data_to_write[5] ),
    .B(net1206),
    .Y(_02471_));
 sg13g2_mux2_1 _07803_ (.A0(net2602),
    .A1(net2610),
    .S(_02456_),
    .X(_02472_));
 sg13g2_nor2b_1 _07804_ (.A(_02472_),
    .B_N(net1206),
    .Y(_02473_));
 sg13g2_nor3_1 _07805_ (.A(net1314),
    .B(_02471_),
    .C(_02473_),
    .Y(_00254_));
 sg13g2_nor2_1 _07806_ (.A(\data_to_write[6] ),
    .B(net1206),
    .Y(_02474_));
 sg13g2_mux2_1 _07807_ (.A0(net1914),
    .A1(net2602),
    .S(_02456_),
    .X(_02475_));
 sg13g2_nor2b_1 _07808_ (.A(_02475_),
    .B_N(net1206),
    .Y(_02476_));
 sg13g2_nor3_1 _07809_ (.A(net1314),
    .B(_02474_),
    .C(_02476_),
    .Y(_00255_));
 sg13g2_nand2_1 _07810_ (.Y(_02477_),
    .A(net1914),
    .B(_02456_));
 sg13g2_o21ai_1 _07811_ (.B1(net1321),
    .Y(_02478_),
    .A1(_00844_),
    .A2(net1206));
 sg13g2_a21oi_1 _07812_ (.A1(net1206),
    .A2(_02477_),
    .Y(_00256_),
    .B1(_02478_));
 sg13g2_or2_1 _07813_ (.X(_02479_),
    .B(_02451_),
    .A(net1319));
 sg13g2_and2_1 _07814_ (.A(net1980),
    .B(_01462_),
    .X(_02480_));
 sg13g2_a21oi_1 _07815_ (.A1(\i_uart_tx.cycle_counter[0] ),
    .A2(_01461_),
    .Y(_02481_),
    .B1(_02480_));
 sg13g2_nor2_1 _07816_ (.A(_02479_),
    .B(net1981),
    .Y(_00257_));
 sg13g2_a21oi_1 _07817_ (.A1(\i_uart_tx.cycle_counter[0] ),
    .A2(_01462_),
    .Y(_02482_),
    .B1(net1968));
 sg13g2_nor2_1 _07818_ (.A(_01461_),
    .B(_02446_),
    .Y(_02483_));
 sg13g2_nor3_1 _07819_ (.A(_02479_),
    .B(net1969),
    .C(_02483_),
    .Y(_00258_));
 sg13g2_nor2_1 _07820_ (.A(net2219),
    .B(_02483_),
    .Y(_02484_));
 sg13g2_and2_1 _07821_ (.A(net2219),
    .B(_02483_),
    .X(_02485_));
 sg13g2_nor3_1 _07822_ (.A(_02479_),
    .B(net2220),
    .C(_02485_),
    .Y(_00259_));
 sg13g2_nor2_1 _07823_ (.A(net2329),
    .B(_02485_),
    .Y(_02486_));
 sg13g2_and2_1 _07824_ (.A(net2329),
    .B(_02485_),
    .X(_02487_));
 sg13g2_nor3_1 _07825_ (.A(net1229),
    .B(_02486_),
    .C(_02487_),
    .Y(_00260_));
 sg13g2_nor2_1 _07826_ (.A(net2334),
    .B(_02487_),
    .Y(_02488_));
 sg13g2_and2_1 _07827_ (.A(net2334),
    .B(_02487_),
    .X(_02489_));
 sg13g2_nor3_1 _07828_ (.A(net1229),
    .B(_02488_),
    .C(_02489_),
    .Y(_00261_));
 sg13g2_nor2_1 _07829_ (.A(net2345),
    .B(_02489_),
    .Y(_02490_));
 sg13g2_and2_1 _07830_ (.A(net2345),
    .B(_02489_),
    .X(_02491_));
 sg13g2_nor3_1 _07831_ (.A(net1229),
    .B(_02490_),
    .C(_02491_),
    .Y(_00262_));
 sg13g2_xnor2_1 _07832_ (.Y(_02492_),
    .A(net2359),
    .B(_02491_));
 sg13g2_nor2_1 _07833_ (.A(net1229),
    .B(_02492_),
    .Y(_00263_));
 sg13g2_a21oi_1 _07834_ (.A1(\i_uart_tx.cycle_counter[6] ),
    .A2(_02491_),
    .Y(_02493_),
    .B1(net2103));
 sg13g2_and3_1 _07835_ (.X(_02494_),
    .A(net2103),
    .B(\i_uart_tx.cycle_counter[6] ),
    .C(_02491_));
 sg13g2_nor3_1 _07836_ (.A(net1229),
    .B(net2104),
    .C(_02494_),
    .Y(_00264_));
 sg13g2_nor2_1 _07837_ (.A(net2343),
    .B(_02494_),
    .Y(_02495_));
 sg13g2_and2_1 _07838_ (.A(net2343),
    .B(_02494_),
    .X(_02496_));
 sg13g2_nor3_1 _07839_ (.A(net1229),
    .B(net2344),
    .C(_02496_),
    .Y(_00265_));
 sg13g2_nor2_1 _07840_ (.A(net2276),
    .B(_02496_),
    .Y(_02497_));
 sg13g2_and2_1 _07841_ (.A(net2276),
    .B(_02496_),
    .X(_02498_));
 sg13g2_nor3_1 _07842_ (.A(net1229),
    .B(net2277),
    .C(_02498_),
    .Y(_00266_));
 sg13g2_a21oi_1 _07843_ (.A1(net2481),
    .A2(_02498_),
    .Y(_02499_),
    .B1(net1229));
 sg13g2_o21ai_1 _07844_ (.B1(_02499_),
    .Y(_02500_),
    .A1(net2481),
    .A2(_02498_));
 sg13g2_inv_1 _07845_ (.Y(_00267_),
    .A(_02500_));
 sg13g2_o21ai_1 _07846_ (.B1(net2549),
    .Y(_02501_),
    .A1(_02447_),
    .A2(_02450_));
 sg13g2_nor2_1 _07847_ (.A(_01461_),
    .B(_02451_),
    .Y(_02502_));
 sg13g2_nor2_1 _07848_ (.A(\i_uart_tx.fsm_state[2] ),
    .B(\i_uart_tx.fsm_state[0] ),
    .Y(_02503_));
 sg13g2_nand3_1 _07849_ (.B(\i_uart_tx.fsm_state[1] ),
    .C(_02503_),
    .A(net2518),
    .Y(_02504_));
 sg13g2_nor2b_1 _07850_ (.A(\i_uart_tx.fsm_state[0] ),
    .B_N(_02504_),
    .Y(_02505_));
 sg13g2_nand2_1 _07851_ (.Y(_02506_),
    .A(_01460_),
    .B(_02505_));
 sg13g2_a21o_1 _07852_ (.A2(_02506_),
    .A1(net1208),
    .B1(_02502_),
    .X(_02507_));
 sg13g2_a21oi_1 _07853_ (.A1(_02501_),
    .A2(_02507_),
    .Y(_00268_),
    .B1(net1314));
 sg13g2_nor2_1 _07854_ (.A(_02502_),
    .B(_02505_),
    .Y(_02508_));
 sg13g2_o21ai_1 _07855_ (.B1(net1321),
    .Y(_02509_),
    .A1(net2397),
    .A2(_02508_));
 sg13g2_a21oi_1 _07856_ (.A1(net2397),
    .A2(_02508_),
    .Y(_00269_),
    .B1(_02509_));
 sg13g2_and2_1 _07857_ (.A(\i_uart_tx.fsm_state[1] ),
    .B(\i_uart_tx.fsm_state[0] ),
    .X(_02510_));
 sg13g2_a21oi_1 _07858_ (.A1(_02451_),
    .A2(_02510_),
    .Y(_02511_),
    .B1(net2365));
 sg13g2_and4_1 _07859_ (.A(net2365),
    .B(net2397),
    .C(\i_uart_tx.fsm_state[0] ),
    .D(_02451_),
    .X(_02512_));
 sg13g2_nor3_1 _07860_ (.A(net1314),
    .B(net2366),
    .C(_02512_),
    .Y(_00270_));
 sg13g2_nand3_1 _07861_ (.B(net2365),
    .C(_02510_),
    .A(net2518),
    .Y(_02513_));
 sg13g2_a21oi_1 _07862_ (.A1(_02504_),
    .A2(_02513_),
    .Y(_02514_),
    .B1(_02502_));
 sg13g2_o21ai_1 _07863_ (.B1(net1321),
    .Y(_02515_),
    .A1(net2518),
    .A2(_02512_));
 sg13g2_nor2_1 _07864_ (.A(_02514_),
    .B(_02515_),
    .Y(_00271_));
 sg13g2_nand2_1 _07865_ (.Y(_02516_),
    .A(\i_uart_rx.cycle_counter[9] ),
    .B(_00815_));
 sg13g2_and2_1 _07866_ (.A(\i_uart_rx.cycle_counter[0] ),
    .B(net2094),
    .X(_02517_));
 sg13g2_nor3_2 _07867_ (.A(net2569),
    .B(net2512),
    .C(net2575),
    .Y(_02518_));
 sg13g2_o21ai_1 _07868_ (.B1(\i_uart_rx.fsm_state[3] ),
    .Y(_02519_),
    .A1(\i_uart_rx.fsm_state[2] ),
    .A2(\i_uart_rx.fsm_state[1] ));
 sg13g2_or4_1 _07869_ (.A(\i_uart_rx.cycle_counter[2] ),
    .B(\i_uart_rx.cycle_counter[4] ),
    .C(\i_uart_rx.cycle_counter[7] ),
    .D(\i_uart_rx.cycle_counter[6] ),
    .X(_02520_));
 sg13g2_nand3_1 _07870_ (.B(\i_uart_rx.cycle_counter[5] ),
    .C(_02517_),
    .A(\i_uart_rx.cycle_counter[3] ),
    .Y(_02521_));
 sg13g2_nor4_2 _07871_ (.A(\i_uart_rx.cycle_counter[10] ),
    .B(_02516_),
    .C(_02520_),
    .Y(_02522_),
    .D(_02521_));
 sg13g2_inv_1 _07872_ (.Y(_02523_),
    .A(_02522_));
 sg13g2_nand3b_1 _07873_ (.B(_02519_),
    .C(_02522_),
    .Y(_02524_),
    .A_N(_02518_));
 sg13g2_mux2_1 _07874_ (.A0(\i_uart_rx.recieved_data[1] ),
    .A1(net2164),
    .S(_02524_),
    .X(_00272_));
 sg13g2_mux2_1 _07875_ (.A0(net2248),
    .A1(\i_uart_rx.recieved_data[1] ),
    .S(_02524_),
    .X(_00273_));
 sg13g2_mux2_1 _07876_ (.A0(net2263),
    .A1(net2248),
    .S(_02524_),
    .X(_00274_));
 sg13g2_mux2_1 _07877_ (.A0(net2309),
    .A1(net2263),
    .S(_02524_),
    .X(_00275_));
 sg13g2_mux2_1 _07878_ (.A0(net2226),
    .A1(\i_uart_rx.recieved_data[4] ),
    .S(_02524_),
    .X(_00276_));
 sg13g2_mux2_1 _07879_ (.A0(net2252),
    .A1(net2226),
    .S(_02524_),
    .X(_00277_));
 sg13g2_mux2_1 _07880_ (.A0(net2264),
    .A1(net2252),
    .S(_02524_),
    .X(_00278_));
 sg13g2_mux2_1 _07881_ (.A0(net2026),
    .A1(\i_uart_rx.recieved_data[7] ),
    .S(_02524_),
    .X(_00279_));
 sg13g2_nor2b_2 _07882_ (.A(net2472),
    .B_N(_02518_),
    .Y(_02525_));
 sg13g2_nor2_2 _07883_ (.A(_02522_),
    .B(_02525_),
    .Y(_02526_));
 sg13g2_nor2_1 _07884_ (.A(net1319),
    .B(_01557_),
    .Y(_02527_));
 sg13g2_nand2_1 _07885_ (.Y(_02528_),
    .A(_02526_),
    .B(_02527_));
 sg13g2_and3_1 _07886_ (.X(_00280_),
    .A(net1816),
    .B(_02526_),
    .C(_02527_));
 sg13g2_nor2_1 _07887_ (.A(\i_uart_rx.cycle_counter[0] ),
    .B(net2094),
    .Y(_02529_));
 sg13g2_nor3_1 _07888_ (.A(_02517_),
    .B(_02528_),
    .C(net2095),
    .Y(_00281_));
 sg13g2_nor2_1 _07889_ (.A(net2332),
    .B(_02517_),
    .Y(_02530_));
 sg13g2_and2_1 _07890_ (.A(net2332),
    .B(_02517_),
    .X(_02531_));
 sg13g2_nor3_1 _07891_ (.A(_02528_),
    .B(net2333),
    .C(_02531_),
    .Y(_00282_));
 sg13g2_nor2_1 _07892_ (.A(net2323),
    .B(_02531_),
    .Y(_02532_));
 sg13g2_and2_1 _07893_ (.A(net2323),
    .B(_02531_),
    .X(_02533_));
 sg13g2_nor3_1 _07894_ (.A(net1228),
    .B(net2324),
    .C(_02533_),
    .Y(_00283_));
 sg13g2_nor2_1 _07895_ (.A(net2281),
    .B(_02533_),
    .Y(_02534_));
 sg13g2_and2_1 _07896_ (.A(net2281),
    .B(_02533_),
    .X(_02535_));
 sg13g2_nor3_1 _07897_ (.A(net1228),
    .B(net2282),
    .C(_02535_),
    .Y(_00284_));
 sg13g2_nor2_1 _07898_ (.A(net2369),
    .B(_02535_),
    .Y(_02536_));
 sg13g2_and2_1 _07899_ (.A(net2369),
    .B(_02535_),
    .X(_02537_));
 sg13g2_nor3_1 _07900_ (.A(net1228),
    .B(_02536_),
    .C(_02537_),
    .Y(_00285_));
 sg13g2_nor2_1 _07901_ (.A(net2357),
    .B(_02537_),
    .Y(_02538_));
 sg13g2_and2_1 _07902_ (.A(net2357),
    .B(_02537_),
    .X(_02539_));
 sg13g2_nor3_1 _07903_ (.A(net1228),
    .B(net2358),
    .C(_02539_),
    .Y(_00286_));
 sg13g2_nor2_1 _07904_ (.A(net2389),
    .B(_02539_),
    .Y(_02540_));
 sg13g2_and2_1 _07905_ (.A(net2389),
    .B(_02539_),
    .X(_02541_));
 sg13g2_nor3_1 _07906_ (.A(net1228),
    .B(_02540_),
    .C(_02541_),
    .Y(_00287_));
 sg13g2_nor2_1 _07907_ (.A(net2303),
    .B(_02541_),
    .Y(_02542_));
 sg13g2_and2_1 _07908_ (.A(net2303),
    .B(_02541_),
    .X(_02543_));
 sg13g2_nor3_1 _07909_ (.A(net1228),
    .B(net2304),
    .C(_02543_),
    .Y(_00288_));
 sg13g2_nor2_1 _07910_ (.A(net2379),
    .B(_02543_),
    .Y(_02544_));
 sg13g2_and2_1 _07911_ (.A(net2379),
    .B(_02543_),
    .X(_02545_));
 sg13g2_nor3_1 _07912_ (.A(net1228),
    .B(_02544_),
    .C(_02545_),
    .Y(_00289_));
 sg13g2_a21oi_1 _07913_ (.A1(net2531),
    .A2(_02545_),
    .Y(_02546_),
    .B1(net1228));
 sg13g2_o21ai_1 _07914_ (.B1(_02546_),
    .Y(_02547_),
    .A1(net2531),
    .A2(_02545_));
 sg13g2_inv_1 _07915_ (.Y(_00290_),
    .A(_02547_));
 sg13g2_nor3_1 _07916_ (.A(\i_uart_rx.cycle_counter[3] ),
    .B(_00814_),
    .C(\i_uart_rx.cycle_counter[5] ),
    .Y(_02548_));
 sg13g2_nor4_1 _07917_ (.A(_00795_),
    .B(\i_uart_rx.cycle_counter[1] ),
    .C(\i_uart_rx.cycle_counter[7] ),
    .D(\i_uart_rx.cycle_counter[6] ),
    .Y(_02549_));
 sg13g2_nand3_1 _07918_ (.B(_02548_),
    .C(_02549_),
    .A(\i_uart_rx.cycle_counter[4] ),
    .Y(_02550_));
 sg13g2_nor4_2 _07919_ (.A(\i_uart_rx.cycle_counter[9] ),
    .B(_00815_),
    .C(\i_uart_rx.cycle_counter[10] ),
    .Y(_02551_),
    .D(_02550_));
 sg13g2_o21ai_1 _07920_ (.B1(net1326),
    .Y(_02552_),
    .A1(\i_uart_rx.bit_sample ),
    .A2(_02551_));
 sg13g2_a21oi_1 _07921_ (.A1(_00781_),
    .A2(_02551_),
    .Y(_00291_),
    .B1(_02552_));
 sg13g2_nand2_1 _07922_ (.Y(_00292_),
    .A(net1326),
    .B(_02518_));
 sg13g2_a21oi_2 _07923_ (.B1(_01558_),
    .Y(_02553_),
    .A2(_01885_),
    .A1(_01474_));
 sg13g2_nor2_1 _07924_ (.A(\i_uart_rx.fsm_state[0] ),
    .B(_01556_),
    .Y(_02554_));
 sg13g2_nor3_1 _07925_ (.A(\i_uart_rx.fsm_state[0] ),
    .B(_00204_),
    .C(_01556_),
    .Y(_02555_));
 sg13g2_a21oi_2 _07926_ (.B1(_02525_),
    .Y(_02556_),
    .A2(_01554_),
    .A1(\i_uart_rx.fsm_state[1] ));
 sg13g2_a22oi_1 _07927_ (.Y(_02557_),
    .B1(_02556_),
    .B2(_00203_),
    .A2(_02555_),
    .A1(_02551_));
 sg13g2_nand2_1 _07928_ (.Y(_02558_),
    .A(_00781_),
    .B(_02525_));
 sg13g2_nand2_2 _07929_ (.Y(_02559_),
    .A(_01556_),
    .B(_02526_));
 sg13g2_nand3_1 _07930_ (.B(_02558_),
    .C(_02559_),
    .A(_02557_),
    .Y(_02560_));
 sg13g2_nor2_1 _07931_ (.A(net2472),
    .B(_02559_),
    .Y(_02561_));
 sg13g2_o21ai_1 _07932_ (.B1(net1326),
    .Y(_02562_),
    .A1(_02553_),
    .A2(_02560_));
 sg13g2_nor2_1 _07933_ (.A(_02561_),
    .B(_02562_),
    .Y(_00293_));
 sg13g2_nand2_1 _07934_ (.Y(_02563_),
    .A(_00204_),
    .B(_02551_));
 sg13g2_a21oi_1 _07935_ (.A1(_02554_),
    .A2(_02563_),
    .Y(_02564_),
    .B1(_02553_));
 sg13g2_nor2b_1 _07936_ (.A(_01554_),
    .B_N(net2575),
    .Y(_02565_));
 sg13g2_nor2_1 _07937_ (.A(net2680),
    .B(_02565_),
    .Y(_02566_));
 sg13g2_o21ai_1 _07938_ (.B1(_02564_),
    .Y(_02567_),
    .A1(_01555_),
    .A2(_02566_));
 sg13g2_a22oi_1 _07939_ (.Y(_02568_),
    .B1(_02567_),
    .B2(_02559_),
    .A2(_02565_),
    .A1(_02526_));
 sg13g2_nor2_1 _07940_ (.A(net1317),
    .B(_02568_),
    .Y(_00294_));
 sg13g2_a21oi_1 _07941_ (.A1(_01555_),
    .A2(_02559_),
    .Y(_02569_),
    .B1(net2512));
 sg13g2_nand2_1 _07942_ (.Y(_02570_),
    .A(\i_uart_rx.fsm_state[2] ),
    .B(_01555_));
 sg13g2_nand3_1 _07943_ (.B(_01555_),
    .C(_02522_),
    .A(net2512),
    .Y(_02571_));
 sg13g2_nand3_1 _07944_ (.B(_02556_),
    .C(_02571_),
    .A(net1325),
    .Y(_02572_));
 sg13g2_nor2_1 _07945_ (.A(net2513),
    .B(_02572_),
    .Y(_00295_));
 sg13g2_xnor2_1 _07946_ (.Y(_02573_),
    .A(\i_uart_rx.fsm_state[3] ),
    .B(_02570_));
 sg13g2_o21ai_1 _07947_ (.B1(_02556_),
    .Y(_02574_),
    .A1(_02523_),
    .A2(_02573_));
 sg13g2_a221oi_1 _07948_ (.B2(_02574_),
    .C1(net1318),
    .B1(_02564_),
    .A1(_00780_),
    .Y(_00296_),
    .A2(_02526_));
 sg13g2_nand2b_1 _07949_ (.Y(_00297_),
    .B(net1326),
    .A_N(net1832));
 sg13g2_nand2b_1 _07950_ (.Y(_00298_),
    .B(net1326),
    .A_N(net8));
 sg13g2_nand2_1 _07951_ (.Y(_02575_),
    .A(net1236),
    .B(_01883_));
 sg13g2_nor2_2 _07952_ (.A(net1454),
    .B(_02575_),
    .Y(_02576_));
 sg13g2_nand2_1 _07953_ (.Y(_02577_),
    .A(net1321),
    .B(_02576_));
 sg13g2_mux2_1 _07954_ (.A0(\data_to_write[8] ),
    .A1(net2201),
    .S(_02577_),
    .X(_00299_));
 sg13g2_nor2_1 _07955_ (.A(net1181),
    .B(net1173),
    .Y(_02578_));
 sg13g2_nand2_2 _07956_ (.Y(_02579_),
    .A(net1176),
    .B(_01833_));
 sg13g2_nand3_1 _07957_ (.B(_01840_),
    .C(net1170),
    .A(net1461),
    .Y(_02580_));
 sg13g2_a21oi_1 _07958_ (.A1(\i_core.cpu.instr_write_offset[2] ),
    .A2(\i_core.cpu.instr_write_offset[1] ),
    .Y(_02581_),
    .B1(_02580_));
 sg13g2_a21oi_1 _07959_ (.A1(_01840_),
    .A2(net1170),
    .Y(_02582_),
    .B1(net1387));
 sg13g2_or2_1 _07960_ (.X(_02583_),
    .B(_02582_),
    .A(_02581_));
 sg13g2_or2_2 _07961_ (.X(_02584_),
    .B(_02581_),
    .A(_02580_));
 sg13g2_nor2_1 _07962_ (.A(\i_core.cpu.instr_data_in[0] ),
    .B(net1129),
    .Y(_02585_));
 sg13g2_a21oi_1 _07963_ (.A1(_00808_),
    .A2(_02583_),
    .Y(_00300_),
    .B1(_02585_));
 sg13g2_nor2_1 _07964_ (.A(\i_core.cpu.instr_data_in[1] ),
    .B(net1129),
    .Y(_02586_));
 sg13g2_a21oi_1 _07965_ (.A1(_00809_),
    .A2(_02583_),
    .Y(_00301_),
    .B1(_02586_));
 sg13g2_nand4_1 _07966_ (.B(_01469_),
    .C(_01473_),
    .A(_01448_),
    .Y(_02587_),
    .D(_01883_));
 sg13g2_nor2_1 _07967_ (.A(\data_to_write[0] ),
    .B(net1205),
    .Y(_02588_));
 sg13g2_nor2_1 _07968_ (.A(\i_debug_uart_tx.cycle_counter[4] ),
    .B(_00779_),
    .Y(_02589_));
 sg13g2_and4_1 _07969_ (.A(\i_debug_uart_tx.cycle_counter[2] ),
    .B(\i_debug_uart_tx.cycle_counter[1] ),
    .C(\i_debug_uart_tx.cycle_counter[0] ),
    .D(_02589_),
    .X(_02590_));
 sg13g2_nand4_1 _07970_ (.B(\i_debug_uart_tx.cycle_counter[1] ),
    .C(\i_debug_uart_tx.cycle_counter[0] ),
    .A(\i_debug_uart_tx.cycle_counter[2] ),
    .Y(_02591_),
    .D(_02589_));
 sg13g2_o21ai_1 _07971_ (.B1(net2395),
    .Y(_02592_),
    .A1(net2292),
    .A2(\i_debug_uart_tx.fsm_state[1] ));
 sg13g2_nand3_1 _07972_ (.B(_02590_),
    .C(_02592_),
    .A(_01468_),
    .Y(_02593_));
 sg13g2_mux2_1 _07973_ (.A0(net2577),
    .A1(net2398),
    .S(_02593_),
    .X(_02594_));
 sg13g2_nor2b_1 _07974_ (.A(_02594_),
    .B_N(net1205),
    .Y(_02595_));
 sg13g2_nor3_1 _07975_ (.A(net1313),
    .B(_02588_),
    .C(_02595_),
    .Y(_00302_));
 sg13g2_nor2_1 _07976_ (.A(\data_to_write[1] ),
    .B(net1203),
    .Y(_02596_));
 sg13g2_mux2_1 _07977_ (.A0(net2589),
    .A1(net2577),
    .S(_02593_),
    .X(_02597_));
 sg13g2_nor2b_1 _07978_ (.A(_02597_),
    .B_N(net1203),
    .Y(_02598_));
 sg13g2_nor3_1 _07979_ (.A(net1313),
    .B(_02596_),
    .C(_02598_),
    .Y(_00303_));
 sg13g2_nor2_1 _07980_ (.A(\data_to_write[2] ),
    .B(net1204),
    .Y(_02599_));
 sg13g2_mux2_1 _07981_ (.A0(net2623),
    .A1(net2589),
    .S(_02593_),
    .X(_02600_));
 sg13g2_nor2b_1 _07982_ (.A(_02600_),
    .B_N(net1204),
    .Y(_02601_));
 sg13g2_nor3_1 _07983_ (.A(net1316),
    .B(_02599_),
    .C(_02601_),
    .Y(_00304_));
 sg13g2_nor2_1 _07984_ (.A(\data_to_write[3] ),
    .B(net1204),
    .Y(_02602_));
 sg13g2_mux2_1 _07985_ (.A0(net2596),
    .A1(\i_debug_uart_tx.data_to_send[3] ),
    .S(_02593_),
    .X(_02603_));
 sg13g2_nor2b_1 _07986_ (.A(net2597),
    .B_N(net1204),
    .Y(_02604_));
 sg13g2_nor3_1 _07987_ (.A(net1313),
    .B(_02602_),
    .C(_02604_),
    .Y(_00305_));
 sg13g2_nor2_1 _07988_ (.A(net2622),
    .B(net1203),
    .Y(_02605_));
 sg13g2_mux2_1 _07989_ (.A0(net2600),
    .A1(net2596),
    .S(_02593_),
    .X(_02606_));
 sg13g2_nor2b_1 _07990_ (.A(_02606_),
    .B_N(net1203),
    .Y(_02607_));
 sg13g2_nor3_1 _07991_ (.A(net1316),
    .B(_02605_),
    .C(_02607_),
    .Y(_00306_));
 sg13g2_nor2_1 _07992_ (.A(\data_to_write[5] ),
    .B(net1203),
    .Y(_02608_));
 sg13g2_mux2_1 _07993_ (.A0(net2565),
    .A1(net2600),
    .S(_02593_),
    .X(_02609_));
 sg13g2_nor2b_1 _07994_ (.A(_02609_),
    .B_N(net1203),
    .Y(_02610_));
 sg13g2_nor3_1 _07995_ (.A(net1313),
    .B(_02608_),
    .C(_02610_),
    .Y(_00307_));
 sg13g2_nor2_1 _07996_ (.A(\data_to_write[6] ),
    .B(net1203),
    .Y(_02611_));
 sg13g2_mux2_1 _07997_ (.A0(net1935),
    .A1(net2565),
    .S(_02593_),
    .X(_02612_));
 sg13g2_nor2b_1 _07998_ (.A(_02612_),
    .B_N(net1203),
    .Y(_02613_));
 sg13g2_nor3_1 _07999_ (.A(net1313),
    .B(_02611_),
    .C(_02613_),
    .Y(_00308_));
 sg13g2_nand2_1 _08000_ (.Y(_02614_),
    .A(net1935),
    .B(_02593_));
 sg13g2_o21ai_1 _08001_ (.B1(net1320),
    .Y(_02615_),
    .A1(_00844_),
    .A2(net1205));
 sg13g2_a21oi_1 _08002_ (.A1(net1205),
    .A2(_02614_),
    .Y(_00309_),
    .B1(_02615_));
 sg13g2_nor2_1 _08003_ (.A(net1871),
    .B(_01469_),
    .Y(_02616_));
 sg13g2_nand2b_1 _08004_ (.Y(_02617_),
    .B(_02591_),
    .A_N(net1319));
 sg13g2_nor2_1 _08005_ (.A(\i_debug_uart_tx.cycle_counter[0] ),
    .B(_01470_),
    .Y(_02618_));
 sg13g2_nor3_1 _08006_ (.A(net1872),
    .B(_02617_),
    .C(_02618_),
    .Y(_00310_));
 sg13g2_a21oi_1 _08007_ (.A1(\i_debug_uart_tx.cycle_counter[0] ),
    .A2(_01470_),
    .Y(_02619_),
    .B1(net2223));
 sg13g2_nand3_1 _08008_ (.B(\i_debug_uart_tx.cycle_counter[0] ),
    .C(_01470_),
    .A(net2223),
    .Y(_02620_));
 sg13g2_nand2b_1 _08009_ (.Y(_02621_),
    .B(_02620_),
    .A_N(_02617_));
 sg13g2_nor2_1 _08010_ (.A(net2224),
    .B(_02621_),
    .Y(_00311_));
 sg13g2_nand4_1 _08011_ (.B(net2223),
    .C(\i_debug_uart_tx.cycle_counter[0] ),
    .A(net2447),
    .Y(_02622_),
    .D(_01470_));
 sg13g2_xor2_1 _08012_ (.B(_02620_),
    .A(net2447),
    .X(_02623_));
 sg13g2_nor2_1 _08013_ (.A(_02617_),
    .B(net2448),
    .Y(_00312_));
 sg13g2_xnor2_1 _08014_ (.Y(_02624_),
    .A(_00779_),
    .B(_02622_));
 sg13g2_nor2_1 _08015_ (.A(_02617_),
    .B(net2536),
    .Y(_00313_));
 sg13g2_o21ai_1 _08016_ (.B1(net1881),
    .Y(_02625_),
    .A1(_00779_),
    .A2(_02622_));
 sg13g2_nor2_1 _08017_ (.A(net1319),
    .B(net1882),
    .Y(_00314_));
 sg13g2_nand2_1 _08018_ (.Y(_02626_),
    .A(_01470_),
    .B(_02591_));
 sg13g2_nor2b_1 _08019_ (.A(\i_debug_uart_tx.fsm_state[2] ),
    .B_N(\i_debug_uart_tx.fsm_state[3] ),
    .Y(_02627_));
 sg13g2_nor2b_1 _08020_ (.A(\i_debug_uart_tx.fsm_state[0] ),
    .B_N(\i_debug_uart_tx.fsm_state[1] ),
    .Y(_02628_));
 sg13g2_a21oi_1 _08021_ (.A1(\i_debug_uart_tx.fsm_state[1] ),
    .A2(_02627_),
    .Y(_02629_),
    .B1(\i_debug_uart_tx.fsm_state[0] ));
 sg13g2_nand2_1 _08022_ (.Y(_02630_),
    .A(_01468_),
    .B(_02629_));
 sg13g2_nand2_1 _08023_ (.Y(_02631_),
    .A(net1205),
    .B(_02630_));
 sg13g2_a22oi_1 _08024_ (.Y(_02632_),
    .B1(_02626_),
    .B2(_02631_),
    .A2(_02591_),
    .A1(net2545));
 sg13g2_nor2_1 _08025_ (.A(net1313),
    .B(net2546),
    .Y(_00315_));
 sg13g2_a21oi_1 _08026_ (.A1(_01470_),
    .A2(_02591_),
    .Y(_02633_),
    .B1(_02629_));
 sg13g2_nor2_1 _08027_ (.A(net2496),
    .B(_02633_),
    .Y(_02634_));
 sg13g2_a21oi_1 _08028_ (.A1(net2496),
    .A2(_02633_),
    .Y(_02635_),
    .B1(net1313));
 sg13g2_nor2b_1 _08029_ (.A(net2497),
    .B_N(_02635_),
    .Y(_00316_));
 sg13g2_and3_1 _08030_ (.X(_02636_),
    .A(\i_debug_uart_tx.fsm_state[1] ),
    .B(\i_debug_uart_tx.fsm_state[0] ),
    .C(_02590_));
 sg13g2_nand3_1 _08031_ (.B(\i_debug_uart_tx.fsm_state[1] ),
    .C(\i_debug_uart_tx.fsm_state[0] ),
    .A(\i_debug_uart_tx.fsm_state[2] ),
    .Y(_02637_));
 sg13g2_o21ai_1 _08032_ (.B1(net1321),
    .Y(_02638_),
    .A1(net2292),
    .A2(_02636_));
 sg13g2_a21oi_1 _08033_ (.A1(net2292),
    .A2(_02636_),
    .Y(_00317_),
    .B1(_02638_));
 sg13g2_xor2_1 _08034_ (.B(_02637_),
    .A(net2395),
    .X(_02639_));
 sg13g2_a21oi_1 _08035_ (.A1(_02627_),
    .A2(_02628_),
    .Y(_02640_),
    .B1(_02639_));
 sg13g2_a22oi_1 _08036_ (.Y(_02641_),
    .B1(_02626_),
    .B2(_02640_),
    .A2(_02591_),
    .A1(net2395));
 sg13g2_nor2_1 _08037_ (.A(net1313),
    .B(net2396),
    .Y(_00318_));
 sg13g2_nand2b_1 _08038_ (.Y(_02642_),
    .B(net1434),
    .A_N(net2687));
 sg13g2_a21oi_1 _08039_ (.A1(_01865_),
    .A2(_02642_),
    .Y(_02643_),
    .B1(net2123));
 sg13g2_and2_1 _08040_ (.A(net1323),
    .B(_01865_),
    .X(_00570_));
 sg13g2_and2_1 _08041_ (.A(_02643_),
    .B(_00570_),
    .X(_00319_));
 sg13g2_xnor2_1 _08042_ (.Y(_02644_),
    .A(\i_spi.clock_divider[0] ),
    .B(\i_spi.clock_count[0] ));
 sg13g2_xnor2_1 _08043_ (.Y(_02645_),
    .A(\i_spi.clock_divider[1] ),
    .B(\i_spi.clock_count[1] ));
 sg13g2_nand2_2 _08044_ (.Y(_02646_),
    .A(_02644_),
    .B(_02645_));
 sg13g2_a21oi_1 _08045_ (.A1(net1455),
    .A2(_02646_),
    .Y(_02647_),
    .B1(net2154));
 sg13g2_and2_1 _08046_ (.A(net1455),
    .B(net2154),
    .X(_02648_));
 sg13g2_nor3_1 _08047_ (.A(net1317),
    .B(_02647_),
    .C(_02648_),
    .Y(_00320_));
 sg13g2_nor2_2 _08048_ (.A(_00778_),
    .B(_02646_),
    .Y(_02649_));
 sg13g2_o21ai_1 _08049_ (.B1(net1325),
    .Y(_02650_),
    .A1(net2484),
    .A2(_02648_));
 sg13g2_a21oi_1 _08050_ (.A1(net2484),
    .A2(_02648_),
    .Y(_02651_),
    .B1(_02650_));
 sg13g2_nor2b_1 _08051_ (.A(_02649_),
    .B_N(_02651_),
    .Y(_00321_));
 sg13g2_a22oi_1 _08052_ (.Y(_02652_),
    .B1(_02646_),
    .B2(net1455),
    .A2(_02575_),
    .A1(_00156_));
 sg13g2_nand2b_1 _08053_ (.Y(_02653_),
    .B(net1454),
    .A_N(\i_spi.spi_clk_out ));
 sg13g2_a21oi_1 _08054_ (.A1(net1965),
    .A2(_00776_),
    .Y(_02654_),
    .B1(_02653_));
 sg13g2_nand3b_1 _08055_ (.B(_02652_),
    .C(net1325),
    .Y(_02655_),
    .A_N(_02654_));
 sg13g2_nand2_1 _08056_ (.Y(_02656_),
    .A(net1455),
    .B(net4));
 sg13g2_o21ai_1 _08057_ (.B1(_02656_),
    .Y(_02657_),
    .A1(_00775_),
    .A2(net1455));
 sg13g2_mux2_1 _08058_ (.A0(_02657_),
    .A1(net2432),
    .S(_02655_),
    .X(_00322_));
 sg13g2_nand2_1 _08059_ (.Y(_02658_),
    .A(_00155_),
    .B(_02649_));
 sg13g2_nand2_1 _08060_ (.Y(_02659_),
    .A(_02652_),
    .B(_02658_));
 sg13g2_nor2_1 _08061_ (.A(net1916),
    .B(\i_spi.bits_remaining[0] ),
    .Y(_02660_));
 sg13g2_nand2b_1 _08062_ (.Y(_02661_),
    .B(_02660_),
    .A_N(\i_spi.bits_remaining[2] ));
 sg13g2_nor2_2 _08063_ (.A(net2315),
    .B(_02661_),
    .Y(_02662_));
 sg13g2_nand3_1 _08064_ (.B(net1455),
    .C(_02662_),
    .A(\i_spi.spi_clk_out ),
    .Y(_02663_));
 sg13g2_nor2b_1 _08065_ (.A(_02659_),
    .B_N(_02663_),
    .Y(_02664_));
 sg13g2_and2_1 _08066_ (.A(net1455),
    .B(_02664_),
    .X(_02665_));
 sg13g2_o21ai_1 _08067_ (.B1(net1321),
    .Y(_02666_),
    .A1(net1978),
    .A2(_02665_));
 sg13g2_a21oi_1 _08068_ (.A1(net1978),
    .A2(_02664_),
    .Y(_00323_),
    .B1(_02666_));
 sg13g2_o21ai_1 _08069_ (.B1(_02664_),
    .Y(_02667_),
    .A1(_00777_),
    .A2(_00778_));
 sg13g2_a22oi_1 _08070_ (.Y(_02668_),
    .B1(_02667_),
    .B2(net1916),
    .A2(_02665_),
    .A1(_02660_));
 sg13g2_nor2_1 _08071_ (.A(net1315),
    .B(net1917),
    .Y(_00324_));
 sg13g2_xor2_1 _08072_ (.B(_02660_),
    .A(net2211),
    .X(_02669_));
 sg13g2_a22oi_1 _08073_ (.Y(_02670_),
    .B1(_02665_),
    .B2(_02669_),
    .A2(_02659_),
    .A1(net2211));
 sg13g2_nor2_1 _08074_ (.A(net1314),
    .B(net2212),
    .Y(_00325_));
 sg13g2_o21ai_1 _08075_ (.B1(_02664_),
    .Y(_02671_),
    .A1(_00156_),
    .A2(_02662_));
 sg13g2_o21ai_1 _08076_ (.B1(net2315),
    .Y(_02672_),
    .A1(_02659_),
    .A2(_02661_));
 sg13g2_a21oi_1 _08077_ (.A1(_02671_),
    .A2(net2316),
    .Y(_00326_),
    .B1(net1317));
 sg13g2_a21oi_1 _08078_ (.A1(net1236),
    .A2(_01883_),
    .Y(_02673_),
    .B1(net1454));
 sg13g2_nand3b_1 _08079_ (.B(_02649_),
    .C(_02662_),
    .Y(_02674_),
    .A_N(\i_spi.spi_clk_out ));
 sg13g2_inv_1 _08080_ (.Y(_02675_),
    .A(_02674_));
 sg13g2_nor3_1 _08081_ (.A(net1317),
    .B(_02673_),
    .C(_02675_),
    .Y(_00327_));
 sg13g2_mux2_1 _08082_ (.A0(\data_to_write[9] ),
    .A1(net2155),
    .S(_02577_),
    .X(_00328_));
 sg13g2_nand2_1 _08083_ (.Y(_02676_),
    .A(net2134),
    .B(_02674_));
 sg13g2_a21oi_1 _08084_ (.A1(\i_spi.end_txn_reg ),
    .A2(_02675_),
    .Y(_02677_),
    .B1(net1314));
 sg13g2_o21ai_1 _08085_ (.B1(_02677_),
    .Y(_00329_),
    .A1(_02576_),
    .A2(_02676_));
 sg13g2_or2_1 _08086_ (.X(_02678_),
    .B(_02649_),
    .A(_02576_));
 sg13g2_o21ai_1 _08087_ (.B1(_02678_),
    .Y(_02679_),
    .A1(_02653_),
    .A2(_02662_));
 sg13g2_o21ai_1 _08088_ (.B1(_02679_),
    .Y(_02680_),
    .A1(net2562),
    .A2(_02678_));
 sg13g2_nor2_1 _08089_ (.A(net1317),
    .B(_02680_),
    .Y(_00330_));
 sg13g2_nand2_1 _08090_ (.Y(_02681_),
    .A(net2398),
    .B(_01468_));
 sg13g2_nand4_1 _08091_ (.B(_01470_),
    .C(_02592_),
    .A(net1320),
    .Y(_00331_),
    .D(net2399));
 sg13g2_or4_2 _08092_ (.A(net1450),
    .B(_01449_),
    .C(_01450_),
    .D(_01884_),
    .X(_02682_));
 sg13g2_nor2_1 _08093_ (.A(net2688),
    .B(_02682_),
    .Y(_02683_));
 sg13g2_nor2b_1 _08094_ (.A(net1965),
    .B_N(_02682_),
    .Y(_02684_));
 sg13g2_nor3_1 _08095_ (.A(net1317),
    .B(_02683_),
    .C(_02684_),
    .Y(_00332_));
 sg13g2_a21oi_1 _08096_ (.A1(net2314),
    .A2(_02682_),
    .Y(_02685_),
    .B1(net1317));
 sg13g2_o21ai_1 _08097_ (.B1(_02685_),
    .Y(_00333_),
    .A1(_00775_),
    .A2(_02682_));
 sg13g2_nor2_1 _08098_ (.A(\data_to_write[1] ),
    .B(_02682_),
    .Y(_02686_));
 sg13g2_nor2b_1 _08099_ (.A(net2042),
    .B_N(_02682_),
    .Y(_02687_));
 sg13g2_nor3_1 _08100_ (.A(net1317),
    .B(_02686_),
    .C(_02687_),
    .Y(_00334_));
 sg13g2_nand4_1 _08101_ (.B(_01237_),
    .C(_01238_),
    .A(_01231_),
    .Y(_02688_),
    .D(_01242_));
 sg13g2_and2_1 _08102_ (.A(net1379),
    .B(_02688_),
    .X(_02689_));
 sg13g2_and2_2 _08103_ (.A(_01231_),
    .B(_01251_),
    .X(_02690_));
 sg13g2_inv_1 _08104_ (.Y(_02691_),
    .A(_02690_));
 sg13g2_nor4_1 _08105_ (.A(net1410),
    .B(_00084_),
    .C(_02689_),
    .D(_02690_),
    .Y(_02692_));
 sg13g2_nand2_1 _08106_ (.Y(_02693_),
    .A(_01234_),
    .B(_02360_));
 sg13g2_o21ai_1 _08107_ (.B1(_02692_),
    .Y(_02694_),
    .A1(_01051_),
    .A2(_02693_));
 sg13g2_nand2_1 _08108_ (.Y(_02695_),
    .A(_01051_),
    .B(_02380_));
 sg13g2_a21oi_2 _08109_ (.B1(_01234_),
    .Y(_02696_),
    .A2(_00841_),
    .A1(\i_core.cpu.i_core.interrupt_req[1] ));
 sg13g2_a22oi_1 _08110_ (.Y(_02697_),
    .B1(_02696_),
    .B2(_00774_),
    .A2(_02695_),
    .A1(_01234_));
 sg13g2_o21ai_1 _08111_ (.B1(_02353_),
    .Y(_02698_),
    .A1(_02694_),
    .A2(_02697_));
 sg13g2_a21oi_1 _08112_ (.A1(_00774_),
    .A2(_02694_),
    .Y(_00335_),
    .B1(_02698_));
 sg13g2_nor2_1 _08113_ (.A(_01090_),
    .B(_02693_),
    .Y(_02699_));
 sg13g2_nor2b_1 _08114_ (.A(_02699_),
    .B_N(_02692_),
    .Y(_02700_));
 sg13g2_nor2b_2 _08115_ (.A(\i_core.cpu.i_core.last_interrupt_req[0] ),
    .B_N(\i_core.cpu.i_core.interrupt_req[0] ),
    .Y(_02701_));
 sg13g2_o21ai_1 _08116_ (.B1(_02700_),
    .Y(_02702_),
    .A1(_01234_),
    .A2(_02701_));
 sg13g2_a21oi_1 _08117_ (.A1(_01090_),
    .A2(_02380_),
    .Y(_02703_),
    .B1(_01235_));
 sg13g2_a221oi_1 _08118_ (.B2(_02700_),
    .C1(_02354_),
    .B1(_02703_),
    .A1(_00773_),
    .Y(_00336_),
    .A2(_02702_));
 sg13g2_o21ai_1 _08119_ (.B1(_02690_),
    .Y(_02704_),
    .A1(_00926_),
    .A2(_02359_));
 sg13g2_a22oi_1 _08120_ (.Y(_02705_),
    .B1(_02704_),
    .B2(net2168),
    .A2(_02381_),
    .A1(_01251_));
 sg13g2_nor2_1 _08121_ (.A(_02354_),
    .B(_02705_),
    .Y(_00337_));
 sg13g2_nand2_1 _08122_ (.Y(_02706_),
    .A(net2683),
    .B(_02360_));
 sg13g2_nand3_1 _08123_ (.B(_02690_),
    .C(_02706_),
    .A(_01003_),
    .Y(_02707_));
 sg13g2_o21ai_1 _08124_ (.B1(_02690_),
    .Y(_02708_),
    .A1(_01003_),
    .A2(_02359_));
 sg13g2_nand2_1 _08125_ (.Y(_02709_),
    .A(net2313),
    .B(_02708_));
 sg13g2_a21oi_1 _08126_ (.A1(_02707_),
    .A2(_02709_),
    .Y(_00338_),
    .B1(_02354_));
 sg13g2_o21ai_1 _08127_ (.B1(_02690_),
    .Y(_02710_),
    .A1(_01051_),
    .A2(_02693_));
 sg13g2_nand2_1 _08128_ (.Y(_02711_),
    .A(net2283),
    .B(_02710_));
 sg13g2_nand3_1 _08129_ (.B(_01251_),
    .C(_02380_),
    .A(_01051_),
    .Y(_02712_));
 sg13g2_a21oi_1 _08130_ (.A1(_02711_),
    .A2(_02712_),
    .Y(_00339_),
    .B1(_02354_));
 sg13g2_nand3_1 _08131_ (.B(_01251_),
    .C(_02380_),
    .A(_01090_),
    .Y(_02713_));
 sg13g2_o21ai_1 _08132_ (.B1(net2326),
    .Y(_02714_),
    .A1(_02691_),
    .A2(_02699_));
 sg13g2_a21oi_1 _08133_ (.A1(_02713_),
    .A2(_02714_),
    .Y(_00340_),
    .B1(_02354_));
 sg13g2_nand2_1 _08134_ (.Y(_02715_),
    .A(net2386),
    .B(_01460_));
 sg13g2_nand4_1 _08135_ (.B(_01462_),
    .C(_02452_),
    .A(net1322),
    .Y(_00341_),
    .D(_02715_));
 sg13g2_nor2b_1 _08136_ (.A(_01167_),
    .B_N(_01370_),
    .Y(_02716_));
 sg13g2_o21ai_1 _08137_ (.B1(_01370_),
    .Y(_02717_),
    .A1(_01163_),
    .A2(net1306));
 sg13g2_mux2_1 _08138_ (.A0(net2543),
    .A1(\i_core.cpu.i_core.i_shift.a[4] ),
    .S(net1267),
    .X(_00342_));
 sg13g2_mux2_1 _08139_ (.A0(net2467),
    .A1(\i_core.cpu.i_core.i_shift.a[5] ),
    .S(net1267),
    .X(_00343_));
 sg13g2_mux2_1 _08140_ (.A0(net2527),
    .A1(\i_core.cpu.i_core.i_shift.a[6] ),
    .S(_02717_),
    .X(_00344_));
 sg13g2_mux2_1 _08141_ (.A0(net2474),
    .A1(\i_core.cpu.i_core.i_shift.a[7] ),
    .S(_02717_),
    .X(_00345_));
 sg13g2_mux2_1 _08142_ (.A0(net2649),
    .A1(net2616),
    .S(net1266),
    .X(_00346_));
 sg13g2_mux2_1 _08143_ (.A0(net2646),
    .A1(\i_core.cpu.i_core.i_shift.a[9] ),
    .S(net1266),
    .X(_00347_));
 sg13g2_mux2_1 _08144_ (.A0(net2629),
    .A1(net2615),
    .S(net1266),
    .X(_00348_));
 sg13g2_mux2_1 _08145_ (.A0(net2636),
    .A1(net2612),
    .S(net1264),
    .X(_00349_));
 sg13g2_mux2_1 _08146_ (.A0(net2616),
    .A1(net2351),
    .S(net1266),
    .X(_00350_));
 sg13g2_mux2_1 _08147_ (.A0(\i_core.cpu.i_core.i_shift.a[9] ),
    .A1(net2632),
    .S(net1266),
    .X(_00351_));
 sg13g2_mux2_1 _08148_ (.A0(net2615),
    .A1(net2255),
    .S(net1266),
    .X(_00352_));
 sg13g2_mux2_1 _08149_ (.A0(net2612),
    .A1(net2409),
    .S(net1266),
    .X(_00353_));
 sg13g2_mux2_1 _08150_ (.A0(net2351),
    .A1(net2325),
    .S(net1265),
    .X(_00354_));
 sg13g2_mux2_1 _08151_ (.A0(\i_core.cpu.i_core.i_shift.a[13] ),
    .A1(net2216),
    .S(net1264),
    .X(_00355_));
 sg13g2_mux2_1 _08152_ (.A0(net2255),
    .A1(net2149),
    .S(net1264),
    .X(_00356_));
 sg13g2_mux2_1 _08153_ (.A0(net2409),
    .A1(net2337),
    .S(net1265),
    .X(_00357_));
 sg13g2_mux2_1 _08154_ (.A0(net2325),
    .A1(net2278),
    .S(net1264),
    .X(_00358_));
 sg13g2_mux2_1 _08155_ (.A0(\i_core.cpu.i_core.i_shift.a[17] ),
    .A1(net2145),
    .S(net1264),
    .X(_00359_));
 sg13g2_mux2_1 _08156_ (.A0(net2149),
    .A1(\i_core.cpu.i_core.i_shift.a[22] ),
    .S(net1264),
    .X(_00360_));
 sg13g2_mux2_1 _08157_ (.A0(net2337),
    .A1(net2273),
    .S(net1264),
    .X(_00361_));
 sg13g2_mux2_1 _08158_ (.A0(net2278),
    .A1(\i_core.cpu.i_core.i_shift.a[24] ),
    .S(net1264),
    .X(_00362_));
 sg13g2_mux2_1 _08159_ (.A0(net2145),
    .A1(net2178),
    .S(net1265),
    .X(_00363_));
 sg13g2_mux2_1 _08160_ (.A0(net2271),
    .A1(\i_core.cpu.i_core.i_shift.a[26] ),
    .S(net1265),
    .X(_00364_));
 sg13g2_mux2_1 _08161_ (.A0(net2273),
    .A1(\i_core.cpu.i_core.i_shift.a[27] ),
    .S(net1265),
    .X(_00365_));
 sg13g2_mux2_1 _08162_ (.A0(net2476),
    .A1(net2301),
    .S(net1267),
    .X(_00366_));
 sg13g2_mux2_1 _08163_ (.A0(net2178),
    .A1(net2250),
    .S(net1265),
    .X(_00367_));
 sg13g2_mux2_1 _08164_ (.A0(net2299),
    .A1(\i_core.cpu.i_core.i_shift.a[30] ),
    .S(net1265),
    .X(_00368_));
 sg13g2_mux2_1 _08165_ (.A0(net2377),
    .A1(\i_core.cpu.i_core.i_shift.a[31] ),
    .S(net1267),
    .X(_00369_));
 sg13g2_nand2_2 _08166_ (.Y(_02718_),
    .A(_01735_),
    .B(net1267));
 sg13g2_nand2_2 _08167_ (.Y(_02719_),
    .A(_01164_),
    .B(_02067_));
 sg13g2_inv_1 _08168_ (.Y(_02720_),
    .A(_02719_));
 sg13g2_nand2b_1 _08169_ (.Y(_02721_),
    .B(_02720_),
    .A_N(_01646_));
 sg13g2_a21oi_1 _08170_ (.A1(_01030_),
    .A2(_02719_),
    .Y(_02722_),
    .B1(net1307));
 sg13g2_a22oi_1 _08171_ (.Y(_02723_),
    .B1(_02721_),
    .B2(_02722_),
    .A2(net1306),
    .A1(_01003_));
 sg13g2_nand2_1 _08172_ (.Y(_02724_),
    .A(_01688_),
    .B(net1267));
 sg13g2_nor2_1 _08173_ (.A(_01734_),
    .B(_02724_),
    .Y(_02725_));
 sg13g2_a21oi_1 _08174_ (.A1(net2542),
    .A2(_02716_),
    .Y(_02726_),
    .B1(_02725_));
 sg13g2_o21ai_1 _08175_ (.B1(_02726_),
    .Y(_00370_),
    .A1(_02718_),
    .A2(_02723_));
 sg13g2_nor2_1 _08176_ (.A(_01928_),
    .B(_02719_),
    .Y(_02727_));
 sg13g2_nand2b_1 _08177_ (.Y(_02728_),
    .B(_02719_),
    .A_N(_00965_));
 sg13g2_nor2_1 _08178_ (.A(net1307),
    .B(_02727_),
    .Y(_02729_));
 sg13g2_a22oi_1 _08179_ (.Y(_02730_),
    .B1(_02728_),
    .B2(_02729_),
    .A2(net1306),
    .A1(_00926_));
 sg13g2_nand2b_1 _08180_ (.Y(_02731_),
    .B(net1267),
    .A_N(_02337_));
 sg13g2_o21ai_1 _08181_ (.B1(_02731_),
    .Y(_02732_),
    .A1(net2655),
    .A2(net1267));
 sg13g2_o21ai_1 _08182_ (.B1(_02732_),
    .Y(_00371_),
    .A1(_02718_),
    .A2(_02730_));
 sg13g2_nand3b_1 _08183_ (.B(_00793_),
    .C(\i_core.cpu.instr_write_offset[1] ),
    .Y(_02733_),
    .A_N(_02580_));
 sg13g2_inv_1 _08184_ (.Y(_02734_),
    .A(net1154));
 sg13g2_nor3_1 _08185_ (.A(net2438),
    .B(net1457),
    .C(_02734_),
    .Y(_02735_));
 sg13g2_a21oi_1 _08186_ (.A1(_00825_),
    .A2(_02734_),
    .Y(_00372_),
    .B1(_02735_));
 sg13g2_nor3_1 _08187_ (.A(net2341),
    .B(net1457),
    .C(_02734_),
    .Y(_02736_));
 sg13g2_a21oi_1 _08188_ (.A1(_00831_),
    .A2(_02734_),
    .Y(_00373_),
    .B1(_02736_));
 sg13g2_nor3_1 _08189_ (.A(\i_core.cpu.instr_write_offset[2] ),
    .B(\i_core.cpu.instr_write_offset[1] ),
    .C(_02580_),
    .Y(_02737_));
 sg13g2_mux2_1 _08190_ (.A0(net2158),
    .A1(\i_core.cpu.instr_data_in[2] ),
    .S(net1151),
    .X(_00374_));
 sg13g2_mux2_1 _08191_ (.A0(net2112),
    .A1(\i_core.cpu.instr_data_in[3] ),
    .S(net1148),
    .X(_00375_));
 sg13g2_mux2_1 _08192_ (.A0(net1931),
    .A1(\i_core.cpu.instr_data_in[4] ),
    .S(net1151),
    .X(_00376_));
 sg13g2_mux2_1 _08193_ (.A0(net1941),
    .A1(\i_core.cpu.instr_data_in[5] ),
    .S(net1149),
    .X(_00377_));
 sg13g2_mux2_1 _08194_ (.A0(net1912),
    .A1(\i_core.cpu.instr_data_in[6] ),
    .S(net1148),
    .X(_00378_));
 sg13g2_mux2_1 _08195_ (.A0(net1939),
    .A1(\i_core.cpu.instr_data_in[7] ),
    .S(net1149),
    .X(_00379_));
 sg13g2_nor2_1 _08196_ (.A(net1933),
    .B(net1148),
    .Y(_02738_));
 sg13g2_a21oi_1 _08197_ (.A1(_00208_),
    .A2(net1148),
    .Y(_00380_),
    .B1(_02738_));
 sg13g2_nor2_1 _08198_ (.A(net1948),
    .B(net1148),
    .Y(_02739_));
 sg13g2_a21oi_1 _08199_ (.A1(_00209_),
    .A2(net1148),
    .Y(_00381_),
    .B1(_02739_));
 sg13g2_nor2_1 _08200_ (.A(net1961),
    .B(net1150),
    .Y(_02740_));
 sg13g2_a21oi_1 _08201_ (.A1(_00210_),
    .A2(net1150),
    .Y(_00382_),
    .B1(_02740_));
 sg13g2_nor2_1 _08202_ (.A(net1899),
    .B(net1148),
    .Y(_02741_));
 sg13g2_a21oi_1 _08203_ (.A1(_00211_),
    .A2(net1149),
    .Y(_00383_),
    .B1(_02741_));
 sg13g2_nor2_1 _08204_ (.A(net1910),
    .B(net1150),
    .Y(_02742_));
 sg13g2_a21oi_1 _08205_ (.A1(_00205_),
    .A2(net1150),
    .Y(_00384_),
    .B1(_02742_));
 sg13g2_nor2_1 _08206_ (.A(net1950),
    .B(net1150),
    .Y(_02743_));
 sg13g2_a21oi_1 _08207_ (.A1(_00206_),
    .A2(net1151),
    .Y(_00385_),
    .B1(_02743_));
 sg13g2_nor2_1 _08208_ (.A(net1922),
    .B(net1149),
    .Y(_02744_));
 sg13g2_a21oi_1 _08209_ (.A1(_00212_),
    .A2(net1149),
    .Y(_00386_),
    .B1(_02744_));
 sg13g2_nor2_1 _08210_ (.A(net1954),
    .B(net1148),
    .Y(_02745_));
 sg13g2_a21oi_1 _08211_ (.A1(_00207_),
    .A2(net1149),
    .Y(_00387_),
    .B1(_02745_));
 sg13g2_or3_2 _08212_ (.A(_00793_),
    .B(\i_core.cpu.instr_write_offset[1] ),
    .C(_02580_),
    .X(_02746_));
 sg13g2_inv_1 _08213_ (.Y(_02747_),
    .A(net1146));
 sg13g2_mux2_1 _08214_ (.A0(\i_core.cpu.instr_data_in[2] ),
    .A1(net2318),
    .S(net1147),
    .X(_00388_));
 sg13g2_mux2_1 _08215_ (.A0(\i_core.cpu.instr_data_in[3] ),
    .A1(net2349),
    .S(net1145),
    .X(_00389_));
 sg13g2_mux2_1 _08216_ (.A0(\i_core.cpu.instr_data_in[4] ),
    .A1(net2012),
    .S(net1147),
    .X(_00390_));
 sg13g2_mux2_1 _08217_ (.A0(\i_core.cpu.instr_data_in[5] ),
    .A1(net2108),
    .S(net1146),
    .X(_00391_));
 sg13g2_mux2_1 _08218_ (.A0(\i_core.cpu.instr_data_in[6] ),
    .A1(net2021),
    .S(net1145),
    .X(_00392_));
 sg13g2_mux2_1 _08219_ (.A0(\i_core.cpu.instr_data_in[7] ),
    .A1(net2049),
    .S(net1146),
    .X(_00393_));
 sg13g2_nand2_1 _08220_ (.Y(_02748_),
    .A(net1867),
    .B(net1145));
 sg13g2_o21ai_1 _08221_ (.B1(_02748_),
    .Y(_00394_),
    .A1(_00208_),
    .A2(net1145));
 sg13g2_nand2_1 _08222_ (.Y(_02749_),
    .A(net1855),
    .B(net1145));
 sg13g2_o21ai_1 _08223_ (.B1(_02749_),
    .Y(_00395_),
    .A1(_00209_),
    .A2(net1145));
 sg13g2_nand2_1 _08224_ (.Y(_02750_),
    .A(net1849),
    .B(net1147));
 sg13g2_o21ai_1 _08225_ (.B1(_02750_),
    .Y(_00396_),
    .A1(_00210_),
    .A2(_02746_));
 sg13g2_nand2_1 _08226_ (.Y(_02751_),
    .A(net1869),
    .B(net1145));
 sg13g2_o21ai_1 _08227_ (.B1(_02751_),
    .Y(_00397_),
    .A1(_00211_),
    .A2(net1145));
 sg13g2_nand2_1 _08228_ (.Y(_02752_),
    .A(net1845),
    .B(net1147));
 sg13g2_o21ai_1 _08229_ (.B1(_02752_),
    .Y(_00398_),
    .A1(_00205_),
    .A2(net1147));
 sg13g2_nand2_1 _08230_ (.Y(_02753_),
    .A(net1828),
    .B(net1147));
 sg13g2_o21ai_1 _08231_ (.B1(_02753_),
    .Y(_00399_),
    .A1(_00206_),
    .A2(net1147));
 sg13g2_nand2_1 _08232_ (.Y(_02754_),
    .A(net1876),
    .B(net1146));
 sg13g2_o21ai_1 _08233_ (.B1(_02754_),
    .Y(_00400_),
    .A1(_00212_),
    .A2(net1146));
 sg13g2_nand2_1 _08234_ (.Y(_02755_),
    .A(net1843),
    .B(net1146));
 sg13g2_o21ai_1 _08235_ (.B1(_02755_),
    .Y(_00401_),
    .A1(_00207_),
    .A2(net1146));
 sg13g2_mux2_1 _08236_ (.A0(\i_core.cpu.instr_data_in[2] ),
    .A1(net2372),
    .S(net1130),
    .X(_00402_));
 sg13g2_mux2_1 _08237_ (.A0(\i_core.cpu.instr_data_in[3] ),
    .A1(net2288),
    .S(net1129),
    .X(_00403_));
 sg13g2_mux2_1 _08238_ (.A0(\i_core.cpu.instr_data_in[4] ),
    .A1(net2073),
    .S(net1130),
    .X(_00404_));
 sg13g2_mux2_1 _08239_ (.A0(\i_core.cpu.instr_data_in[5] ),
    .A1(net2017),
    .S(net1128),
    .X(_00405_));
 sg13g2_mux2_1 _08240_ (.A0(\i_core.cpu.instr_data_in[6] ),
    .A1(net2079),
    .S(net1128),
    .X(_00406_));
 sg13g2_mux2_1 _08241_ (.A0(\i_core.cpu.instr_data_in[7] ),
    .A1(net2019),
    .S(net1128),
    .X(_00407_));
 sg13g2_nand2_1 _08242_ (.Y(_02756_),
    .A(net1863),
    .B(net1128));
 sg13g2_o21ai_1 _08243_ (.B1(_02756_),
    .Y(_00408_),
    .A1(_00208_),
    .A2(net1128));
 sg13g2_nand2_1 _08244_ (.Y(_02757_),
    .A(net1865),
    .B(net1128));
 sg13g2_o21ai_1 _08245_ (.B1(_02757_),
    .Y(_00409_),
    .A1(_00209_),
    .A2(net1128));
 sg13g2_nand2_1 _08246_ (.Y(_02758_),
    .A(net1853),
    .B(_02584_));
 sg13g2_o21ai_1 _08247_ (.B1(_02758_),
    .Y(_00410_),
    .A1(_00210_),
    .A2(_02584_));
 sg13g2_nand2_1 _08248_ (.Y(_02759_),
    .A(net1857),
    .B(net1130));
 sg13g2_o21ai_1 _08249_ (.B1(_02759_),
    .Y(_00411_),
    .A1(_00211_),
    .A2(net1129));
 sg13g2_nand2_1 _08250_ (.Y(_02760_),
    .A(net1885),
    .B(net1130));
 sg13g2_o21ai_1 _08251_ (.B1(_02760_),
    .Y(_00412_),
    .A1(_00205_),
    .A2(net1130));
 sg13g2_nand2_1 _08252_ (.Y(_02761_),
    .A(net1833),
    .B(net1130));
 sg13g2_o21ai_1 _08253_ (.B1(_02761_),
    .Y(_00413_),
    .A1(_00206_),
    .A2(net1130));
 sg13g2_nand2_1 _08254_ (.Y(_02762_),
    .A(net1839),
    .B(net1128));
 sg13g2_o21ai_1 _08255_ (.B1(_02762_),
    .Y(_00414_),
    .A1(_00212_),
    .A2(net1129));
 sg13g2_nand2_1 _08256_ (.Y(_02763_),
    .A(net1883),
    .B(net1129));
 sg13g2_o21ai_1 _08257_ (.B1(_02763_),
    .Y(_00415_),
    .A1(_00207_),
    .A2(net1129));
 sg13g2_nand3b_1 _08258_ (.B(_02658_),
    .C(_02678_),
    .Y(_02764_),
    .A_N(net1319));
 sg13g2_nand2b_1 _08259_ (.Y(_02765_),
    .B(net1454),
    .A_N(\i_spi.data[0] ));
 sg13g2_o21ai_1 _08260_ (.B1(_02765_),
    .Y(_02766_),
    .A1(\data_to_write[1] ),
    .A2(net1454));
 sg13g2_nand2_1 _08261_ (.Y(_02767_),
    .A(net2001),
    .B(net1183));
 sg13g2_o21ai_1 _08262_ (.B1(_02767_),
    .Y(_00416_),
    .A1(net1183),
    .A2(_02766_));
 sg13g2_nand2b_1 _08263_ (.Y(_02768_),
    .B(net1454),
    .A_N(net2001));
 sg13g2_o21ai_1 _08264_ (.B1(_02768_),
    .Y(_02769_),
    .A1(\data_to_write[2] ),
    .A2(net1454));
 sg13g2_nand2_1 _08265_ (.Y(_02770_),
    .A(net2039),
    .B(net1183));
 sg13g2_o21ai_1 _08266_ (.B1(_02770_),
    .Y(_00417_),
    .A1(net1183),
    .A2(_02769_));
 sg13g2_nand2b_1 _08267_ (.Y(_02771_),
    .B(net1456),
    .A_N(\i_spi.data[2] ));
 sg13g2_o21ai_1 _08268_ (.B1(_02771_),
    .Y(_02772_),
    .A1(net1453),
    .A2(\data_to_write[3] ));
 sg13g2_nand2_1 _08269_ (.Y(_02773_),
    .A(net1997),
    .B(net1182));
 sg13g2_o21ai_1 _08270_ (.B1(_02773_),
    .Y(_00418_),
    .A1(net1182),
    .A2(_02772_));
 sg13g2_nand2b_1 _08271_ (.Y(_02774_),
    .B(net1453),
    .A_N(\i_spi.data[3] ));
 sg13g2_o21ai_1 _08272_ (.B1(_02774_),
    .Y(_02775_),
    .A1(net1453),
    .A2(\data_to_write[4] ));
 sg13g2_nand2_1 _08273_ (.Y(_02776_),
    .A(net1952),
    .B(net1182));
 sg13g2_o21ai_1 _08274_ (.B1(_02776_),
    .Y(_00419_),
    .A1(net1182),
    .A2(_02775_));
 sg13g2_nand2b_1 _08275_ (.Y(_02777_),
    .B(net1453),
    .A_N(net1952));
 sg13g2_o21ai_1 _08276_ (.B1(_02777_),
    .Y(_02778_),
    .A1(net1453),
    .A2(\data_to_write[5] ));
 sg13g2_nand2_1 _08277_ (.Y(_02779_),
    .A(net2005),
    .B(net1182));
 sg13g2_o21ai_1 _08278_ (.B1(_02779_),
    .Y(_00420_),
    .A1(net1182),
    .A2(_02778_));
 sg13g2_nand2b_1 _08279_ (.Y(_02780_),
    .B(net1453),
    .A_N(\i_spi.data[5] ));
 sg13g2_o21ai_1 _08280_ (.B1(_02780_),
    .Y(_02781_),
    .A1(net1453),
    .A2(\data_to_write[6] ));
 sg13g2_nand2_1 _08281_ (.Y(_02782_),
    .A(net1993),
    .B(net1183));
 sg13g2_o21ai_1 _08282_ (.B1(_02782_),
    .Y(_00421_),
    .A1(net1183),
    .A2(_02781_));
 sg13g2_nand2b_1 _08283_ (.Y(_02783_),
    .B(net1456),
    .A_N(\i_spi.data[6] ));
 sg13g2_o21ai_1 _08284_ (.B1(_02783_),
    .Y(_02784_),
    .A1(net1453),
    .A2(\data_to_write[7] ));
 sg13g2_nand2_1 _08285_ (.Y(_02785_),
    .A(net1959),
    .B(net1182));
 sg13g2_o21ai_1 _08286_ (.B1(_02785_),
    .Y(_00422_),
    .A1(net1182),
    .A2(_02784_));
 sg13g2_nor2_1 _08287_ (.A(net1457),
    .B(net1247),
    .Y(_02786_));
 sg13g2_nor2_1 _08288_ (.A(net2233),
    .B(net1224),
    .Y(_02787_));
 sg13g2_nand2b_1 _08289_ (.Y(_02788_),
    .B(net1298),
    .A_N(\i_core.cpu.i_core.i_shift.a[4] ));
 sg13g2_o21ai_1 _08290_ (.B1(_02788_),
    .Y(_02789_),
    .A1(\i_core.cpu.i_core.mepc[0] ),
    .A2(net1298));
 sg13g2_a21oi_1 _08291_ (.A1(net1224),
    .A2(_02789_),
    .Y(_00423_),
    .B1(_02787_));
 sg13g2_and2_1 _08292_ (.A(\i_core.cpu.i_core.i_shift.a[5] ),
    .B(net1299),
    .X(_02790_));
 sg13g2_a21oi_2 _08293_ (.B1(_02790_),
    .Y(_02791_),
    .A2(net1274),
    .A1(\i_core.cpu.i_core.mepc[1] ));
 sg13g2_nor2_1 _08294_ (.A(net2051),
    .B(net1227),
    .Y(_02792_));
 sg13g2_a21oi_1 _08295_ (.A1(net1224),
    .A2(_02791_),
    .Y(_00424_),
    .B1(_02792_));
 sg13g2_and2_1 _08296_ (.A(\i_core.cpu.i_core.i_shift.a[6] ),
    .B(net1299),
    .X(_02793_));
 sg13g2_a21oi_2 _08297_ (.B1(_02793_),
    .Y(_02794_),
    .A2(net1274),
    .A1(\i_core.cpu.i_core.mepc[2] ));
 sg13g2_nor2_1 _08298_ (.A(net1452),
    .B(net1223),
    .Y(_02795_));
 sg13g2_a21oi_1 _08299_ (.A1(net1223),
    .A2(_02794_),
    .Y(_00425_),
    .B1(_02795_));
 sg13g2_and2_1 _08300_ (.A(\i_core.cpu.i_core.i_shift.a[7] ),
    .B(net1299),
    .X(_02796_));
 sg13g2_a21oi_2 _08301_ (.B1(_02796_),
    .Y(_02797_),
    .A2(net1274),
    .A1(\i_core.cpu.i_core.mepc[3] ));
 sg13g2_nor2_1 _08302_ (.A(net2098),
    .B(net1224),
    .Y(_02798_));
 sg13g2_a21oi_1 _08303_ (.A1(net1224),
    .A2(_02797_),
    .Y(_00426_),
    .B1(_02798_));
 sg13g2_and2_1 _08304_ (.A(\i_core.cpu.i_core.i_shift.a[8] ),
    .B(net1295),
    .X(_02799_));
 sg13g2_a21oi_2 _08305_ (.B1(_02799_),
    .Y(_02800_),
    .A2(net1275),
    .A1(net2335));
 sg13g2_nor2_1 _08306_ (.A(net2449),
    .B(net1225),
    .Y(_02801_));
 sg13g2_a21oi_1 _08307_ (.A1(net1225),
    .A2(_02800_),
    .Y(_00427_),
    .B1(_02801_));
 sg13g2_and2_1 _08308_ (.A(\i_core.cpu.i_core.i_shift.a[9] ),
    .B(net1295),
    .X(_02802_));
 sg13g2_a21oi_2 _08309_ (.B1(_02802_),
    .Y(_02803_),
    .A2(net1275),
    .A1(net2346));
 sg13g2_nor2_1 _08310_ (.A(net2444),
    .B(net1225),
    .Y(_02804_));
 sg13g2_a21oi_1 _08311_ (.A1(net1226),
    .A2(_02803_),
    .Y(_00428_),
    .B1(_02804_));
 sg13g2_nor2_1 _08312_ (.A(net2136),
    .B(net1227),
    .Y(_02805_));
 sg13g2_nand2b_1 _08313_ (.Y(_02806_),
    .B(net1297),
    .A_N(\i_core.cpu.i_core.i_shift.a[10] ));
 sg13g2_o21ai_1 _08314_ (.B1(_02806_),
    .Y(_02807_),
    .A1(\i_core.cpu.i_core.mepc[6] ),
    .A2(net1298));
 sg13g2_a21oi_1 _08315_ (.A1(net1224),
    .A2(_02807_),
    .Y(_00429_),
    .B1(_02805_));
 sg13g2_nor2_1 _08316_ (.A(net2153),
    .B(net1224),
    .Y(_02808_));
 sg13g2_nand2b_1 _08317_ (.Y(_02809_),
    .B(net1297),
    .A_N(\i_core.cpu.i_core.i_shift.a[11] ));
 sg13g2_o21ai_1 _08318_ (.B1(_02809_),
    .Y(_02810_),
    .A1(\i_core.cpu.i_core.mepc[7] ),
    .A2(net1297));
 sg13g2_a21oi_1 _08319_ (.A1(net1224),
    .A2(_02810_),
    .Y(_00430_),
    .B1(_02808_));
 sg13g2_nor2_1 _08320_ (.A(net2434),
    .B(net1225),
    .Y(_02811_));
 sg13g2_nand2b_1 _08321_ (.Y(_02812_),
    .B(net1295),
    .A_N(\i_core.cpu.i_core.i_shift.a[12] ));
 sg13g2_o21ai_1 _08322_ (.B1(_02812_),
    .Y(_02813_),
    .A1(\i_core.cpu.i_core.mepc[8] ),
    .A2(net1295));
 sg13g2_a21oi_1 _08323_ (.A1(net1225),
    .A2(_02813_),
    .Y(_00431_),
    .B1(_02811_));
 sg13g2_and2_1 _08324_ (.A(\i_core.cpu.i_core.i_shift.a[13] ),
    .B(net1296),
    .X(_02814_));
 sg13g2_a21oi_2 _08325_ (.B1(_02814_),
    .Y(_02815_),
    .A2(net1275),
    .A1(net2269));
 sg13g2_nor2_1 _08326_ (.A(net2388),
    .B(net1225),
    .Y(_02816_));
 sg13g2_a21oi_1 _08327_ (.A1(net1225),
    .A2(_02815_),
    .Y(_00432_),
    .B1(_02816_));
 sg13g2_nor2_1 _08328_ (.A(net2429),
    .B(net1226),
    .Y(_02817_));
 sg13g2_nand2b_1 _08329_ (.Y(_02818_),
    .B(net1297),
    .A_N(\i_core.cpu.i_core.i_shift.a[14] ));
 sg13g2_o21ai_1 _08330_ (.B1(_02818_),
    .Y(_02819_),
    .A1(\i_core.cpu.i_core.mepc[10] ),
    .A2(net1297));
 sg13g2_a21oi_1 _08331_ (.A1(net1225),
    .A2(_02819_),
    .Y(_00433_),
    .B1(_02817_));
 sg13g2_and2_1 _08332_ (.A(\i_core.cpu.i_core.i_shift.a[15] ),
    .B(net1297),
    .X(_02820_));
 sg13g2_a21oi_2 _08333_ (.B1(_02820_),
    .Y(_02821_),
    .A2(net1275),
    .A1(net2043));
 sg13g2_nor2_1 _08334_ (.A(net2391),
    .B(net1226),
    .Y(_02822_));
 sg13g2_a21oi_1 _08335_ (.A1(net1226),
    .A2(_02821_),
    .Y(_00434_),
    .B1(_02822_));
 sg13g2_nor2_1 _08336_ (.A(net2302),
    .B(net1226),
    .Y(_02823_));
 sg13g2_nand2b_1 _08337_ (.Y(_02824_),
    .B(net1295),
    .A_N(\i_core.cpu.i_core.i_shift.a[16] ));
 sg13g2_o21ai_1 _08338_ (.B1(_02824_),
    .Y(_02825_),
    .A1(\i_core.cpu.i_core.mepc[12] ),
    .A2(net1295));
 sg13g2_a21oi_1 _08339_ (.A1(net1226),
    .A2(_02825_),
    .Y(_00435_),
    .B1(_02823_));
 sg13g2_and2_1 _08340_ (.A(net2216),
    .B(net1296),
    .X(_02826_));
 sg13g2_a21oi_2 _08341_ (.B1(_02826_),
    .Y(_02827_),
    .A2(net1275),
    .A1(net2208));
 sg13g2_nor2_1 _08342_ (.A(net2267),
    .B(net1221),
    .Y(_02828_));
 sg13g2_a21oi_1 _08343_ (.A1(net1221),
    .A2(_02827_),
    .Y(_00436_),
    .B1(_02828_));
 sg13g2_nor2_1 _08344_ (.A(net2186),
    .B(net1226),
    .Y(_02829_));
 sg13g2_nand2b_1 _08345_ (.Y(_02830_),
    .B(net1297),
    .A_N(\i_core.cpu.i_core.i_shift.a[18] ));
 sg13g2_o21ai_1 _08346_ (.B1(_02830_),
    .Y(_02831_),
    .A1(\i_core.cpu.i_core.mepc[14] ),
    .A2(net1297));
 sg13g2_a21oi_1 _08347_ (.A1(net1222),
    .A2(_02831_),
    .Y(_00437_),
    .B1(_02829_));
 sg13g2_and2_1 _08348_ (.A(\i_core.cpu.i_core.i_shift.a[19] ),
    .B(net1296),
    .X(_02832_));
 sg13g2_a21oi_2 _08349_ (.B1(_02832_),
    .Y(_02833_),
    .A2(net1274),
    .A1(\i_core.cpu.i_core.mepc[15] ));
 sg13g2_nor2_1 _08350_ (.A(net2230),
    .B(net1221),
    .Y(_02834_));
 sg13g2_a21oi_1 _08351_ (.A1(net1221),
    .A2(_02833_),
    .Y(_00438_),
    .B1(_02834_));
 sg13g2_nor2_1 _08352_ (.A(net2256),
    .B(net1221),
    .Y(_02835_));
 sg13g2_nand2b_1 _08353_ (.Y(_02836_),
    .B(net1295),
    .A_N(\i_core.cpu.i_core.i_shift.a[20] ));
 sg13g2_o21ai_1 _08354_ (.B1(_02836_),
    .Y(_02837_),
    .A1(\i_core.cpu.i_core.mepc[16] ),
    .A2(net1295));
 sg13g2_a21oi_1 _08355_ (.A1(net1221),
    .A2(_02837_),
    .Y(_00439_),
    .B1(_02835_));
 sg13g2_and2_1 _08356_ (.A(net2145),
    .B(net1298),
    .X(_02838_));
 sg13g2_a21oi_2 _08357_ (.B1(_02838_),
    .Y(_02839_),
    .A2(net1275),
    .A1(net2235));
 sg13g2_nor2_1 _08358_ (.A(net2244),
    .B(net1221),
    .Y(_02840_));
 sg13g2_a21oi_1 _08359_ (.A1(net1221),
    .A2(_02839_),
    .Y(_00440_),
    .B1(_02840_));
 sg13g2_nor2_1 _08360_ (.A(net2140),
    .B(net1222),
    .Y(_02841_));
 sg13g2_nand2b_1 _08361_ (.Y(_02842_),
    .B(net1298),
    .A_N(\i_core.cpu.i_core.i_shift.a[22] ));
 sg13g2_o21ai_1 _08362_ (.B1(_02842_),
    .Y(_02843_),
    .A1(\i_core.cpu.i_core.mepc[18] ),
    .A2(net1298));
 sg13g2_a21oi_1 _08363_ (.A1(net1222),
    .A2(_02843_),
    .Y(_00441_),
    .B1(_02841_));
 sg13g2_nor2_1 _08364_ (.A(net2382),
    .B(net1222),
    .Y(_02844_));
 sg13g2_nand2b_1 _08365_ (.Y(_02845_),
    .B(net1298),
    .A_N(\i_core.cpu.i_core.i_shift.a[23] ));
 sg13g2_o21ai_1 _08366_ (.B1(_02845_),
    .Y(_02846_),
    .A1(\i_core.cpu.i_core.mepc[19] ),
    .A2(net1298));
 sg13g2_a21oi_1 _08367_ (.A1(net1222),
    .A2(_02846_),
    .Y(_00442_),
    .B1(_02844_));
 sg13g2_and2_1 _08368_ (.A(\i_core.cpu.i_core.i_shift.a[24] ),
    .B(net1299),
    .X(_02847_));
 sg13g2_a21oi_2 _08369_ (.B1(_02847_),
    .Y(_02848_),
    .A2(net1274),
    .A1(net2686));
 sg13g2_nor2_1 _08370_ (.A(net2172),
    .B(net1220),
    .Y(_02849_));
 sg13g2_a21oi_1 _08371_ (.A1(net1220),
    .A2(_02848_),
    .Y(_00443_),
    .B1(_02849_));
 sg13g2_and2_1 _08372_ (.A(net2178),
    .B(net1299),
    .X(_02850_));
 sg13g2_a21oi_2 _08373_ (.B1(_02850_),
    .Y(_02851_),
    .A2(net1275),
    .A1(\i_core.cpu.i_core.mepc[21] ));
 sg13g2_nor2_1 _08374_ (.A(net2205),
    .B(net1220),
    .Y(_02852_));
 sg13g2_a21oi_1 _08375_ (.A1(net1220),
    .A2(_02851_),
    .Y(_00444_),
    .B1(_02852_));
 sg13g2_and2_1 _08376_ (.A(\i_core.cpu.i_core.i_shift.a[26] ),
    .B(net1299),
    .X(_02853_));
 sg13g2_a21oi_2 _08377_ (.B1(_02853_),
    .Y(_02854_),
    .A2(net1274),
    .A1(\i_core.cpu.i_core.mepc[22] ));
 sg13g2_nor2_1 _08378_ (.A(net2198),
    .B(net1220),
    .Y(_02855_));
 sg13g2_a21oi_1 _08379_ (.A1(net1220),
    .A2(_02854_),
    .Y(_00445_),
    .B1(_02855_));
 sg13g2_and2_1 _08380_ (.A(\i_core.cpu.i_core.i_shift.a[27] ),
    .B(net1299),
    .X(_02856_));
 sg13g2_a21oi_2 _08381_ (.B1(_02856_),
    .Y(_02857_),
    .A2(net1274),
    .A1(\i_core.cpu.i_core.mepc[23] ));
 sg13g2_nor2_1 _08382_ (.A(net2110),
    .B(net1220),
    .Y(_02858_));
 sg13g2_a21oi_1 _08383_ (.A1(net1220),
    .A2(_02857_),
    .Y(_00446_),
    .B1(_02858_));
 sg13g2_nor2_2 _08384_ (.A(net1274),
    .B(_02069_),
    .Y(_02859_));
 sg13g2_a22oi_1 _08385_ (.Y(_02860_),
    .B1(_02859_),
    .B2(net2301),
    .A2(net1247),
    .A1(net2415));
 sg13g2_nor2_1 _08386_ (.A(net1386),
    .B(_02860_),
    .Y(_00447_));
 sg13g2_a22oi_1 _08387_ (.Y(_02861_),
    .B1(_02859_),
    .B2(net2250),
    .A2(net1247),
    .A1(net2331));
 sg13g2_nor2_1 _08388_ (.A(net1386),
    .B(_02861_),
    .Y(_00448_));
 sg13g2_a22oi_1 _08389_ (.Y(_02862_),
    .B1(_02859_),
    .B2(\i_core.cpu.i_core.i_shift.a[30] ),
    .A2(net1247),
    .A1(net2430));
 sg13g2_nor2_1 _08390_ (.A(net1386),
    .B(net2431),
    .Y(_00449_));
 sg13g2_a22oi_1 _08391_ (.Y(_02863_),
    .B1(_02859_),
    .B2(\i_core.cpu.i_core.i_shift.a[31] ),
    .A2(net1247),
    .A1(net2405));
 sg13g2_nor2_1 _08392_ (.A(net1385),
    .B(net2406),
    .Y(_00450_));
 sg13g2_mux2_1 _08393_ (.A0(\i_core.cpu.instr_data_in[2] ),
    .A1(net2265),
    .S(net1154),
    .X(_00451_));
 sg13g2_mux2_1 _08394_ (.A0(\i_core.cpu.instr_data_in[3] ),
    .A1(net2221),
    .S(net1152),
    .X(_00452_));
 sg13g2_mux2_1 _08395_ (.A0(\i_core.cpu.instr_data_in[4] ),
    .A1(net2077),
    .S(net1154),
    .X(_00453_));
 sg13g2_mux2_1 _08396_ (.A0(\i_core.cpu.instr_data_in[5] ),
    .A1(net2056),
    .S(net1153),
    .X(_00454_));
 sg13g2_mux2_1 _08397_ (.A0(\i_core.cpu.instr_data_in[6] ),
    .A1(net2117),
    .S(net1152),
    .X(_00455_));
 sg13g2_mux2_1 _08398_ (.A0(\i_core.cpu.instr_data_in[7] ),
    .A1(net2075),
    .S(net1153),
    .X(_00456_));
 sg13g2_nand2_1 _08399_ (.Y(_02864_),
    .A(net1837),
    .B(net1152));
 sg13g2_o21ai_1 _08400_ (.B1(_02864_),
    .Y(_00457_),
    .A1(_00208_),
    .A2(net1152));
 sg13g2_nand2_1 _08401_ (.Y(_02865_),
    .A(net1851),
    .B(net1152));
 sg13g2_o21ai_1 _08402_ (.B1(_02865_),
    .Y(_00458_),
    .A1(_00209_),
    .A2(net1152));
 sg13g2_nand2_1 _08403_ (.Y(_02866_),
    .A(net1859),
    .B(_02733_));
 sg13g2_o21ai_1 _08404_ (.B1(_02866_),
    .Y(_00459_),
    .A1(_00210_),
    .A2(net1154));
 sg13g2_nand2_1 _08405_ (.Y(_02867_),
    .A(net1878),
    .B(net1153));
 sg13g2_o21ai_1 _08406_ (.B1(_02867_),
    .Y(_00460_),
    .A1(_00211_),
    .A2(net1152));
 sg13g2_nand2_1 _08407_ (.Y(_02868_),
    .A(net1847),
    .B(net1154));
 sg13g2_o21ai_1 _08408_ (.B1(_02868_),
    .Y(_00461_),
    .A1(_00205_),
    .A2(net1154));
 sg13g2_nand2_1 _08409_ (.Y(_02869_),
    .A(net1835),
    .B(net1154));
 sg13g2_o21ai_1 _08410_ (.B1(_02869_),
    .Y(_00462_),
    .A1(_00206_),
    .A2(net1154));
 sg13g2_nand2_1 _08411_ (.Y(_02870_),
    .A(net1841),
    .B(net1153));
 sg13g2_o21ai_1 _08412_ (.B1(_02870_),
    .Y(_00463_),
    .A1(_00212_),
    .A2(net1153));
 sg13g2_nand2_1 _08413_ (.Y(_02871_),
    .A(net1861),
    .B(net1153));
 sg13g2_o21ai_1 _08414_ (.B1(_02871_),
    .Y(_00464_),
    .A1(_00207_),
    .A2(net1152));
 sg13g2_mux2_1 _08415_ (.A0(\i_core.cpu.i_core.mepc[0] ),
    .A1(net2335),
    .S(net1350),
    .X(_00465_));
 sg13g2_mux2_1 _08416_ (.A0(\i_core.cpu.i_core.mepc[1] ),
    .A1(net2346),
    .S(net1353),
    .X(_00466_));
 sg13g2_mux2_1 _08417_ (.A0(net2364),
    .A1(net2355),
    .S(net1351),
    .X(_00467_));
 sg13g2_mux2_1 _08418_ (.A0(\i_core.cpu.i_core.mepc[3] ),
    .A1(net2352),
    .S(net1351),
    .X(_00468_));
 sg13g2_mux2_1 _08419_ (.A0(\i_core.cpu.i_core.mepc[4] ),
    .A1(net2228),
    .S(net1350),
    .X(_00469_));
 sg13g2_mux2_1 _08420_ (.A0(\i_core.cpu.i_core.mepc[5] ),
    .A1(net2269),
    .S(net1350),
    .X(_00470_));
 sg13g2_mux2_1 _08421_ (.A0(net2355),
    .A1(\i_core.cpu.i_core.mepc[10] ),
    .S(net1351),
    .X(_00471_));
 sg13g2_mux2_1 _08422_ (.A0(\i_core.cpu.i_core.mepc[7] ),
    .A1(net2043),
    .S(net1351),
    .X(_00472_));
 sg13g2_mux2_1 _08423_ (.A0(\i_core.cpu.i_core.mepc[8] ),
    .A1(net2151),
    .S(net1350),
    .X(_00473_));
 sg13g2_mux2_1 _08424_ (.A0(\i_core.cpu.i_core.mepc[9] ),
    .A1(net2208),
    .S(net1351),
    .X(_00474_));
 sg13g2_mux2_1 _08425_ (.A0(\i_core.cpu.i_core.mepc[10] ),
    .A1(net2260),
    .S(net1351),
    .X(_00475_));
 sg13g2_mux2_1 _08426_ (.A0(net2043),
    .A1(net2251),
    .S(net1350),
    .X(_00476_));
 sg13g2_mux2_1 _08427_ (.A0(net2151),
    .A1(net2173),
    .S(net1350),
    .X(_00477_));
 sg13g2_mux2_1 _08428_ (.A0(net2208),
    .A1(net2235),
    .S(net1350),
    .X(_00478_));
 sg13g2_mux2_1 _08429_ (.A0(\i_core.cpu.i_core.mepc[14] ),
    .A1(net2166),
    .S(net1351),
    .X(_00479_));
 sg13g2_mux2_1 _08430_ (.A0(net2251),
    .A1(net2126),
    .S(net1352),
    .X(_00480_));
 sg13g2_mux2_1 _08431_ (.A0(net2173),
    .A1(\i_core.cpu.i_core.mepc[20] ),
    .S(net1350),
    .X(_00481_));
 sg13g2_nor2_1 _08432_ (.A(net2235),
    .B(net1352),
    .Y(_02872_));
 sg13g2_a21oi_1 _08433_ (.A1(_00842_),
    .A2(net1352),
    .Y(_00482_),
    .B1(_02872_));
 sg13g2_mux2_1 _08434_ (.A0(net2166),
    .A1(net2259),
    .S(net1352),
    .X(_00483_));
 sg13g2_nor2_1 _08435_ (.A(net2126),
    .B(net1352),
    .Y(_02873_));
 sg13g2_a21oi_1 _08436_ (.A1(_00843_),
    .A2(net1352),
    .Y(_00484_),
    .B1(_02873_));
 sg13g2_nand2_2 _08437_ (.Y(_02874_),
    .A(net1278),
    .B(_02067_));
 sg13g2_mux2_2 _08438_ (.A0(_01102_),
    .A1(_01122_),
    .S(_01170_),
    .X(_02875_));
 sg13g2_mux2_1 _08439_ (.A0(_02875_),
    .A1(net1444),
    .S(_02874_),
    .X(_00485_));
 sg13g2_nor2_1 _08440_ (.A(_01071_),
    .B(_01170_),
    .Y(_02876_));
 sg13g2_a21oi_2 _08441_ (.B1(_02876_),
    .Y(_02877_),
    .A2(_01170_),
    .A1(_01065_));
 sg13g2_nor2_1 _08442_ (.A(_02874_),
    .B(_02877_),
    .Y(_02878_));
 sg13g2_a21oi_1 _08443_ (.A1(net1370),
    .A2(_02874_),
    .Y(_00486_),
    .B1(_02878_));
 sg13g2_o21ai_1 _08444_ (.B1(_01170_),
    .Y(_02879_),
    .A1(_01027_),
    .A2(_01029_));
 sg13g2_o21ai_1 _08445_ (.B1(_02879_),
    .Y(_02880_),
    .A1(_01013_),
    .A2(_01170_));
 sg13g2_mux2_1 _08446_ (.A0(_02880_),
    .A1(net2576),
    .S(_02874_),
    .X(_00487_));
 sg13g2_nor2b_1 _08447_ (.A(_00965_),
    .B_N(_01170_),
    .Y(_02881_));
 sg13g2_a21oi_2 _08448_ (.B1(_01170_),
    .Y(_02882_),
    .A2(_00973_),
    .A1(_00969_));
 sg13g2_nor3_2 _08449_ (.A(_02874_),
    .B(_02881_),
    .C(_02882_),
    .Y(_02883_));
 sg13g2_a21o_1 _08450_ (.A2(_02874_),
    .A1(net2268),
    .B1(_02883_),
    .X(_00488_));
 sg13g2_nor3_1 _08451_ (.A(net2451),
    .B(net1457),
    .C(net1150),
    .Y(_02884_));
 sg13g2_a21oi_1 _08452_ (.A1(_00825_),
    .A2(net1149),
    .Y(_00489_),
    .B1(_02884_));
 sg13g2_nor3_1 _08453_ (.A(net2403),
    .B(net1457),
    .C(net1150),
    .Y(_02885_));
 sg13g2_a21oi_1 _08454_ (.A1(_00831_),
    .A2(net1150),
    .Y(_00490_),
    .B1(_02885_));
 sg13g2_a21oi_1 _08455_ (.A1(_01482_),
    .A2(_01490_),
    .Y(_02886_),
    .B1(net1319));
 sg13g2_nand2_1 _08456_ (.Y(_02887_),
    .A(\data_to_write[0] ),
    .B(net1324));
 sg13g2_o21ai_1 _08457_ (.B1(_02887_),
    .Y(_02888_),
    .A1(net1324),
    .A2(_00837_));
 sg13g2_mux2_1 _08458_ (.A0(_02888_),
    .A1(net2620),
    .S(_02886_),
    .X(_00491_));
 sg13g2_nor2_1 _08459_ (.A(\i_core.mem.qspi_data_byte_idx[1] ),
    .B(\i_core.mem.qspi_data_byte_idx[0] ),
    .Y(_02889_));
 sg13g2_nand3_1 _08460_ (.B(_01856_),
    .C(_02889_),
    .A(_01430_),
    .Y(_02890_));
 sg13g2_xor2_1 _08461_ (.B(_01190_),
    .A(net1437),
    .X(_02891_));
 sg13g2_xor2_1 _08462_ (.B(net1437),
    .A(\i_core.mem.qspi_data_byte_idx[1] ),
    .X(_02892_));
 sg13g2_xor2_1 _08463_ (.B(_02892_),
    .A(_01187_),
    .X(_02893_));
 sg13g2_and2_1 _08464_ (.A(\i_core.mem.q_ctrl.data_req ),
    .B(_02893_),
    .X(_02894_));
 sg13g2_a22oi_1 _08465_ (.Y(_02895_),
    .B1(_02891_),
    .B2(_02894_),
    .A2(_02890_),
    .A1(\i_core.mem.data_stall ));
 sg13g2_a21oi_1 _08466_ (.A1(_01428_),
    .A2(_02895_),
    .Y(_00492_),
    .B1(_00822_));
 sg13g2_nand2_1 _08467_ (.Y(_02896_),
    .A(\i_core.cpu.i_core.i_shift.a[15] ),
    .B(net1217));
 sg13g2_o21ai_1 _08468_ (.B1(_02309_),
    .Y(_02897_),
    .A1(_02286_),
    .A2(_02307_));
 sg13g2_and2_1 _08469_ (.A(\i_core.cpu.i_core.i_shift.a[14] ),
    .B(net1232),
    .X(_02898_));
 sg13g2_nand2b_1 _08470_ (.Y(_02899_),
    .B(_02898_),
    .A_N(_02306_));
 sg13g2_xnor2_1 _08471_ (.Y(_02900_),
    .A(_02306_),
    .B(_02898_));
 sg13g2_and2_1 _08472_ (.A(_02897_),
    .B(_02900_),
    .X(_02901_));
 sg13g2_xor2_1 _08473_ (.B(_02900_),
    .A(_02897_),
    .X(_02902_));
 sg13g2_nor2b_1 _08474_ (.A(_02896_),
    .B_N(_02902_),
    .Y(_02903_));
 sg13g2_xnor2_1 _08475_ (.Y(_02904_),
    .A(_02896_),
    .B(_02902_));
 sg13g2_o21ai_1 _08476_ (.B1(_02311_),
    .Y(_02905_),
    .A1(_00872_),
    .A2(_02312_));
 sg13g2_nand2_1 _08477_ (.Y(_02906_),
    .A(_02904_),
    .B(_02905_));
 sg13g2_xor2_1 _08478_ (.B(_02905_),
    .A(_02904_),
    .X(_02907_));
 sg13g2_o21ai_1 _08479_ (.B1(_02314_),
    .Y(_02908_),
    .A1(_02302_),
    .A2(_02315_));
 sg13g2_nand2_1 _08480_ (.Y(_02909_),
    .A(_02907_),
    .B(_02908_));
 sg13g2_xor2_1 _08481_ (.B(_02908_),
    .A(_02907_),
    .X(_02910_));
 sg13g2_a21oi_1 _08482_ (.A1(_02299_),
    .A2(_02301_),
    .Y(_02911_),
    .B1(_02318_));
 sg13g2_o21ai_1 _08483_ (.B1(_02910_),
    .Y(_02912_),
    .A1(_02319_),
    .A2(_02911_));
 sg13g2_or3_1 _08484_ (.A(_02319_),
    .B(_02910_),
    .C(_02911_),
    .X(_02913_));
 sg13g2_and2_1 _08485_ (.A(_02912_),
    .B(_02913_),
    .X(_00493_));
 sg13g2_nand2_1 _08486_ (.Y(_02914_),
    .A(\i_core.cpu.i_core.i_shift.a[15] ),
    .B(net1232));
 sg13g2_nand3_1 _08487_ (.B(net1230),
    .C(_02307_),
    .A(\i_core.cpu.i_core.i_shift.a[14] ),
    .Y(_02915_));
 sg13g2_nand2_1 _08488_ (.Y(_02916_),
    .A(net2409),
    .B(net1230));
 sg13g2_xor2_1 _08489_ (.B(_02915_),
    .A(_02914_),
    .X(_02917_));
 sg13g2_o21ai_1 _08490_ (.B1(_02917_),
    .Y(_02918_),
    .A1(_02901_),
    .A2(_02903_));
 sg13g2_or3_1 _08491_ (.A(_02901_),
    .B(_02903_),
    .C(_02917_),
    .X(_02919_));
 sg13g2_and2_1 _08492_ (.A(_02918_),
    .B(_02919_),
    .X(_02920_));
 sg13g2_nor2b_1 _08493_ (.A(_02906_),
    .B_N(_02920_),
    .Y(_02921_));
 sg13g2_xor2_1 _08494_ (.B(_02920_),
    .A(_02906_),
    .X(_02922_));
 sg13g2_a21oi_1 _08495_ (.A1(_02909_),
    .A2(_02912_),
    .Y(_02923_),
    .B1(_02922_));
 sg13g2_nand3_1 _08496_ (.B(_02912_),
    .C(_02922_),
    .A(_02909_),
    .Y(_02924_));
 sg13g2_nor2b_1 _08497_ (.A(_02923_),
    .B_N(_02924_),
    .Y(_00494_));
 sg13g2_nor2_1 _08498_ (.A(_02898_),
    .B(_02916_),
    .Y(_02925_));
 sg13g2_o21ai_1 _08499_ (.B1(_02918_),
    .Y(_02926_),
    .A1(\i_core.cpu.i_core.i_shift.a[15] ),
    .A2(_02899_));
 sg13g2_xor2_1 _08500_ (.B(_02926_),
    .A(_02925_),
    .X(_02927_));
 sg13g2_o21ai_1 _08501_ (.B1(_02927_),
    .Y(_02928_),
    .A1(_02921_),
    .A2(_02923_));
 sg13g2_or3_1 _08502_ (.A(_02921_),
    .B(_02923_),
    .C(_02927_),
    .X(_02929_));
 sg13g2_and2_1 _08503_ (.A(_02928_),
    .B(_02929_),
    .X(_00495_));
 sg13g2_nor2b_1 _08504_ (.A(_02898_),
    .B_N(_02918_),
    .Y(_02930_));
 sg13g2_o21ai_1 _08505_ (.B1(_02928_),
    .Y(_00496_),
    .A1(_02916_),
    .A2(_02930_));
 sg13g2_nand3_1 _08506_ (.B(_01853_),
    .C(_01860_),
    .A(net2501),
    .Y(_02931_));
 sg13g2_nand2_1 _08507_ (.Y(_02932_),
    .A(_01835_),
    .B(_01855_));
 sg13g2_nor2_1 _08508_ (.A(_02931_),
    .B(_02932_),
    .Y(_02933_));
 sg13g2_nor2_2 _08509_ (.A(_00813_),
    .B(_02933_),
    .Y(_02934_));
 sg13g2_o21ai_1 _08510_ (.B1(_00089_),
    .Y(_02935_),
    .A1(_02931_),
    .A2(_02932_));
 sg13g2_nor3_1 _08511_ (.A(_01188_),
    .B(_02891_),
    .C(_02935_),
    .Y(_02936_));
 sg13g2_a21oi_1 _08512_ (.A1(_01837_),
    .A2(_02935_),
    .Y(_02937_),
    .B1(_02936_));
 sg13g2_nor2b_1 _08513_ (.A(_01862_),
    .B_N(net2537),
    .Y(_02938_));
 sg13g2_a22oi_1 _08514_ (.Y(_02939_),
    .B1(_02937_),
    .B2(_02938_),
    .A2(_01862_),
    .A1(net1437));
 sg13g2_nand2_1 _08515_ (.Y(_02940_),
    .A(_01853_),
    .B(_02932_));
 sg13g2_nand3_1 _08516_ (.B(_01860_),
    .C(_02940_),
    .A(_00151_),
    .Y(_02941_));
 sg13g2_or2_1 _08517_ (.X(_02942_),
    .B(_02931_),
    .A(_01855_));
 sg13g2_and2_2 _08518_ (.A(_02941_),
    .B(_02942_),
    .X(_02943_));
 sg13g2_nand2_1 _08519_ (.Y(_02944_),
    .A(_02941_),
    .B(_02942_));
 sg13g2_nor3_1 _08520_ (.A(_00154_),
    .B(net2538),
    .C(net1125),
    .Y(_00497_));
 sg13g2_nor2b_1 _08521_ (.A(_01862_),
    .B_N(_02892_),
    .Y(_02945_));
 sg13g2_a22oi_1 _08522_ (.Y(_02946_),
    .B1(_02937_),
    .B2(_02945_),
    .A2(_01862_),
    .A1(net2654));
 sg13g2_nor3_1 _08523_ (.A(_00154_),
    .B(net1125),
    .C(_02946_),
    .Y(_00498_));
 sg13g2_nand2_1 _08524_ (.Y(_02947_),
    .A(\i_core.mem.q_ctrl.data_ready ),
    .B(_02889_));
 sg13g2_nor2_1 _08525_ (.A(net2483),
    .B(net1286),
    .Y(_02948_));
 sg13g2_a21oi_1 _08526_ (.A1(_00825_),
    .A2(net1285),
    .Y(_00499_),
    .B1(_02948_));
 sg13g2_nor2_1 _08527_ (.A(net2374),
    .B(net1286),
    .Y(_02949_));
 sg13g2_a21oi_1 _08528_ (.A1(_00831_),
    .A2(net1285),
    .Y(_00500_),
    .B1(_02949_));
 sg13g2_mux2_1 _08529_ (.A0(\i_core.cpu.instr_data_in[10] ),
    .A1(net2626),
    .S(net1285),
    .X(_00501_));
 sg13g2_mux2_1 _08530_ (.A0(net2370),
    .A1(net2564),
    .S(net1287),
    .X(_00502_));
 sg13g2_nand2_1 _08531_ (.Y(_02950_),
    .A(net2552),
    .B(net1285));
 sg13g2_o21ai_1 _08532_ (.B1(_02950_),
    .Y(_00503_),
    .A1(_00827_),
    .A2(net1285));
 sg13g2_nand2_1 _08533_ (.Y(_02951_),
    .A(\i_core.cpu.instr_data_in[5] ),
    .B(net1286));
 sg13g2_o21ai_1 _08534_ (.B1(_02951_),
    .Y(_00504_),
    .A1(_00833_),
    .A2(net1285));
 sg13g2_nand2_1 _08535_ (.Y(_02952_),
    .A(net2411),
    .B(net1285));
 sg13g2_o21ai_1 _08536_ (.B1(_02952_),
    .Y(_00505_),
    .A1(_00835_),
    .A2(net1285));
 sg13g2_nand2_1 _08537_ (.Y(_02953_),
    .A(\i_core.cpu.instr_data_in[7] ),
    .B(net1287));
 sg13g2_o21ai_1 _08538_ (.B1(_02953_),
    .Y(_00506_),
    .A1(_00838_),
    .A2(net1287));
 sg13g2_nand2_2 _08539_ (.Y(_02954_),
    .A(\i_core.mem.q_ctrl.data_ready ),
    .B(_02892_));
 sg13g2_or2_1 _08540_ (.X(_02955_),
    .B(_02889_),
    .A(_00157_));
 sg13g2_nor2_1 _08541_ (.A(_00208_),
    .B(net1282),
    .Y(_02956_));
 sg13g2_nor3_1 _08542_ (.A(_00208_),
    .B(_02954_),
    .C(net1282),
    .Y(_02957_));
 sg13g2_a21o_1 _08543_ (.A2(net1288),
    .A1(net2085),
    .B1(_02957_),
    .X(_00507_));
 sg13g2_nor2_1 _08544_ (.A(_00209_),
    .B(net1282),
    .Y(_02958_));
 sg13g2_nor3_1 _08545_ (.A(_00209_),
    .B(_02954_),
    .C(net1282),
    .Y(_02959_));
 sg13g2_a21o_1 _08546_ (.A2(net1288),
    .A1(net2099),
    .B1(_02959_),
    .X(_00508_));
 sg13g2_nor2_1 _08547_ (.A(_00210_),
    .B(net1283),
    .Y(_02960_));
 sg13g2_nor3_1 _08548_ (.A(_00210_),
    .B(_02954_),
    .C(net1283),
    .Y(_02961_));
 sg13g2_a21o_1 _08549_ (.A2(net1288),
    .A1(net2081),
    .B1(_02961_),
    .X(_00509_));
 sg13g2_nor2_1 _08550_ (.A(_00211_),
    .B(net1284),
    .Y(_02962_));
 sg13g2_nor3_1 _08551_ (.A(_00211_),
    .B(_02954_),
    .C(net1284),
    .Y(_02963_));
 sg13g2_a21o_1 _08552_ (.A2(_01838_),
    .A1(net2124),
    .B1(_02963_),
    .X(_00510_));
 sg13g2_nor2_1 _08553_ (.A(_00205_),
    .B(net1283),
    .Y(_02964_));
 sg13g2_nor3_1 _08554_ (.A(_00205_),
    .B(_02954_),
    .C(net1282),
    .Y(_02965_));
 sg13g2_a21o_1 _08555_ (.A2(net1288),
    .A1(net2058),
    .B1(_02965_),
    .X(_00511_));
 sg13g2_nor2_1 _08556_ (.A(_00206_),
    .B(net1283),
    .Y(_02966_));
 sg13g2_nor3_1 _08557_ (.A(_00206_),
    .B(_02954_),
    .C(net1282),
    .Y(_02967_));
 sg13g2_a21o_1 _08558_ (.A2(net1288),
    .A1(net2055),
    .B1(_02967_),
    .X(_00512_));
 sg13g2_nor2_1 _08559_ (.A(_00212_),
    .B(net1282),
    .Y(_02968_));
 sg13g2_nor3_1 _08560_ (.A(_00212_),
    .B(_02954_),
    .C(net1282),
    .Y(_02969_));
 sg13g2_a21o_1 _08561_ (.A2(net1288),
    .A1(net2053),
    .B1(_02969_),
    .X(_00513_));
 sg13g2_nor2_1 _08562_ (.A(_00207_),
    .B(net1284),
    .Y(_02970_));
 sg13g2_nor3_1 _08563_ (.A(_00207_),
    .B(_02954_),
    .C(net1284),
    .Y(_02971_));
 sg13g2_a21o_1 _08564_ (.A2(_01838_),
    .A1(net2003),
    .B1(_02971_),
    .X(_00514_));
 sg13g2_nand3b_1 _08565_ (.B(\i_core.mem.q_ctrl.data_ready ),
    .C(\i_core.mem.qspi_data_byte_idx[1] ),
    .Y(_02972_),
    .A_N(net1437));
 sg13g2_nand2_1 _08566_ (.Y(_02973_),
    .A(net1888),
    .B(net1331));
 sg13g2_o21ai_1 _08567_ (.B1(_02973_),
    .Y(_00515_),
    .A1(_00208_),
    .A2(net1331));
 sg13g2_nand2_1 _08568_ (.Y(_02974_),
    .A(net1918),
    .B(net1331));
 sg13g2_o21ai_1 _08569_ (.B1(_02974_),
    .Y(_00516_),
    .A1(_00209_),
    .A2(net1331));
 sg13g2_nand2_1 _08570_ (.Y(_02975_),
    .A(net1893),
    .B(net1332));
 sg13g2_o21ai_1 _08571_ (.B1(_02975_),
    .Y(_00517_),
    .A1(_00210_),
    .A2(_02972_));
 sg13g2_nand2_1 _08572_ (.Y(_02976_),
    .A(net1895),
    .B(net1332));
 sg13g2_o21ai_1 _08573_ (.B1(_02976_),
    .Y(_00518_),
    .A1(_00211_),
    .A2(net1332));
 sg13g2_nand2_1 _08574_ (.Y(_02977_),
    .A(net1971),
    .B(net1331));
 sg13g2_o21ai_1 _08575_ (.B1(_02977_),
    .Y(_00519_),
    .A1(_00205_),
    .A2(net1331));
 sg13g2_nand2_1 _08576_ (.Y(_02978_),
    .A(net1904),
    .B(net1331));
 sg13g2_o21ai_1 _08577_ (.B1(_02978_),
    .Y(_00520_),
    .A1(_00206_),
    .A2(net1331));
 sg13g2_nand2_1 _08578_ (.Y(_02979_),
    .A(net1907),
    .B(net1332));
 sg13g2_o21ai_1 _08579_ (.B1(_02979_),
    .Y(_00521_),
    .A1(_00212_),
    .A2(net1332));
 sg13g2_nand2_1 _08580_ (.Y(_02980_),
    .A(net1891),
    .B(net1332));
 sg13g2_o21ai_1 _08581_ (.B1(_02980_),
    .Y(_00522_),
    .A1(_00207_),
    .A2(net1332));
 sg13g2_nand3_1 _08582_ (.B(net1437),
    .C(\i_core.mem.q_ctrl.data_ready ),
    .A(\i_core.mem.qspi_data_byte_idx[1] ),
    .Y(_02981_));
 sg13g2_nor2_2 _08583_ (.A(_00794_),
    .B(_02892_),
    .Y(_02982_));
 sg13g2_a22oi_1 _08584_ (.Y(_02983_),
    .B1(_02982_),
    .B2(_02956_),
    .A2(_02981_),
    .A1(net1963));
 sg13g2_inv_1 _08585_ (.Y(_00523_),
    .A(net1964));
 sg13g2_a22oi_1 _08586_ (.Y(_02984_),
    .B1(_02982_),
    .B2(_02958_),
    .A2(_02981_),
    .A1(net2121));
 sg13g2_inv_1 _08587_ (.Y(_00524_),
    .A(net2122));
 sg13g2_a22oi_1 _08588_ (.Y(_02985_),
    .B1(_02982_),
    .B2(_02960_),
    .A2(_02981_),
    .A1(net2047));
 sg13g2_inv_1 _08589_ (.Y(_00525_),
    .A(net2048));
 sg13g2_a22oi_1 _08590_ (.Y(_02986_),
    .B1(_02982_),
    .B2(_02962_),
    .A2(_02981_),
    .A1(net1984));
 sg13g2_inv_1 _08591_ (.Y(_00526_),
    .A(net1985));
 sg13g2_a22oi_1 _08592_ (.Y(_02987_),
    .B1(_02982_),
    .B2(_02964_),
    .A2(_02981_),
    .A1(net2025));
 sg13g2_inv_1 _08593_ (.Y(_00527_),
    .A(_02987_));
 sg13g2_a22oi_1 _08594_ (.Y(_02988_),
    .B1(_02982_),
    .B2(_02966_),
    .A2(_02981_),
    .A1(net2006));
 sg13g2_inv_1 _08595_ (.Y(_00528_),
    .A(_02988_));
 sg13g2_a22oi_1 _08596_ (.Y(_02989_),
    .B1(_02982_),
    .B2(_02968_),
    .A2(_02981_),
    .A1(net2059));
 sg13g2_inv_1 _08597_ (.Y(_00529_),
    .A(net2060));
 sg13g2_a22oi_1 _08598_ (.Y(_02990_),
    .B1(_02982_),
    .B2(_02970_),
    .A2(_02981_),
    .A1(net1982));
 sg13g2_inv_1 _08599_ (.Y(_00530_),
    .A(net1983));
 sg13g2_nor3_1 _08600_ (.A(net1318),
    .B(_02931_),
    .C(_02932_),
    .Y(_00531_));
 sg13g2_a21oi_1 _08601_ (.A1(net2464),
    .A2(_01861_),
    .Y(_02991_),
    .B1(_02933_));
 sg13g2_nor3_1 _08602_ (.A(net1319),
    .B(_01865_),
    .C(net2465),
    .Y(_00532_));
 sg13g2_nand2b_1 _08603_ (.Y(_02992_),
    .B(_02643_),
    .A_N(net1319));
 sg13g2_nor2_2 _08604_ (.A(_01860_),
    .B(net1123),
    .Y(_02993_));
 sg13g2_nor2_1 _08605_ (.A(net1436),
    .B(\i_core.mem.q_ctrl.read_cycles_count[0] ),
    .Y(_02994_));
 sg13g2_nor3_2 _08606_ (.A(\i_core.mem.q_ctrl.read_cycles_count[1] ),
    .B(\i_core.mem.q_ctrl.read_cycles_count[0] ),
    .C(\i_core.mem.q_ctrl.read_cycles_count[2] ),
    .Y(_02995_));
 sg13g2_nor2_1 _08607_ (.A(net2203),
    .B(_02995_),
    .Y(_02996_));
 sg13g2_and2_2 _08608_ (.A(\i_core.mem.q_ctrl.fsm_state[2] ),
    .B(_02016_),
    .X(_02997_));
 sg13g2_nand2_2 _08609_ (.Y(_02998_),
    .A(net1430),
    .B(_02016_));
 sg13g2_nor2_1 _08610_ (.A(\i_core.mem.q_ctrl.nibbles_remaining[1] ),
    .B(\i_core.mem.q_ctrl.nibbles_remaining[0] ),
    .Y(_02999_));
 sg13g2_nor3_2 _08611_ (.A(net2433),
    .B(net2554),
    .C(net2613),
    .Y(_03000_));
 sg13g2_nand2_2 _08612_ (.Y(_03001_),
    .A(_00769_),
    .B(_02999_));
 sg13g2_nand2_1 _08613_ (.Y(_03002_),
    .A(\i_core.mem.q_ctrl.fsm_state[1] ),
    .B(\i_core.mem.q_ctrl.fsm_state[0] ));
 sg13g2_nand2_1 _08614_ (.Y(_03003_),
    .A(net1431),
    .B(_02023_));
 sg13g2_nand3_1 _08615_ (.B(\i_core.mem.q_ctrl.delay_cycles_cfg[2] ),
    .C(_02023_),
    .A(net1431),
    .Y(_03004_));
 sg13g2_nand2_2 _08616_ (.Y(_03005_),
    .A(_03001_),
    .B(_03004_));
 sg13g2_o21ai_1 _08617_ (.B1(_02023_),
    .Y(_03006_),
    .A1(net1431),
    .A2(_00159_));
 sg13g2_nor2_1 _08618_ (.A(_02995_),
    .B(_03006_),
    .Y(_03007_));
 sg13g2_a21oi_2 _08619_ (.B1(_03007_),
    .Y(_03008_),
    .A2(_03006_),
    .A1(net2617));
 sg13g2_inv_1 _08620_ (.Y(_03009_),
    .A(_03008_));
 sg13g2_nand2_2 _08621_ (.Y(_03010_),
    .A(_03005_),
    .B(_03008_));
 sg13g2_nand2_2 _08622_ (.Y(_03011_),
    .A(net1430),
    .B(_01859_));
 sg13g2_nor2_1 _08623_ (.A(_03010_),
    .B(_03011_),
    .Y(_03012_));
 sg13g2_nor2_1 _08624_ (.A(_02996_),
    .B(_03012_),
    .Y(_03013_));
 sg13g2_nand3_1 _08625_ (.B(\i_core.mem.q_ctrl.delay_cycles_cfg[0] ),
    .C(_01859_),
    .A(net1430),
    .Y(_03014_));
 sg13g2_a21oi_1 _08626_ (.A1(net1333),
    .A2(_03014_),
    .Y(_03015_),
    .B1(_03010_));
 sg13g2_o21ai_1 _08627_ (.B1(_02998_),
    .Y(_03016_),
    .A1(_03013_),
    .A2(_03015_));
 sg13g2_nand2b_2 _08628_ (.Y(_03017_),
    .B(_01850_),
    .A_N(\i_core.mem.data_stall ));
 sg13g2_nor3_2 _08629_ (.A(net1436),
    .B(\i_core.mem.q_ctrl.read_cycles_count[2] ),
    .C(_03017_),
    .Y(_03018_));
 sg13g2_nand2b_1 _08630_ (.Y(_03019_),
    .B(_02997_),
    .A_N(_03018_));
 sg13g2_nand3b_1 _08631_ (.B(net2093),
    .C(_03018_),
    .Y(_03020_),
    .A_N(net1434));
 sg13g2_or2_1 _08632_ (.X(_03021_),
    .B(_03017_),
    .A(net1333));
 sg13g2_nor2_1 _08633_ (.A(_03010_),
    .B(_03021_),
    .Y(_03022_));
 sg13g2_a21oi_1 _08634_ (.A1(_02996_),
    .A2(_03022_),
    .Y(_03023_),
    .B1(_03016_));
 sg13g2_o21ai_1 _08635_ (.B1(_03020_),
    .Y(_03024_),
    .A1(_02996_),
    .A2(_03018_));
 sg13g2_a21oi_1 _08636_ (.A1(_02997_),
    .A2(_03024_),
    .Y(_03025_),
    .B1(_03023_));
 sg13g2_nor2_1 _08637_ (.A(net2510),
    .B(_02993_),
    .Y(_03026_));
 sg13g2_a21oi_1 _08638_ (.A1(_02993_),
    .A2(_03025_),
    .Y(_00533_),
    .B1(_03026_));
 sg13g2_xnor2_1 _08639_ (.Y(_03027_),
    .A(net1436),
    .B(\i_core.mem.q_ctrl.read_cycles_count[0] ));
 sg13g2_o21ai_1 _08640_ (.B1(_03027_),
    .Y(_03028_),
    .A1(net1436),
    .A2(\i_core.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_mux2_1 _08641_ (.A0(_03028_),
    .A1(_00851_),
    .S(_03017_),
    .X(_03029_));
 sg13g2_nor2_1 _08642_ (.A(net1333),
    .B(_03029_),
    .Y(_03030_));
 sg13g2_o21ai_1 _08643_ (.B1(net1333),
    .Y(_03031_),
    .A1(\i_core.mem.q_ctrl.delay_cycles_cfg[1] ),
    .A2(_03011_));
 sg13g2_a21oi_1 _08644_ (.A1(_03011_),
    .A2(_03028_),
    .Y(_03032_),
    .B1(_03031_));
 sg13g2_nor3_1 _08645_ (.A(_03010_),
    .B(_03030_),
    .C(_03032_),
    .Y(_03033_));
 sg13g2_a21o_1 _08646_ (.A2(_03028_),
    .A1(_03010_),
    .B1(_03033_),
    .X(_03034_));
 sg13g2_nor2b_1 _08647_ (.A(net1434),
    .B_N(\i_core.mem.q_ctrl.delay_cycles_cfg[2] ),
    .Y(_03035_));
 sg13g2_a21oi_1 _08648_ (.A1(_03018_),
    .A2(_03035_),
    .Y(_03036_),
    .B1(_02998_));
 sg13g2_a22oi_1 _08649_ (.Y(_03037_),
    .B1(_03036_),
    .B2(_03028_),
    .A2(_03034_),
    .A1(_02998_));
 sg13g2_mux2_1 _08650_ (.A0(net1436),
    .A1(_03037_),
    .S(_02993_),
    .X(_00534_));
 sg13g2_nor2b_1 _08651_ (.A(_02994_),
    .B_N(\i_core.mem.q_ctrl.read_cycles_count[2] ),
    .Y(_03038_));
 sg13g2_a21oi_1 _08652_ (.A1(_03005_),
    .A2(_03008_),
    .Y(_03039_),
    .B1(_03038_));
 sg13g2_or2_1 _08653_ (.X(_03040_),
    .B(_03039_),
    .A(_02997_));
 sg13g2_o21ai_1 _08654_ (.B1(_03019_),
    .Y(_03041_),
    .A1(_03021_),
    .A2(_03040_));
 sg13g2_nand3_1 _08655_ (.B(_02023_),
    .C(_03017_),
    .A(net2551),
    .Y(_03042_));
 sg13g2_mux2_1 _08656_ (.A0(\i_core.mem.q_ctrl.delay_cycles_cfg[2] ),
    .A1(_03038_),
    .S(_03011_),
    .X(_03043_));
 sg13g2_a21oi_1 _08657_ (.A1(net1333),
    .A2(_03043_),
    .Y(_03044_),
    .B1(_03010_));
 sg13g2_a21oi_1 _08658_ (.A1(_03042_),
    .A2(_03044_),
    .Y(_03045_),
    .B1(_03040_));
 sg13g2_a21oi_1 _08659_ (.A1(_03038_),
    .A2(_03041_),
    .Y(_03046_),
    .B1(_03045_));
 sg13g2_nor2_1 _08660_ (.A(net2573),
    .B(_02993_),
    .Y(_03047_));
 sg13g2_a21oi_1 _08661_ (.A1(_02993_),
    .A2(_03046_),
    .Y(_00535_),
    .B1(_03047_));
 sg13g2_nor2_1 _08662_ (.A(_01860_),
    .B(_02997_),
    .Y(_03048_));
 sg13g2_nand2_2 _08663_ (.Y(_03049_),
    .A(_01861_),
    .B(_02998_));
 sg13g2_nor2_1 _08664_ (.A(_03008_),
    .B(_03049_),
    .Y(_03050_));
 sg13g2_nand4_1 _08665_ (.B(_02025_),
    .C(_03000_),
    .A(net1434),
    .Y(_03051_),
    .D(_03050_));
 sg13g2_nor2_1 _08666_ (.A(net1124),
    .B(_03051_),
    .Y(_00536_));
 sg13g2_nand2_1 _08667_ (.Y(_03052_),
    .A(\addr[24] ),
    .B(_02934_));
 sg13g2_nand3_1 _08668_ (.B(_00161_),
    .C(_02934_),
    .A(\addr[24] ),
    .Y(_03053_));
 sg13g2_nor2_1 _08669_ (.A(net2348),
    .B(_03052_),
    .Y(_03054_));
 sg13g2_a21oi_1 _08670_ (.A1(_00821_),
    .A2(_03054_),
    .Y(_03055_),
    .B1(_02943_));
 sg13g2_o21ai_1 _08671_ (.B1(_03055_),
    .Y(_03056_),
    .A1(net2668),
    .A2(_03053_));
 sg13g2_nand2_1 _08672_ (.Y(_03057_),
    .A(_02998_),
    .B(_03005_));
 sg13g2_nor3_1 _08673_ (.A(net1430),
    .B(net1429),
    .C(_03001_),
    .Y(_03058_));
 sg13g2_or2_1 _08674_ (.X(_03059_),
    .B(_03058_),
    .A(_03050_));
 sg13g2_a21oi_2 _08675_ (.B1(_03059_),
    .Y(_03060_),
    .A2(net1112),
    .A1(_03049_));
 sg13g2_nand4_1 _08676_ (.B(_01861_),
    .C(_03004_),
    .A(net2613),
    .Y(_03061_),
    .D(_03060_));
 sg13g2_o21ai_1 _08677_ (.B1(_03061_),
    .Y(_03062_),
    .A1(net2613),
    .A2(_03060_));
 sg13g2_nor2_1 _08678_ (.A(net1124),
    .B(_03062_),
    .Y(_00537_));
 sg13g2_nand2b_1 _08679_ (.Y(_03063_),
    .B(_03004_),
    .A_N(_02999_));
 sg13g2_a21oi_1 _08680_ (.A1(\i_core.mem.q_ctrl.nibbles_remaining[1] ),
    .A2(\i_core.mem.q_ctrl.nibbles_remaining[0] ),
    .Y(_03064_),
    .B1(_03063_));
 sg13g2_o21ai_1 _08681_ (.B1(_02026_),
    .Y(_03065_),
    .A1(_00767_),
    .A2(net1435));
 sg13g2_nand4_1 _08682_ (.B(net1429),
    .C(net1333),
    .A(net1431),
    .Y(_03066_),
    .D(_03065_));
 sg13g2_a21o_1 _08683_ (.A2(_03066_),
    .A1(_03005_),
    .B1(_03064_),
    .X(_03067_));
 sg13g2_o21ai_1 _08684_ (.B1(_03060_),
    .Y(_03068_),
    .A1(_01860_),
    .A2(_03067_));
 sg13g2_o21ai_1 _08685_ (.B1(_03068_),
    .Y(_03069_),
    .A1(net2554),
    .A2(_03060_));
 sg13g2_nor2_1 _08686_ (.A(net1123),
    .B(_03069_),
    .Y(_00538_));
 sg13g2_nand4_1 _08687_ (.B(net1429),
    .C(_02017_),
    .A(_00768_),
    .Y(_03070_),
    .D(_03000_));
 sg13g2_o21ai_1 _08688_ (.B1(_03070_),
    .Y(_03071_),
    .A1(_00769_),
    .A2(_03063_));
 sg13g2_a21oi_2 _08689_ (.B1(_01861_),
    .Y(_03072_),
    .A2(_02934_),
    .A1(\addr[24] ));
 sg13g2_a21oi_1 _08690_ (.A1(_01861_),
    .A2(_03071_),
    .Y(_03073_),
    .B1(_03072_));
 sg13g2_nand2_1 _08691_ (.Y(_03074_),
    .A(_03060_),
    .B(_03073_));
 sg13g2_o21ai_1 _08692_ (.B1(_03074_),
    .Y(_03075_),
    .A1(net2433),
    .A2(_03060_));
 sg13g2_nor2_1 _08693_ (.A(net1123),
    .B(_03075_),
    .Y(_00539_));
 sg13g2_nor2_1 _08694_ (.A(_03052_),
    .B(_03056_),
    .Y(_03076_));
 sg13g2_a22oi_1 _08695_ (.Y(_03077_),
    .B1(_03076_),
    .B2(_02941_),
    .A2(_03056_),
    .A1(net1434));
 sg13g2_nor2_1 _08696_ (.A(net1124),
    .B(net2669),
    .Y(_00540_));
 sg13g2_nand2_1 _08697_ (.Y(_03078_),
    .A(_01861_),
    .B(_03019_));
 sg13g2_o21ai_1 _08698_ (.B1(net2393),
    .Y(_03079_),
    .A1(_02997_),
    .A2(_03022_));
 sg13g2_nor3_1 _08699_ (.A(net1123),
    .B(_03078_),
    .C(net2394),
    .Y(_00541_));
 sg13g2_nand2_1 _08700_ (.Y(_03080_),
    .A(net1112),
    .B(_03078_));
 sg13g2_a21oi_1 _08701_ (.A1(_03001_),
    .A2(_03003_),
    .Y(_03081_),
    .B1(_03009_));
 sg13g2_nor2_2 _08702_ (.A(_02997_),
    .B(_03000_),
    .Y(_03082_));
 sg13g2_nand2_2 _08703_ (.Y(_03083_),
    .A(_02998_),
    .B(_03001_));
 sg13g2_o21ai_1 _08704_ (.B1(_03080_),
    .Y(_03084_),
    .A1(_03049_),
    .A2(_03081_));
 sg13g2_o21ai_1 _08705_ (.B1(_03065_),
    .Y(_03085_),
    .A1(_00850_),
    .A2(_02026_));
 sg13g2_a221oi_1 _08706_ (.B2(net1333),
    .C1(_03049_),
    .B1(_03085_),
    .A1(_03001_),
    .Y(_03086_),
    .A2(_03004_));
 sg13g2_a21oi_1 _08707_ (.A1(_03021_),
    .A2(_03086_),
    .Y(_03087_),
    .B1(_03072_));
 sg13g2_mux2_1 _08708_ (.A0(_03087_),
    .A1(net2679),
    .S(_03084_),
    .X(_03088_));
 sg13g2_nor2b_1 _08709_ (.A(net1123),
    .B_N(_03088_),
    .Y(_00542_));
 sg13g2_nor2b_1 _08710_ (.A(net1431),
    .B_N(_03084_),
    .Y(_03089_));
 sg13g2_o21ai_1 _08711_ (.B1(_00159_),
    .Y(_03090_),
    .A1(\i_core.mem.q_ctrl.delay_cycles_cfg[2] ),
    .A2(\i_core.mem.q_ctrl.delay_cycles_cfg[1] ));
 sg13g2_o21ai_1 _08712_ (.B1(_02026_),
    .Y(_03091_),
    .A1(\i_core.mem.q_ctrl.spi_flash_select ),
    .A2(net1434));
 sg13g2_o21ai_1 _08713_ (.B1(_03091_),
    .Y(_03092_),
    .A1(_02016_),
    .A2(_02017_));
 sg13g2_a21oi_1 _08714_ (.A1(net1334),
    .A2(_03092_),
    .Y(_03093_),
    .B1(_03057_));
 sg13g2_nand2_1 _08715_ (.Y(_03094_),
    .A(_03021_),
    .B(_03093_));
 sg13g2_o21ai_1 _08716_ (.B1(_03094_),
    .Y(_03095_),
    .A1(_02998_),
    .A2(_03090_));
 sg13g2_nor3_1 _08717_ (.A(_03072_),
    .B(_03084_),
    .C(_03095_),
    .Y(_03096_));
 sg13g2_nor3_1 _08718_ (.A(net1123),
    .B(_03089_),
    .C(_03096_),
    .Y(_00543_));
 sg13g2_xnor2_1 _08719_ (.Y(_03097_),
    .A(_00152_),
    .B(_03002_));
 sg13g2_nand3_1 _08720_ (.B(_03091_),
    .C(_03097_),
    .A(net1334),
    .Y(_03098_));
 sg13g2_o21ai_1 _08721_ (.B1(_01861_),
    .Y(_03099_),
    .A1(_03057_),
    .A2(_03098_));
 sg13g2_mux2_1 _08722_ (.A0(_03099_),
    .A1(_00768_),
    .S(_03084_),
    .X(_03100_));
 sg13g2_nor2_1 _08723_ (.A(net1123),
    .B(_03100_),
    .Y(_00544_));
 sg13g2_a21oi_1 _08724_ (.A1(net1906),
    .A2(net1112),
    .Y(_03101_),
    .B1(net1124));
 sg13g2_o21ai_1 _08725_ (.B1(_03101_),
    .Y(_00545_),
    .A1(_03054_),
    .A2(net1112));
 sg13g2_a22oi_1 _08726_ (.Y(_03102_),
    .B1(net1112),
    .B2(net1937),
    .A2(_03055_),
    .A1(_03053_));
 sg13g2_nand2b_1 _08727_ (.Y(_00546_),
    .B(net2328),
    .A_N(net1124));
 sg13g2_a21oi_1 _08728_ (.A1(net2540),
    .A2(net1112),
    .Y(_03103_),
    .B1(net1124));
 sg13g2_nand2b_1 _08729_ (.Y(_00547_),
    .B(_03103_),
    .A_N(_03076_));
 sg13g2_nand2b_1 _08730_ (.Y(_03104_),
    .B(_03048_),
    .A_N(net2376));
 sg13g2_nand3_1 _08731_ (.B(_01860_),
    .C(net1112),
    .A(net2376),
    .Y(_03105_));
 sg13g2_a21oi_1 _08732_ (.A1(_03104_),
    .A2(_03105_),
    .Y(_00548_),
    .B1(net1124));
 sg13g2_and4_1 _08733_ (.A(_02020_),
    .B(net1333),
    .C(_03048_),
    .D(_03081_),
    .X(_03106_));
 sg13g2_o21ai_1 _08734_ (.B1(_00159_),
    .Y(_03107_),
    .A1(\i_core.mem.q_ctrl.spi_flash_select ),
    .A2(net1435));
 sg13g2_nor2b_1 _08735_ (.A(_00158_),
    .B_N(_02026_),
    .Y(_03108_));
 sg13g2_nor2_1 _08736_ (.A(net1429),
    .B(_00158_),
    .Y(_03109_));
 sg13g2_a22oi_1 _08737_ (.Y(_03110_),
    .B1(_03109_),
    .B2(net1334),
    .A2(_03108_),
    .A1(_03107_));
 sg13g2_or2_1 _08738_ (.X(_03111_),
    .B(_03110_),
    .A(_03057_));
 sg13g2_a221oi_1 _08739_ (.B2(_03111_),
    .C1(net1123),
    .B1(_03106_),
    .A1(_00766_),
    .Y(_00549_),
    .A2(net1112));
 sg13g2_o21ai_1 _08740_ (.B1(_01166_),
    .Y(_03112_),
    .A1(_01122_),
    .A2(_02720_));
 sg13g2_a21oi_1 _08741_ (.A1(_01286_),
    .A2(_02720_),
    .Y(_03113_),
    .B1(_03112_));
 sg13g2_a21oi_1 _08742_ (.A1(_01090_),
    .A2(net1306),
    .Y(_03114_),
    .B1(_03113_));
 sg13g2_nand2_1 _08743_ (.Y(_03115_),
    .A(net2301),
    .B(_02716_));
 sg13g2_o21ai_1 _08744_ (.B1(_03115_),
    .Y(_00550_),
    .A1(_02718_),
    .A2(_03114_));
 sg13g2_o21ai_1 _08745_ (.B1(_01166_),
    .Y(_03116_),
    .A1(_01580_),
    .A2(_02719_));
 sg13g2_a21oi_1 _08746_ (.A1(_01065_),
    .A2(_02719_),
    .Y(_03117_),
    .B1(_03116_));
 sg13g2_a21oi_1 _08747_ (.A1(_01051_),
    .A2(net1306),
    .Y(_03118_),
    .B1(_03117_));
 sg13g2_nand2_1 _08748_ (.Y(_03119_),
    .A(net2250),
    .B(_02716_));
 sg13g2_o21ai_1 _08749_ (.B1(_03119_),
    .Y(_00551_),
    .A1(_02718_),
    .A2(_03118_));
 sg13g2_o21ai_1 _08750_ (.B1(_00160_),
    .Y(_03120_),
    .A1(net1436),
    .A2(\i_core.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_nor3_1 _08751_ (.A(net1432),
    .B(_02998_),
    .C(net2204),
    .Y(_03121_));
 sg13g2_nor2_1 _08752_ (.A(net2090),
    .B(net1260),
    .Y(_03122_));
 sg13g2_a21oi_1 _08753_ (.A1(_00853_),
    .A2(net1259),
    .Y(_00552_),
    .B1(net2091));
 sg13g2_nor2_1 _08754_ (.A(net2187),
    .B(net1259),
    .Y(_03123_));
 sg13g2_a21oi_1 _08755_ (.A1(_00854_),
    .A2(net1259),
    .Y(_00553_),
    .B1(_03123_));
 sg13g2_mux2_1 _08756_ (.A0(net1957),
    .A1(net11),
    .S(net1259),
    .X(_00554_));
 sg13g2_nor2_1 _08757_ (.A(net2137),
    .B(net1260),
    .Y(_03124_));
 sg13g2_a21oi_1 _08758_ (.A1(_00856_),
    .A2(net1259),
    .Y(_00555_),
    .B1(net2138));
 sg13g2_mux2_1 _08759_ (.A0(net2030),
    .A1(\i_core.mem.q_ctrl.spi_in_buffer[0] ),
    .S(net1260),
    .X(_00556_));
 sg13g2_mux2_1 _08760_ (.A0(net1999),
    .A1(\i_core.mem.q_ctrl.spi_in_buffer[1] ),
    .S(net1259),
    .X(_00557_));
 sg13g2_nand2_1 _08761_ (.Y(_03125_),
    .A(net1957),
    .B(net1259));
 sg13g2_o21ai_1 _08762_ (.B1(_03125_),
    .Y(_00558_),
    .A1(_00855_),
    .A2(net1259));
 sg13g2_mux2_1 _08763_ (.A0(net1995),
    .A1(\i_core.mem.q_ctrl.spi_in_buffer[3] ),
    .S(net1260),
    .X(_00559_));
 sg13g2_and2_1 _08764_ (.A(_02025_),
    .B(_02995_),
    .X(_03126_));
 sg13g2_nor3_2 _08765_ (.A(\i_core.mem.q_ctrl.read_cycles_count[0] ),
    .B(\i_core.mem.q_ctrl.read_cycles_count[2] ),
    .C(_03003_),
    .Y(_03127_));
 sg13g2_nor3_1 _08766_ (.A(net1433),
    .B(_03126_),
    .C(_03127_),
    .Y(_03128_));
 sg13g2_o21ai_1 _08767_ (.B1(net2685),
    .Y(_03129_),
    .A1(_02025_),
    .A2(_03000_));
 sg13g2_nor2_1 _08768_ (.A(_00159_),
    .B(_02997_),
    .Y(_03130_));
 sg13g2_a21oi_2 _08769_ (.B1(_03128_),
    .Y(_03131_),
    .A2(_03130_),
    .A1(_03129_));
 sg13g2_a21o_1 _08770_ (.A2(_03130_),
    .A1(_03129_),
    .B1(_03128_),
    .X(_03132_));
 sg13g2_nand2_1 _08771_ (.Y(_03133_),
    .A(net1437),
    .B(\i_core.mem.q_ctrl.data_req ));
 sg13g2_xor2_1 _08772_ (.B(\i_core.mem.q_ctrl.data_req ),
    .A(net1437),
    .X(_03134_));
 sg13g2_xnor2_1 _08773_ (.Y(_03135_),
    .A(net1437),
    .B(\i_core.mem.q_ctrl.data_req ));
 sg13g2_xor2_1 _08774_ (.B(_03133_),
    .A(\i_core.mem.qspi_data_byte_idx[1] ),
    .X(_03136_));
 sg13g2_mux4_1 _08775_ (.S0(net1329),
    .A0(\data_to_write[24] ),
    .A1(\data_to_write[16] ),
    .A2(\data_to_write[8] ),
    .A3(\data_to_write[0] ),
    .S1(net1281),
    .X(_03137_));
 sg13g2_o21ai_1 _08776_ (.B1(net1432),
    .Y(_03138_),
    .A1(_03082_),
    .A2(_03137_));
 sg13g2_a21oi_1 _08777_ (.A1(_00853_),
    .A2(_03082_),
    .Y(_03139_),
    .B1(_03138_));
 sg13g2_and2_2 _08778_ (.A(net1436),
    .B(_03127_),
    .X(_03140_));
 sg13g2_nand2_1 _08779_ (.Y(_03141_),
    .A(net1436),
    .B(_03127_));
 sg13g2_nand2_1 _08780_ (.Y(_03142_),
    .A(net2030),
    .B(_03140_));
 sg13g2_a21oi_1 _08781_ (.A1(\i_core.mem.q_ctrl.spi_in_buffer[0] ),
    .A2(_03141_),
    .Y(_03143_),
    .B1(net1258));
 sg13g2_a221oi_1 _08782_ (.B2(_03143_),
    .C1(net1432),
    .B1(_03142_),
    .A1(_00853_),
    .Y(_03144_),
    .A2(net1258));
 sg13g2_nor3_2 _08783_ (.A(net1219),
    .B(_03139_),
    .C(_03144_),
    .Y(_03145_));
 sg13g2_a21oi_1 _08784_ (.A1(_00826_),
    .A2(net1218),
    .Y(_00560_),
    .B1(_03145_));
 sg13g2_nand2_1 _08785_ (.Y(_03146_),
    .A(\i_core.mem.q_ctrl.spi_in_buffer[5] ),
    .B(_03140_));
 sg13g2_a21oi_1 _08786_ (.A1(\i_core.mem.q_ctrl.spi_in_buffer[1] ),
    .A2(_03141_),
    .Y(_03147_),
    .B1(net1258));
 sg13g2_a22oi_1 _08787_ (.Y(_03148_),
    .B1(_03146_),
    .B2(_03147_),
    .A2(net1258),
    .A1(_00854_));
 sg13g2_mux4_1 _08788_ (.S0(net1329),
    .A0(\data_to_write[25] ),
    .A1(\data_to_write[17] ),
    .A2(\data_to_write[9] ),
    .A3(\data_to_write[1] ),
    .S1(net1281),
    .X(_03149_));
 sg13g2_and2_1 _08789_ (.A(_03083_),
    .B(_03149_),
    .X(_03150_));
 sg13g2_a21oi_1 _08790_ (.A1(net10),
    .A2(_03082_),
    .Y(_03151_),
    .B1(_03150_));
 sg13g2_a21oi_1 _08791_ (.A1(net1433),
    .A2(_03151_),
    .Y(_03152_),
    .B1(net1219));
 sg13g2_o21ai_1 _08792_ (.B1(_03152_),
    .Y(_03153_),
    .A1(net1432),
    .A2(_03148_));
 sg13g2_o21ai_1 _08793_ (.B1(_03153_),
    .Y(_00561_),
    .A1(_00832_),
    .A2(_03131_));
 sg13g2_a21oi_1 _08794_ (.A1(_00855_),
    .A2(_03140_),
    .Y(_03154_),
    .B1(net1258));
 sg13g2_o21ai_1 _08795_ (.B1(_03154_),
    .Y(_03155_),
    .A1(net1957),
    .A2(_03140_));
 sg13g2_a21oi_1 _08796_ (.A1(net11),
    .A2(net1258),
    .Y(_03156_),
    .B1(net1432));
 sg13g2_nand2_1 _08797_ (.Y(_03157_),
    .A(\data_to_write[2] ),
    .B(net1329));
 sg13g2_nand2_1 _08798_ (.Y(_03158_),
    .A(\data_to_write[10] ),
    .B(net1330));
 sg13g2_nand3_1 _08799_ (.B(_03157_),
    .C(_03158_),
    .A(net1281),
    .Y(_03159_));
 sg13g2_nand2_1 _08800_ (.Y(_03160_),
    .A(\data_to_write[18] ),
    .B(net1329));
 sg13g2_a21oi_1 _08801_ (.A1(\data_to_write[26] ),
    .A2(net1330),
    .Y(_03161_),
    .B1(net1281));
 sg13g2_a21oi_1 _08802_ (.A1(_03160_),
    .A2(_03161_),
    .Y(_03162_),
    .B1(_03082_));
 sg13g2_a22oi_1 _08803_ (.Y(_03163_),
    .B1(_03159_),
    .B2(_03162_),
    .A2(_03082_),
    .A1(net11));
 sg13g2_a221oi_1 _08804_ (.B2(net1432),
    .C1(net1219),
    .B1(_03163_),
    .A1(_03155_),
    .Y(_03164_),
    .A2(_03156_));
 sg13g2_a21o_1 _08805_ (.A2(net1219),
    .A1(net2630),
    .B1(_03164_),
    .X(_00562_));
 sg13g2_nand2_1 _08806_ (.Y(_03165_),
    .A(net2370),
    .B(net1218));
 sg13g2_mux4_1 _08807_ (.S0(net1328),
    .A0(\data_to_write[27] ),
    .A1(\data_to_write[19] ),
    .A2(\data_to_write[11] ),
    .A3(\data_to_write[3] ),
    .S1(net1280),
    .X(_03166_));
 sg13g2_o21ai_1 _08808_ (.B1(net1432),
    .Y(_03167_),
    .A1(_00856_),
    .A2(_03083_));
 sg13g2_a21oi_1 _08809_ (.A1(_03083_),
    .A2(_03166_),
    .Y(_03168_),
    .B1(_03167_));
 sg13g2_nand2_1 _08810_ (.Y(_03169_),
    .A(net1995),
    .B(_03140_));
 sg13g2_a21oi_1 _08811_ (.A1(\i_core.mem.q_ctrl.spi_in_buffer[3] ),
    .A2(_03141_),
    .Y(_03170_),
    .B1(net1258));
 sg13g2_a22oi_1 _08812_ (.Y(_03171_),
    .B1(_03169_),
    .B2(_03170_),
    .A2(net1258),
    .A1(_00856_));
 sg13g2_o21ai_1 _08813_ (.B1(_03131_),
    .Y(_03172_),
    .A1(net1432),
    .A2(_03171_));
 sg13g2_o21ai_1 _08814_ (.B1(_03165_),
    .Y(_00563_),
    .A1(_03168_),
    .A2(_03172_));
 sg13g2_nand2_2 _08815_ (.Y(_03173_),
    .A(net1433),
    .B(_03083_));
 sg13g2_nand2_1 _08816_ (.Y(_03174_),
    .A(net2133),
    .B(net1330));
 sg13g2_nand2_1 _08817_ (.Y(_03175_),
    .A(\data_to_write[4] ),
    .B(net1328));
 sg13g2_nand3_1 _08818_ (.B(_03174_),
    .C(_03175_),
    .A(net1280),
    .Y(_03176_));
 sg13g2_nand2_1 _08819_ (.Y(_03177_),
    .A(net2191),
    .B(net1328));
 sg13g2_a21oi_1 _08820_ (.A1(net1903),
    .A2(net1330),
    .Y(_03178_),
    .B1(net1280));
 sg13g2_a21oi_1 _08821_ (.A1(_03177_),
    .A2(_03178_),
    .Y(_03179_),
    .B1(_03173_));
 sg13g2_a221oi_1 _08822_ (.B2(_03179_),
    .C1(net1218),
    .B1(_03176_),
    .A1(\i_core.cpu.instr_data_in[8] ),
    .Y(_03180_),
    .A2(_03173_));
 sg13g2_a21oi_1 _08823_ (.A1(_00827_),
    .A2(net1218),
    .Y(_00564_),
    .B1(_03180_));
 sg13g2_mux2_1 _08824_ (.A0(net1880),
    .A1(net2184),
    .S(net1328),
    .X(_03181_));
 sg13g2_and2_1 _08825_ (.A(\data_to_write[13] ),
    .B(net1330),
    .X(_03182_));
 sg13g2_a21oi_1 _08826_ (.A1(\data_to_write[5] ),
    .A2(net1328),
    .Y(_03183_),
    .B1(_03182_));
 sg13g2_a21oi_1 _08827_ (.A1(net1280),
    .A2(_03183_),
    .Y(_03184_),
    .B1(_03173_));
 sg13g2_o21ai_1 _08828_ (.B1(_03184_),
    .Y(_03185_),
    .A1(net1280),
    .A2(_03181_));
 sg13g2_a21oi_1 _08829_ (.A1(net2374),
    .A2(_03173_),
    .Y(_03186_),
    .B1(net1218));
 sg13g2_a22oi_1 _08830_ (.Y(_00565_),
    .B1(_03185_),
    .B2(_03186_),
    .A2(net1218),
    .A1(_00833_));
 sg13g2_nand2_1 _08831_ (.Y(_03187_),
    .A(net2183),
    .B(net1330));
 sg13g2_nand2_1 _08832_ (.Y(_03188_),
    .A(\data_to_write[6] ),
    .B(net1328));
 sg13g2_nand3_1 _08833_ (.B(_03187_),
    .C(_03188_),
    .A(net1280),
    .Y(_03189_));
 sg13g2_nand2_1 _08834_ (.Y(_03190_),
    .A(net2181),
    .B(net1328));
 sg13g2_a21oi_1 _08835_ (.A1(net1890),
    .A2(net1330),
    .Y(_03191_),
    .B1(net1280));
 sg13g2_a21oi_1 _08836_ (.A1(_03190_),
    .A2(_03191_),
    .Y(_03192_),
    .B1(_03173_));
 sg13g2_a221oi_1 _08837_ (.B2(_03192_),
    .C1(net1218),
    .B1(_03189_),
    .A1(net2630),
    .Y(_03193_),
    .A2(_03173_));
 sg13g2_a21oi_1 _08838_ (.A1(_00835_),
    .A2(net1218),
    .Y(_00566_),
    .B1(_03193_));
 sg13g2_nand2_1 _08839_ (.Y(_03194_),
    .A(net2188),
    .B(net1330));
 sg13g2_nand2_1 _08840_ (.Y(_03195_),
    .A(\data_to_write[7] ),
    .B(net1329));
 sg13g2_nand3_1 _08841_ (.B(_03194_),
    .C(_03195_),
    .A(net1280),
    .Y(_03196_));
 sg13g2_nand2_1 _08842_ (.Y(_03197_),
    .A(net2175),
    .B(net1328));
 sg13g2_a21oi_1 _08843_ (.A1(net1909),
    .A2(_03134_),
    .Y(_03198_),
    .B1(net1281));
 sg13g2_a21oi_1 _08844_ (.A1(_03197_),
    .A2(_03198_),
    .Y(_03199_),
    .B1(_03173_));
 sg13g2_a221oi_1 _08845_ (.B2(_03199_),
    .C1(net1219),
    .B1(_03196_),
    .A1(net2370),
    .Y(_03200_),
    .A2(_03173_));
 sg13g2_a21oi_1 _08846_ (.A1(_00838_),
    .A2(net1219),
    .Y(_00567_),
    .B1(_03200_));
 sg13g2_nand2b_1 _08847_ (.Y(_00568_),
    .B(net1322),
    .A_N(net1906));
 sg13g2_nand2b_1 _08848_ (.Y(_00569_),
    .B(net1320),
    .A_N(net1937));
 sg13g2_nor3_1 _08849_ (.A(net2498),
    .B(net1457),
    .C(_02747_),
    .Y(_03201_));
 sg13g2_a21oi_1 _08850_ (.A1(_00825_),
    .A2(_02747_),
    .Y(_00571_),
    .B1(_03201_));
 sg13g2_nor3_1 _08851_ (.A(net2307),
    .B(net1457),
    .C(_02747_),
    .Y(_03202_));
 sg13g2_a21oi_1 _08852_ (.A1(_00831_),
    .A2(_02747_),
    .Y(_00572_),
    .B1(_03202_));
 sg13g2_nand2_1 _08853_ (.Y(_03203_),
    .A(net1320),
    .B(net2093));
 sg13g2_o21ai_1 _08854_ (.B1(_03203_),
    .Y(_00573_),
    .A1(net1320),
    .A2(_00853_));
 sg13g2_nor2_1 _08855_ (.A(net1320),
    .B(net10),
    .Y(_03204_));
 sg13g2_a21oi_1 _08856_ (.A1(net1320),
    .A2(_00851_),
    .Y(_00574_),
    .B1(_03204_));
 sg13g2_mux2_1 _08857_ (.A0(net11),
    .A1(net2551),
    .S(net1320),
    .X(_00575_));
 sg13g2_nand2_1 _08858_ (.Y(_03205_),
    .A(\i_core.cpu.pc[1] ),
    .B(\i_core.cpu.i_core.imm_lo[1] ));
 sg13g2_xnor2_1 _08859_ (.Y(_03206_),
    .A(\i_core.cpu.pc[1] ),
    .B(\i_core.cpu.i_core.imm_lo[1] ));
 sg13g2_or2_1 _08860_ (.X(_03207_),
    .B(_03206_),
    .A(net1344));
 sg13g2_o21ai_1 _08861_ (.B1(_03207_),
    .Y(_03208_),
    .A1(net1348),
    .A2(_02791_));
 sg13g2_a22oi_1 _08862_ (.Y(_03209_),
    .B1(_03208_),
    .B2(net1180),
    .A2(net1172),
    .A1(net1825));
 sg13g2_nand2_1 _08863_ (.Y(_03210_),
    .A(_01846_),
    .B(net1170));
 sg13g2_a21oi_1 _08864_ (.A1(_03209_),
    .A2(_03210_),
    .Y(_00576_),
    .B1(net1385));
 sg13g2_nand2_1 _08865_ (.Y(_03211_),
    .A(\i_core.cpu.pc[2] ),
    .B(\i_core.cpu.i_core.imm_lo[2] ));
 sg13g2_xnor2_1 _08866_ (.Y(_03212_),
    .A(\i_core.cpu.pc[2] ),
    .B(\i_core.cpu.i_core.imm_lo[2] ));
 sg13g2_xnor2_1 _08867_ (.Y(_03213_),
    .A(_03205_),
    .B(_03212_));
 sg13g2_nand2_1 _08868_ (.Y(_03214_),
    .A(net1346),
    .B(_03213_));
 sg13g2_a21oi_1 _08869_ (.A1(net1344),
    .A2(_02794_),
    .Y(_03215_),
    .B1(net1176));
 sg13g2_a22oi_1 _08870_ (.Y(_03216_),
    .B1(_03214_),
    .B2(_03215_),
    .A2(net1172),
    .A1(net1826));
 sg13g2_o21ai_1 _08871_ (.B1(_03216_),
    .Y(_03217_),
    .A1(_01845_),
    .A2(_02579_));
 sg13g2_and2_1 _08872_ (.A(net1464),
    .B(_03217_),
    .X(_00577_));
 sg13g2_nor2_1 _08873_ (.A(_02935_),
    .B(_02943_),
    .Y(_03218_));
 sg13g2_nand2_2 _08874_ (.Y(_03219_),
    .A(_02934_),
    .B(net1125));
 sg13g2_nor2_1 _08875_ (.A(net1125),
    .B(net1263),
    .Y(_03220_));
 sg13g2_nor2_2 _08876_ (.A(_02934_),
    .B(_02943_),
    .Y(_03221_));
 sg13g2_nand2_2 _08877_ (.Y(_03222_),
    .A(_02935_),
    .B(_02944_));
 sg13g2_nor2_1 _08878_ (.A(net1422),
    .B(\i_core.cpu.instr_write_offset[1] ),
    .Y(_03223_));
 sg13g2_a21oi_2 _08879_ (.B1(_03223_),
    .Y(_03224_),
    .A2(_03206_),
    .A1(net1422));
 sg13g2_a22oi_1 _08880_ (.Y(_03225_),
    .B1(net1113),
    .B2(_03224_),
    .A2(net1117),
    .A1(net2143));
 sg13g2_o21ai_1 _08881_ (.B1(_03225_),
    .Y(_00578_),
    .A1(_00816_),
    .A2(_03219_));
 sg13g2_nor2_1 _08882_ (.A(net1389),
    .B(_03213_),
    .Y(_03226_));
 sg13g2_a21oi_1 _08883_ (.A1(net1389),
    .A2(\i_core.cpu.instr_write_offset[2] ),
    .Y(_03227_),
    .B1(_03226_));
 sg13g2_a22oi_1 _08884_ (.Y(_03228_),
    .B1(net1118),
    .B2(net2088),
    .A2(net1120),
    .A1(net1452));
 sg13g2_o21ai_1 _08885_ (.B1(net2089),
    .Y(_00579_),
    .A1(_03222_),
    .A2(_03227_));
 sg13g2_or2_1 _08886_ (.X(_03229_),
    .B(\i_core.cpu.i_core.imm_lo[3] ),
    .A(net1428));
 sg13g2_and2_1 _08887_ (.A(net1428),
    .B(\i_core.cpu.i_core.imm_lo[3] ),
    .X(_03230_));
 sg13g2_xnor2_1 _08888_ (.Y(_03231_),
    .A(net1428),
    .B(\i_core.cpu.i_core.imm_lo[3] ));
 sg13g2_o21ai_1 _08889_ (.B1(_03211_),
    .Y(_03232_),
    .A1(_03205_),
    .A2(_03212_));
 sg13g2_xnor2_1 _08890_ (.Y(_03233_),
    .A(_03231_),
    .B(_03232_));
 sg13g2_nand2_2 _08891_ (.Y(_03234_),
    .A(net1428),
    .B(\i_core.cpu.instr_write_offset[3] ));
 sg13g2_nor2_1 _08892_ (.A(net1428),
    .B(\i_core.cpu.instr_write_offset[3] ),
    .Y(_03235_));
 sg13g2_nor2_1 _08893_ (.A(net1422),
    .B(_03235_),
    .Y(_03236_));
 sg13g2_a22oi_1 _08894_ (.Y(_03237_),
    .B1(_03234_),
    .B2(_03236_),
    .A2(_03233_),
    .A1(net1422));
 sg13g2_a22oi_1 _08895_ (.Y(_03238_),
    .B1(net1118),
    .B2(net2033),
    .A2(net1121),
    .A1(net2098));
 sg13g2_o21ai_1 _08896_ (.B1(_03238_),
    .Y(_00580_),
    .A1(_03222_),
    .A2(_03237_));
 sg13g2_o21ai_1 _08897_ (.B1(net1170),
    .Y(_03239_),
    .A1(_01526_),
    .A2(net1189));
 sg13g2_and2_1 _08898_ (.A(net1188),
    .B(net1167),
    .X(_03240_));
 sg13g2_nand2_1 _08899_ (.Y(_03241_),
    .A(net1188),
    .B(net1167));
 sg13g2_o21ai_1 _08900_ (.B1(net1464),
    .Y(_03242_),
    .A1(net2638),
    .A2(net1160));
 sg13g2_a21oi_1 _08901_ (.A1(_03209_),
    .A2(_03239_),
    .Y(_00581_),
    .B1(_03242_));
 sg13g2_o21ai_1 _08902_ (.B1(net1168),
    .Y(_03243_),
    .A1(_01675_),
    .A2(net1189));
 sg13g2_o21ai_1 _08903_ (.B1(net1464),
    .Y(_03244_),
    .A1(net2644),
    .A2(net1160));
 sg13g2_a21oi_1 _08904_ (.A1(_03216_),
    .A2(_03243_),
    .Y(_00582_),
    .B1(_03244_));
 sg13g2_nor2_1 _08905_ (.A(net1344),
    .B(_03233_),
    .Y(_03245_));
 sg13g2_a21oi_1 _08906_ (.A1(net1344),
    .A2(_02797_),
    .Y(_03246_),
    .B1(_03245_));
 sg13g2_a22oi_1 _08907_ (.Y(_03247_),
    .B1(_03246_),
    .B2(net1180),
    .A2(net1172),
    .A1(net1827));
 sg13g2_o21ai_1 _08908_ (.B1(net1168),
    .Y(_03248_),
    .A1(net1189),
    .A2(_01979_));
 sg13g2_o21ai_1 _08909_ (.B1(net1465),
    .Y(_03249_),
    .A1(net1428),
    .A2(net1160));
 sg13g2_a21oi_1 _08910_ (.A1(_03247_),
    .A2(_03248_),
    .Y(_00583_),
    .B1(_03249_));
 sg13g2_nand2_1 _08911_ (.Y(_03250_),
    .A(\i_core.cpu.instr_data_start[4] ),
    .B(\i_core.cpu.i_core.imm_lo[4] ));
 sg13g2_xnor2_1 _08912_ (.Y(_03251_),
    .A(\i_core.cpu.instr_data_start[4] ),
    .B(\i_core.cpu.i_core.imm_lo[4] ));
 sg13g2_a21oi_2 _08913_ (.B1(_03230_),
    .Y(_03252_),
    .A2(_03232_),
    .A1(_03229_));
 sg13g2_xnor2_1 _08914_ (.Y(_03253_),
    .A(_03251_),
    .B(_03252_));
 sg13g2_mux2_1 _08915_ (.A0(_02800_),
    .A1(_03253_),
    .S(net1348),
    .X(_03254_));
 sg13g2_a22oi_1 _08916_ (.Y(_03255_),
    .B1(_03254_),
    .B2(net1180),
    .A2(net1172),
    .A1(_00857_));
 sg13g2_o21ai_1 _08917_ (.B1(_03255_),
    .Y(_03256_),
    .A1(_01217_),
    .A2(_02579_));
 sg13g2_o21ai_1 _08918_ (.B1(net1465),
    .Y(_03257_),
    .A1(net2578),
    .A2(net1160));
 sg13g2_a21oi_1 _08919_ (.A1(net1160),
    .A2(_03256_),
    .Y(_00584_),
    .B1(_03257_));
 sg13g2_or2_1 _08920_ (.X(_03258_),
    .B(\i_core.cpu.i_core.imm_lo[5] ),
    .A(\i_core.cpu.instr_data_start[5] ));
 sg13g2_and2_1 _08921_ (.A(\i_core.cpu.instr_data_start[5] ),
    .B(\i_core.cpu.i_core.imm_lo[5] ),
    .X(_03259_));
 sg13g2_xnor2_1 _08922_ (.Y(_03260_),
    .A(\i_core.cpu.instr_data_start[5] ),
    .B(\i_core.cpu.i_core.imm_lo[5] ));
 sg13g2_o21ai_1 _08923_ (.B1(_03250_),
    .Y(_03261_),
    .A1(_03251_),
    .A2(_03252_));
 sg13g2_xnor2_1 _08924_ (.Y(_03262_),
    .A(_03260_),
    .B(_03261_));
 sg13g2_nor2_1 _08925_ (.A(net1344),
    .B(_03262_),
    .Y(_03263_));
 sg13g2_a21oi_1 _08926_ (.A1(net1345),
    .A2(_02803_),
    .Y(_03264_),
    .B1(_03263_));
 sg13g2_a22oi_1 _08927_ (.Y(_03265_),
    .B1(_03264_),
    .B2(net1181),
    .A2(net1172),
    .A1(net1810));
 sg13g2_o21ai_1 _08928_ (.B1(net1168),
    .Y(_03266_),
    .A1(_01524_),
    .A2(_01773_));
 sg13g2_a221oi_1 _08929_ (.B2(_03266_),
    .C1(net1385),
    .B1(_03265_),
    .A1(_00765_),
    .Y(_00585_),
    .A2(net1163));
 sg13g2_nand2_1 _08930_ (.Y(_03267_),
    .A(\i_core.cpu.instr_data_start[6] ),
    .B(\i_core.cpu.i_core.imm_lo[6] ));
 sg13g2_xnor2_1 _08931_ (.Y(_03268_),
    .A(\i_core.cpu.instr_data_start[6] ),
    .B(\i_core.cpu.i_core.imm_lo[6] ));
 sg13g2_a21oi_1 _08932_ (.A1(_03258_),
    .A2(_03261_),
    .Y(_03269_),
    .B1(_03259_));
 sg13g2_xor2_1 _08933_ (.B(_03269_),
    .A(_03268_),
    .X(_03270_));
 sg13g2_o21ai_1 _08934_ (.B1(net1180),
    .Y(_03271_),
    .A1(net1347),
    .A2(_02807_));
 sg13g2_a21oi_1 _08935_ (.A1(net1348),
    .A2(_03270_),
    .Y(_03272_),
    .B1(_03271_));
 sg13g2_a221oi_1 _08936_ (.B2(_01673_),
    .C1(_03272_),
    .B1(net1168),
    .A1(_00858_),
    .Y(_03273_),
    .A2(net1172));
 sg13g2_o21ai_1 _08937_ (.B1(net1466),
    .Y(_03274_),
    .A1(net1163),
    .A2(_03273_));
 sg13g2_a21oi_1 _08938_ (.A1(_00764_),
    .A2(net1163),
    .Y(_00586_),
    .B1(_03274_));
 sg13g2_and2_1 _08939_ (.A(net1427),
    .B(\i_core.cpu.i_core.imm_lo[7] ),
    .X(_03275_));
 sg13g2_xor2_1 _08940_ (.B(\i_core.cpu.i_core.imm_lo[7] ),
    .A(net1427),
    .X(_03276_));
 sg13g2_o21ai_1 _08941_ (.B1(_03267_),
    .Y(_03277_),
    .A1(_03268_),
    .A2(_03269_));
 sg13g2_xnor2_1 _08942_ (.Y(_03278_),
    .A(_03276_),
    .B(_03277_));
 sg13g2_nand2_1 _08943_ (.Y(_03279_),
    .A(net1347),
    .B(_03278_));
 sg13g2_a21oi_1 _08944_ (.A1(net1345),
    .A2(_02810_),
    .Y(_03280_),
    .B1(net1177));
 sg13g2_a22oi_1 _08945_ (.Y(_03281_),
    .B1(_03279_),
    .B2(_03280_),
    .A2(net1169),
    .A1(_01977_));
 sg13g2_a21oi_1 _08946_ (.A1(net1812),
    .A2(net1174),
    .Y(_03282_),
    .B1(_03240_));
 sg13g2_o21ai_1 _08947_ (.B1(net1466),
    .Y(_03283_),
    .A1(net2435),
    .A2(net1162));
 sg13g2_a21oi_1 _08948_ (.A1(_03281_),
    .A2(_03282_),
    .Y(_00587_),
    .B1(_03283_));
 sg13g2_nor2_1 _08949_ (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .B(net1171),
    .Y(_03284_));
 sg13g2_a21oi_2 _08950_ (.B1(_03284_),
    .Y(_03285_),
    .A2(_01833_),
    .A1(_01216_));
 sg13g2_nand2_1 _08951_ (.Y(_03286_),
    .A(\i_core.cpu.instr_data_start[8] ),
    .B(\i_core.cpu.i_core.imm_lo[8] ));
 sg13g2_xnor2_1 _08952_ (.Y(_03287_),
    .A(\i_core.cpu.instr_data_start[8] ),
    .B(\i_core.cpu.i_core.imm_lo[8] ));
 sg13g2_a21oi_1 _08953_ (.A1(_03276_),
    .A2(_03277_),
    .Y(_03288_),
    .B1(_03275_));
 sg13g2_xnor2_1 _08954_ (.Y(_03289_),
    .A(_03287_),
    .B(_03288_));
 sg13g2_mux2_1 _08955_ (.A0(_02813_),
    .A1(_03289_),
    .S(net1347),
    .X(_03290_));
 sg13g2_nand2_1 _08956_ (.Y(_03291_),
    .A(net1181),
    .B(_03290_));
 sg13g2_o21ai_1 _08957_ (.B1(_03291_),
    .Y(_03292_),
    .A1(net1181),
    .A2(_03285_));
 sg13g2_o21ai_1 _08958_ (.B1(net1466),
    .Y(_03293_),
    .A1(net2651),
    .A2(net1162));
 sg13g2_a21oi_1 _08959_ (.A1(net1162),
    .A2(_03292_),
    .Y(_00588_),
    .B1(_03293_));
 sg13g2_o21ai_1 _08960_ (.B1(_03286_),
    .Y(_03294_),
    .A1(_03287_),
    .A2(_03288_));
 sg13g2_and2_1 _08961_ (.A(\i_core.cpu.instr_data_start[9] ),
    .B(\i_core.cpu.i_core.imm_lo[9] ),
    .X(_03295_));
 sg13g2_xor2_1 _08962_ (.B(\i_core.cpu.i_core.imm_lo[9] ),
    .A(\i_core.cpu.instr_data_start[9] ),
    .X(_03296_));
 sg13g2_xnor2_1 _08963_ (.Y(_03297_),
    .A(_03294_),
    .B(_03296_));
 sg13g2_nand2_1 _08964_ (.Y(_03298_),
    .A(net1347),
    .B(_03297_));
 sg13g2_a21oi_1 _08965_ (.A1(net1345),
    .A2(_02815_),
    .Y(_03299_),
    .B1(net1177));
 sg13g2_a22oi_1 _08966_ (.Y(_03300_),
    .B1(_03298_),
    .B2(_03299_),
    .A2(net1172),
    .A1(net1797));
 sg13g2_o21ai_1 _08967_ (.B1(net1168),
    .Y(_03301_),
    .A1(_01528_),
    .A2(net1189));
 sg13g2_a221oi_1 _08968_ (.B2(_03301_),
    .C1(net1385),
    .B1(_03300_),
    .A1(_00763_),
    .Y(_00589_),
    .A2(net1163));
 sg13g2_a21oi_1 _08969_ (.A1(_03294_),
    .A2(_03296_),
    .Y(_03302_),
    .B1(_03295_));
 sg13g2_nor2_1 _08970_ (.A(\i_core.cpu.instr_data_start[10] ),
    .B(\i_core.cpu.i_core.imm_lo[10] ),
    .Y(_03303_));
 sg13g2_xnor2_1 _08971_ (.Y(_03304_),
    .A(\i_core.cpu.instr_data_start[10] ),
    .B(\i_core.cpu.i_core.imm_lo[10] ));
 sg13g2_xnor2_1 _08972_ (.Y(_03305_),
    .A(_03302_),
    .B(_03304_));
 sg13g2_mux2_1 _08973_ (.A0(_02819_),
    .A1(_03305_),
    .S(net1347),
    .X(_03306_));
 sg13g2_nor2_1 _08974_ (.A(net1791),
    .B(net1171),
    .Y(_03307_));
 sg13g2_a221oi_1 _08975_ (.B2(net1180),
    .C1(_03307_),
    .B1(_03306_),
    .A1(_01671_),
    .Y(_03308_),
    .A2(net1169));
 sg13g2_o21ai_1 _08976_ (.B1(net1466),
    .Y(_03309_),
    .A1(net1163),
    .A2(_03308_));
 sg13g2_a21oi_1 _08977_ (.A1(_00762_),
    .A2(net1163),
    .Y(_00590_),
    .B1(_03309_));
 sg13g2_mux2_1 _08978_ (.A0(net1724),
    .A1(_01976_),
    .S(net1171),
    .X(_03310_));
 sg13g2_xnor2_1 _08979_ (.Y(_03311_),
    .A(\i_core.cpu.instr_data_start[11] ),
    .B(\i_core.cpu.i_core.imm_lo[11] ));
 sg13g2_a221oi_1 _08980_ (.B2(_03296_),
    .C1(_03295_),
    .B1(_03294_),
    .A1(\i_core.cpu.instr_data_start[10] ),
    .Y(_03312_),
    .A2(\i_core.cpu.i_core.imm_lo[10] ));
 sg13g2_nor3_1 _08981_ (.A(_03303_),
    .B(_03311_),
    .C(_03312_),
    .Y(_03313_));
 sg13g2_o21ai_1 _08982_ (.B1(_03311_),
    .Y(_03314_),
    .A1(_03303_),
    .A2(_03312_));
 sg13g2_nand2b_1 _08983_ (.Y(_03315_),
    .B(_03314_),
    .A_N(_03313_));
 sg13g2_nand2_1 _08984_ (.Y(_03316_),
    .A(net1347),
    .B(_03315_));
 sg13g2_a21oi_1 _08985_ (.A1(net1344),
    .A2(_02821_),
    .Y(_03317_),
    .B1(net1177));
 sg13g2_a22oi_1 _08986_ (.Y(_03318_),
    .B1(_03316_),
    .B2(_03317_),
    .A2(_03310_),
    .A1(net1177));
 sg13g2_o21ai_1 _08987_ (.B1(net1466),
    .Y(_03319_),
    .A1(net2648),
    .A2(net1160));
 sg13g2_a21oi_1 _08988_ (.A1(net1160),
    .A2(_03318_),
    .Y(_00591_),
    .B1(_03319_));
 sg13g2_a21oi_1 _08989_ (.A1(\i_core.cpu.instr_data_start[11] ),
    .A2(\i_core.cpu.i_core.imm_lo[11] ),
    .Y(_03320_),
    .B1(_03313_));
 sg13g2_nor2_1 _08990_ (.A(\i_core.cpu.instr_data_start[12] ),
    .B(\i_core.cpu.imm[12] ),
    .Y(_03321_));
 sg13g2_nand2_1 _08991_ (.Y(_03322_),
    .A(\i_core.cpu.instr_data_start[12] ),
    .B(\i_core.cpu.imm[12] ));
 sg13g2_nor2b_1 _08992_ (.A(_03321_),
    .B_N(_03322_),
    .Y(_03323_));
 sg13g2_xnor2_1 _08993_ (.Y(_03324_),
    .A(_03320_),
    .B(_03323_));
 sg13g2_o21ai_1 _08994_ (.B1(net1180),
    .Y(_03325_),
    .A1(net1347),
    .A2(_02825_));
 sg13g2_a21oi_1 _08995_ (.A1(net1347),
    .A2(_03324_),
    .Y(_03326_),
    .B1(_03325_));
 sg13g2_a221oi_1 _08996_ (.B2(_01213_),
    .C1(_03326_),
    .B1(net1168),
    .A1(_00859_),
    .Y(_03327_),
    .A2(net1174));
 sg13g2_o21ai_1 _08997_ (.B1(net1466),
    .Y(_03328_),
    .A1(net1163),
    .A2(_03327_));
 sg13g2_a21oi_1 _08998_ (.A1(_00761_),
    .A2(net1163),
    .Y(_00592_),
    .B1(_03328_));
 sg13g2_nand2b_1 _08999_ (.Y(_03329_),
    .B(net1168),
    .A_N(_01522_));
 sg13g2_and2_1 _09000_ (.A(\i_core.cpu.instr_data_start[13] ),
    .B(\i_core.cpu.imm[13] ),
    .X(_03330_));
 sg13g2_xor2_1 _09001_ (.B(\i_core.cpu.imm[13] ),
    .A(\i_core.cpu.instr_data_start[13] ),
    .X(_03331_));
 sg13g2_o21ai_1 _09002_ (.B1(_03322_),
    .Y(_03332_),
    .A1(_03320_),
    .A2(_03321_));
 sg13g2_xnor2_1 _09003_ (.Y(_03333_),
    .A(_03331_),
    .B(_03332_));
 sg13g2_nand2_1 _09004_ (.Y(_03334_),
    .A(net1346),
    .B(_03333_));
 sg13g2_a21oi_1 _09005_ (.A1(net1344),
    .A2(_02827_),
    .Y(_03335_),
    .B1(net1176));
 sg13g2_a221oi_1 _09006_ (.B2(_03335_),
    .C1(_03240_),
    .B1(_03334_),
    .A1(net1773),
    .Y(_03336_),
    .A2(net1174));
 sg13g2_a221oi_1 _09007_ (.B2(_03336_),
    .C1(net1385),
    .B1(_03329_),
    .A1(_00760_),
    .Y(_00593_),
    .A2(net1164));
 sg13g2_a21oi_1 _09008_ (.A1(_03331_),
    .A2(_03332_),
    .Y(_03337_),
    .B1(_03330_));
 sg13g2_nor2_1 _09009_ (.A(net1426),
    .B(\i_core.cpu.imm[14] ),
    .Y(_03338_));
 sg13g2_xor2_1 _09010_ (.B(\i_core.cpu.imm[14] ),
    .A(net1426),
    .X(_03339_));
 sg13g2_xnor2_1 _09011_ (.Y(_03340_),
    .A(_03337_),
    .B(_03339_));
 sg13g2_o21ai_1 _09012_ (.B1(net1180),
    .Y(_03341_),
    .A1(net1346),
    .A2(_02831_));
 sg13g2_a21o_1 _09013_ (.A2(_03340_),
    .A1(net1349),
    .B1(_03341_),
    .X(_03342_));
 sg13g2_o21ai_1 _09014_ (.B1(_03342_),
    .Y(_03343_),
    .A1(net1766),
    .A2(net1171));
 sg13g2_a21o_1 _09015_ (.A2(net1169),
    .A1(_01669_),
    .B1(_03343_),
    .X(_03344_));
 sg13g2_o21ai_1 _09016_ (.B1(net1463),
    .Y(_03345_),
    .A1(net2456),
    .A2(net1160));
 sg13g2_a21oi_1 _09017_ (.A1(net1161),
    .A2(_03344_),
    .Y(_00594_),
    .B1(_03345_));
 sg13g2_a21oi_1 _09018_ (.A1(net1794),
    .A2(net1173),
    .Y(_03346_),
    .B1(net1164));
 sg13g2_xnor2_1 _09019_ (.Y(_03347_),
    .A(net1425),
    .B(\i_core.cpu.imm[15] ));
 sg13g2_a221oi_1 _09020_ (.B2(_03332_),
    .C1(_03330_),
    .B1(_03331_),
    .A1(net1426),
    .Y(_03348_),
    .A2(\i_core.cpu.imm[14] ));
 sg13g2_nor3_1 _09021_ (.A(_03338_),
    .B(_03347_),
    .C(_03348_),
    .Y(_03349_));
 sg13g2_o21ai_1 _09022_ (.B1(_03347_),
    .Y(_03350_),
    .A1(_03338_),
    .A2(_03348_));
 sg13g2_nand2b_1 _09023_ (.Y(_03351_),
    .B(_03350_),
    .A_N(_03349_));
 sg13g2_nand2_1 _09024_ (.Y(_03352_),
    .A(net1344),
    .B(_02833_));
 sg13g2_a21oi_1 _09025_ (.A1(net1346),
    .A2(_03351_),
    .Y(_03353_),
    .B1(net1176));
 sg13g2_a22oi_1 _09026_ (.Y(_03354_),
    .B1(_03352_),
    .B2(_03353_),
    .A2(net1168),
    .A1(_01974_));
 sg13g2_o21ai_1 _09027_ (.B1(net1463),
    .Y(_03355_),
    .A1(net1425),
    .A2(net1161));
 sg13g2_a21oi_1 _09028_ (.A1(_03346_),
    .A2(_03354_),
    .Y(_00595_),
    .B1(_03355_));
 sg13g2_a21o_1 _09029_ (.A2(\i_core.cpu.imm[15] ),
    .A1(net1425),
    .B1(_03349_),
    .X(_03356_));
 sg13g2_or2_1 _09030_ (.X(_03357_),
    .B(\i_core.cpu.imm[16] ),
    .A(net1424));
 sg13g2_and2_1 _09031_ (.A(net1424),
    .B(\i_core.cpu.imm[16] ),
    .X(_03358_));
 sg13g2_xnor2_1 _09032_ (.Y(_03359_),
    .A(net1424),
    .B(\i_core.cpu.imm[16] ));
 sg13g2_xnor2_1 _09033_ (.Y(_03360_),
    .A(_03356_),
    .B(_03359_));
 sg13g2_o21ai_1 _09034_ (.B1(net1179),
    .Y(_03361_),
    .A1(net1346),
    .A2(_02837_));
 sg13g2_a21oi_1 _09035_ (.A1(net1349),
    .A2(_03360_),
    .Y(_03362_),
    .B1(_03361_));
 sg13g2_a221oi_1 _09036_ (.B2(_01228_),
    .C1(_03362_),
    .B1(net1167),
    .A1(_00860_),
    .Y(_03363_),
    .A2(net1172));
 sg13g2_o21ai_1 _09037_ (.B1(net1463),
    .Y(_03364_),
    .A1(net1164),
    .A2(_03363_));
 sg13g2_a21oi_1 _09038_ (.A1(_00759_),
    .A2(net1164),
    .Y(_00596_),
    .B1(_03364_));
 sg13g2_nor2_1 _09039_ (.A(\i_core.cpu.instr_data_start[17] ),
    .B(\i_core.cpu.imm[17] ),
    .Y(_03365_));
 sg13g2_nand2_1 _09040_ (.Y(_03366_),
    .A(\i_core.cpu.instr_data_start[17] ),
    .B(\i_core.cpu.imm[17] ));
 sg13g2_nor2b_1 _09041_ (.A(_03365_),
    .B_N(_03366_),
    .Y(_03367_));
 sg13g2_a21oi_1 _09042_ (.A1(_03356_),
    .A2(_03357_),
    .Y(_03368_),
    .B1(_03358_));
 sg13g2_xnor2_1 _09043_ (.Y(_03369_),
    .A(_03367_),
    .B(_03368_));
 sg13g2_o21ai_1 _09044_ (.B1(net1179),
    .Y(_03370_),
    .A1(net1345),
    .A2(_03369_));
 sg13g2_a21oi_1 _09045_ (.A1(net1343),
    .A2(_02839_),
    .Y(_03371_),
    .B1(_03370_));
 sg13g2_or2_1 _09046_ (.X(_03372_),
    .B(_01773_),
    .A(_01519_));
 sg13g2_a221oi_1 _09047_ (.B2(_03372_),
    .C1(_03371_),
    .B1(net1169),
    .A1(net1787),
    .Y(_03373_),
    .A2(net1173));
 sg13g2_o21ai_1 _09048_ (.B1(net1463),
    .Y(_03374_),
    .A1(net2522),
    .A2(net1161));
 sg13g2_nor2_1 _09049_ (.A(_03373_),
    .B(_03374_),
    .Y(_00597_));
 sg13g2_o21ai_1 _09050_ (.B1(_03366_),
    .Y(_03375_),
    .A1(_03365_),
    .A2(_03368_));
 sg13g2_xor2_1 _09051_ (.B(\i_core.cpu.imm[18] ),
    .A(\i_core.cpu.instr_data_start[18] ),
    .X(_03376_));
 sg13g2_xnor2_1 _09052_ (.Y(_03377_),
    .A(_03375_),
    .B(_03376_));
 sg13g2_mux2_1 _09053_ (.A0(_02843_),
    .A1(_03377_),
    .S(net1346),
    .X(_03378_));
 sg13g2_nor2_1 _09054_ (.A(net1749),
    .B(net1171),
    .Y(_03379_));
 sg13g2_a221oi_1 _09055_ (.B2(net1181),
    .C1(_03379_),
    .B1(_03378_),
    .A1(_01681_),
    .Y(_03380_),
    .A2(net1167));
 sg13g2_o21ai_1 _09056_ (.B1(net1463),
    .Y(_03381_),
    .A1(net1164),
    .A2(_03380_));
 sg13g2_a21oi_1 _09057_ (.A1(_00758_),
    .A2(net1164),
    .Y(_00598_),
    .B1(_03381_));
 sg13g2_nand2_1 _09058_ (.Y(_03382_),
    .A(\i_core.cpu.instr_data_start[19] ),
    .B(\i_core.cpu.imm[19] ));
 sg13g2_xnor2_1 _09059_ (.Y(_03383_),
    .A(\i_core.cpu.instr_data_start[19] ),
    .B(\i_core.cpu.imm[19] ));
 sg13g2_a21o_1 _09060_ (.A2(\i_core.cpu.imm[18] ),
    .A1(\i_core.cpu.instr_data_start[18] ),
    .B1(_03375_),
    .X(_03384_));
 sg13g2_o21ai_1 _09061_ (.B1(_03384_),
    .Y(_03385_),
    .A1(\i_core.cpu.instr_data_start[18] ),
    .A2(\i_core.cpu.imm[18] ));
 sg13g2_xnor2_1 _09062_ (.Y(_03386_),
    .A(_03383_),
    .B(_03385_));
 sg13g2_mux2_1 _09063_ (.A0(_02846_),
    .A1(_03386_),
    .S(net1346),
    .X(_03387_));
 sg13g2_o21ai_1 _09064_ (.B1(net1161),
    .Y(_03388_),
    .A1(net1750),
    .A2(net1171));
 sg13g2_a221oi_1 _09065_ (.B2(net1179),
    .C1(_03388_),
    .B1(_03387_),
    .A1(_01969_),
    .Y(_03389_),
    .A2(net1167));
 sg13g2_a21oi_1 _09066_ (.A1(net2599),
    .A2(net1164),
    .Y(_03390_),
    .B1(_03389_));
 sg13g2_nor2_1 _09067_ (.A(net1385),
    .B(_03390_),
    .Y(_00599_));
 sg13g2_o21ai_1 _09068_ (.B1(_03382_),
    .Y(_03391_),
    .A1(_03383_),
    .A2(_03385_));
 sg13g2_or2_1 _09069_ (.X(_03392_),
    .B(\i_core.cpu.imm[20] ),
    .A(net1423));
 sg13g2_and2_1 _09070_ (.A(net1423),
    .B(\i_core.cpu.imm[20] ),
    .X(_03393_));
 sg13g2_xor2_1 _09071_ (.B(\i_core.cpu.imm[20] ),
    .A(net1423),
    .X(_03394_));
 sg13g2_xnor2_1 _09072_ (.Y(_03395_),
    .A(_03391_),
    .B(_03394_));
 sg13g2_a21o_1 _09073_ (.A2(_03395_),
    .A1(net1346),
    .B1(net1178),
    .X(_03396_));
 sg13g2_a21oi_1 _09074_ (.A1(net1343),
    .A2(_02848_),
    .Y(_03397_),
    .B1(_03396_));
 sg13g2_nand2b_1 _09075_ (.Y(_03398_),
    .B(_01225_),
    .A_N(net1188));
 sg13g2_a221oi_1 _09076_ (.B2(_03398_),
    .C1(_03397_),
    .B1(net1167),
    .A1(net1887),
    .Y(_03399_),
    .A2(net1173));
 sg13g2_o21ai_1 _09077_ (.B1(net1462),
    .Y(_03400_),
    .A1(net1423),
    .A2(net1161));
 sg13g2_nor2_1 _09078_ (.A(_03399_),
    .B(_03400_),
    .Y(_00600_));
 sg13g2_nor2_1 _09079_ (.A(\i_core.cpu.instr_data_start[21] ),
    .B(\i_core.cpu.imm[21] ),
    .Y(_03401_));
 sg13g2_nand2_1 _09080_ (.Y(_03402_),
    .A(\i_core.cpu.instr_data_start[21] ),
    .B(\i_core.cpu.imm[21] ));
 sg13g2_nor2b_1 _09081_ (.A(_03401_),
    .B_N(_03402_),
    .Y(_03403_));
 sg13g2_a21oi_1 _09082_ (.A1(_03391_),
    .A2(_03392_),
    .Y(_03404_),
    .B1(_03393_));
 sg13g2_xnor2_1 _09083_ (.Y(_03405_),
    .A(_03403_),
    .B(_03404_));
 sg13g2_o21ai_1 _09084_ (.B1(net1179),
    .Y(_03406_),
    .A1(net1343),
    .A2(_03405_));
 sg13g2_a21oi_1 _09085_ (.A1(net1343),
    .A2(_02851_),
    .Y(_03407_),
    .B1(_03406_));
 sg13g2_nand2b_1 _09086_ (.Y(_03408_),
    .B(_01517_),
    .A_N(net1188));
 sg13g2_a221oi_1 _09087_ (.B2(_03408_),
    .C1(_03407_),
    .B1(net1169),
    .A1(net2016),
    .Y(_03409_),
    .A2(net1173));
 sg13g2_o21ai_1 _09088_ (.B1(net1462),
    .Y(_03410_),
    .A1(net2657),
    .A2(net1161));
 sg13g2_nor2_1 _09089_ (.A(_03409_),
    .B(_03410_),
    .Y(_00601_));
 sg13g2_o21ai_1 _09090_ (.B1(_03402_),
    .Y(_03411_),
    .A1(_03401_),
    .A2(_03404_));
 sg13g2_or2_1 _09091_ (.X(_03412_),
    .B(\i_core.cpu.imm[22] ),
    .A(\i_core.cpu.instr_data_start[22] ));
 sg13g2_and2_1 _09092_ (.A(\i_core.cpu.instr_data_start[22] ),
    .B(\i_core.cpu.imm[22] ),
    .X(_03413_));
 sg13g2_xor2_1 _09093_ (.B(\i_core.cpu.imm[22] ),
    .A(\i_core.cpu.instr_data_start[22] ),
    .X(_03414_));
 sg13g2_xnor2_1 _09094_ (.Y(_03415_),
    .A(_03411_),
    .B(_03414_));
 sg13g2_inv_1 _09095_ (.Y(_03416_),
    .A(_03415_));
 sg13g2_o21ai_1 _09096_ (.B1(net1179),
    .Y(_03417_),
    .A1(net1343),
    .A2(_03416_));
 sg13g2_a21oi_1 _09097_ (.A1(net1343),
    .A2(_02854_),
    .Y(_03418_),
    .B1(_03417_));
 sg13g2_nand2b_1 _09098_ (.Y(_03419_),
    .B(_01680_),
    .A_N(net1189));
 sg13g2_a221oi_1 _09099_ (.B2(_03419_),
    .C1(_03418_),
    .B1(net1167),
    .A1(net2092),
    .Y(_03420_),
    .A2(net1173));
 sg13g2_o21ai_1 _09100_ (.B1(net1462),
    .Y(_03421_),
    .A1(net2650),
    .A2(net1161));
 sg13g2_nor2_1 _09101_ (.A(_03420_),
    .B(_03421_),
    .Y(_00602_));
 sg13g2_a21oi_1 _09102_ (.A1(_03411_),
    .A2(_03412_),
    .Y(_03422_),
    .B1(_03413_));
 sg13g2_xor2_1 _09103_ (.B(\i_core.cpu.imm[23] ),
    .A(\i_core.cpu.instr_data_start[23] ),
    .X(_03423_));
 sg13g2_xnor2_1 _09104_ (.Y(_03424_),
    .A(_03422_),
    .B(_03423_));
 sg13g2_o21ai_1 _09105_ (.B1(net1179),
    .Y(_03425_),
    .A1(net1343),
    .A2(_03424_));
 sg13g2_a21oi_1 _09106_ (.A1(net1343),
    .A2(_02857_),
    .Y(_03426_),
    .B1(_03425_));
 sg13g2_or2_1 _09107_ (.X(_03427_),
    .B(_01966_),
    .A(net1188));
 sg13g2_a221oi_1 _09108_ (.B2(_03427_),
    .C1(_03426_),
    .B1(net1167),
    .A1(net1898),
    .Y(_03428_),
    .A2(net1173));
 sg13g2_o21ai_1 _09109_ (.B1(net1462),
    .Y(_03429_),
    .A1(net2515),
    .A2(net1161));
 sg13g2_nor2_1 _09110_ (.A(_03428_),
    .B(_03429_),
    .Y(_00603_));
 sg13g2_a21o_1 _09111_ (.A2(_00819_),
    .A1(net2640),
    .B1(\i_core.cpu.instr_fetch_started ),
    .X(_03430_));
 sg13g2_nand3_1 _09112_ (.B(net1171),
    .C(net2641),
    .A(_01799_),
    .Y(_03431_));
 sg13g2_o21ai_1 _09113_ (.B1(net1462),
    .Y(_03432_),
    .A1(net1417),
    .A2(net1178));
 sg13g2_a21oi_1 _09114_ (.A1(net1178),
    .A2(_03431_),
    .Y(_00604_),
    .B1(_03432_));
 sg13g2_o21ai_1 _09115_ (.B1(net1464),
    .Y(_03433_),
    .A1(net1419),
    .A2(net1310));
 sg13g2_a21oi_1 _09116_ (.A1(net1310),
    .A2(_01799_),
    .Y(_00605_),
    .B1(_03433_));
 sg13g2_nor2_1 _09117_ (.A(\i_core.cpu.i_core.mem_op[0] ),
    .B(_02072_),
    .Y(_03434_));
 sg13g2_nand3_1 _09118_ (.B(_01430_),
    .C(_02072_),
    .A(_01185_),
    .Y(_03435_));
 sg13g2_nor2_1 _09119_ (.A(net2532),
    .B(_03435_),
    .Y(_03436_));
 sg13g2_o21ai_1 _09120_ (.B1(net1462),
    .Y(_00606_),
    .A1(_03434_),
    .A2(_03436_));
 sg13g2_nor2_1 _09121_ (.A(\i_core.cpu.i_core.mem_op[1] ),
    .B(_02072_),
    .Y(_03437_));
 sg13g2_nor2_1 _09122_ (.A(net2489),
    .B(_03435_),
    .Y(_03438_));
 sg13g2_o21ai_1 _09123_ (.B1(net1462),
    .Y(_00607_),
    .A1(_03437_),
    .A2(_03438_));
 sg13g2_a21oi_1 _09124_ (.A1(net1920),
    .A2(_01882_),
    .Y(_03439_),
    .B1(_02070_));
 sg13g2_nand2_1 _09125_ (.Y(_03440_),
    .A(\i_core.cpu.i_core.mem_op[0] ),
    .B(_02068_));
 sg13g2_nand2_1 _09126_ (.Y(_03441_),
    .A(net2491),
    .B(net1247));
 sg13g2_nand3_1 _09127_ (.B(_03440_),
    .C(_03441_),
    .A(_03439_),
    .Y(_00608_));
 sg13g2_nand2_1 _09128_ (.Y(_03442_),
    .A(\i_core.cpu.i_core.mem_op[1] ),
    .B(_02068_));
 sg13g2_nand2_1 _09129_ (.Y(_03443_),
    .A(net2533),
    .B(net1247));
 sg13g2_nand3_1 _09130_ (.B(_03442_),
    .C(_03443_),
    .A(_03439_),
    .Y(_00609_));
 sg13g2_nor2_1 _09131_ (.A(net1202),
    .B(_01855_),
    .Y(_03444_));
 sg13g2_nand2_1 _09132_ (.Y(_03445_),
    .A(net1310),
    .B(_02072_));
 sg13g2_a21oi_1 _09133_ (.A1(net2392),
    .A2(net1309),
    .Y(_03446_),
    .B1(net1385));
 sg13g2_o21ai_1 _09134_ (.B1(_03446_),
    .Y(_00610_),
    .A1(_03444_),
    .A2(_03445_));
 sg13g2_a21oi_1 _09135_ (.A1(_00754_),
    .A2(net1247),
    .Y(_00611_),
    .B1(_02070_));
 sg13g2_nor2_2 _09136_ (.A(_00875_),
    .B(_01174_),
    .Y(_03447_));
 sg13g2_nor2_1 _09137_ (.A(net1312),
    .B(_01174_),
    .Y(_03448_));
 sg13g2_nand2_1 _09138_ (.Y(_03449_),
    .A(net1279),
    .B(net1336));
 sg13g2_nand2_2 _09139_ (.Y(_03450_),
    .A(net2503),
    .B(_03448_));
 sg13g2_a22oi_1 _09140_ (.Y(_03451_),
    .B1(_03450_),
    .B2(\data_to_write[0] ),
    .A2(_03448_),
    .A1(_01122_));
 sg13g2_inv_1 _09141_ (.Y(_00612_),
    .A(_03451_));
 sg13g2_nand2_1 _09142_ (.Y(_03452_),
    .A(\data_to_write[1] ),
    .B(_03450_));
 sg13g2_o21ai_1 _09143_ (.B1(_03452_),
    .Y(_00613_),
    .A1(_01065_),
    .A2(_03449_));
 sg13g2_nand2_1 _09144_ (.Y(_03453_),
    .A(net2678),
    .B(_03450_));
 sg13g2_o21ai_1 _09145_ (.B1(_03453_),
    .Y(_00614_),
    .A1(_01030_),
    .A2(_03449_));
 sg13g2_a22oi_1 _09146_ (.Y(_03454_),
    .B1(_03450_),
    .B2(net2674),
    .A2(_03448_),
    .A1(_00965_));
 sg13g2_inv_1 _09147_ (.Y(_00615_),
    .A(_03454_));
 sg13g2_xnor2_1 _09148_ (.Y(_03455_),
    .A(net1404),
    .B(net1368));
 sg13g2_nand2_2 _09149_ (.Y(_03456_),
    .A(net1336),
    .B(_03455_));
 sg13g2_a21oi_2 _09150_ (.B1(_00218_),
    .Y(_03457_),
    .A2(_00882_),
    .A1(_00880_));
 sg13g2_nand2b_2 _09151_ (.Y(_03458_),
    .B(_03457_),
    .A_N(_03456_));
 sg13g2_nor2_1 _09152_ (.A(net1279),
    .B(_01497_),
    .Y(_03459_));
 sg13g2_and2_2 _09153_ (.A(_01122_),
    .B(_03459_),
    .X(_03460_));
 sg13g2_mux2_1 _09154_ (.A0(_03460_),
    .A1(net2622),
    .S(_03458_),
    .X(_00616_));
 sg13g2_nor2b_2 _09155_ (.A(_01065_),
    .B_N(_03459_),
    .Y(_03461_));
 sg13g2_mux2_1 _09156_ (.A0(_03461_),
    .A1(net2682),
    .S(_03458_),
    .X(_00617_));
 sg13g2_nor2b_2 _09157_ (.A(_01030_),
    .B_N(_03459_),
    .Y(_03462_));
 sg13g2_mux2_1 _09158_ (.A0(_03462_),
    .A1(\data_to_write[6] ),
    .S(_03458_),
    .X(_00618_));
 sg13g2_and2_2 _09159_ (.A(_00965_),
    .B(_03459_),
    .X(_03463_));
 sg13g2_mux2_1 _09160_ (.A0(_03463_),
    .A1(net2471),
    .S(_03458_),
    .X(_00619_));
 sg13g2_nand2_1 _09161_ (.Y(_03464_),
    .A(net1357),
    .B(_03460_));
 sg13g2_nand2_2 _09162_ (.Y(_03465_),
    .A(_00995_),
    .B(net1336));
 sg13g2_nand2_1 _09163_ (.Y(_03466_),
    .A(net2458),
    .B(_03465_));
 sg13g2_o21ai_1 _09164_ (.B1(_03466_),
    .Y(_00620_),
    .A1(_03456_),
    .A2(_03464_));
 sg13g2_nand2_1 _09165_ (.Y(_03467_),
    .A(net1357),
    .B(_03461_));
 sg13g2_nand2_1 _09166_ (.Y(_03468_),
    .A(net2461),
    .B(_03465_));
 sg13g2_o21ai_1 _09167_ (.B1(_03468_),
    .Y(_00621_),
    .A1(_03456_),
    .A2(_03467_));
 sg13g2_nand2_1 _09168_ (.Y(_03469_),
    .A(net1357),
    .B(_03462_));
 sg13g2_nand2_1 _09169_ (.Y(_03470_),
    .A(net1901),
    .B(_03465_));
 sg13g2_o21ai_1 _09170_ (.B1(_03470_),
    .Y(_00622_),
    .A1(_03456_),
    .A2(_03469_));
 sg13g2_nand2_1 _09171_ (.Y(_03471_),
    .A(net1357),
    .B(_03463_));
 sg13g2_nand2_1 _09172_ (.Y(_03472_),
    .A(net1924),
    .B(_03465_));
 sg13g2_o21ai_1 _09173_ (.B1(_03472_),
    .Y(_00623_),
    .A1(_03456_),
    .A2(_03471_));
 sg13g2_nor3_2 _09174_ (.A(_00218_),
    .B(net1360),
    .C(net1357),
    .Y(_03473_));
 sg13g2_nand3_1 _09175_ (.B(_03455_),
    .C(_03473_),
    .A(net1336),
    .Y(_03474_));
 sg13g2_mux2_1 _09176_ (.A0(_03460_),
    .A1(net2133),
    .S(_03474_),
    .X(_00624_));
 sg13g2_mux2_1 _09177_ (.A0(_03461_),
    .A1(net2132),
    .S(_03474_),
    .X(_00625_));
 sg13g2_mux2_1 _09178_ (.A0(_03462_),
    .A1(net2183),
    .S(_03474_),
    .X(_00626_));
 sg13g2_mux2_1 _09179_ (.A0(_03463_),
    .A1(net2188),
    .S(_03474_),
    .X(_00627_));
 sg13g2_nand2_2 _09180_ (.Y(_03475_),
    .A(net1404),
    .B(_03447_));
 sg13g2_a22oi_1 _09181_ (.Y(_03476_),
    .B1(_03475_),
    .B2(net1990),
    .A2(_03460_),
    .A1(_03447_));
 sg13g2_inv_1 _09182_ (.Y(_00628_),
    .A(net1991));
 sg13g2_a22oi_1 _09183_ (.Y(_03477_),
    .B1(_03475_),
    .B2(net1974),
    .A2(_03461_),
    .A1(_03447_));
 sg13g2_inv_1 _09184_ (.Y(_00629_),
    .A(net1975));
 sg13g2_a22oi_1 _09185_ (.Y(_03478_),
    .B1(_03475_),
    .B2(net2037),
    .A2(_03462_),
    .A1(_03447_));
 sg13g2_inv_1 _09186_ (.Y(_00630_),
    .A(net2038));
 sg13g2_a22oi_1 _09187_ (.Y(_03479_),
    .B1(_03475_),
    .B2(net1927),
    .A2(_03463_),
    .A1(_03447_));
 sg13g2_inv_1 _09188_ (.Y(_00631_),
    .A(net1928));
 sg13g2_nor2_1 _09189_ (.A(_01174_),
    .B(_03455_),
    .Y(_03480_));
 sg13g2_nand2b_2 _09190_ (.Y(_03481_),
    .B(net1336),
    .A_N(_03455_));
 sg13g2_nand2_2 _09191_ (.Y(_03482_),
    .A(_03457_),
    .B(_03480_));
 sg13g2_mux2_1 _09192_ (.A0(_03460_),
    .A1(net2191),
    .S(_03482_),
    .X(_00632_));
 sg13g2_mux2_1 _09193_ (.A0(_03461_),
    .A1(net2184),
    .S(_03482_),
    .X(_00633_));
 sg13g2_mux2_1 _09194_ (.A0(_03462_),
    .A1(net2181),
    .S(_03482_),
    .X(_00634_));
 sg13g2_mux2_1 _09195_ (.A0(_03463_),
    .A1(net2175),
    .S(_03482_),
    .X(_00635_));
 sg13g2_nand3_1 _09196_ (.B(net1354),
    .C(net1336),
    .A(net1378),
    .Y(_03483_));
 sg13g2_nand2_1 _09197_ (.Y(_03484_),
    .A(net1938),
    .B(_03483_));
 sg13g2_o21ai_1 _09198_ (.B1(_03484_),
    .Y(_00636_),
    .A1(_03464_),
    .A2(_03481_));
 sg13g2_nand2_1 _09199_ (.Y(_03485_),
    .A(net2087),
    .B(_03483_));
 sg13g2_o21ai_1 _09200_ (.B1(_03485_),
    .Y(_00637_),
    .A1(_03467_),
    .A2(_03481_));
 sg13g2_nand2_1 _09201_ (.Y(_03486_),
    .A(net1897),
    .B(_03483_));
 sg13g2_o21ai_1 _09202_ (.B1(_03486_),
    .Y(_00638_),
    .A1(_03469_),
    .A2(_03481_));
 sg13g2_nand2_1 _09203_ (.Y(_03487_),
    .A(net1902),
    .B(_03483_));
 sg13g2_o21ai_1 _09204_ (.B1(_03487_),
    .Y(_00639_),
    .A1(_03471_),
    .A2(_03481_));
 sg13g2_and2_2 _09205_ (.A(_03473_),
    .B(_03480_),
    .X(_03488_));
 sg13g2_nand4_1 _09206_ (.B(_00820_),
    .C(net1354),
    .A(net1414),
    .Y(_03489_),
    .D(net1336));
 sg13g2_a22oi_1 _09207_ (.Y(_03490_),
    .B1(_03489_),
    .B2(net1903),
    .A2(_03488_),
    .A1(_03460_));
 sg13g2_inv_1 _09208_ (.Y(_00640_),
    .A(_03490_));
 sg13g2_a22oi_1 _09209_ (.Y(_03491_),
    .B1(_03489_),
    .B2(net1880),
    .A2(_03488_),
    .A1(_03461_));
 sg13g2_inv_1 _09210_ (.Y(_00641_),
    .A(_03491_));
 sg13g2_a22oi_1 _09211_ (.Y(_03492_),
    .B1(_03489_),
    .B2(net1890),
    .A2(_03488_),
    .A1(_03462_));
 sg13g2_inv_1 _09212_ (.Y(_00642_),
    .A(_03492_));
 sg13g2_a22oi_1 _09213_ (.Y(_03493_),
    .B1(_03489_),
    .B2(net1909),
    .A2(_03488_),
    .A1(_03463_));
 sg13g2_inv_1 _09214_ (.Y(_00643_),
    .A(_03493_));
 sg13g2_nor2_1 _09215_ (.A(net1385),
    .B(_00820_),
    .Y(_00644_));
 sg13g2_o21ai_1 _09216_ (.B1(net1462),
    .Y(_03494_),
    .A1(net1360),
    .A2(net1357));
 sg13g2_inv_1 _09217_ (.Y(_00645_),
    .A(_03494_));
 sg13g2_o21ai_1 _09218_ (.B1(net1464),
    .Y(_03495_),
    .A1(net1404),
    .A2(net1365));
 sg13g2_a21oi_1 _09219_ (.A1(net1414),
    .A2(net1354),
    .Y(_00646_),
    .B1(_03495_));
 sg13g2_nor2_1 _09220_ (.A(net2176),
    .B(_01882_),
    .Y(_03496_));
 sg13g2_o21ai_1 _09221_ (.B1(net1464),
    .Y(_03497_),
    .A1(net2401),
    .A2(net1310));
 sg13g2_a21oi_1 _09222_ (.A1(net1310),
    .A2(_03496_),
    .Y(_00647_),
    .B1(_03497_));
 sg13g2_nor3_1 _09223_ (.A(net1458),
    .B(net1310),
    .C(_03496_),
    .Y(_00648_));
 sg13g2_nand2_1 _09224_ (.Y(_03498_),
    .A(net1185),
    .B(_02388_));
 sg13g2_and2_1 _09225_ (.A(net1185),
    .B(_02389_),
    .X(_03499_));
 sg13g2_nand2_1 _09226_ (.Y(_03500_),
    .A(net1185),
    .B(_02389_));
 sg13g2_mux4_1 _09227_ (.S0(net1289),
    .A0(_00148_),
    .A1(_00147_),
    .A2(_00150_),
    .A3(_00149_),
    .S1(net1269),
    .X(_03501_));
 sg13g2_nor3_2 _09228_ (.A(net1215),
    .B(_01801_),
    .C(_01803_),
    .Y(_03502_));
 sg13g2_inv_1 _09229_ (.Y(_03503_),
    .A(_03502_));
 sg13g2_a21oi_1 _09230_ (.A1(_01752_),
    .A2(_01780_),
    .Y(_03504_),
    .B1(_01800_));
 sg13g2_and2_1 _09231_ (.A(_02399_),
    .B(_03504_),
    .X(_03505_));
 sg13g2_a221oi_1 _09232_ (.B2(_03502_),
    .C1(_03505_),
    .B1(net1246),
    .A1(net1200),
    .Y(_03506_),
    .A2(_01810_));
 sg13g2_o21ai_1 _09233_ (.B1(net1460),
    .Y(_03507_),
    .A1(net2676),
    .A2(net1159));
 sg13g2_a21oi_1 _09234_ (.A1(net1159),
    .A2(_03506_),
    .Y(_00649_),
    .B1(_03507_));
 sg13g2_or2_1 _09235_ (.X(_03508_),
    .B(_03501_),
    .A(_01817_));
 sg13g2_inv_1 _09236_ (.Y(_03509_),
    .A(_03508_));
 sg13g2_nand2_2 _09237_ (.Y(_03510_),
    .A(net1213),
    .B(_03509_));
 sg13g2_inv_1 _09238_ (.Y(_03511_),
    .A(_03510_));
 sg13g2_nand2_1 _09239_ (.Y(_03512_),
    .A(_02398_),
    .B(_02401_));
 sg13g2_a21oi_1 _09240_ (.A1(_02395_),
    .A2(_03510_),
    .Y(_03513_),
    .B1(_03512_));
 sg13g2_nor3_1 _09241_ (.A(_01790_),
    .B(net1252),
    .C(net1251),
    .Y(_03514_));
 sg13g2_nand4_1 _09242_ (.B(net1255),
    .C(net1253),
    .A(net1200),
    .Y(_03515_),
    .D(_03514_));
 sg13g2_nand3_1 _09243_ (.B(_01819_),
    .C(net1248),
    .A(_01817_),
    .Y(_03516_));
 sg13g2_nor2_2 _09244_ (.A(net1249),
    .B(_03516_),
    .Y(_03517_));
 sg13g2_nand2_2 _09245_ (.Y(_03518_),
    .A(_02405_),
    .B(_03517_));
 sg13g2_inv_1 _09246_ (.Y(_03519_),
    .A(_03518_));
 sg13g2_nand4_1 _09247_ (.B(_03513_),
    .C(_03515_),
    .A(net1158),
    .Y(_03520_),
    .D(_03518_));
 sg13g2_o21ai_1 _09248_ (.B1(_03520_),
    .Y(_03521_),
    .A1(net2628),
    .A2(net1158));
 sg13g2_nor2_1 _09249_ (.A(net1383),
    .B(_03521_),
    .Y(_00650_));
 sg13g2_nand2_1 _09250_ (.Y(_03522_),
    .A(net2210),
    .B(net1157));
 sg13g2_nor2_2 _09251_ (.A(net1199),
    .B(net1157),
    .Y(_03523_));
 sg13g2_nor3_2 _09252_ (.A(_01790_),
    .B(_01793_),
    .C(net1250),
    .Y(_03524_));
 sg13g2_and2_1 _09253_ (.A(net1253),
    .B(_03524_),
    .X(_03525_));
 sg13g2_nand2_2 _09254_ (.Y(_03526_),
    .A(_01788_),
    .B(_03524_));
 sg13g2_nand3_1 _09255_ (.B(_03523_),
    .C(net1193),
    .A(net1256),
    .Y(_03527_));
 sg13g2_a21oi_1 _09256_ (.A1(_03522_),
    .A2(_03527_),
    .Y(_00651_),
    .B1(net1384));
 sg13g2_nor2_1 _09257_ (.A(net1246),
    .B(_03503_),
    .Y(_03528_));
 sg13g2_nor2_2 _09258_ (.A(net1257),
    .B(_01803_),
    .Y(_03529_));
 sg13g2_nor3_1 _09259_ (.A(net1201),
    .B(_03528_),
    .C(_03529_),
    .Y(_03530_));
 sg13g2_nor2_2 _09260_ (.A(net1255),
    .B(_01807_),
    .Y(_03531_));
 sg13g2_or2_2 _09261_ (.X(_03532_),
    .B(_01807_),
    .A(net1255));
 sg13g2_nand2_2 _09262_ (.Y(_03533_),
    .A(net1254),
    .B(_03531_));
 sg13g2_o21ai_1 _09263_ (.B1(net1461),
    .Y(_03534_),
    .A1(net2618),
    .A2(net1158));
 sg13g2_a221oi_1 _09264_ (.B2(_03523_),
    .C1(_03534_),
    .B1(_03533_),
    .A1(net1158),
    .Y(_00652_),
    .A2(_03530_));
 sg13g2_a221oi_1 _09265_ (.B2(_03511_),
    .C1(net1200),
    .B1(_02395_),
    .A1(_01783_),
    .Y(_03535_),
    .A2(_01804_));
 sg13g2_o21ai_1 _09266_ (.B1(_03535_),
    .Y(_03536_),
    .A1(_01806_),
    .A2(_01810_));
 sg13g2_nand3b_1 _09267_ (.B(net1253),
    .C(_03514_),
    .Y(_03537_),
    .A_N(net1255));
 sg13g2_o21ai_1 _09268_ (.B1(net1459),
    .Y(_03538_),
    .A1(net1156),
    .A2(_03536_));
 sg13g2_a221oi_1 _09269_ (.B2(_03537_),
    .C1(_03538_),
    .B1(_03523_),
    .A1(_00752_),
    .Y(_00653_),
    .A2(net1156));
 sg13g2_nor2_1 _09270_ (.A(_02406_),
    .B(_03517_),
    .Y(_03539_));
 sg13g2_nor3_1 _09271_ (.A(net1198),
    .B(net1256),
    .C(net1191),
    .Y(_03540_));
 sg13g2_nor3_1 _09272_ (.A(net1156),
    .B(_03539_),
    .C(_03540_),
    .Y(_03541_));
 sg13g2_o21ai_1 _09273_ (.B1(net1460),
    .Y(_03542_),
    .A1(net2568),
    .A2(net1159));
 sg13g2_nor2_1 _09274_ (.A(_03541_),
    .B(_03542_),
    .Y(_00654_));
 sg13g2_nor2_2 _09275_ (.A(net1254),
    .B(_03532_),
    .Y(_03543_));
 sg13g2_nor2_2 _09276_ (.A(net1257),
    .B(_02394_),
    .Y(_03544_));
 sg13g2_nand2b_2 _09277_ (.Y(_03545_),
    .B(_01782_),
    .A_N(_02394_));
 sg13g2_nor2_1 _09278_ (.A(net1156),
    .B(_03545_),
    .Y(_03546_));
 sg13g2_a221oi_1 _09279_ (.B2(_03543_),
    .C1(_03546_),
    .B1(_03523_),
    .A1(net2667),
    .Y(_03547_),
    .A2(net1156));
 sg13g2_nor2_1 _09280_ (.A(net1383),
    .B(_03547_),
    .Y(_00655_));
 sg13g2_nor2_1 _09281_ (.A(_01794_),
    .B(net1250),
    .Y(_03548_));
 sg13g2_nand2_1 _09282_ (.Y(_03549_),
    .A(net1249),
    .B(net1246));
 sg13g2_nor2_1 _09283_ (.A(_03516_),
    .B(_03549_),
    .Y(_03550_));
 sg13g2_nor3_1 _09284_ (.A(_01812_),
    .B(net1156),
    .C(_03550_),
    .Y(_03551_));
 sg13g2_a221oi_1 _09285_ (.B2(_03548_),
    .C1(_03551_),
    .B1(_03523_),
    .A1(net2660),
    .Y(_03552_),
    .A2(net1156));
 sg13g2_nor2_1 _09286_ (.A(net1383),
    .B(_03552_),
    .Y(_00656_));
 sg13g2_o21ai_1 _09287_ (.B1(net1465),
    .Y(_03553_),
    .A1(_01798_),
    .A2(net1157));
 sg13g2_a21oi_1 _09288_ (.A1(_00750_),
    .A2(net1157),
    .Y(_00657_),
    .B1(_03553_));
 sg13g2_nand2_2 _09289_ (.Y(_03554_),
    .A(_02396_),
    .B(_02403_));
 sg13g2_nand2_2 _09290_ (.Y(_03555_),
    .A(_01786_),
    .B(_03545_));
 sg13g2_nor2_1 _09291_ (.A(_03554_),
    .B(_03555_),
    .Y(_03556_));
 sg13g2_nor2_2 _09292_ (.A(net1215),
    .B(_02401_),
    .Y(_03557_));
 sg13g2_nor2_1 _09293_ (.A(_01803_),
    .B(_02404_),
    .Y(_03558_));
 sg13g2_nor3_2 _09294_ (.A(net1215),
    .B(_01803_),
    .C(_02404_),
    .Y(_03559_));
 sg13g2_nand2_2 _09295_ (.Y(_03560_),
    .A(_01752_),
    .B(_03558_));
 sg13g2_and2_1 _09296_ (.A(net1215),
    .B(_03529_),
    .X(_03561_));
 sg13g2_nand2_1 _09297_ (.Y(_03562_),
    .A(net1215),
    .B(_03529_));
 sg13g2_nor3_2 _09298_ (.A(_03557_),
    .B(_03559_),
    .C(_03561_),
    .Y(_03563_));
 sg13g2_nor4_2 _09299_ (.A(_01746_),
    .B(net1215),
    .C(_01780_),
    .Y(_03564_),
    .D(net1257));
 sg13g2_nor2_1 _09300_ (.A(_03502_),
    .B(_03564_),
    .Y(_03565_));
 sg13g2_nand4_1 _09301_ (.B(_02414_),
    .C(_03563_),
    .A(_02406_),
    .Y(_03566_),
    .D(_03565_));
 sg13g2_nor3_1 _09302_ (.A(_03554_),
    .B(_03555_),
    .C(_03566_),
    .Y(_03567_));
 sg13g2_nand3_1 _09303_ (.B(_01789_),
    .C(_03514_),
    .A(net1200),
    .Y(_03568_));
 sg13g2_a22oi_1 _09304_ (.Y(_03569_),
    .B1(_03567_),
    .B2(_01752_),
    .A2(_03550_),
    .A1(_01811_));
 sg13g2_nand3_1 _09305_ (.B(_03568_),
    .C(_03569_),
    .A(net1158),
    .Y(_03570_));
 sg13g2_o21ai_1 _09306_ (.B1(_03570_),
    .Y(_03571_),
    .A1(net2591),
    .A2(net1158));
 sg13g2_nor2_1 _09307_ (.A(net1383),
    .B(_03571_),
    .Y(_00658_));
 sg13g2_nor2_1 _09308_ (.A(net2381),
    .B(net1158),
    .Y(_03572_));
 sg13g2_nor3_1 _09309_ (.A(net1387),
    .B(_03523_),
    .C(_03572_),
    .Y(_00659_));
 sg13g2_nand2_1 _09310_ (.Y(_03573_),
    .A(net2493),
    .B(net1157));
 sg13g2_nand3b_1 _09311_ (.B(_03573_),
    .C(net1464),
    .Y(_00660_),
    .A_N(_03523_));
 sg13g2_nor2_1 _09312_ (.A(net1458),
    .B(net1157),
    .Y(_03574_));
 sg13g2_nand2b_1 _09313_ (.Y(_03575_),
    .B(net1159),
    .A_N(net1458));
 sg13g2_nor2_1 _09314_ (.A(net1198),
    .B(net1193),
    .Y(_03576_));
 sg13g2_nand2_2 _09315_ (.Y(_03577_),
    .A(net1201),
    .B(net1191));
 sg13g2_nor2_1 _09316_ (.A(net1268),
    .B(net1292),
    .Y(_03578_));
 sg13g2_nor2_1 _09317_ (.A(_01741_),
    .B(net1290),
    .Y(_03579_));
 sg13g2_a22oi_1 _09318_ (.Y(_03580_),
    .B1(net1294),
    .B2(_00105_),
    .A2(net1271),
    .A1(_00106_));
 sg13g2_a22oi_1 _09319_ (.Y(_03581_),
    .B1(net1242),
    .B2(_00103_),
    .A2(net1245),
    .A1(_00104_));
 sg13g2_o21ai_1 _09320_ (.B1(_03581_),
    .Y(_03582_),
    .A1(net1242),
    .A2(_03580_));
 sg13g2_nand3b_1 _09321_ (.B(_03532_),
    .C(_01797_),
    .Y(_03583_),
    .A_N(_03582_));
 sg13g2_o21ai_1 _09322_ (.B1(_03583_),
    .Y(_03584_),
    .A1(net1248),
    .A2(_03533_));
 sg13g2_nor2_1 _09323_ (.A(net1253),
    .B(_01818_),
    .Y(_03585_));
 sg13g2_a22oi_1 _09324_ (.Y(_03586_),
    .B1(_03585_),
    .B2(_03502_),
    .A2(_03550_),
    .A1(_01805_));
 sg13g2_nor2_1 _09325_ (.A(net1214),
    .B(_02396_),
    .Y(_03587_));
 sg13g2_nand2_2 _09326_ (.Y(_03588_),
    .A(_03509_),
    .B(_03587_));
 sg13g2_nand2_1 _09327_ (.Y(_03589_),
    .A(_03586_),
    .B(_03588_));
 sg13g2_nor2_1 _09328_ (.A(net1213),
    .B(_03508_),
    .Y(_03590_));
 sg13g2_a221oi_1 _09329_ (.B2(_03584_),
    .C1(_03589_),
    .B1(_03576_),
    .A1(net1252),
    .Y(_03591_),
    .A2(_03554_));
 sg13g2_nor2_1 _09330_ (.A(net2529),
    .B(net1141),
    .Y(_03592_));
 sg13g2_a21oi_1 _09331_ (.A1(net1141),
    .A2(_03591_),
    .Y(_00661_),
    .B1(_03592_));
 sg13g2_o21ai_1 _09332_ (.B1(_03588_),
    .Y(_03593_),
    .A1(net1255),
    .A2(_03503_));
 sg13g2_o21ai_1 _09333_ (.B1(net1197),
    .Y(_03594_),
    .A1(_03567_),
    .A2(_03593_));
 sg13g2_a22oi_1 _09334_ (.Y(_03595_),
    .B1(net1293),
    .B2(_00109_),
    .A2(net1270),
    .A1(_00110_));
 sg13g2_a22oi_1 _09335_ (.Y(_03596_),
    .B1(net1243),
    .B2(_00107_),
    .A2(net1244),
    .A1(_00108_));
 sg13g2_o21ai_1 _09336_ (.B1(_03596_),
    .Y(_03597_),
    .A1(net1240),
    .A2(_03595_));
 sg13g2_nand2_1 _09337_ (.Y(_03598_),
    .A(net1249),
    .B(_03531_));
 sg13g2_a21oi_1 _09338_ (.A1(_03532_),
    .A2(_03597_),
    .Y(_03599_),
    .B1(_03577_));
 sg13g2_o21ai_1 _09339_ (.B1(_03594_),
    .Y(_03600_),
    .A1(_02426_),
    .A2(_03556_));
 sg13g2_a21oi_2 _09340_ (.B1(_03600_),
    .Y(_03601_),
    .A2(_03599_),
    .A1(_03598_));
 sg13g2_nor2_1 _09341_ (.A(net2593),
    .B(net1140),
    .Y(_03602_));
 sg13g2_a21oi_1 _09342_ (.A1(net1141),
    .A2(_03601_),
    .Y(_00662_),
    .B1(_03602_));
 sg13g2_a21oi_1 _09343_ (.A1(_01790_),
    .A2(_03588_),
    .Y(_03603_),
    .B1(_03556_));
 sg13g2_nor2_1 _09344_ (.A(_03557_),
    .B(_03564_),
    .Y(_03604_));
 sg13g2_nand2_1 _09345_ (.Y(_03605_),
    .A(_01791_),
    .B(_02408_));
 sg13g2_nor2_1 _09346_ (.A(_01819_),
    .B(_03562_),
    .Y(_03606_));
 sg13g2_a22oi_1 _09347_ (.Y(_03607_),
    .B1(net1292),
    .B2(_00113_),
    .A2(net1268),
    .A1(_00114_));
 sg13g2_a22oi_1 _09348_ (.Y(_03608_),
    .B1(net1239),
    .B2(_00111_),
    .A2(net1244),
    .A1(_00112_));
 sg13g2_o21ai_1 _09349_ (.B1(_03608_),
    .Y(_03609_),
    .A1(net1239),
    .A2(_03607_));
 sg13g2_a21o_1 _09350_ (.A2(_03531_),
    .A1(_01819_),
    .B1(_03577_),
    .X(_03610_));
 sg13g2_a21oi_1 _09351_ (.A1(_03532_),
    .A2(_03609_),
    .Y(_03611_),
    .B1(_03610_));
 sg13g2_o21ai_1 _09352_ (.B1(_03605_),
    .Y(_03612_),
    .A1(net1254),
    .A2(_03604_));
 sg13g2_nor4_2 _09353_ (.A(_03603_),
    .B(_03606_),
    .C(_03611_),
    .Y(_03613_),
    .D(_03612_));
 sg13g2_nor2_1 _09354_ (.A(net2604),
    .B(net1142),
    .Y(_03614_));
 sg13g2_a21oi_1 _09355_ (.A1(net1142),
    .A2(_03613_),
    .Y(_00663_),
    .B1(_03614_));
 sg13g2_nor2_1 _09356_ (.A(_01785_),
    .B(_03557_),
    .Y(_03615_));
 sg13g2_nor2_1 _09357_ (.A(_02408_),
    .B(_03554_),
    .Y(_03616_));
 sg13g2_a21oi_1 _09358_ (.A1(_03615_),
    .A2(_03616_),
    .Y(_03617_),
    .B1(net1256));
 sg13g2_or3_1 _09359_ (.A(_03544_),
    .B(_03561_),
    .C(_03564_),
    .X(_03618_));
 sg13g2_a22oi_1 _09360_ (.Y(_03619_),
    .B1(net1293),
    .B2(_00129_),
    .A2(net1270),
    .A1(_00130_));
 sg13g2_a22oi_1 _09361_ (.Y(_03620_),
    .B1(net1241),
    .B2(_00127_),
    .A2(net1245),
    .A1(_00128_));
 sg13g2_o21ai_1 _09362_ (.B1(_03620_),
    .Y(_03621_),
    .A1(net1241),
    .A2(_03619_));
 sg13g2_nand2_1 _09363_ (.Y(_03622_),
    .A(_01817_),
    .B(_03531_));
 sg13g2_a21oi_1 _09364_ (.A1(_03532_),
    .A2(_03621_),
    .Y(_03623_),
    .B1(_03577_));
 sg13g2_a22oi_1 _09365_ (.Y(_03624_),
    .B1(_03622_),
    .B2(_03623_),
    .A2(_03618_),
    .A1(_01818_));
 sg13g2_nand2_1 _09366_ (.Y(_03625_),
    .A(_03588_),
    .B(_03624_));
 sg13g2_nor3_1 _09367_ (.A(net1135),
    .B(_03617_),
    .C(_03625_),
    .Y(_03626_));
 sg13g2_a21oi_1 _09368_ (.A1(_00797_),
    .A2(net1135),
    .Y(_00664_),
    .B1(_03626_));
 sg13g2_nand2_1 _09369_ (.Y(_03627_),
    .A(net1254),
    .B(_03588_));
 sg13g2_and2_1 _09370_ (.A(_01801_),
    .B(_02400_),
    .X(_03628_));
 sg13g2_nor2_1 _09371_ (.A(_03554_),
    .B(_03628_),
    .Y(_03629_));
 sg13g2_o21ai_1 _09372_ (.B1(_03629_),
    .Y(_03630_),
    .A1(net1254),
    .A2(_03518_));
 sg13g2_nor4_1 _09373_ (.A(_01785_),
    .B(_03557_),
    .C(_03559_),
    .D(_03618_),
    .Y(_03631_));
 sg13g2_a22oi_1 _09374_ (.Y(_03632_),
    .B1(net1292),
    .B2(_00133_),
    .A2(net1268),
    .A1(_00134_));
 sg13g2_a22oi_1 _09375_ (.Y(_03633_),
    .B1(net1239),
    .B2(_00131_),
    .A2(net1244),
    .A1(_00132_));
 sg13g2_o21ai_1 _09376_ (.B1(_03633_),
    .Y(_03634_),
    .A1(net1239),
    .A2(_03632_));
 sg13g2_nand2_1 _09377_ (.Y(_03635_),
    .A(_03532_),
    .B(_03634_));
 sg13g2_a21oi_1 _09378_ (.A1(net1246),
    .A2(_03531_),
    .Y(_03636_),
    .B1(_03577_));
 sg13g2_a22oi_1 _09379_ (.Y(_03637_),
    .B1(_03635_),
    .B2(_03636_),
    .A2(_03630_),
    .A1(_03627_));
 sg13g2_o21ai_1 _09380_ (.B1(_03637_),
    .Y(_03638_),
    .A1(net1246),
    .A2(_03631_));
 sg13g2_mux2_1 _09381_ (.A0(net2560),
    .A1(_03638_),
    .S(net1141),
    .X(_00665_));
 sg13g2_nand3_1 _09382_ (.B(_03604_),
    .C(_03616_),
    .A(_03562_),
    .Y(_03639_));
 sg13g2_nand2_1 _09383_ (.Y(_03640_),
    .A(net1184),
    .B(_03518_));
 sg13g2_o21ai_1 _09384_ (.B1(_01792_),
    .Y(_03641_),
    .A1(_03555_),
    .A2(_03640_));
 sg13g2_a22oi_1 _09385_ (.Y(_03642_),
    .B1(net1292),
    .B2(_00137_),
    .A2(net1268),
    .A1(_00138_));
 sg13g2_a22oi_1 _09386_ (.Y(_03643_),
    .B1(net1239),
    .B2(_00135_),
    .A2(net1244),
    .A1(_00136_));
 sg13g2_o21ai_1 _09387_ (.B1(_03643_),
    .Y(_03644_),
    .A1(net1239),
    .A2(_03642_));
 sg13g2_nor2_2 _09388_ (.A(net1196),
    .B(_03644_),
    .Y(_03645_));
 sg13g2_o21ai_1 _09389_ (.B1(_03641_),
    .Y(_03646_),
    .A1(_01817_),
    .A2(_03560_));
 sg13g2_a221oi_1 _09390_ (.B2(_03526_),
    .C1(_03646_),
    .B1(_03645_),
    .A1(_01828_),
    .Y(_03647_),
    .A2(_03639_));
 sg13g2_nor2_1 _09391_ (.A(net2625),
    .B(net1141),
    .Y(_03648_));
 sg13g2_a21oi_1 _09392_ (.A1(net1140),
    .A2(_03647_),
    .Y(_00666_),
    .B1(_03648_));
 sg13g2_nor3_1 _09393_ (.A(_03544_),
    .B(_03564_),
    .C(_03640_),
    .Y(_03649_));
 sg13g2_a21oi_1 _09394_ (.A1(_01786_),
    .A2(_03563_),
    .Y(_03650_),
    .B1(net1248));
 sg13g2_a21oi_2 _09395_ (.B1(net1214),
    .Y(_03651_),
    .A2(_02403_),
    .A1(_02396_));
 sg13g2_a22oi_1 _09396_ (.Y(_03652_),
    .B1(net1294),
    .B2(_00141_),
    .A2(net1272),
    .A1(_00142_));
 sg13g2_a22oi_1 _09397_ (.Y(_03653_),
    .B1(net1242),
    .B2(_00139_),
    .A2(net1245),
    .A1(_00140_));
 sg13g2_o21ai_1 _09398_ (.B1(_03653_),
    .Y(_03654_),
    .A1(net1242),
    .A2(_03652_));
 sg13g2_nor2_1 _09399_ (.A(_03577_),
    .B(_03654_),
    .Y(_03655_));
 sg13g2_a21oi_1 _09400_ (.A1(_01792_),
    .A2(_02408_),
    .Y(_03656_),
    .B1(_03651_));
 sg13g2_o21ai_1 _09401_ (.B1(_03656_),
    .Y(_03657_),
    .A1(net1256),
    .A2(_03649_));
 sg13g2_nor4_2 _09402_ (.A(net1135),
    .B(_03650_),
    .C(_03655_),
    .Y(_03658_),
    .D(_03657_));
 sg13g2_a21oi_1 _09403_ (.A1(_00801_),
    .A2(net1135),
    .Y(_00667_),
    .B1(_03658_));
 sg13g2_o21ai_1 _09404_ (.B1(net1251),
    .Y(_03659_),
    .A1(_03519_),
    .A2(_03628_));
 sg13g2_o21ai_1 _09405_ (.B1(_03659_),
    .Y(_03660_),
    .A1(net1249),
    .A2(_03563_));
 sg13g2_a22oi_1 _09406_ (.Y(_03661_),
    .B1(net1292),
    .B2(_00149_),
    .A2(net1269),
    .A1(_00150_));
 sg13g2_a22oi_1 _09407_ (.Y(_03662_),
    .B1(net1240),
    .B2(_00147_),
    .A2(net1244),
    .A1(_00148_));
 sg13g2_o21ai_1 _09408_ (.B1(_03662_),
    .Y(_03663_),
    .A1(net1239),
    .A2(_03661_));
 sg13g2_nand2b_1 _09409_ (.Y(_03664_),
    .B(_03555_),
    .A_N(net1254));
 sg13g2_o21ai_1 _09410_ (.B1(_03664_),
    .Y(_03665_),
    .A1(_03577_),
    .A2(_03663_));
 sg13g2_nor4_2 _09411_ (.A(net1135),
    .B(_03651_),
    .C(_03660_),
    .Y(_03666_),
    .D(_03665_));
 sg13g2_a21oi_1 _09412_ (.A1(_00798_),
    .A2(net1135),
    .Y(_00668_),
    .B1(_03666_));
 sg13g2_a21o_1 _09413_ (.A2(_03545_),
    .A1(_02403_),
    .B1(net1213),
    .X(_03667_));
 sg13g2_nor2_1 _09414_ (.A(_03508_),
    .B(_03524_),
    .Y(_03668_));
 sg13g2_nor3_2 _09415_ (.A(net1214),
    .B(_02396_),
    .C(_03668_),
    .Y(_03669_));
 sg13g2_a21oi_1 _09416_ (.A1(net1251),
    .A2(_03587_),
    .Y(_03670_),
    .B1(_03669_));
 sg13g2_nand2_1 _09417_ (.Y(_03671_),
    .A(_03667_),
    .B(_03670_));
 sg13g2_a21oi_1 _09418_ (.A1(net1184),
    .A2(_03518_),
    .Y(_03672_),
    .B1(_01790_));
 sg13g2_a22oi_1 _09419_ (.Y(_03673_),
    .B1(net1294),
    .B2(_00145_),
    .A2(net1272),
    .A1(_00146_));
 sg13g2_a22oi_1 _09420_ (.Y(_03674_),
    .B1(net1241),
    .B2(_00143_),
    .A2(net1245),
    .A1(_00144_));
 sg13g2_o21ai_1 _09421_ (.B1(_03674_),
    .Y(_03675_),
    .A1(net1241),
    .A2(_03673_));
 sg13g2_nor2_1 _09422_ (.A(_03577_),
    .B(_03675_),
    .Y(_03676_));
 sg13g2_a21oi_1 _09423_ (.A1(_03560_),
    .A2(_03615_),
    .Y(_03677_),
    .B1(_01819_));
 sg13g2_nor4_2 _09424_ (.A(_03671_),
    .B(_03672_),
    .C(_03676_),
    .Y(_03678_),
    .D(_03677_));
 sg13g2_nor2_1 _09425_ (.A(net2653),
    .B(net1142),
    .Y(_03679_));
 sg13g2_a21oi_1 _09426_ (.A1(net1142),
    .A2(_03678_),
    .Y(_00669_),
    .B1(_03679_));
 sg13g2_a21oi_1 _09427_ (.A1(_03518_),
    .A2(_03560_),
    .Y(_03680_),
    .B1(net1213));
 sg13g2_o21ai_1 _09428_ (.B1(_03667_),
    .Y(_03681_),
    .A1(net1214),
    .A2(net1184));
 sg13g2_nor2_1 _09429_ (.A(_03680_),
    .B(_03681_),
    .Y(_03682_));
 sg13g2_nand2_1 _09430_ (.Y(_03683_),
    .A(_03670_),
    .B(_03682_));
 sg13g2_a22oi_1 _09431_ (.Y(_03684_),
    .B1(net1294),
    .B2(_00117_),
    .A2(net1271),
    .A1(_00118_));
 sg13g2_nand2b_1 _09432_ (.Y(_03685_),
    .B(_03684_),
    .A_N(net1241));
 sg13g2_nand2b_1 _09433_ (.Y(_03686_),
    .B(net1241),
    .A_N(_00115_));
 sg13g2_a221oi_1 _09434_ (.B2(_03686_),
    .C1(net1196),
    .B1(_03685_),
    .A1(_00116_),
    .Y(_03687_),
    .A2(net1245));
 sg13g2_a21oi_1 _09435_ (.A1(_03526_),
    .A2(_03687_),
    .Y(_03688_),
    .B1(_03683_));
 sg13g2_o21ai_1 _09436_ (.B1(_03688_),
    .Y(_03689_),
    .A1(_01817_),
    .A2(_03615_));
 sg13g2_mux2_1 _09437_ (.A0(net2643),
    .A1(_03689_),
    .S(net1141),
    .X(_00670_));
 sg13g2_a22oi_1 _09438_ (.Y(_03690_),
    .B1(net1293),
    .B2(_00121_),
    .A2(net1270),
    .A1(_00122_));
 sg13g2_nor2_1 _09439_ (.A(net1240),
    .B(_03690_),
    .Y(_03691_));
 sg13g2_a221oi_1 _09440_ (.B2(_00119_),
    .C1(_03691_),
    .B1(net1240),
    .A1(_00120_),
    .Y(_03692_),
    .A2(net1244));
 sg13g2_a221oi_1 _09441_ (.B2(_03692_),
    .C1(_03683_),
    .B1(_03576_),
    .A1(_01785_),
    .Y(_03693_),
    .A2(_01822_));
 sg13g2_nor2_1 _09442_ (.A(net2658),
    .B(net1142),
    .Y(_03694_));
 sg13g2_a21oi_1 _09443_ (.A1(net1142),
    .A2(_03693_),
    .Y(_00671_),
    .B1(_03694_));
 sg13g2_nor2_1 _09444_ (.A(_01786_),
    .B(net1213),
    .Y(_03695_));
 sg13g2_nor2_1 _09445_ (.A(_03683_),
    .B(_03695_),
    .Y(_03696_));
 sg13g2_a22oi_1 _09446_ (.Y(_03697_),
    .B1(net1292),
    .B2(_00125_),
    .A2(net1269),
    .A1(_00126_));
 sg13g2_a22oi_1 _09447_ (.Y(_03698_),
    .B1(net1240),
    .B2(_00123_),
    .A2(net1244),
    .A1(_00124_));
 sg13g2_o21ai_1 _09448_ (.B1(_03698_),
    .Y(_03699_),
    .A1(net1240),
    .A2(_03697_));
 sg13g2_nor2_1 _09449_ (.A(_01796_),
    .B(_03699_),
    .Y(_03700_));
 sg13g2_nor2_1 _09450_ (.A(_01797_),
    .B(_03582_),
    .Y(_03701_));
 sg13g2_nor3_1 _09451_ (.A(_03543_),
    .B(_03700_),
    .C(_03701_),
    .Y(_03702_));
 sg13g2_a21o_1 _09452_ (.A2(_03543_),
    .A1(net1248),
    .B1(_03702_),
    .X(_03703_));
 sg13g2_o21ai_1 _09453_ (.B1(_03696_),
    .Y(_03704_),
    .A1(_03577_),
    .A2(_03703_));
 sg13g2_mux2_1 _09454_ (.A0(net2637),
    .A1(_03704_),
    .S(net1141),
    .X(_00672_));
 sg13g2_nand2_1 _09455_ (.Y(_03705_),
    .A(net1194),
    .B(_03696_));
 sg13g2_nor2_2 _09456_ (.A(_01796_),
    .B(net1192),
    .Y(_03706_));
 sg13g2_nor2_2 _09457_ (.A(net1194),
    .B(_03706_),
    .Y(_03707_));
 sg13g2_a21oi_1 _09458_ (.A1(net1191),
    .A2(_03700_),
    .Y(_03708_),
    .B1(net1195));
 sg13g2_a21oi_1 _09459_ (.A1(net1195),
    .A2(_03696_),
    .Y(_03709_),
    .B1(_03708_));
 sg13g2_a221oi_1 _09460_ (.B2(_01828_),
    .C1(_03709_),
    .B1(_03707_),
    .A1(net1252),
    .Y(_03710_),
    .A2(_03539_));
 sg13g2_nor2_1 _09461_ (.A(net2428),
    .B(net1140),
    .Y(_03711_));
 sg13g2_a21oi_1 _09462_ (.A1(net1140),
    .A2(_03710_),
    .Y(_00673_),
    .B1(_03711_));
 sg13g2_a221oi_1 _09463_ (.B2(_01780_),
    .C1(_03709_),
    .B1(_03707_),
    .A1(net1250),
    .Y(_03712_),
    .A2(_03539_));
 sg13g2_nor2_1 _09464_ (.A(net2520),
    .B(net1140),
    .Y(_03713_));
 sg13g2_a21oi_1 _09465_ (.A1(net1140),
    .A2(_03712_),
    .Y(_00674_),
    .B1(_03713_));
 sg13g2_nor2_1 _09466_ (.A(net1197),
    .B(_01781_),
    .Y(_03714_));
 sg13g2_a221oi_1 _09467_ (.B2(_01782_),
    .C1(_03709_),
    .B1(_03707_),
    .A1(_01791_),
    .Y(_03715_),
    .A2(_03539_));
 sg13g2_nor2_1 _09468_ (.A(net2553),
    .B(net1140),
    .Y(_03716_));
 sg13g2_a21oi_1 _09469_ (.A1(net1140),
    .A2(_03715_),
    .Y(_00675_),
    .B1(_03716_));
 sg13g2_nor3_1 _09470_ (.A(net1256),
    .B(_02406_),
    .C(_03517_),
    .Y(_03717_));
 sg13g2_o21ai_1 _09471_ (.B1(_03708_),
    .Y(_03718_),
    .A1(_01802_),
    .A2(_03706_));
 sg13g2_o21ai_1 _09472_ (.B1(_03718_),
    .Y(_03719_),
    .A1(_03705_),
    .A2(_03717_));
 sg13g2_nand2_1 _09473_ (.Y(_03720_),
    .A(net2459),
    .B(net1133));
 sg13g2_o21ai_1 _09474_ (.B1(_03720_),
    .Y(_00676_),
    .A1(net1133),
    .A2(_03719_));
 sg13g2_a22oi_1 _09475_ (.Y(_03721_),
    .B1(net1292),
    .B2(\i_core.cpu.instr_data[2][0] ),
    .A2(net1270),
    .A1(\i_core.cpu.instr_data[3][0] ));
 sg13g2_a22oi_1 _09476_ (.Y(_03722_),
    .B1(net1241),
    .B2(\i_core.cpu.instr_data[0][0] ),
    .A2(net1245),
    .A1(\i_core.cpu.instr_data[1][0] ));
 sg13g2_o21ai_1 _09477_ (.B1(_03722_),
    .Y(_03723_),
    .A1(net1241),
    .A2(_03721_));
 sg13g2_o21ai_1 _09478_ (.B1(_03723_),
    .Y(_03724_),
    .A1(_01796_),
    .A2(net1192));
 sg13g2_nor3_1 _09479_ (.A(_03669_),
    .B(_03681_),
    .C(_03695_),
    .Y(_03725_));
 sg13g2_nor3_1 _09480_ (.A(net1254),
    .B(_02406_),
    .C(_03517_),
    .Y(_03726_));
 sg13g2_nor3_1 _09481_ (.A(net1201),
    .B(_03680_),
    .C(_03726_),
    .Y(_03727_));
 sg13g2_a221oi_1 _09482_ (.B2(_03727_),
    .C1(net1134),
    .B1(_03725_),
    .A1(_03708_),
    .Y(_03728_),
    .A2(_03724_));
 sg13g2_a21o_1 _09483_ (.A2(net1134),
    .A1(net2504),
    .B1(_03728_),
    .X(_00677_));
 sg13g2_o21ai_1 _09484_ (.B1(_01828_),
    .Y(_03729_),
    .A1(_02405_),
    .A2(_03559_));
 sg13g2_nand2_1 _09485_ (.Y(_03730_),
    .A(_03725_),
    .B(_03729_));
 sg13g2_nor2_1 _09486_ (.A(net1194),
    .B(_03699_),
    .Y(_03731_));
 sg13g2_a21oi_1 _09487_ (.A1(_03706_),
    .A2(_03731_),
    .Y(_03732_),
    .B1(_03730_));
 sg13g2_inv_1 _09488_ (.Y(_03733_),
    .A(_03732_));
 sg13g2_mux4_1 _09489_ (.S0(_01741_),
    .A0(\i_core.cpu.instr_data[0][1] ),
    .A1(\i_core.cpu.instr_data[2][1] ),
    .A2(\i_core.cpu.instr_data[3][1] ),
    .A3(\i_core.cpu.instr_data[1][1] ),
    .S1(net1290),
    .X(_03734_));
 sg13g2_nand2_1 _09490_ (.Y(_03735_),
    .A(net1201),
    .B(_03734_));
 sg13g2_o21ai_1 _09491_ (.B1(_03732_),
    .Y(_03736_),
    .A1(_03706_),
    .A2(_03735_));
 sg13g2_mux2_1 _09492_ (.A0(net2517),
    .A1(_03736_),
    .S(net1137),
    .X(_00678_));
 sg13g2_mux4_1 _09493_ (.S0(net1271),
    .A0(\i_core.cpu.instr_data[1][2] ),
    .A1(\i_core.cpu.instr_data[3][2] ),
    .A2(\i_core.cpu.instr_data[2][2] ),
    .A3(\i_core.cpu.instr_data[0][2] ),
    .S1(net1294),
    .X(_03737_));
 sg13g2_nand2_2 _09494_ (.Y(_03738_),
    .A(net1201),
    .B(_03737_));
 sg13g2_o21ai_1 _09495_ (.B1(_03732_),
    .Y(_03739_),
    .A1(_03706_),
    .A2(_03738_));
 sg13g2_mux2_1 _09496_ (.A0(net2580),
    .A1(_03739_),
    .S(net1139),
    .X(_00679_));
 sg13g2_a22oi_1 _09497_ (.Y(_03740_),
    .B1(net1292),
    .B2(\i_core.cpu.instr_data[2][3] ),
    .A2(net1268),
    .A1(\i_core.cpu.instr_data[3][3] ));
 sg13g2_a22oi_1 _09498_ (.Y(_03741_),
    .B1(net1239),
    .B2(\i_core.cpu.instr_data[0][3] ),
    .A2(net1244),
    .A1(\i_core.cpu.instr_data[1][3] ));
 sg13g2_o21ai_1 _09499_ (.B1(_03741_),
    .Y(_03742_),
    .A1(net1240),
    .A2(_03740_));
 sg13g2_a21oi_1 _09500_ (.A1(_03707_),
    .A2(_03742_),
    .Y(_03743_),
    .B1(_03733_));
 sg13g2_nor2_1 _09501_ (.A(net2500),
    .B(net1139),
    .Y(_03744_));
 sg13g2_a21oi_1 _09502_ (.A1(net1139),
    .A2(_03743_),
    .Y(_00680_),
    .B1(_03744_));
 sg13g2_a21o_1 _09503_ (.A2(_03731_),
    .A1(net1191),
    .B1(_03730_),
    .X(_03745_));
 sg13g2_nor2_2 _09504_ (.A(net1195),
    .B(_03582_),
    .Y(_03746_));
 sg13g2_a21oi_1 _09505_ (.A1(net1192),
    .A2(_03746_),
    .Y(_03747_),
    .B1(net1175));
 sg13g2_nor2_1 _09506_ (.A(net2526),
    .B(net1138),
    .Y(_03748_));
 sg13g2_a21oi_1 _09507_ (.A1(net1138),
    .A2(_03747_),
    .Y(_00681_),
    .B1(_03748_));
 sg13g2_nor2_1 _09508_ (.A(net1195),
    .B(_03597_),
    .Y(_03749_));
 sg13g2_a21oi_1 _09509_ (.A1(net1192),
    .A2(_03749_),
    .Y(_03750_),
    .B1(net1175));
 sg13g2_nor2_1 _09510_ (.A(net2594),
    .B(net1137),
    .Y(_03751_));
 sg13g2_a21oi_1 _09511_ (.A1(net1138),
    .A2(_03750_),
    .Y(_00682_),
    .B1(_03751_));
 sg13g2_nor2_2 _09512_ (.A(net1194),
    .B(_03609_),
    .Y(_03752_));
 sg13g2_a21oi_1 _09513_ (.A1(net1193),
    .A2(_03752_),
    .Y(_03753_),
    .B1(net1175));
 sg13g2_nor2_1 _09514_ (.A(net2516),
    .B(net1137),
    .Y(_03754_));
 sg13g2_a21oi_1 _09515_ (.A1(net1137),
    .A2(_03753_),
    .Y(_00683_),
    .B1(_03754_));
 sg13g2_nor2_2 _09516_ (.A(net1196),
    .B(_03621_),
    .Y(_03755_));
 sg13g2_a21oi_1 _09517_ (.A1(net1192),
    .A2(_03755_),
    .Y(_03756_),
    .B1(net1175));
 sg13g2_nor2_1 _09518_ (.A(net2466),
    .B(net1137),
    .Y(_03757_));
 sg13g2_a21oi_1 _09519_ (.A1(net1137),
    .A2(_03756_),
    .Y(_00684_),
    .B1(_03757_));
 sg13g2_nor3_1 _09520_ (.A(net1194),
    .B(net1191),
    .C(_03634_),
    .Y(_03758_));
 sg13g2_nor3_1 _09521_ (.A(net1133),
    .B(_03745_),
    .C(_03758_),
    .Y(_03759_));
 sg13g2_a21oi_1 _09522_ (.A1(_00804_),
    .A2(net1134),
    .Y(_00685_),
    .B1(_03759_));
 sg13g2_a21oi_1 _09523_ (.A1(net1192),
    .A2(_03645_),
    .Y(_03760_),
    .B1(_03745_));
 sg13g2_nor2_1 _09524_ (.A(net2032),
    .B(net1138),
    .Y(_03761_));
 sg13g2_a21oi_1 _09525_ (.A1(net1138),
    .A2(_03760_),
    .Y(_00686_),
    .B1(_03761_));
 sg13g2_nor3_1 _09526_ (.A(net1194),
    .B(net1191),
    .C(_03654_),
    .Y(_03762_));
 sg13g2_nor3_1 _09527_ (.A(net1133),
    .B(net1175),
    .C(_03762_),
    .Y(_03763_));
 sg13g2_a21oi_1 _09528_ (.A1(_00802_),
    .A2(net1134),
    .Y(_00687_),
    .B1(_03763_));
 sg13g2_nor3_1 _09529_ (.A(net1194),
    .B(net1191),
    .C(_03663_),
    .Y(_03764_));
 sg13g2_nor3_1 _09530_ (.A(net1133),
    .B(net1175),
    .C(_03764_),
    .Y(_03765_));
 sg13g2_a21oi_1 _09531_ (.A1(_00799_),
    .A2(net1133),
    .Y(_00688_),
    .B1(_03765_));
 sg13g2_nor3_1 _09532_ (.A(net1194),
    .B(net1191),
    .C(_03675_),
    .Y(_03766_));
 sg13g2_nor3_1 _09533_ (.A(net1133),
    .B(_03745_),
    .C(_03766_),
    .Y(_03767_));
 sg13g2_a21oi_1 _09534_ (.A1(_00805_),
    .A2(net1134),
    .Y(_00689_),
    .B1(_03767_));
 sg13g2_a21oi_1 _09535_ (.A1(net1192),
    .A2(_03687_),
    .Y(_03768_),
    .B1(net1175));
 sg13g2_nor2_1 _09536_ (.A(net2125),
    .B(net1137),
    .Y(_03769_));
 sg13g2_a21oi_1 _09537_ (.A1(net1137),
    .A2(_03768_),
    .Y(_00690_),
    .B1(_03769_));
 sg13g2_nand3_1 _09538_ (.B(net1192),
    .C(_03692_),
    .A(net1201),
    .Y(_03770_));
 sg13g2_nor2b_1 _09539_ (.A(net1175),
    .B_N(_03770_),
    .Y(_03771_));
 sg13g2_nor2_1 _09540_ (.A(net2097),
    .B(net1138),
    .Y(_03772_));
 sg13g2_a21oi_1 _09541_ (.A1(net1138),
    .A2(_03771_),
    .Y(_00691_),
    .B1(_03772_));
 sg13g2_nor3_1 _09542_ (.A(net1133),
    .B(_03730_),
    .C(_03731_),
    .Y(_03773_));
 sg13g2_a21oi_1 _09543_ (.A1(_00800_),
    .A2(net1134),
    .Y(_00692_),
    .B1(_03773_));
 sg13g2_nand2_1 _09544_ (.Y(_03774_),
    .A(net1200),
    .B(_01794_));
 sg13g2_a221oi_1 _09545_ (.B2(net1255),
    .C1(_03774_),
    .B1(net1193),
    .A1(_01788_),
    .Y(_03775_),
    .A2(_01808_));
 sg13g2_nor2_1 _09546_ (.A(_03537_),
    .B(_03654_),
    .Y(_03776_));
 sg13g2_or2_1 _09547_ (.X(_03777_),
    .B(_03776_),
    .A(_03543_));
 sg13g2_inv_1 _09548_ (.Y(_03778_),
    .A(_03777_));
 sg13g2_nand2_1 _09549_ (.Y(_03779_),
    .A(_01780_),
    .B(_03543_));
 sg13g2_o21ai_1 _09550_ (.B1(_03779_),
    .Y(_03780_),
    .A1(net1213),
    .A2(_03777_));
 sg13g2_nand2_1 _09551_ (.Y(_03781_),
    .A(_03775_),
    .B(_03780_));
 sg13g2_a21oi_1 _09552_ (.A1(_03524_),
    .A2(_03590_),
    .Y(_03782_),
    .B1(_02396_));
 sg13g2_o21ai_1 _09553_ (.B1(_03782_),
    .Y(_03783_),
    .A1(_01789_),
    .A2(_03510_));
 sg13g2_and4_2 _09554_ (.A(_02402_),
    .B(net1142),
    .C(_03781_),
    .D(_03783_),
    .X(_03784_));
 sg13g2_a21oi_1 _09555_ (.A1(_00792_),
    .A2(net1136),
    .Y(_00693_),
    .B1(_03784_));
 sg13g2_nand2_1 _09556_ (.Y(_03785_),
    .A(_01781_),
    .B(_03543_));
 sg13g2_a22oi_1 _09557_ (.Y(_03786_),
    .B1(_03778_),
    .B2(_01779_),
    .A2(_03543_),
    .A1(net1257));
 sg13g2_a21oi_1 _09558_ (.A1(net1253),
    .A2(_03511_),
    .Y(_03787_),
    .B1(net1246));
 sg13g2_a22oi_1 _09559_ (.Y(_03788_),
    .B1(_03787_),
    .B2(_03782_),
    .A2(_03786_),
    .A1(_03775_));
 sg13g2_and3_2 _09560_ (.X(_03789_),
    .A(_02407_),
    .B(net1142),
    .C(_03788_));
 sg13g2_a21oi_1 _09561_ (.A1(net1374),
    .A2(net1136),
    .Y(_00694_),
    .B1(_03789_));
 sg13g2_o21ai_1 _09562_ (.B1(_03785_),
    .Y(_03790_),
    .A1(net1257),
    .A2(_03777_));
 sg13g2_nor2_1 _09563_ (.A(_01809_),
    .B(_03510_),
    .Y(_03791_));
 sg13g2_o21ai_1 _09564_ (.B1(_03545_),
    .Y(_03792_),
    .A1(_02396_),
    .A2(_03791_));
 sg13g2_a21oi_2 _09565_ (.B1(_03792_),
    .Y(_03793_),
    .A2(_03790_),
    .A1(_03775_));
 sg13g2_nor2_1 _09566_ (.A(net1394),
    .B(net1143),
    .Y(_03794_));
 sg13g2_a21oi_1 _09567_ (.A1(net1143),
    .A2(_03793_),
    .Y(_00695_),
    .B1(_03794_));
 sg13g2_o21ai_1 _09568_ (.B1(net1255),
    .Y(_03795_),
    .A1(_01780_),
    .A2(net1213));
 sg13g2_a21oi_1 _09569_ (.A1(_03692_),
    .A2(_03795_),
    .Y(_03796_),
    .B1(_03776_));
 sg13g2_nor2_1 _09570_ (.A(_03543_),
    .B(_03796_),
    .Y(_03797_));
 sg13g2_a21oi_1 _09571_ (.A1(_01818_),
    .A2(net1246),
    .Y(_03798_),
    .B1(_03791_));
 sg13g2_o21ai_1 _09572_ (.B1(_02407_),
    .Y(_03799_),
    .A1(_02396_),
    .A2(_03798_));
 sg13g2_a21oi_2 _09573_ (.B1(_03799_),
    .Y(_03800_),
    .A2(_03797_),
    .A1(_03775_));
 sg13g2_nor2_1 _09574_ (.A(net2666),
    .B(net1143),
    .Y(_03801_));
 sg13g2_a21oi_1 _09575_ (.A1(net1143),
    .A2(_03800_),
    .Y(_00696_),
    .B1(_03801_));
 sg13g2_and4_1 _09576_ (.A(_01780_),
    .B(net1253),
    .C(_01808_),
    .D(_01828_),
    .X(_03802_));
 sg13g2_nor3_1 _09577_ (.A(net1196),
    .B(_01827_),
    .C(_03802_),
    .Y(_03803_));
 sg13g2_nor2_1 _09578_ (.A(_03505_),
    .B(_03529_),
    .Y(_03804_));
 sg13g2_nand3_1 _09579_ (.B(_03545_),
    .C(_03804_),
    .A(_01818_),
    .Y(_03805_));
 sg13g2_o21ai_1 _09580_ (.B1(_03805_),
    .Y(_03806_),
    .A1(_02394_),
    .A2(_02404_));
 sg13g2_a21oi_1 _09581_ (.A1(net1196),
    .A2(_03806_),
    .Y(_03807_),
    .B1(_03803_));
 sg13g2_nor2_1 _09582_ (.A(net2665),
    .B(net1139),
    .Y(_03808_));
 sg13g2_a21oi_1 _09583_ (.A1(net1139),
    .A2(_03807_),
    .Y(_00697_),
    .B1(_03808_));
 sg13g2_o21ai_1 _09584_ (.B1(_03804_),
    .Y(_03809_),
    .A1(net1196),
    .A2(_01779_));
 sg13g2_mux2_1 _09585_ (.A0(net2588),
    .A1(_03809_),
    .S(net1139),
    .X(_00698_));
 sg13g2_nand2b_1 _09586_ (.Y(_03810_),
    .B(_01818_),
    .A_N(net1254));
 sg13g2_nand3_1 _09587_ (.B(net1246),
    .C(_03810_),
    .A(net1196),
    .Y(_03811_));
 sg13g2_nor4_2 _09588_ (.A(_03505_),
    .B(_03529_),
    .C(_03544_),
    .Y(_03812_),
    .D(_03811_));
 sg13g2_nor3_1 _09589_ (.A(_01828_),
    .B(_02404_),
    .C(_03533_),
    .Y(_03813_));
 sg13g2_nor2_1 _09590_ (.A(_03802_),
    .B(_03813_),
    .Y(_03814_));
 sg13g2_inv_1 _09591_ (.Y(_03815_),
    .A(_03814_));
 sg13g2_a21oi_2 _09592_ (.B1(_03812_),
    .Y(_03816_),
    .A2(_03814_),
    .A1(_03714_));
 sg13g2_nor2_1 _09593_ (.A(net2287),
    .B(net1139),
    .Y(_03817_));
 sg13g2_a21oi_1 _09594_ (.A1(net1139),
    .A2(_03816_),
    .Y(_00699_),
    .B1(_03817_));
 sg13g2_o21ai_1 _09595_ (.B1(_03565_),
    .Y(_03818_),
    .A1(_01783_),
    .A2(_02394_));
 sg13g2_o21ai_1 _09596_ (.B1(_02417_),
    .Y(_03819_),
    .A1(_01782_),
    .A2(_02398_));
 sg13g2_nand3_1 _09597_ (.B(_02402_),
    .C(_02407_),
    .A(_01812_),
    .Y(_03820_));
 sg13g2_nor3_2 _09598_ (.A(_03818_),
    .B(_03819_),
    .C(_03820_),
    .Y(_03821_));
 sg13g2_nor2_1 _09599_ (.A(net1248),
    .B(_03821_),
    .Y(_03822_));
 sg13g2_nor2_1 _09600_ (.A(net1198),
    .B(_01802_),
    .Y(_03823_));
 sg13g2_nand2_1 _09601_ (.Y(_03824_),
    .A(net1184),
    .B(_03560_));
 sg13g2_nor4_2 _09602_ (.A(net1135),
    .B(_03822_),
    .C(_03823_),
    .Y(_03825_),
    .D(_03824_));
 sg13g2_a21oi_1 _09603_ (.A1(_00796_),
    .A2(net1136),
    .Y(_00700_),
    .B1(_03825_));
 sg13g2_o21ai_1 _09604_ (.B1(_01779_),
    .Y(_03826_),
    .A1(_02408_),
    .A2(_03561_));
 sg13g2_nor4_1 _09605_ (.A(net1201),
    .B(_02405_),
    .C(_03557_),
    .D(_03824_),
    .Y(_03827_));
 sg13g2_and2_1 _09606_ (.A(_03826_),
    .B(_03827_),
    .X(_03828_));
 sg13g2_o21ai_1 _09607_ (.B1(_03828_),
    .Y(_03829_),
    .A1(net1249),
    .A2(_03821_));
 sg13g2_o21ai_1 _09608_ (.B1(_03829_),
    .Y(_03830_),
    .A1(net1198),
    .A2(_03723_));
 sg13g2_nand2_1 _09609_ (.Y(_03831_),
    .A(net2450),
    .B(net1136));
 sg13g2_o21ai_1 _09610_ (.B1(_03831_),
    .Y(_00701_),
    .A1(net1136),
    .A2(_03830_));
 sg13g2_nor2_1 _09611_ (.A(_01819_),
    .B(_03821_),
    .Y(_03832_));
 sg13g2_nor2_1 _09612_ (.A(_01752_),
    .B(_02404_),
    .Y(_03833_));
 sg13g2_o21ai_1 _09613_ (.B1(net1195),
    .Y(_03834_),
    .A1(_03832_),
    .A2(_03833_));
 sg13g2_a21oi_2 _09614_ (.B1(net1134),
    .Y(_03835_),
    .A2(_03834_),
    .A1(_03735_));
 sg13g2_a21o_1 _09615_ (.A2(net1136),
    .A1(net2509),
    .B1(_03835_),
    .X(_00702_));
 sg13g2_o21ai_1 _09616_ (.B1(net1197),
    .Y(_03836_),
    .A1(_01818_),
    .A2(_03818_));
 sg13g2_o21ai_1 _09617_ (.B1(_03738_),
    .Y(_03837_),
    .A1(_03821_),
    .A2(_03836_));
 sg13g2_mux2_1 _09618_ (.A0(net2550),
    .A1(_03837_),
    .S(net1143),
    .X(_00703_));
 sg13g2_xnor2_1 _09619_ (.Y(_03838_),
    .A(\i_core.cpu.i_core.i_registers.rs2[0] ),
    .B(\i_core.cpu.mem_op_increment_reg ));
 sg13g2_nand2_1 _09620_ (.Y(_03839_),
    .A(net1197),
    .B(_03545_));
 sg13g2_a21o_1 _09621_ (.A2(_03560_),
    .A1(_01793_),
    .B1(_03839_),
    .X(_03840_));
 sg13g2_nor2_1 _09622_ (.A(_01775_),
    .B(_03746_),
    .Y(_03841_));
 sg13g2_a22oi_1 _09623_ (.Y(_03842_),
    .B1(_03840_),
    .B2(_03841_),
    .A2(_03838_),
    .A1(net1186));
 sg13g2_mux2_1 _09624_ (.A0(net2606),
    .A1(_03842_),
    .S(_02391_),
    .X(_00704_));
 sg13g2_nor3_1 _09625_ (.A(_02426_),
    .B(_03544_),
    .C(_03559_),
    .Y(_03843_));
 sg13g2_o21ai_1 _09626_ (.B1(net1185),
    .Y(_03844_),
    .A1(_03749_),
    .A2(_03843_));
 sg13g2_a21oi_1 _09627_ (.A1(\i_core.cpu.i_core.i_registers.rs2[0] ),
    .A2(\i_core.cpu.mem_op_increment_reg ),
    .Y(_03845_),
    .B1(\i_core.cpu.i_core.i_registers.rs2[1] ));
 sg13g2_nand2_1 _09628_ (.Y(_03846_),
    .A(\i_core.cpu.mem_op_increment_reg ),
    .B(net1337));
 sg13g2_nand2b_1 _09629_ (.Y(_03847_),
    .B(_03846_),
    .A_N(_03845_));
 sg13g2_o21ai_1 _09630_ (.B1(_03844_),
    .Y(_03848_),
    .A1(net1185),
    .A2(_03847_));
 sg13g2_mux2_1 _09631_ (.A0(net2521),
    .A1(_03848_),
    .S(_02391_),
    .X(_00705_));
 sg13g2_nand3_1 _09632_ (.B(\i_core.cpu.mem_op_increment_reg ),
    .C(net1337),
    .A(\i_core.cpu.i_core.i_registers.rs2[2] ),
    .Y(_03849_));
 sg13g2_xor2_1 _09633_ (.B(_03846_),
    .A(\i_core.cpu.i_core.i_registers.rs2[2] ),
    .X(_03850_));
 sg13g2_nor3_1 _09634_ (.A(_01790_),
    .B(_03559_),
    .C(_03839_),
    .Y(_03851_));
 sg13g2_nor3_2 _09635_ (.A(net1187),
    .B(_03752_),
    .C(_03851_),
    .Y(_03852_));
 sg13g2_a21oi_1 _09636_ (.A1(net1186),
    .A2(_03850_),
    .Y(_03853_),
    .B1(_03852_));
 sg13g2_mux2_1 _09637_ (.A0(net2595),
    .A1(_03853_),
    .S(net1155),
    .X(_00706_));
 sg13g2_o21ai_1 _09638_ (.B1(net1256),
    .Y(_03854_),
    .A1(_01804_),
    .A2(_03558_));
 sg13g2_nor2b_1 _09639_ (.A(_03839_),
    .B_N(_03854_),
    .Y(_03855_));
 sg13g2_nor3_2 _09640_ (.A(net1187),
    .B(_03755_),
    .C(_03855_),
    .Y(_03856_));
 sg13g2_xor2_1 _09641_ (.B(_03849_),
    .A(\i_core.cpu.i_core.i_registers.rs2[3] ),
    .X(_03857_));
 sg13g2_a21oi_1 _09642_ (.A1(net1186),
    .A2(_03857_),
    .Y(_03858_),
    .B1(_03856_));
 sg13g2_mux2_1 _09643_ (.A0(net2585),
    .A1(_03858_),
    .S(net1155),
    .X(_00707_));
 sg13g2_nor2_1 _09644_ (.A(net1248),
    .B(net1184),
    .Y(_03859_));
 sg13g2_a221oi_1 _09645_ (.B2(net1200),
    .C1(_03859_),
    .B1(_03815_),
    .A1(net1252),
    .Y(_03860_),
    .A2(_03559_));
 sg13g2_a22oi_1 _09646_ (.Y(_03861_),
    .B1(_02390_),
    .B2(\i_core.cpu.additional_mem_ops[0] ),
    .A2(net1187),
    .A1(net2407));
 sg13g2_o21ai_1 _09647_ (.B1(net2408),
    .Y(_03862_),
    .A1(net1156),
    .A2(_03860_));
 sg13g2_and2_1 _09648_ (.A(net1460),
    .B(_03862_),
    .X(_00708_));
 sg13g2_o21ai_1 _09649_ (.B1(net1185),
    .Y(_03863_),
    .A1(net1249),
    .A2(net1184));
 sg13g2_a221oi_1 _09650_ (.B2(_03815_),
    .C1(_03863_),
    .B1(_03714_),
    .A1(net1251),
    .Y(_03864_),
    .A2(_03559_));
 sg13g2_nand2_1 _09651_ (.Y(_03865_),
    .A(net2320),
    .B(\i_core.cpu.additional_mem_ops[0] ));
 sg13g2_a21oi_1 _09652_ (.A1(_00748_),
    .A2(_00749_),
    .Y(_03866_),
    .B1(_01184_));
 sg13g2_a21oi_1 _09653_ (.A1(_03865_),
    .A2(_03866_),
    .Y(_03867_),
    .B1(_03864_));
 sg13g2_o21ai_1 _09654_ (.B1(net1459),
    .Y(_03868_),
    .A1(_02390_),
    .A2(_03867_));
 sg13g2_a21oi_1 _09655_ (.A1(_00748_),
    .A2(_02390_),
    .Y(_00709_),
    .B1(_03868_));
 sg13g2_nand2_1 _09656_ (.Y(_03869_),
    .A(_01791_),
    .B(_03559_));
 sg13g2_o21ai_1 _09657_ (.B1(_03869_),
    .Y(_03870_),
    .A1(_01819_),
    .A2(net1184));
 sg13g2_nand2_1 _09658_ (.Y(_03871_),
    .A(net1158),
    .B(_03870_));
 sg13g2_o21ai_1 _09659_ (.B1(net2200),
    .Y(_03872_),
    .A1(_02390_),
    .A2(_03866_));
 sg13g2_a21oi_1 _09660_ (.A1(_03871_),
    .A2(_03872_),
    .Y(_00710_),
    .B1(net1383));
 sg13g2_nor2_1 _09661_ (.A(net2460),
    .B(net1143),
    .Y(_03873_));
 sg13g2_and2_1 _09662_ (.A(net1200),
    .B(_03813_),
    .X(_03874_));
 sg13g2_a21oi_1 _09663_ (.A1(net1143),
    .A2(_03874_),
    .Y(_00711_),
    .B1(_03873_));
 sg13g2_a22oi_1 _09664_ (.Y(_03875_),
    .B1(_03498_),
    .B2(net2139),
    .A2(net1185),
    .A1(_01769_));
 sg13g2_nor2_1 _09665_ (.A(net1386),
    .B(_03875_),
    .Y(_00712_));
 sg13g2_o21ai_1 _09666_ (.B1(_03498_),
    .Y(_03876_),
    .A1(_01770_),
    .A2(net1187));
 sg13g2_nand2b_1 _09667_ (.Y(_03877_),
    .B(_01771_),
    .A_N(_01831_));
 sg13g2_o21ai_1 _09668_ (.B1(_03876_),
    .Y(_03878_),
    .A1(net1180),
    .A2(_03877_));
 sg13g2_o21ai_1 _09669_ (.B1(net1465),
    .Y(_03879_),
    .A1(net1392),
    .A2(_03876_));
 sg13g2_nor2b_1 _09670_ (.A(_03879_),
    .B_N(_03878_),
    .Y(_00713_));
 sg13g2_a22oi_1 _09671_ (.Y(_03880_),
    .B1(net1118),
    .B2(net1874),
    .A2(net1122),
    .A1(\addr[0] ));
 sg13g2_inv_1 _09672_ (.Y(_00714_),
    .A(net1875));
 sg13g2_nor3_1 _09673_ (.A(net1457),
    .B(_01844_),
    .C(_02579_),
    .Y(_00715_));
 sg13g2_xnor2_1 _09674_ (.Y(_03881_),
    .A(\i_core.cpu.instr_data_start[4] ),
    .B(_03234_));
 sg13g2_nor2_1 _09675_ (.A(net1422),
    .B(_03881_),
    .Y(_03882_));
 sg13g2_a21oi_2 _09676_ (.B1(_03882_),
    .Y(_03883_),
    .A2(_03253_),
    .A1(net1422));
 sg13g2_a22oi_1 _09677_ (.Y(_03884_),
    .B1(net1113),
    .B2(_03883_),
    .A2(net1262),
    .A1(net1874));
 sg13g2_a22oi_1 _09678_ (.Y(_03885_),
    .B1(net1117),
    .B2(net2035),
    .A2(net1121),
    .A1(\addr[4] ));
 sg13g2_nand2_1 _09679_ (.Y(_00716_),
    .A(_03884_),
    .B(net2036));
 sg13g2_nand2_1 _09680_ (.Y(_03886_),
    .A(net1929),
    .B(net1117));
 sg13g2_nor3_2 _09681_ (.A(_00765_),
    .B(_00163_),
    .C(_03234_),
    .Y(_03887_));
 sg13g2_o21ai_1 _09682_ (.B1(_00765_),
    .Y(_03888_),
    .A1(_00163_),
    .A2(_03234_));
 sg13g2_nand2_1 _09683_ (.Y(_03889_),
    .A(net1388),
    .B(_03888_));
 sg13g2_o21ai_1 _09684_ (.B1(_03221_),
    .Y(_03890_),
    .A1(_03887_),
    .A2(_03889_));
 sg13g2_a21oi_1 _09685_ (.A1(net1420),
    .A2(_03262_),
    .Y(_03891_),
    .B1(_03890_));
 sg13g2_a21o_1 _09686_ (.A2(net1261),
    .A1(\i_core.mem.q_ctrl.addr[1] ),
    .B1(net1125),
    .X(_03892_));
 sg13g2_o21ai_1 _09687_ (.B1(_03892_),
    .Y(_03893_),
    .A1(\addr[5] ),
    .A2(_03219_));
 sg13g2_o21ai_1 _09688_ (.B1(_03886_),
    .Y(_00717_),
    .A1(_03891_),
    .A2(_03893_));
 sg13g2_a21oi_1 _09689_ (.A1(\i_core.mem.q_ctrl.addr[2] ),
    .A2(net1261),
    .Y(_03894_),
    .B1(net1125));
 sg13g2_and2_1 _09690_ (.A(\i_core.cpu.instr_data_start[6] ),
    .B(_03887_),
    .X(_03895_));
 sg13g2_o21ai_1 _09691_ (.B1(net1388),
    .Y(_03896_),
    .A1(\i_core.cpu.instr_data_start[6] ),
    .A2(_03887_));
 sg13g2_nor2_1 _09692_ (.A(_03895_),
    .B(_03896_),
    .Y(_03897_));
 sg13g2_a21oi_2 _09693_ (.B1(_03897_),
    .Y(_03898_),
    .A2(_03270_),
    .A1(net1420));
 sg13g2_a221oi_1 _09694_ (.B2(_03898_),
    .C1(_03894_),
    .B1(net1113),
    .A1(_00817_),
    .Y(_03899_),
    .A2(net1121));
 sg13g2_a21o_1 _09695_ (.A2(net1117),
    .A1(net2061),
    .B1(_03899_),
    .X(_00718_));
 sg13g2_xor2_1 _09696_ (.B(_03895_),
    .A(\i_core.cpu.instr_data_start[7] ),
    .X(_03900_));
 sg13g2_nand2_1 _09697_ (.Y(_03901_),
    .A(net1420),
    .B(_03278_));
 sg13g2_o21ai_1 _09698_ (.B1(_03901_),
    .Y(_03902_),
    .A1(net1420),
    .A2(_03900_));
 sg13g2_nand2b_1 _09699_ (.Y(_03903_),
    .B(net1117),
    .A_N(\i_core.mem.q_ctrl.addr[7] ));
 sg13g2_o21ai_1 _09700_ (.B1(_03903_),
    .Y(_03904_),
    .A1(\addr[7] ),
    .A2(_03219_));
 sg13g2_a221oi_1 _09701_ (.B2(_03902_),
    .C1(_03904_),
    .B1(net1113),
    .A1(_00852_),
    .Y(_00719_),
    .A2(net1263));
 sg13g2_nand3_1 _09702_ (.B(net1427),
    .C(_03895_),
    .A(\i_core.cpu.instr_data_start[8] ),
    .Y(_03905_));
 sg13g2_a21o_1 _09703_ (.A2(_03895_),
    .A1(net1427),
    .B1(\i_core.cpu.instr_data_start[8] ),
    .X(_03906_));
 sg13g2_nand3_1 _09704_ (.B(_03905_),
    .C(_03906_),
    .A(net1388),
    .Y(_03907_));
 sg13g2_o21ai_1 _09705_ (.B1(_03907_),
    .Y(_03908_),
    .A1(net1388),
    .A2(_03289_));
 sg13g2_a22oi_1 _09706_ (.Y(_03909_),
    .B1(net1113),
    .B2(_03908_),
    .A2(net1262),
    .A1(net2035));
 sg13g2_a22oi_1 _09707_ (.Y(_03910_),
    .B1(net1117),
    .B2(net2141),
    .A2(net1122),
    .A1(\addr[8] ));
 sg13g2_nand2_1 _09708_ (.Y(_00720_),
    .A(_03909_),
    .B(net2142));
 sg13g2_or2_1 _09709_ (.X(_03911_),
    .B(_03905_),
    .A(_00763_));
 sg13g2_a21oi_1 _09710_ (.A1(_00763_),
    .A2(_03905_),
    .Y(_03912_),
    .B1(net1421));
 sg13g2_nor2_1 _09711_ (.A(net1389),
    .B(_03297_),
    .Y(_03913_));
 sg13g2_a21o_1 _09712_ (.A2(_03912_),
    .A1(_03911_),
    .B1(_03913_),
    .X(_03914_));
 sg13g2_a22oi_1 _09713_ (.Y(_03915_),
    .B1(net1114),
    .B2(_03914_),
    .A2(net1261),
    .A1(net1929));
 sg13g2_a22oi_1 _09714_ (.Y(_03916_),
    .B1(net1119),
    .B2(net2082),
    .A2(net1121),
    .A1(\addr[9] ));
 sg13g2_nand2_1 _09715_ (.Y(_00721_),
    .A(_03915_),
    .B(net2083));
 sg13g2_nor2_1 _09716_ (.A(_00762_),
    .B(_03911_),
    .Y(_03917_));
 sg13g2_xnor2_1 _09717_ (.Y(_03918_),
    .A(\i_core.cpu.instr_data_start[10] ),
    .B(_03911_));
 sg13g2_nand2_1 _09718_ (.Y(_03919_),
    .A(net1388),
    .B(_03918_));
 sg13g2_o21ai_1 _09719_ (.B1(_03919_),
    .Y(_03920_),
    .A1(net1388),
    .A2(_03305_));
 sg13g2_a22oi_1 _09720_ (.Y(_03921_),
    .B1(net1114),
    .B2(_03920_),
    .A2(net1262),
    .A1(net2061));
 sg13g2_a22oi_1 _09721_ (.Y(_03922_),
    .B1(net1117),
    .B2(net2106),
    .A2(net1121),
    .A1(\addr[10] ));
 sg13g2_nand2_1 _09722_ (.Y(_00722_),
    .A(_03921_),
    .B(net2107));
 sg13g2_xnor2_1 _09723_ (.Y(_03923_),
    .A(_00201_),
    .B(_03917_));
 sg13g2_nor2_1 _09724_ (.A(net1420),
    .B(_03923_),
    .Y(_03924_));
 sg13g2_a21oi_1 _09725_ (.A1(net1420),
    .A2(_03315_),
    .Y(_03925_),
    .B1(_03924_));
 sg13g2_a22oi_1 _09726_ (.Y(_03926_),
    .B1(net1113),
    .B2(_03925_),
    .A2(net1262),
    .A1(\i_core.mem.q_ctrl.addr[7] ));
 sg13g2_a22oi_1 _09727_ (.Y(_03927_),
    .B1(net1118),
    .B2(net2161),
    .A2(net1121),
    .A1(\addr[11] ));
 sg13g2_nand2_1 _09728_ (.Y(_00723_),
    .A(_03926_),
    .B(net2162));
 sg13g2_and3_1 _09729_ (.X(_03928_),
    .A(\i_core.cpu.instr_data_start[12] ),
    .B(\i_core.cpu.instr_data_start[11] ),
    .C(_03917_));
 sg13g2_a21oi_1 _09730_ (.A1(\i_core.cpu.instr_data_start[11] ),
    .A2(_03917_),
    .Y(_03929_),
    .B1(\i_core.cpu.instr_data_start[12] ));
 sg13g2_nor3_1 _09731_ (.A(net1420),
    .B(_03928_),
    .C(_03929_),
    .Y(_03930_));
 sg13g2_a21o_1 _09732_ (.A2(_03324_),
    .A1(net1420),
    .B1(_03930_),
    .X(_03931_));
 sg13g2_a22oi_1 _09733_ (.Y(_03932_),
    .B1(net1114),
    .B2(_03931_),
    .A2(net1261),
    .A1(net2141));
 sg13g2_a22oi_1 _09734_ (.Y(_03933_),
    .B1(net1117),
    .B2(net2240),
    .A2(net1121),
    .A1(\addr[12] ));
 sg13g2_nand2_1 _09735_ (.Y(_00724_),
    .A(_03932_),
    .B(net2241));
 sg13g2_o21ai_1 _09736_ (.B1(net1388),
    .Y(_03934_),
    .A1(\i_core.cpu.instr_data_start[13] ),
    .A2(_03928_));
 sg13g2_a21o_1 _09737_ (.A2(_03928_),
    .A1(\i_core.cpu.instr_data_start[13] ),
    .B1(_03934_),
    .X(_03935_));
 sg13g2_o21ai_1 _09738_ (.B1(_03935_),
    .Y(_03936_),
    .A1(net1388),
    .A2(_03333_));
 sg13g2_a22oi_1 _09739_ (.Y(_03937_),
    .B1(net1113),
    .B2(_03936_),
    .A2(net1261),
    .A1(\i_core.mem.q_ctrl.addr[9] ));
 sg13g2_a22oi_1 _09740_ (.Y(_03938_),
    .B1(net1118),
    .B2(net2068),
    .A2(net1122),
    .A1(\addr[13] ));
 sg13g2_nand2_1 _09741_ (.Y(_00725_),
    .A(_03937_),
    .B(net2069));
 sg13g2_and3_1 _09742_ (.X(_03939_),
    .A(net1426),
    .B(\i_core.cpu.instr_data_start[13] ),
    .C(_03928_));
 sg13g2_a21oi_1 _09743_ (.A1(\i_core.cpu.instr_data_start[13] ),
    .A2(_03928_),
    .Y(_03940_),
    .B1(net1426));
 sg13g2_nor3_1 _09744_ (.A(net1421),
    .B(_03939_),
    .C(_03940_),
    .Y(_03941_));
 sg13g2_a21o_1 _09745_ (.A2(_03340_),
    .A1(net1421),
    .B1(_03941_),
    .X(_03942_));
 sg13g2_a22oi_1 _09746_ (.Y(_03943_),
    .B1(net1113),
    .B2(_03942_),
    .A2(net1261),
    .A1(net2106));
 sg13g2_a22oi_1 _09747_ (.Y(_03944_),
    .B1(net1118),
    .B2(net2119),
    .A2(net1121),
    .A1(\addr[14] ));
 sg13g2_nand2_1 _09748_ (.Y(_00726_),
    .A(_03943_),
    .B(net2120));
 sg13g2_xor2_1 _09749_ (.B(_03939_),
    .A(net1425),
    .X(_03945_));
 sg13g2_nor2_1 _09750_ (.A(net1421),
    .B(_03945_),
    .Y(_03946_));
 sg13g2_a21oi_2 _09751_ (.B1(_03946_),
    .Y(_03947_),
    .A2(_03351_),
    .A1(net1421));
 sg13g2_a22oi_1 _09752_ (.Y(_03948_),
    .B1(_03947_),
    .B2(net1125),
    .A2(net1261),
    .A1(\i_core.mem.q_ctrl.addr[11] ));
 sg13g2_a22oi_1 _09753_ (.Y(_03949_),
    .B1(net1118),
    .B2(net2114),
    .A2(net1120),
    .A1(\addr[15] ));
 sg13g2_o21ai_1 _09754_ (.B1(net2115),
    .Y(_00727_),
    .A1(net1120),
    .A2(_03948_));
 sg13g2_a22oi_1 _09755_ (.Y(_03950_),
    .B1(net1120),
    .B2(\addr[16] ),
    .A2(net1261),
    .A1(\i_core.mem.q_ctrl.addr[12] ));
 sg13g2_and3_1 _09756_ (.X(_03951_),
    .A(net1424),
    .B(net1425),
    .C(_03939_));
 sg13g2_a21oi_1 _09757_ (.A1(net1425),
    .A2(_03939_),
    .Y(_03952_),
    .B1(net1424));
 sg13g2_nor3_1 _09758_ (.A(net1418),
    .B(_03951_),
    .C(_03952_),
    .Y(_03953_));
 sg13g2_a21o_1 _09759_ (.A2(_03360_),
    .A1(net1418),
    .B1(_03953_),
    .X(_03954_));
 sg13g2_a22oi_1 _09760_ (.Y(_03955_),
    .B1(net1114),
    .B2(_03954_),
    .A2(net1115),
    .A1(net2170));
 sg13g2_nand2_1 _09761_ (.Y(_00728_),
    .A(_03950_),
    .B(_03955_));
 sg13g2_a22oi_1 _09762_ (.Y(_03956_),
    .B1(net1116),
    .B2(net2071),
    .A2(net1263),
    .A1(net2068));
 sg13g2_and2_1 _09763_ (.A(\i_core.cpu.instr_data_start[17] ),
    .B(_03951_),
    .X(_03957_));
 sg13g2_o21ai_1 _09764_ (.B1(net1389),
    .Y(_03958_),
    .A1(\i_core.cpu.instr_data_start[17] ),
    .A2(_03951_));
 sg13g2_nand2_1 _09765_ (.Y(_03959_),
    .A(net1418),
    .B(_03369_));
 sg13g2_o21ai_1 _09766_ (.B1(_03959_),
    .Y(_03960_),
    .A1(_03957_),
    .A2(_03958_));
 sg13g2_a22oi_1 _09767_ (.Y(_03961_),
    .B1(net1114),
    .B2(_03960_),
    .A2(net1120),
    .A1(\addr[17] ));
 sg13g2_nand2_1 _09768_ (.Y(_00729_),
    .A(_03956_),
    .B(_03961_));
 sg13g2_or2_1 _09769_ (.X(_03962_),
    .B(_03957_),
    .A(\i_core.cpu.instr_data_start[18] ));
 sg13g2_nand2_1 _09770_ (.Y(_03963_),
    .A(\i_core.cpu.instr_data_start[18] ),
    .B(_03957_));
 sg13g2_a21oi_1 _09771_ (.A1(_03962_),
    .A2(_03963_),
    .Y(_03964_),
    .B1(net1417));
 sg13g2_a21oi_2 _09772_ (.B1(_03964_),
    .Y(_03965_),
    .A2(_03377_),
    .A1(net1418));
 sg13g2_a22oi_1 _09773_ (.Y(_03966_),
    .B1(net1116),
    .B2(net2182),
    .A2(net1120),
    .A1(net2140));
 sg13g2_a22oi_1 _09774_ (.Y(_03967_),
    .B1(net1114),
    .B2(_03965_),
    .A2(net1263),
    .A1(net2119));
 sg13g2_nand2_1 _09775_ (.Y(_00730_),
    .A(_03966_),
    .B(_03967_));
 sg13g2_and3_1 _09776_ (.X(_03968_),
    .A(\i_core.cpu.instr_data_start[19] ),
    .B(\i_core.cpu.instr_data_start[18] ),
    .C(_03957_));
 sg13g2_xnor2_1 _09777_ (.Y(_03969_),
    .A(\i_core.cpu.instr_data_start[19] ),
    .B(_03963_));
 sg13g2_o21ai_1 _09778_ (.B1(_03221_),
    .Y(_03970_),
    .A1(net1417),
    .A2(_03969_));
 sg13g2_a21oi_1 _09779_ (.A1(net1418),
    .A2(_03386_),
    .Y(_03971_),
    .B1(_03970_));
 sg13g2_a221oi_1 _09780_ (.B2(\addr[19] ),
    .C1(_03971_),
    .B1(net1120),
    .A1(\i_core.mem.q_ctrl.addr[15] ),
    .Y(_03972_),
    .A2(_02943_));
 sg13g2_nand2_1 _09781_ (.Y(_03973_),
    .A(net1976),
    .B(net1115));
 sg13g2_o21ai_1 _09782_ (.B1(_03973_),
    .Y(_00731_),
    .A1(net1115),
    .A2(_03972_));
 sg13g2_nor2_1 _09783_ (.A(_00165_),
    .B(_03963_),
    .Y(_03974_));
 sg13g2_xnor2_1 _09784_ (.Y(_03975_),
    .A(_00757_),
    .B(_03974_));
 sg13g2_nand2_1 _09785_ (.Y(_03976_),
    .A(net1418),
    .B(_03395_));
 sg13g2_o21ai_1 _09786_ (.B1(_03976_),
    .Y(_03977_),
    .A1(net1417),
    .A2(_03975_));
 sg13g2_nand2b_1 _09787_ (.Y(_03978_),
    .B(net1263),
    .A_N(net2170));
 sg13g2_o21ai_1 _09788_ (.B1(_03978_),
    .Y(_03979_),
    .A1(net2172),
    .A2(_03219_));
 sg13g2_a221oi_1 _09789_ (.B2(_03977_),
    .C1(_03979_),
    .B1(net1114),
    .A1(_00846_),
    .Y(_00732_),
    .A2(net1116));
 sg13g2_and3_1 _09790_ (.X(_03980_),
    .A(\i_core.cpu.instr_data_start[21] ),
    .B(net1423),
    .C(_03968_));
 sg13g2_a21oi_1 _09791_ (.A1(net1423),
    .A2(_03968_),
    .Y(_03981_),
    .B1(\i_core.cpu.instr_data_start[21] ));
 sg13g2_o21ai_1 _09792_ (.B1(net1389),
    .Y(_03982_),
    .A1(_03980_),
    .A2(_03981_));
 sg13g2_o21ai_1 _09793_ (.B1(_03982_),
    .Y(_03983_),
    .A1(net1389),
    .A2(_03405_));
 sg13g2_a22oi_1 _09794_ (.Y(_03984_),
    .B1(net1120),
    .B2(net2205),
    .A2(_02943_),
    .A1(net2071));
 sg13g2_nor2_1 _09795_ (.A(net1116),
    .B(_03984_),
    .Y(_03985_));
 sg13g2_a21oi_1 _09796_ (.A1(net2368),
    .A2(net1115),
    .Y(_03986_),
    .B1(_03985_));
 sg13g2_o21ai_1 _09797_ (.B1(_03986_),
    .Y(_00733_),
    .A1(_03222_),
    .A2(_03983_));
 sg13g2_nand2_1 _09798_ (.Y(_03987_),
    .A(\i_core.cpu.instr_data_start[22] ),
    .B(_03980_));
 sg13g2_nor2_1 _09799_ (.A(\i_core.cpu.instr_data_start[22] ),
    .B(_03980_),
    .Y(_03988_));
 sg13g2_nor2_1 _09800_ (.A(net1417),
    .B(_03988_),
    .Y(_03989_));
 sg13g2_a221oi_1 _09801_ (.B2(_03989_),
    .C1(_02934_),
    .B1(_03987_),
    .A1(net1417),
    .Y(_03990_),
    .A2(_03416_));
 sg13g2_o21ai_1 _09802_ (.B1(net1125),
    .Y(_03991_),
    .A1(net2198),
    .A2(_02935_));
 sg13g2_or2_1 _09803_ (.X(_03992_),
    .B(_03991_),
    .A(_03990_));
 sg13g2_a21oi_1 _09804_ (.A1(net2182),
    .A2(_02943_),
    .Y(_03993_),
    .B1(net1115));
 sg13g2_a22oi_1 _09805_ (.Y(_00734_),
    .B1(_03992_),
    .B2(_03993_),
    .A2(net1115),
    .A1(_00847_));
 sg13g2_xnor2_1 _09806_ (.Y(_03994_),
    .A(_00162_),
    .B(_03987_));
 sg13g2_a21oi_1 _09807_ (.A1(net1417),
    .A2(_03424_),
    .Y(_03995_),
    .B1(_02934_));
 sg13g2_o21ai_1 _09808_ (.B1(_03995_),
    .Y(_03996_),
    .A1(net1417),
    .A2(_03994_));
 sg13g2_a21oi_1 _09809_ (.A1(_00161_),
    .A2(_02934_),
    .Y(_03997_),
    .B1(_02943_));
 sg13g2_a221oi_1 _09810_ (.B2(_03997_),
    .C1(net1115),
    .B1(_03996_),
    .A1(net1976),
    .Y(_03998_),
    .A2(_02943_));
 sg13g2_a21oi_1 _09811_ (.A1(_00849_),
    .A2(net1115),
    .Y(_00735_),
    .B1(_03998_));
 sg13g2_nor3_1 _09812_ (.A(\i_core.cpu.i_core.i_cycles.cy ),
    .B(net2523),
    .C(net1278),
    .Y(_03999_));
 sg13g2_nand2_1 _09813_ (.Y(_04000_),
    .A(net1459),
    .B(_02343_));
 sg13g2_nor2_1 _09814_ (.A(net2524),
    .B(_04000_),
    .Y(_00736_));
 sg13g2_a21oi_1 _09815_ (.A1(_00823_),
    .A2(_02343_),
    .Y(_04001_),
    .B1(net1384));
 sg13g2_nor2b_1 _09816_ (.A(_02344_),
    .B_N(_04001_),
    .Y(_00737_));
 sg13g2_o21ai_1 _09817_ (.B1(net1459),
    .Y(_04002_),
    .A1(net2487),
    .A2(_02344_));
 sg13g2_nor2_1 _09818_ (.A(_02345_),
    .B(net2488),
    .Y(_00738_));
 sg13g2_o21ai_1 _09819_ (.B1(net1459),
    .Y(_04003_),
    .A1(net2413),
    .A2(_02345_));
 sg13g2_nor2b_1 _09820_ (.A(_04003_),
    .B_N(_02346_),
    .Y(_00739_));
 sg13g2_mux2_2 _09821_ (.A0(_00216_),
    .A1(net2213),
    .S(net1311),
    .X(_04004_));
 sg13g2_nor2_1 _09822_ (.A(_00824_),
    .B(_04004_),
    .Y(_04005_));
 sg13g2_nor3_1 _09823_ (.A(_00824_),
    .B(_00199_),
    .C(net2214),
    .Y(_04006_));
 sg13g2_nand2_1 _09824_ (.Y(_04007_),
    .A(net2571),
    .B(_04006_));
 sg13g2_nor3_1 _09825_ (.A(net1383),
    .B(_00836_),
    .C(_04007_),
    .Y(_00740_));
 sg13g2_nand3_1 _09826_ (.B(net1362),
    .C(_02067_),
    .A(net1382),
    .Y(_04008_));
 sg13g2_mux2_1 _09827_ (.A0(_02875_),
    .A1(net2478),
    .S(_04008_),
    .X(_00741_));
 sg13g2_nor2_1 _09828_ (.A(net1383),
    .B(net2414),
    .Y(_00742_));
 sg13g2_o21ai_1 _09829_ (.B1(net1459),
    .Y(_04009_),
    .A1(_00164_),
    .A2(net2214));
 sg13g2_a21oi_2 _09830_ (.B1(_04009_),
    .Y(_00743_),
    .A2(net2214),
    .A1(_00164_));
 sg13g2_o21ai_1 _09831_ (.B1(net1459),
    .Y(_04010_),
    .A1(net1830),
    .A2(_04005_));
 sg13g2_a21oi_1 _09832_ (.A1(net1830),
    .A2(_04005_),
    .Y(_00744_),
    .B1(_04010_));
 sg13g2_o21ai_1 _09833_ (.B1(net1459),
    .Y(_04011_),
    .A1(net2571),
    .A2(_04006_));
 sg13g2_nor2b_1 _09834_ (.A(net2572),
    .B_N(_04007_),
    .Y(_00745_));
 sg13g2_xnor2_1 _09835_ (.Y(_04012_),
    .A(_00836_),
    .B(_04007_));
 sg13g2_nor2_1 _09836_ (.A(net1383),
    .B(_04012_),
    .Y(_00746_));
 sg13g2_dfrbp_1 _09837_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net1037),
    .D(net1657),
    .Q_N(_04405_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[15][0] ));
 sg13g2_dfrbp_1 _09838_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net1038),
    .D(net1644),
    .Q_N(_00094_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[15][1] ));
 sg13g2_dfrbp_1 _09839_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net1039),
    .D(net1697),
    .Q_N(_00093_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[15][2] ));
 sg13g2_dfrbp_1 _09840_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net1040),
    .D(net1084),
    .Q_N(_00091_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[15][3] ));
 sg13g2_dfrbp_1 _09841_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net1041),
    .D(net1716),
    .Q_N(_04406_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _09842_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net1042),
    .D(net1472),
    .Q_N(_04407_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _09843_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net1043),
    .D(net1068),
    .Q_N(_04408_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _09844_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net1044),
    .D(net1589),
    .Q_N(_04409_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _09845_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net1045),
    .D(net1714),
    .Q_N(_04410_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _09846_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net1046),
    .D(net1731),
    .Q_N(_04411_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _09847_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net1047),
    .D(net1584),
    .Q_N(_04412_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _09848_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net1048),
    .D(net1727),
    .Q_N(_04413_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _09849_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net13),
    .D(net1561),
    .Q_N(_04414_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _09850_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net14),
    .D(net1571),
    .Q_N(_04415_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _09851_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net15),
    .D(net1732),
    .Q_N(_04416_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _09852_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net16),
    .D(net1070),
    .Q_N(_04417_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _09853_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net17),
    .D(net1640),
    .Q_N(_04418_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _09854_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net18),
    .D(net1069),
    .Q_N(_04419_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _09855_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net19),
    .D(net1515),
    .Q_N(_04420_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _09856_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net20),
    .D(net1588),
    .Q_N(_04421_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _09857_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net21),
    .D(net1680),
    .Q_N(_04422_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _09858_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net22),
    .D(net1583),
    .Q_N(_04423_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _09859_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net23),
    .D(net1610),
    .Q_N(_04424_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _09860_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net24),
    .D(net1499),
    .Q_N(_04425_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _09861_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net25),
    .D(net1702),
    .Q_N(_04426_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _09862_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net26),
    .D(net1652),
    .Q_N(_04427_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _09863_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net27),
    .D(net1676),
    .Q_N(_04428_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _09864_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net28),
    .D(net1658),
    .Q_N(_04429_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _09865_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net29),
    .D(_00050_),
    .Q_N(_04430_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _09866_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net30),
    .D(_00051_),
    .Q_N(_04431_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _09867_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net31),
    .D(_00052_),
    .Q_N(_04432_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _09868_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net32),
    .D(_00053_),
    .Q_N(_04433_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _09869_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net33),
    .D(net1772),
    .Q_N(_04434_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[14][0] ));
 sg13g2_dfrbp_1 _09870_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net34),
    .D(net1711),
    .Q_N(_04435_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[14][1] ));
 sg13g2_dfrbp_1 _09871_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net35),
    .D(net1701),
    .Q_N(_04436_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[14][2] ));
 sg13g2_dfrbp_1 _09872_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net36),
    .D(net1799),
    .Q_N(_04437_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[14][3] ));
 sg13g2_dfrbp_1 _09873_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net37),
    .D(net1067),
    .Q_N(_04438_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _09874_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net38),
    .D(net1756),
    .Q_N(_04439_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _09875_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net39),
    .D(net1101),
    .Q_N(_04440_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _09876_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net40),
    .D(net1077),
    .Q_N(_04441_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _09877_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net41),
    .D(net1484),
    .Q_N(_04442_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _09878_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net42),
    .D(net1591),
    .Q_N(_04443_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _09879_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net43),
    .D(net1628),
    .Q_N(_04444_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _09880_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net44),
    .D(net1604),
    .Q_N(_04445_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _09881_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net45),
    .D(net1485),
    .Q_N(_04446_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _09882_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net46),
    .D(net1627),
    .Q_N(_04447_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _09883_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net47),
    .D(net1679),
    .Q_N(_04448_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _09884_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net48),
    .D(net1546),
    .Q_N(_04449_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _09885_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net49),
    .D(net1488),
    .Q_N(_04450_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _09886_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net50),
    .D(net1504),
    .Q_N(_04451_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _09887_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net51),
    .D(net1771),
    .Q_N(_04452_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _09888_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net52),
    .D(net1550),
    .Q_N(_04453_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _09889_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net53),
    .D(net1757),
    .Q_N(_04454_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _09890_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net54),
    .D(net1719),
    .Q_N(_04455_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _09891_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net55),
    .D(net1107),
    .Q_N(_04456_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _09892_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net56),
    .D(net1603),
    .Q_N(_04457_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _09893_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net57),
    .D(net1763),
    .Q_N(_04458_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _09894_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net58),
    .D(net1104),
    .Q_N(_04459_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _09895_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net59),
    .D(net1598),
    .Q_N(_04460_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _09896_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net60),
    .D(net1807),
    .Q_N(_04461_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _09897_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net61),
    .D(_00046_),
    .Q_N(_04462_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _09898_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net62),
    .D(_00047_),
    .Q_N(_04463_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _09899_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net63),
    .D(_00048_),
    .Q_N(_04464_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _09900_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net64),
    .D(_00049_),
    .Q_N(_04465_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _09901_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net65),
    .D(net1803),
    .Q_N(_04466_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[13][0] ));
 sg13g2_dfrbp_1 _09902_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net66),
    .D(net1802),
    .Q_N(_04467_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[13][1] ));
 sg13g2_dfrbp_1 _09903_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net67),
    .D(net1705),
    .Q_N(_04468_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[13][2] ));
 sg13g2_dfrbp_1 _09904_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net68),
    .D(net1097),
    .Q_N(_04469_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[13][3] ));
 sg13g2_dfrbp_1 _09905_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net69),
    .D(net1693),
    .Q_N(_04470_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _09906_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net70),
    .D(net1681),
    .Q_N(_04471_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _09907_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net71),
    .D(net1663),
    .Q_N(_04472_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _09908_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net72),
    .D(net1491),
    .Q_N(_04473_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _09909_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net73),
    .D(net1768),
    .Q_N(_04474_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _09910_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net74),
    .D(net1526),
    .Q_N(_04475_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _09911_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net75),
    .D(net1083),
    .Q_N(_04476_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _09912_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net76),
    .D(net1473),
    .Q_N(_04477_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _09913_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net77),
    .D(net1088),
    .Q_N(_04478_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _09914_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net78),
    .D(net1527),
    .Q_N(_04479_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _09915_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net79),
    .D(net1492),
    .Q_N(_04480_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _09916_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net80),
    .D(net1494),
    .Q_N(_04481_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _09917_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net81),
    .D(net1624),
    .Q_N(_04482_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _09918_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net82),
    .D(net1552),
    .Q_N(_04483_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _09919_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net83),
    .D(net1493),
    .Q_N(_04484_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _09920_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net84),
    .D(net1513),
    .Q_N(_04485_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _09921_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net85),
    .D(net1551),
    .Q_N(_04486_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _09922_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net86),
    .D(net1778),
    .Q_N(_04487_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _09923_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net87),
    .D(net1708),
    .Q_N(_04488_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _09924_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net88),
    .D(net1808),
    .Q_N(_04489_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _09925_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net89),
    .D(net1059),
    .Q_N(_04490_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _09926_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net90),
    .D(net1102),
    .Q_N(_04491_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _09927_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net91),
    .D(net1078),
    .Q_N(_04492_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _09928_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net92),
    .D(net1575),
    .Q_N(_04493_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _09929_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net93),
    .D(_00042_),
    .Q_N(_04494_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _09930_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net94),
    .D(_00043_),
    .Q_N(_04495_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _09931_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net95),
    .D(_00044_),
    .Q_N(_04496_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _09932_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net96),
    .D(_00045_),
    .Q_N(_04497_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _09933_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net97),
    .D(net1675),
    .Q_N(_04498_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[12][0] ));
 sg13g2_dfrbp_1 _09934_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net98),
    .D(net1684),
    .Q_N(_04499_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[12][1] ));
 sg13g2_dfrbp_1 _09935_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net99),
    .D(net1668),
    .Q_N(_04500_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[12][2] ));
 sg13g2_dfrbp_1 _09936_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net100),
    .D(net1747),
    .Q_N(_04501_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[12][3] ));
 sg13g2_dfrbp_1 _09937_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net101),
    .D(net1721),
    .Q_N(_04502_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _09938_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net102),
    .D(net1788),
    .Q_N(_04503_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _09939_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net103),
    .D(net1801),
    .Q_N(_04504_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _09940_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net104),
    .D(net1670),
    .Q_N(_04505_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _09941_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net105),
    .D(net1786),
    .Q_N(_04506_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _09942_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net106),
    .D(net1547),
    .Q_N(_04507_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _09943_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net107),
    .D(net1572),
    .Q_N(_04508_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _09944_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net108),
    .D(net1081),
    .Q_N(_04509_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _09945_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net109),
    .D(net1545),
    .Q_N(_04510_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _09946_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net110),
    .D(net1717),
    .Q_N(_04511_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _09947_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net111),
    .D(net1065),
    .Q_N(_04512_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _09948_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net112),
    .D(net1592),
    .Q_N(_04513_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _09949_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net113),
    .D(net1718),
    .Q_N(_04514_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _09950_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net114),
    .D(net1082),
    .Q_N(_04515_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _09951_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net115),
    .D(net1556),
    .Q_N(_04516_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _09952_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net116),
    .D(net1619),
    .Q_N(_04517_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _09953_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net117),
    .D(net1564),
    .Q_N(_04518_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _09954_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net118),
    .D(net1689),
    .Q_N(_04519_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _09955_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net119),
    .D(net1742),
    .Q_N(_04520_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _09956_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net120),
    .D(net1483),
    .Q_N(_04521_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _09957_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net121),
    .D(net1631),
    .Q_N(_04522_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _09958_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net122),
    .D(net1098),
    .Q_N(_04523_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _09959_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net123),
    .D(net1567),
    .Q_N(_04524_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _09960_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net124),
    .D(net1800),
    .Q_N(_04525_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _09961_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net125),
    .D(_00038_),
    .Q_N(_04526_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _09962_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net126),
    .D(_00039_),
    .Q_N(_04527_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _09963_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net127),
    .D(_00040_),
    .Q_N(_04528_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _09964_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net128),
    .D(_00041_),
    .Q_N(_04529_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _09965_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net129),
    .D(net1822),
    .Q_N(_04530_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[11][0] ));
 sg13g2_dfrbp_1 _09966_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net130),
    .D(net1815),
    .Q_N(_04531_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[11][1] ));
 sg13g2_dfrbp_1 _09967_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net131),
    .D(net1798),
    .Q_N(_04532_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[11][2] ));
 sg13g2_dfrbp_1 _09968_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net132),
    .D(net1767),
    .Q_N(_04533_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[11][3] ));
 sg13g2_dfrbp_1 _09969_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net133),
    .D(net1608),
    .Q_N(_04534_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _09970_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net134),
    .D(net1690),
    .Q_N(_04535_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _09971_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net135),
    .D(net1506),
    .Q_N(_04536_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _09972_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net136),
    .D(net1478),
    .Q_N(_04537_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _09973_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net137),
    .D(net1540),
    .Q_N(_04538_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _09974_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net138),
    .D(net1064),
    .Q_N(_04539_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _09975_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net139),
    .D(net1060),
    .Q_N(_04540_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _09976_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net140),
    .D(net1653),
    .Q_N(_04541_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _09977_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net141),
    .D(net1538),
    .Q_N(_04542_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _09978_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net142),
    .D(net1489),
    .Q_N(_04543_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _09979_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net143),
    .D(net1576),
    .Q_N(_04544_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _09980_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net144),
    .D(net1751),
    .Q_N(_04545_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _09981_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net145),
    .D(net1051),
    .Q_N(_04546_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _09982_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net146),
    .D(net1713),
    .Q_N(_04547_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _09983_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net147),
    .D(net1475),
    .Q_N(_04548_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _09984_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net148),
    .D(net1662),
    .Q_N(_04549_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _09985_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net149),
    .D(net1497),
    .Q_N(_04550_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _09986_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net150),
    .D(net1637),
    .Q_N(_04551_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _09987_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net151),
    .D(net1646),
    .Q_N(_04552_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _09988_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net152),
    .D(net1094),
    .Q_N(_04553_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _09989_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net153),
    .D(net1476),
    .Q_N(_04554_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _09990_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net154),
    .D(net1055),
    .Q_N(_04555_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _09991_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net155),
    .D(net1741),
    .Q_N(_04556_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _09992_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net156),
    .D(net1748),
    .Q_N(_04557_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _09993_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net157),
    .D(_00034_),
    .Q_N(_04558_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _09994_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net158),
    .D(_00035_),
    .Q_N(_04559_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _09995_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net159),
    .D(_00036_),
    .Q_N(_04560_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _09996_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net160),
    .D(_00037_),
    .Q_N(_04561_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _09997_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net161),
    .D(net1761),
    .Q_N(_04562_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[10][0] ));
 sg13g2_dfrbp_1 _09998_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net162),
    .D(net1085),
    .Q_N(_04563_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[10][1] ));
 sg13g2_dfrbp_1 _09999_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net163),
    .D(net1568),
    .Q_N(_04564_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[10][2] ));
 sg13g2_dfrbp_1 _10000_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net164),
    .D(net1783),
    .Q_N(_04565_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[10][3] ));
 sg13g2_dfrbp_1 _10001_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net165),
    .D(net1720),
    .Q_N(_04566_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10002_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net166),
    .D(net1743),
    .Q_N(_04567_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10003_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net167),
    .D(net1481),
    .Q_N(_04568_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10004_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net168),
    .D(net1660),
    .Q_N(_04569_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10005_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net169),
    .D(net1753),
    .Q_N(_04570_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10006_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net170),
    .D(net1080),
    .Q_N(_04571_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10007_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net171),
    .D(net1587),
    .Q_N(_04572_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10008_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net172),
    .D(net1549),
    .Q_N(_04573_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10009_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net173),
    .D(net1534),
    .Q_N(_04574_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10010_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net174),
    .D(net1733),
    .Q_N(_04575_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10011_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net175),
    .D(net1715),
    .Q_N(_04576_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10012_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net176),
    .D(net1052),
    .Q_N(_04577_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10013_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net177),
    .D(net1569),
    .Q_N(_04578_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10014_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net178),
    .D(net1516),
    .Q_N(_04579_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10015_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net179),
    .D(net1654),
    .Q_N(_04580_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10016_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net180),
    .D(net1487),
    .Q_N(_04581_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10017_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net181),
    .D(net1503),
    .Q_N(_04582_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10018_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net182),
    .D(net1651),
    .Q_N(_04583_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10019_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net183),
    .D(net1754),
    .Q_N(_04584_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10020_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net184),
    .D(net1746),
    .Q_N(_04585_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10021_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net185),
    .D(net1667),
    .Q_N(_04586_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10022_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net186),
    .D(net1664),
    .Q_N(_04587_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10023_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net187),
    .D(net1537),
    .Q_N(_04588_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10024_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net188),
    .D(net1774),
    .Q_N(_04589_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10025_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net189),
    .D(_00030_),
    .Q_N(_04590_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10026_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net190),
    .D(_00031_),
    .Q_N(_04591_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10027_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net191),
    .D(_00032_),
    .Q_N(_04592_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10028_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net192),
    .D(_00033_),
    .Q_N(_04593_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _10029_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net193),
    .D(net1824),
    .Q_N(_04594_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[9][0] ));
 sg13g2_dfrbp_1 _10030_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net194),
    .D(net1784),
    .Q_N(_04595_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[9][1] ));
 sg13g2_dfrbp_1 _10031_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net195),
    .D(net1820),
    .Q_N(_04596_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[9][2] ));
 sg13g2_dfrbp_1 _10032_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net196),
    .D(net1821),
    .Q_N(_04597_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[9][3] ));
 sg13g2_dfrbp_1 _10033_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net197),
    .D(net1704),
    .Q_N(_04598_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10034_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net198),
    .D(net1486),
    .Q_N(_04599_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10035_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net199),
    .D(net1573),
    .Q_N(_04600_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10036_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net200),
    .D(net1066),
    .Q_N(_04601_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10037_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net201),
    .D(net1536),
    .Q_N(_04602_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10038_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net202),
    .D(net1722),
    .Q_N(_04603_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10039_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net203),
    .D(net1585),
    .Q_N(_04604_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10040_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net204),
    .D(net1581),
    .Q_N(_04605_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10041_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net205),
    .D(net1605),
    .Q_N(_04606_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10042_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net206),
    .D(net1630),
    .Q_N(_04607_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10043_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net207),
    .D(net1100),
    .Q_N(_04608_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10044_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net208),
    .D(net1730),
    .Q_N(_04609_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10045_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net209),
    .D(net1099),
    .Q_N(_04610_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10046_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net210),
    .D(net1518),
    .Q_N(_04611_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10047_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net211),
    .D(net1586),
    .Q_N(_04612_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10048_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net212),
    .D(net1517),
    .Q_N(_04613_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10049_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net213),
    .D(net1594),
    .Q_N(_04614_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10050_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net214),
    .D(net1519),
    .Q_N(_04615_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10051_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net215),
    .D(net1505),
    .Q_N(_04616_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10052_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net216),
    .D(net1531),
    .Q_N(_04617_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10053_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net217),
    .D(net1053),
    .Q_N(_04618_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10054_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net218),
    .D(net1647),
    .Q_N(_04619_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10055_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net219),
    .D(net1056),
    .Q_N(_04620_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10056_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net220),
    .D(net1073),
    .Q_N(_04621_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10057_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net221),
    .D(_00078_),
    .Q_N(_04622_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10058_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net222),
    .D(_00079_),
    .Q_N(_04623_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10059_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net223),
    .D(_00080_),
    .Q_N(_04624_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10060_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net224),
    .D(_00081_),
    .Q_N(_04625_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _10061_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net225),
    .D(net1795),
    .Q_N(_04626_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[8][0] ));
 sg13g2_dfrbp_1 _10062_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net226),
    .D(net1108),
    .Q_N(_04627_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[8][1] ));
 sg13g2_dfrbp_1 _10063_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net227),
    .D(net1813),
    .Q_N(_04628_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[8][2] ));
 sg13g2_dfrbp_1 _10064_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net228),
    .D(net1776),
    .Q_N(_04629_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[8][3] ));
 sg13g2_dfrbp_1 _10065_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net229),
    .D(net1699),
    .Q_N(_04630_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10066_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net230),
    .D(net1796),
    .Q_N(_04631_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10067_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net231),
    .D(net1523),
    .Q_N(_04632_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10068_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net232),
    .D(net1600),
    .Q_N(_04633_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10069_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net233),
    .D(net1105),
    .Q_N(_04634_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10070_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net234),
    .D(net1548),
    .Q_N(_04635_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10071_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net235),
    .D(net1635),
    .Q_N(_04636_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10072_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net236),
    .D(net1641),
    .Q_N(_04637_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10073_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net237),
    .D(net1530),
    .Q_N(_04638_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10074_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net238),
    .D(net1520),
    .Q_N(_04639_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10075_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net239),
    .D(net1541),
    .Q_N(_04640_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10076_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net240),
    .D(net1095),
    .Q_N(_04641_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10077_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net241),
    .D(net1613),
    .Q_N(_04642_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10078_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net242),
    .D(net1694),
    .Q_N(_04643_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10079_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net243),
    .D(net1500),
    .Q_N(_04644_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10080_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net244),
    .D(net1599),
    .Q_N(_04645_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10081_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net245),
    .D(net1687),
    .Q_N(_04646_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10082_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net246),
    .D(net1554),
    .Q_N(_04647_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10083_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net247),
    .D(net1597),
    .Q_N(_04648_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10084_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net248),
    .D(net1521),
    .Q_N(_04649_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10085_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net249),
    .D(net1745),
    .Q_N(_04650_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10086_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net250),
    .D(net1691),
    .Q_N(_04651_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10087_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net251),
    .D(net1764),
    .Q_N(_04652_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10088_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net252),
    .D(net1765),
    .Q_N(_04653_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10089_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net253),
    .D(_00074_),
    .Q_N(_04654_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10090_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net254),
    .D(_00075_),
    .Q_N(_04655_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10091_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net255),
    .D(_00076_),
    .Q_N(_04656_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10092_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net256),
    .D(_00077_),
    .Q_N(_04657_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _10093_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net257),
    .D(net1805),
    .Q_N(_04658_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_dfrbp_1 _10094_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net258),
    .D(net1809),
    .Q_N(_04659_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[7][1] ));
 sg13g2_dfrbp_1 _10095_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net259),
    .D(net1804),
    .Q_N(_04660_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[7][2] ));
 sg13g2_dfrbp_1 _10096_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net260),
    .D(net1823),
    .Q_N(_04661_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[7][3] ));
 sg13g2_dfrbp_1 _10097_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net261),
    .D(net1723),
    .Q_N(_04662_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10098_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net262),
    .D(net1779),
    .Q_N(_04663_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10099_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net263),
    .D(net1785),
    .Q_N(_04664_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10100_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net264),
    .D(net1087),
    .Q_N(_04665_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10101_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net265),
    .D(net1710),
    .Q_N(_04666_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10102_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net266),
    .D(net1477),
    .Q_N(_04667_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10103_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net267),
    .D(net1557),
    .Q_N(_04668_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10104_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net268),
    .D(net1502),
    .Q_N(_04669_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10105_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net269),
    .D(net1507),
    .Q_N(_04670_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10106_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net270),
    .D(net1063),
    .Q_N(_04671_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10107_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net271),
    .D(net1086),
    .Q_N(_04672_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10108_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net272),
    .D(net1058),
    .Q_N(_04673_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10109_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net273),
    .D(net1645),
    .Q_N(_04674_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10110_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net274),
    .D(net1563),
    .Q_N(_04675_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10111_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net275),
    .D(net1590),
    .Q_N(_04676_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10112_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net276),
    .D(net1565),
    .Q_N(_04677_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10113_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net277),
    .D(net1793),
    .Q_N(_04678_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10114_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net278),
    .D(net1050),
    .Q_N(_04679_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10115_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net279),
    .D(net1062),
    .Q_N(_04680_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10116_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net280),
    .D(net1093),
    .Q_N(_04681_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10117_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net281),
    .D(net1709),
    .Q_N(_04682_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10118_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net282),
    .D(net1480),
    .Q_N(_04683_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10119_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net283),
    .D(net1054),
    .Q_N(_04684_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10120_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net284),
    .D(net1498),
    .Q_N(_04685_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10121_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net285),
    .D(_00070_),
    .Q_N(_04686_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10122_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net286),
    .D(_00071_),
    .Q_N(_04687_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10123_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net287),
    .D(_00072_),
    .Q_N(_04688_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10124_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net288),
    .D(_00073_),
    .Q_N(_04689_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _10125_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net289),
    .D(net1642),
    .Q_N(_04690_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[6][0] ));
 sg13g2_dfrbp_1 _10126_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net290),
    .D(net1512),
    .Q_N(_04691_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[6][1] ));
 sg13g2_dfrbp_1 _10127_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net291),
    .D(net1578),
    .Q_N(_04692_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[6][2] ));
 sg13g2_dfrbp_1 _10128_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net292),
    .D(net1759),
    .Q_N(_04693_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[6][3] ));
 sg13g2_dfrbp_1 _10129_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net293),
    .D(net1075),
    .Q_N(_04694_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10130_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net294),
    .D(net1655),
    .Q_N(_04695_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10131_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net295),
    .D(net1671),
    .Q_N(_04696_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10132_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net296),
    .D(net1074),
    .Q_N(_04697_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10133_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net297),
    .D(net1683),
    .Q_N(_04698_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10134_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net298),
    .D(net1726),
    .Q_N(_04699_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10135_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net299),
    .D(net1103),
    .Q_N(_04700_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10136_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net300),
    .D(net1471),
    .Q_N(_04701_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10137_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net301),
    .D(net1535),
    .Q_N(_04702_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10138_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net302),
    .D(net1522),
    .Q_N(_04703_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10139_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net303),
    .D(net1533),
    .Q_N(_04704_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10140_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net304),
    .D(net1482),
    .Q_N(_04705_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10141_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net305),
    .D(net1539),
    .Q_N(_04706_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10142_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net306),
    .D(net1524),
    .Q_N(_04707_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10143_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net307),
    .D(net1560),
    .Q_N(_04708_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10144_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net308),
    .D(net1510),
    .Q_N(_04709_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10145_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net309),
    .D(net1661),
    .Q_N(_04710_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10146_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net310),
    .D(net1525),
    .Q_N(_04711_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10147_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net311),
    .D(net1703),
    .Q_N(_04712_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10148_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net312),
    .D(net1558),
    .Q_N(_04713_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10149_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net313),
    .D(net1579),
    .Q_N(_04714_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10150_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net314),
    .D(net1792),
    .Q_N(_04715_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10151_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net315),
    .D(net1508),
    .Q_N(_04716_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10152_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net316),
    .D(net1806),
    .Q_N(_04717_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10153_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net317),
    .D(_00066_),
    .Q_N(_04718_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10154_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net318),
    .D(_00067_),
    .Q_N(_04719_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10155_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net319),
    .D(_00068_),
    .Q_N(_04720_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10156_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net320),
    .D(_00069_),
    .Q_N(_04721_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _10157_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net321),
    .D(net1769),
    .Q_N(_04722_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[5][0] ));
 sg13g2_dfrbp_1 _10158_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net322),
    .D(net1712),
    .Q_N(_04723_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[5][1] ));
 sg13g2_dfrbp_1 _10159_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net323),
    .D(net1076),
    .Q_N(_04724_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[5][2] ));
 sg13g2_dfrbp_1 _10160_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net324),
    .D(net1606),
    .Q_N(_04725_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[5][3] ));
 sg13g2_dfrbp_1 _10161_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net325),
    .D(net1780),
    .Q_N(_04726_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10162_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net326),
    .D(net1781),
    .Q_N(_04727_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10163_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net327),
    .D(net1725),
    .Q_N(_04728_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10164_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net328),
    .D(net1739),
    .Q_N(_04729_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10165_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net329),
    .D(net1495),
    .Q_N(_04730_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10166_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net330),
    .D(net1496),
    .Q_N(_04731_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10167_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net331),
    .D(net1601),
    .Q_N(_04732_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10168_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net332),
    .D(net1562),
    .Q_N(_04733_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10169_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net333),
    .D(net1595),
    .Q_N(_04734_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10170_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net334),
    .D(net1071),
    .Q_N(_04735_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10171_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net335),
    .D(net1695),
    .Q_N(_04736_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10172_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net336),
    .D(net1582),
    .Q_N(_04737_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10173_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net337),
    .D(net1639),
    .Q_N(_04738_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10174_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net338),
    .D(net1672),
    .Q_N(_04739_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10175_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net339),
    .D(net1474),
    .Q_N(_04740_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10176_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net340),
    .D(net1682),
    .Q_N(_04741_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10177_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net341),
    .D(net1061),
    .Q_N(_04742_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10178_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net342),
    .D(net1096),
    .Q_N(_04743_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10179_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net343),
    .D(net1643),
    .Q_N(_04744_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10180_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net344),
    .D(net1514),
    .Q_N(_04745_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10181_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net345),
    .D(net1629),
    .Q_N(_04746_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10182_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net346),
    .D(net1602),
    .Q_N(_04747_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10183_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net347),
    .D(net1650),
    .Q_N(_04748_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10184_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net348),
    .D(net1593),
    .Q_N(_04749_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10185_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net349),
    .D(_00062_),
    .Q_N(_04750_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10186_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net350),
    .D(_00063_),
    .Q_N(_04751_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10187_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net351),
    .D(_00064_),
    .Q_N(_04752_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10188_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net352),
    .D(_00065_),
    .Q_N(_04753_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _10189_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net353),
    .D(net1782),
    .Q_N(_04754_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[2][0] ));
 sg13g2_dfrbp_1 _10190_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net354),
    .D(net1760),
    .Q_N(_04755_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[2][1] ));
 sg13g2_dfrbp_1 _10191_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net355),
    .D(net1729),
    .Q_N(_04756_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[2][2] ));
 sg13g2_dfrbp_1 _10192_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net356),
    .D(net1775),
    .Q_N(_04757_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[2][3] ));
 sg13g2_dfrbp_1 _10193_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net357),
    .D(net1666),
    .Q_N(_04758_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10194_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net358),
    .D(net1706),
    .Q_N(_04759_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10195_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net359),
    .D(net1509),
    .Q_N(_04760_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10196_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net360),
    .D(net1685),
    .Q_N(_04761_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10197_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net361),
    .D(net1542),
    .Q_N(_04762_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10198_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net362),
    .D(net1091),
    .Q_N(_04763_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10199_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net363),
    .D(net1057),
    .Q_N(_04764_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10200_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net364),
    .D(net1544),
    .Q_N(_04765_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10201_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net365),
    .D(net1090),
    .Q_N(_04766_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10202_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net366),
    .D(net1634),
    .Q_N(_04767_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10203_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net367),
    .D(net1744),
    .Q_N(_04768_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10204_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net368),
    .D(net1543),
    .Q_N(_04769_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10205_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net369),
    .D(net1490),
    .Q_N(_04770_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10206_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net370),
    .D(net1656),
    .Q_N(_04771_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10207_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net371),
    .D(net1632),
    .Q_N(_04772_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10208_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net372),
    .D(net1106),
    .Q_N(_04773_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10209_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net373),
    .D(net1636),
    .Q_N(_04774_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10210_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net374),
    .D(net1740),
    .Q_N(_04775_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10211_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net375),
    .D(net1737),
    .Q_N(_04776_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10212_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net376),
    .D(net1659),
    .Q_N(_04777_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10213_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net377),
    .D(net1762),
    .Q_N(_04778_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10214_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net378),
    .D(net1501),
    .Q_N(_04779_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10215_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net379),
    .D(net1696),
    .Q_N(_04780_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10216_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net380),
    .D(net1777),
    .Q_N(_04781_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10217_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net381),
    .D(_00058_),
    .Q_N(_04782_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10218_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net382),
    .D(_00059_),
    .Q_N(_04783_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10219_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net383),
    .D(_00060_),
    .Q_N(_04784_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10220_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net384),
    .D(_00061_),
    .Q_N(_04785_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _10221_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net385),
    .D(net1700),
    .Q_N(_04786_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[1][0] ));
 sg13g2_dfrbp_1 _10222_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net386),
    .D(net1825),
    .Q_N(_04787_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[1][1] ));
 sg13g2_dfrbp_1 _10223_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net387),
    .D(net1826),
    .Q_N(_04788_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[1][2] ));
 sg13g2_dfrbp_1 _10224_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net388),
    .D(net1827),
    .Q_N(_04789_),
    .Q(\i_core.cpu.i_core.i_registers.reg_access[1][3] ));
 sg13g2_dfrbp_1 _10225_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net389),
    .D(net1790),
    .Q_N(_04790_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10226_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net390),
    .D(net1810),
    .Q_N(_04791_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10227_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net391),
    .D(net1814),
    .Q_N(_04792_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10228_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net392),
    .D(net1812),
    .Q_N(_04793_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10229_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net393),
    .D(net1818),
    .Q_N(_04794_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10230_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net394),
    .D(net1797),
    .Q_N(_04795_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10231_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net395),
    .D(net1791),
    .Q_N(_04796_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10232_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net396),
    .D(net1724),
    .Q_N(_04797_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10233_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net397),
    .D(net1755),
    .Q_N(_04798_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10234_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net398),
    .D(net1773),
    .Q_N(_04799_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10235_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net399),
    .D(net1766),
    .Q_N(_04800_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10236_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net400),
    .D(net1794),
    .Q_N(_04801_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10237_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net401),
    .D(net1758),
    .Q_N(_04802_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10238_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net402),
    .D(net1787),
    .Q_N(_04803_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10239_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net403),
    .D(net1749),
    .Q_N(_04804_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10240_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net404),
    .D(net1750),
    .Q_N(_04805_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10241_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net405),
    .D(net1887),
    .Q_N(_04806_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10242_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net406),
    .D(net2016),
    .Q_N(_04807_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10243_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net407),
    .D(net2092),
    .Q_N(_04808_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10244_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net408),
    .D(net1898),
    .Q_N(_04809_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10245_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net409),
    .D(net1770),
    .Q_N(_04810_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10246_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net410),
    .D(net1532),
    .Q_N(_04811_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10247_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net411),
    .D(net1698),
    .Q_N(_04812_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10248_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net412),
    .D(net1811),
    .Q_N(_04813_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10249_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net413),
    .D(_00054_),
    .Q_N(_04814_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10250_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net414),
    .D(_00055_),
    .Q_N(_04815_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10251_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net415),
    .D(_00056_),
    .Q_N(_04816_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10252_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net427),
    .D(_00057_),
    .Q_N(_04817_),
    .Q(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _10253_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net1036),
    .D(\i_core.cpu.i_core.cy_out ),
    .Q_N(_00095_),
    .Q(\i_core.cpu.i_core.cy ));
 sg13g2_dfrbp_1 _10254_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net629),
    .D(net2190),
    .Q_N(_04404_),
    .Q(\i_core.cpu.i_core.load_done ));
 sg13g2_dfrbp_1 _10255_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net628),
    .D(_00225_),
    .Q_N(_00085_),
    .Q(\i_core.cpu.i_core.cycle[0] ));
 sg13g2_dfrbp_1 _10256_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net626),
    .D(_00226_),
    .Q_N(_04403_),
    .Q(\i_core.cpu.i_core.cycle[1] ));
 sg13g2_dfrbp_1 _10257_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net624),
    .D(_00227_),
    .Q_N(_04402_),
    .Q(\i_core.cpu.i_core.mcause[0] ));
 sg13g2_dfrbp_1 _10258_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net622),
    .D(net2384),
    .Q_N(_04401_),
    .Q(\i_core.cpu.i_core.mcause[1] ));
 sg13g2_dfrbp_1 _10259_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net620),
    .D(net1967),
    .Q_N(_04400_),
    .Q(\i_core.cpu.i_core.mcause[3] ));
 sg13g2_dfrbp_1 _10260_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net618),
    .D(_00230_),
    .Q_N(_04399_),
    .Q(\i_core.cpu.i_core.mcause[4] ));
 sg13g2_dfrbp_1 _10261_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net616),
    .D(net2286),
    .Q_N(_04398_),
    .Q(\i_core.cpu.i_core.is_double_fault_r ));
 sg13g2_dfrbp_1 _10262_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net615),
    .D(net1945),
    .Q_N(_00222_),
    .Q(\i_core.cpu.i_core.time_hi[0] ));
 sg13g2_dfrbp_1 _10263_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net613),
    .D(net2129),
    .Q_N(_04397_),
    .Q(\i_core.cpu.i_core.time_hi[1] ));
 sg13g2_dfrbp_1 _10264_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net442),
    .D(net2009),
    .Q_N(_04818_),
    .Q(\i_core.cpu.i_core.time_hi[2] ));
 sg13g2_dfrbp_1 _10265_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net611),
    .D(_00029_),
    .Q_N(_00216_),
    .Q(\i_core.cpu.i_core.i_instrret.add ));
 sg13g2_dfrbp_1 _10266_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net609),
    .D(net2131),
    .Q_N(_04396_),
    .Q(\i_core.cpu.i_core.last_interrupt_req[0] ));
 sg13g2_dfrbp_1 _10267_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net608),
    .D(net2148),
    .Q_N(_04395_),
    .Q(\i_core.cpu.i_core.last_interrupt_req[1] ));
 sg13g2_dfrbp_1 _10268_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net607),
    .D(_00237_),
    .Q_N(_04394_),
    .Q(\i_core.cpu.i_core.mepc[20] ));
 sg13g2_dfrbp_1 _10269_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net605),
    .D(_00238_),
    .Q_N(_04393_),
    .Q(\i_core.cpu.i_core.mepc[21] ));
 sg13g2_dfrbp_1 _10270_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net603),
    .D(_00239_),
    .Q_N(_04392_),
    .Q(\i_core.cpu.i_core.mepc[22] ));
 sg13g2_dfrbp_1 _10271_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net601),
    .D(_00240_),
    .Q_N(_04391_),
    .Q(\i_core.cpu.i_core.mepc[23] ));
 sg13g2_dfrbp_1 _10272_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net599),
    .D(net2363),
    .Q_N(_04390_),
    .Q(\i_core.cpu.i_core.mstatus_mpie ));
 sg13g2_dfrbp_1 _10273_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net597),
    .D(net2559),
    .Q_N(_04389_),
    .Q(\i_core.cpu.i_core.mstatus_mie ));
 sg13g2_dfrbp_1 _10274_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net595),
    .D(net2441),
    .Q_N(_04388_),
    .Q(\i_core.cpu.i_core.mstatus_mte ));
 sg13g2_dfrbp_1 _10275_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net593),
    .D(net1926),
    .Q_N(_00215_),
    .Q(\i_core.cpu.i_core.i_registers.rd[0] ));
 sg13g2_dfrbp_1 _10276_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net592),
    .D(_00245_),
    .Q_N(_04387_),
    .Q(\i_core.cpu.i_core.i_registers.rd[1] ));
 sg13g2_dfrbp_1 _10277_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net591),
    .D(_00246_),
    .Q_N(_04386_),
    .Q(\i_core.cpu.i_core.i_registers.rd[2] ));
 sg13g2_dfrbp_1 _10278_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net590),
    .D(_00247_),
    .Q_N(_04385_),
    .Q(\i_core.cpu.i_core.i_registers.rd[3] ));
 sg13g2_dfrbp_1 _10279_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net443),
    .D(_00248_),
    .Q_N(_04819_),
    .Q(\i_core.cpu.i_core.load_top_bit ));
 sg13g2_dfrbp_1 _10280_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net536),
    .D(\i_core.cpu.i_core.cmp_out ),
    .Q_N(_04820_),
    .Q(\i_core.cpu.i_core.cmp ));
 sg13g2_dfrbp_1 _10281_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net589),
    .D(net1323),
    .Q_N(_00153_),
    .Q(\i_core.cpu.i_core.i_cycles.rstn ));
 sg13g2_dfrbp_1 _10282_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net587),
    .D(_00249_),
    .Q_N(_04384_),
    .Q(\i_uart_tx.data_to_send[0] ));
 sg13g2_dfrbp_1 _10283_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net585),
    .D(_00250_),
    .Q_N(_04383_),
    .Q(\i_uart_tx.data_to_send[1] ));
 sg13g2_dfrbp_1 _10284_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net583),
    .D(_00251_),
    .Q_N(_04382_),
    .Q(\i_uart_tx.data_to_send[2] ));
 sg13g2_dfrbp_1 _10285_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net581),
    .D(net2609),
    .Q_N(_04381_),
    .Q(\i_uart_tx.data_to_send[3] ));
 sg13g2_dfrbp_1 _10286_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net579),
    .D(_00253_),
    .Q_N(_04380_),
    .Q(\i_uart_tx.data_to_send[4] ));
 sg13g2_dfrbp_1 _10287_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net577),
    .D(net2611),
    .Q_N(_04379_),
    .Q(\i_uart_tx.data_to_send[5] ));
 sg13g2_dfrbp_1 _10288_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net575),
    .D(net2603),
    .Q_N(_04378_),
    .Q(\i_uart_tx.data_to_send[6] ));
 sg13g2_dfrbp_1 _10289_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net573),
    .D(net1915),
    .Q_N(_04377_),
    .Q(\i_uart_tx.data_to_send[7] ));
 sg13g2_dfrbp_1 _10290_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net571),
    .D(_00257_),
    .Q_N(_00221_),
    .Q(\i_uart_tx.cycle_counter[0] ));
 sg13g2_dfrbp_1 _10291_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net569),
    .D(net1970),
    .Q_N(_04376_),
    .Q(\i_uart_tx.cycle_counter[1] ));
 sg13g2_dfrbp_1 _10292_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net567),
    .D(_00259_),
    .Q_N(_04375_),
    .Q(\i_uart_tx.cycle_counter[2] ));
 sg13g2_dfrbp_1 _10293_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net565),
    .D(_00260_),
    .Q_N(_04374_),
    .Q(\i_uart_tx.cycle_counter[3] ));
 sg13g2_dfrbp_1 _10294_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net563),
    .D(_00261_),
    .Q_N(_04373_),
    .Q(\i_uart_tx.cycle_counter[4] ));
 sg13g2_dfrbp_1 _10295_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net561),
    .D(_00262_),
    .Q_N(_04372_),
    .Q(\i_uart_tx.cycle_counter[5] ));
 sg13g2_dfrbp_1 _10296_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net559),
    .D(_00263_),
    .Q_N(_04371_),
    .Q(\i_uart_tx.cycle_counter[6] ));
 sg13g2_dfrbp_1 _10297_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net535),
    .D(net2105),
    .Q_N(_04370_),
    .Q(\i_uart_tx.cycle_counter[7] ));
 sg13g2_dfrbp_1 _10298_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net533),
    .D(_00265_),
    .Q_N(_04369_),
    .Q(\i_uart_tx.cycle_counter[8] ));
 sg13g2_dfrbp_1 _10299_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net531),
    .D(_00266_),
    .Q_N(_04368_),
    .Q(\i_uart_tx.cycle_counter[9] ));
 sg13g2_dfrbp_1 _10300_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net529),
    .D(_00267_),
    .Q_N(_04367_),
    .Q(\i_uart_tx.cycle_counter[10] ));
 sg13g2_dfrbp_1 _10301_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net527),
    .D(_00268_),
    .Q_N(_04366_),
    .Q(\i_uart_tx.fsm_state[0] ));
 sg13g2_dfrbp_1 _10302_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net525),
    .D(_00269_),
    .Q_N(_04365_),
    .Q(\i_uart_tx.fsm_state[1] ));
 sg13g2_dfrbp_1 _10303_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net523),
    .D(net2367),
    .Q_N(_04364_),
    .Q(\i_uart_tx.fsm_state[2] ));
 sg13g2_dfrbp_1 _10304_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net521),
    .D(net2519),
    .Q_N(_04363_),
    .Q(\i_uart_tx.fsm_state[3] ));
 sg13g2_dfrbp_1 _10305_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net519),
    .D(net2165),
    .Q_N(_04362_),
    .Q(\i_uart_rx.recieved_data[0] ));
 sg13g2_dfrbp_1 _10306_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net518),
    .D(net2249),
    .Q_N(_04361_),
    .Q(\i_uart_rx.recieved_data[1] ));
 sg13g2_dfrbp_1 _10307_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net517),
    .D(_00274_),
    .Q_N(_04360_),
    .Q(\i_uart_rx.recieved_data[2] ));
 sg13g2_dfrbp_1 _10308_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net516),
    .D(_00275_),
    .Q_N(_04359_),
    .Q(\i_uart_rx.recieved_data[3] ));
 sg13g2_dfrbp_1 _10309_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net515),
    .D(net2227),
    .Q_N(_04358_),
    .Q(\i_uart_rx.recieved_data[4] ));
 sg13g2_dfrbp_1 _10310_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net514),
    .D(_00277_),
    .Q_N(_04357_),
    .Q(\i_uart_rx.recieved_data[5] ));
 sg13g2_dfrbp_1 _10311_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net513),
    .D(_00278_),
    .Q_N(_04356_),
    .Q(\i_uart_rx.recieved_data[6] ));
 sg13g2_dfrbp_1 _10312_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net512),
    .D(net2027),
    .Q_N(_04355_),
    .Q(\i_uart_rx.recieved_data[7] ));
 sg13g2_dfrbp_1 _10313_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net511),
    .D(_00280_),
    .Q_N(_00220_),
    .Q(\i_uart_rx.cycle_counter[0] ));
 sg13g2_dfrbp_1 _10314_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net510),
    .D(net2096),
    .Q_N(_04354_),
    .Q(\i_uart_rx.cycle_counter[1] ));
 sg13g2_dfrbp_1 _10315_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net509),
    .D(_00282_),
    .Q_N(_04353_),
    .Q(\i_uart_rx.cycle_counter[2] ));
 sg13g2_dfrbp_1 _10316_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net508),
    .D(_00283_),
    .Q_N(_04352_),
    .Q(\i_uart_rx.cycle_counter[3] ));
 sg13g2_dfrbp_1 _10317_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net507),
    .D(_00284_),
    .Q_N(_04351_),
    .Q(\i_uart_rx.cycle_counter[4] ));
 sg13g2_dfrbp_1 _10318_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net506),
    .D(_00285_),
    .Q_N(_04350_),
    .Q(\i_uart_rx.cycle_counter[5] ));
 sg13g2_dfrbp_1 _10319_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net505),
    .D(_00286_),
    .Q_N(_04349_),
    .Q(\i_uart_rx.cycle_counter[6] ));
 sg13g2_dfrbp_1 _10320_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net504),
    .D(_00287_),
    .Q_N(_04348_),
    .Q(\i_uart_rx.cycle_counter[7] ));
 sg13g2_dfrbp_1 _10321_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net503),
    .D(_00288_),
    .Q_N(_04347_),
    .Q(\i_uart_rx.cycle_counter[8] ));
 sg13g2_dfrbp_1 _10322_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net502),
    .D(_00289_),
    .Q_N(_04346_),
    .Q(\i_uart_rx.cycle_counter[9] ));
 sg13g2_dfrbp_1 _10323_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net501),
    .D(_00290_),
    .Q_N(_04345_),
    .Q(\i_uart_rx.cycle_counter[10] ));
 sg13g2_dfrbp_1 _10324_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net500),
    .D(net2024),
    .Q_N(_04344_),
    .Q(\i_uart_rx.bit_sample ));
 sg13g2_dfrbp_1 _10325_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net498),
    .D(_00292_),
    .Q_N(_04343_),
    .Q(\i_uart_rx.uart_rts ));
 sg13g2_dfrbp_1 _10326_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net497),
    .D(net2473),
    .Q_N(_00203_),
    .Q(\i_uart_rx.fsm_state[0] ));
 sg13g2_dfrbp_1 _10327_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net495),
    .D(_00294_),
    .Q_N(_04342_),
    .Q(\i_uart_rx.fsm_state[1] ));
 sg13g2_dfrbp_1 _10328_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net493),
    .D(net2514),
    .Q_N(_04341_),
    .Q(\i_uart_rx.fsm_state[2] ));
 sg13g2_dfrbp_1 _10329_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net491),
    .D(net2570),
    .Q_N(_04340_),
    .Q(\i_uart_rx.fsm_state[3] ));
 sg13g2_dfrbp_1 _10330_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net489),
    .D(_00297_),
    .Q_N(_00204_),
    .Q(\i_uart_rx.rxd_reg[0] ));
 sg13g2_dfrbp_1 _10331_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net488),
    .D(_00298_),
    .Q_N(_04339_),
    .Q(\i_uart_rx.rxd_reg[1] ));
 sg13g2_dfrbp_1 _10332_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net487),
    .D(net2202),
    .Q_N(_04338_),
    .Q(\i_spi.end_txn_reg ));
 sg13g2_dfrbp_1 _10333_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net486),
    .D(net2046),
    .Q_N(_04337_),
    .Q(\i_core.cpu.instr_data[3][0] ));
 sg13g2_dfrbp_1 _10334_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net485),
    .D(net1947),
    .Q_N(_00102_),
    .Q(\i_core.cpu.instr_data[3][1] ));
 sg13g2_dfrbp_1 _10335_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net484),
    .D(_00302_),
    .Q_N(_04336_),
    .Q(\i_debug_uart_tx.data_to_send[0] ));
 sg13g2_dfrbp_1 _10336_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net482),
    .D(_00303_),
    .Q_N(_04335_),
    .Q(\i_debug_uart_tx.data_to_send[1] ));
 sg13g2_dfrbp_1 _10337_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net480),
    .D(net2624),
    .Q_N(_04334_),
    .Q(\i_debug_uart_tx.data_to_send[2] ));
 sg13g2_dfrbp_1 _10338_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net478),
    .D(net2598),
    .Q_N(_04333_),
    .Q(\i_debug_uart_tx.data_to_send[3] ));
 sg13g2_dfrbp_1 _10339_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net476),
    .D(_00306_),
    .Q_N(_04332_),
    .Q(\i_debug_uart_tx.data_to_send[4] ));
 sg13g2_dfrbp_1 _10340_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net474),
    .D(net2601),
    .Q_N(_04331_),
    .Q(\i_debug_uart_tx.data_to_send[5] ));
 sg13g2_dfrbp_1 _10341_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net472),
    .D(net2566),
    .Q_N(_04330_),
    .Q(\i_debug_uart_tx.data_to_send[6] ));
 sg13g2_dfrbp_1 _10342_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net470),
    .D(net1936),
    .Q_N(_04329_),
    .Q(\i_debug_uart_tx.data_to_send[7] ));
 sg13g2_dfrbp_1 _10343_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net468),
    .D(net1873),
    .Q_N(_00219_),
    .Q(\i_debug_uart_tx.cycle_counter[0] ));
 sg13g2_dfrbp_1 _10344_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net466),
    .D(net2225),
    .Q_N(_04328_),
    .Q(\i_debug_uart_tx.cycle_counter[1] ));
 sg13g2_dfrbp_1 _10345_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net464),
    .D(_00312_),
    .Q_N(_04327_),
    .Q(\i_debug_uart_tx.cycle_counter[2] ));
 sg13g2_dfrbp_1 _10346_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net462),
    .D(_00313_),
    .Q_N(_04326_),
    .Q(\i_debug_uart_tx.cycle_counter[3] ));
 sg13g2_dfrbp_1 _10347_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net460),
    .D(_00314_),
    .Q_N(_04325_),
    .Q(\i_debug_uart_tx.cycle_counter[4] ));
 sg13g2_dfrbp_1 _10348_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net458),
    .D(_00315_),
    .Q_N(_04324_),
    .Q(\i_debug_uart_tx.fsm_state[0] ));
 sg13g2_dfrbp_1 _10349_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net456),
    .D(_00316_),
    .Q_N(_04323_),
    .Q(\i_debug_uart_tx.fsm_state[1] ));
 sg13g2_dfrbp_1 _10350_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net454),
    .D(net2293),
    .Q_N(_04322_),
    .Q(\i_debug_uart_tx.fsm_state[2] ));
 sg13g2_dfrbp_1 _10351_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net452),
    .D(_00318_),
    .Q_N(_04321_),
    .Q(\i_debug_uart_tx.fsm_state[3] ));
 sg13g2_dfrbp_1 _10352_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net450),
    .D(_00319_),
    .Q_N(_04320_),
    .Q(\i_core.mem.q_ctrl.stop_txn_reg ));
 sg13g2_dfrbp_1 _10353_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net449),
    .D(_00320_),
    .Q_N(_04319_),
    .Q(\i_spi.clock_count[0] ));
 sg13g2_dfrbp_1 _10354_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net447),
    .D(net2485),
    .Q_N(_04318_),
    .Q(\i_spi.clock_count[1] ));
 sg13g2_dfrbp_1 _10355_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net445),
    .D(_00322_),
    .Q_N(_04317_),
    .Q(\i_spi.data[0] ));
 sg13g2_dfrbp_1 _10356_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net444),
    .D(net1979),
    .Q_N(_04316_),
    .Q(\i_spi.bits_remaining[0] ));
 sg13g2_dfrbp_1 _10357_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net440),
    .D(_00324_),
    .Q_N(_04315_),
    .Q(\i_spi.bits_remaining[1] ));
 sg13g2_dfrbp_1 _10358_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net438),
    .D(_00325_),
    .Q_N(_04314_),
    .Q(\i_spi.bits_remaining[2] ));
 sg13g2_dfrbp_1 _10359_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net436),
    .D(net2317),
    .Q_N(_04313_),
    .Q(\i_spi.bits_remaining[3] ));
 sg13g2_dfrbp_1 _10360_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net434),
    .D(_00327_),
    .Q_N(_00156_),
    .Q(\i_spi.busy ));
 sg13g2_dfrbp_1 _10361_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net433),
    .D(net2156),
    .Q_N(_04312_),
    .Q(\i_spi.spi_dc ));
 sg13g2_dfrbp_1 _10362_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net432),
    .D(net2135),
    .Q_N(_04311_),
    .Q(\i_spi.spi_select ));
 sg13g2_dfrbp_1 _10363_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net430),
    .D(_00330_),
    .Q_N(_00155_),
    .Q(\i_spi.spi_clk_out ));
 sg13g2_dfrbp_1 _10364_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net428),
    .D(net2400),
    .Q_N(_04310_),
    .Q(debug_uart_txd));
 sg13g2_dfrbp_1 _10365_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net426),
    .D(_00332_),
    .Q_N(_04309_),
    .Q(\i_spi.read_latency ));
 sg13g2_dfrbp_1 _10366_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net424),
    .D(_00333_),
    .Q_N(_04308_),
    .Q(\i_spi.clock_divider[0] ));
 sg13g2_dfrbp_1 _10367_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net422),
    .D(_00334_),
    .Q_N(_04307_),
    .Q(\i_spi.clock_divider[1] ));
 sg13g2_dfrbp_1 _10368_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net420),
    .D(net2421),
    .Q_N(_04306_),
    .Q(\i_core.cpu.i_core.mip[17] ));
 sg13g2_dfrbp_1 _10369_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net418),
    .D(net2339),
    .Q_N(_04305_),
    .Q(\i_core.cpu.i_core.mip[16] ));
 sg13g2_dfrbp_1 _10370_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net416),
    .D(net2169),
    .Q_N(_04304_),
    .Q(\i_core.cpu.i_core.mie[19] ));
 sg13g2_dfrbp_1 _10371_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net1034),
    .D(_00338_),
    .Q_N(_04303_),
    .Q(\i_core.cpu.i_core.mie[18] ));
 sg13g2_dfrbp_1 _10372_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net1032),
    .D(net2284),
    .Q_N(_04302_),
    .Q(\i_core.cpu.i_core.mie[17] ));
 sg13g2_dfrbp_1 _10373_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net537),
    .D(_00340_),
    .Q_N(_04821_),
    .Q(\i_core.cpu.i_core.mie[16] ));
 sg13g2_dfrbp_1 _10374_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net538),
    .D(\debug_rd[0] ),
    .Q_N(_04822_),
    .Q(\debug_rd_r[0] ));
 sg13g2_dfrbp_1 _10375_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net539),
    .D(net1132),
    .Q_N(_04823_),
    .Q(\debug_rd_r[1] ));
 sg13g2_dfrbp_1 _10376_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net541),
    .D(net1127),
    .Q_N(_04824_),
    .Q(\debug_rd_r[2] ));
 sg13g2_dfrbp_1 _10377_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net1030),
    .D(\debug_rd[3] ),
    .Q_N(_04301_),
    .Q(\debug_rd_r[3] ));
 sg13g2_dfrbp_1 _10378_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net542),
    .D(net2387),
    .Q_N(_04825_),
    .Q(\i_uart_tx.txd_reg ));
 sg13g2_dfrbp_1 _10379_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net543),
    .D(_00008_),
    .Q_N(_04826_),
    .Q(\gpio_out_sel[0] ));
 sg13g2_dfrbp_1 _10380_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net544),
    .D(_00009_),
    .Q_N(_04827_),
    .Q(\gpio_out_sel[1] ));
 sg13g2_dfrbp_1 _10381_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net545),
    .D(net2194),
    .Q_N(_04828_),
    .Q(\gpio_out_sel[2] ));
 sg13g2_dfrbp_1 _10382_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net546),
    .D(net2196),
    .Q_N(_04829_),
    .Q(\gpio_out_sel[3] ));
 sg13g2_dfrbp_1 _10383_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net547),
    .D(net2247),
    .Q_N(_04830_),
    .Q(\gpio_out_sel[4] ));
 sg13g2_dfrbp_1 _10384_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net548),
    .D(net2254),
    .Q_N(_04831_),
    .Q(\gpio_out_sel[5] ));
 sg13g2_dfrbp_1 _10385_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net549),
    .D(net2311),
    .Q_N(_04832_),
    .Q(\gpio_out_sel[6] ));
 sg13g2_dfrbp_1 _10386_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net550),
    .D(_00015_),
    .Q_N(_04833_),
    .Q(\gpio_out_sel[7] ));
 sg13g2_dfrbp_1 _10387_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net551),
    .D(_00000_),
    .Q_N(_04834_),
    .Q(\gpio_out[0] ));
 sg13g2_dfrbp_1 _10388_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net552),
    .D(_00001_),
    .Q_N(_04835_),
    .Q(\gpio_out[1] ));
 sg13g2_dfrbp_1 _10389_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net553),
    .D(net2011),
    .Q_N(_04836_),
    .Q(\gpio_out[2] ));
 sg13g2_dfrbp_1 _10390_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net554),
    .D(net2015),
    .Q_N(_04837_),
    .Q(\gpio_out[3] ));
 sg13g2_dfrbp_1 _10391_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net555),
    .D(net1987),
    .Q_N(_04838_),
    .Q(\gpio_out[4] ));
 sg13g2_dfrbp_1 _10392_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net556),
    .D(net2102),
    .Q_N(_04839_),
    .Q(\gpio_out[5] ));
 sg13g2_dfrbp_1 _10393_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net557),
    .D(net2067),
    .Q_N(_04840_),
    .Q(\gpio_out[6] ));
 sg13g2_dfrbp_1 _10394_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net558),
    .D(net1989),
    .Q_N(_04841_),
    .Q(\gpio_out[7] ));
 sg13g2_dfrbp_1 _10395_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net707),
    .D(net2),
    .Q_N(_04842_),
    .Q(\i_core.cpu.i_core.interrupt_req[0] ));
 sg13g2_dfrbp_1 _10396_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1000),
    .D(net3),
    .Q_N(_04300_),
    .Q(\i_core.cpu.i_core.interrupt_req[1] ));
 sg13g2_dfrbp_1 _10397_ (.CLK(net1049),
    .RESET_B(net999),
    .D(net1),
    .Q_N(_00154_),
    .Q(\i_core.mem.q_ctrl.rstn ));
 sg13g2_dfrbp_1 _10398_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net998),
    .D(net2544),
    .Q_N(_00198_),
    .Q(\i_core.cpu.i_core.i_shift.a[0] ));
 sg13g2_dfrbp_1 _10399_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net997),
    .D(net2468),
    .Q_N(_00196_),
    .Q(\i_core.cpu.i_core.i_shift.a[1] ));
 sg13g2_dfrbp_1 _10400_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net996),
    .D(net2528),
    .Q_N(_00194_),
    .Q(\i_core.cpu.i_core.i_shift.a[2] ));
 sg13g2_dfrbp_1 _10401_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net967),
    .D(net2475),
    .Q_N(_00168_),
    .Q(\i_core.cpu.i_core.i_shift.a[3] ));
 sg13g2_dfrbp_1 _10402_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net966),
    .D(_00346_),
    .Q_N(_00169_),
    .Q(\i_core.cpu.i_core.i_shift.a[4] ));
 sg13g2_dfrbp_1 _10403_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net965),
    .D(net2647),
    .Q_N(_00171_),
    .Q(\i_core.cpu.i_core.i_shift.a[5] ));
 sg13g2_dfrbp_1 _10404_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net964),
    .D(_00348_),
    .Q_N(_00173_),
    .Q(\i_core.cpu.i_core.i_shift.a[6] ));
 sg13g2_dfrbp_1 _10405_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net963),
    .D(_00349_),
    .Q_N(_00175_),
    .Q(\i_core.cpu.i_core.i_shift.a[7] ));
 sg13g2_dfrbp_1 _10406_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net962),
    .D(_00350_),
    .Q_N(_00177_),
    .Q(\i_core.cpu.i_core.i_shift.a[8] ));
 sg13g2_dfrbp_1 _10407_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net961),
    .D(net2633),
    .Q_N(_00179_),
    .Q(\i_core.cpu.i_core.i_shift.a[9] ));
 sg13g2_dfrbp_1 _10408_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net960),
    .D(_00352_),
    .Q_N(_00181_),
    .Q(\i_core.cpu.i_core.i_shift.a[10] ));
 sg13g2_dfrbp_1 _10409_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net959),
    .D(_00353_),
    .Q_N(_00183_),
    .Q(\i_core.cpu.i_core.i_shift.a[11] ));
 sg13g2_dfrbp_1 _10410_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net958),
    .D(_00354_),
    .Q_N(_00185_),
    .Q(\i_core.cpu.i_core.i_shift.a[12] ));
 sg13g2_dfrbp_1 _10411_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net957),
    .D(net2217),
    .Q_N(_00187_),
    .Q(\i_core.cpu.i_core.i_shift.a[13] ));
 sg13g2_dfrbp_1 _10412_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net956),
    .D(_00356_),
    .Q_N(_00189_),
    .Q(\i_core.cpu.i_core.i_shift.a[14] ));
 sg13g2_dfrbp_1 _10413_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net955),
    .D(_00357_),
    .Q_N(_00191_),
    .Q(\i_core.cpu.i_core.i_shift.a[15] ));
 sg13g2_dfrbp_1 _10414_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net954),
    .D(_00358_),
    .Q_N(_00192_),
    .Q(\i_core.cpu.i_core.i_shift.a[16] ));
 sg13g2_dfrbp_1 _10415_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net953),
    .D(net2146),
    .Q_N(_00190_),
    .Q(\i_core.cpu.i_core.i_shift.a[17] ));
 sg13g2_dfrbp_1 _10416_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net952),
    .D(net2150),
    .Q_N(_00188_),
    .Q(\i_core.cpu.i_core.i_shift.a[18] ));
 sg13g2_dfrbp_1 _10417_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net951),
    .D(_00361_),
    .Q_N(_00186_),
    .Q(\i_core.cpu.i_core.i_shift.a[19] ));
 sg13g2_dfrbp_1 _10418_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net950),
    .D(net2279),
    .Q_N(_00184_),
    .Q(\i_core.cpu.i_core.i_shift.a[20] ));
 sg13g2_dfrbp_1 _10419_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net949),
    .D(_00363_),
    .Q_N(_00182_),
    .Q(\i_core.cpu.i_core.i_shift.a[21] ));
 sg13g2_dfrbp_1 _10420_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net948),
    .D(net2272),
    .Q_N(_00180_),
    .Q(\i_core.cpu.i_core.i_shift.a[22] ));
 sg13g2_dfrbp_1 _10421_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net947),
    .D(net2274),
    .Q_N(_00178_),
    .Q(\i_core.cpu.i_core.i_shift.a[23] ));
 sg13g2_dfrbp_1 _10422_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net946),
    .D(_00366_),
    .Q_N(_00176_),
    .Q(\i_core.cpu.i_core.i_shift.a[24] ));
 sg13g2_dfrbp_1 _10423_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net945),
    .D(_00367_),
    .Q_N(_00174_),
    .Q(\i_core.cpu.i_core.i_shift.a[25] ));
 sg13g2_dfrbp_1 _10424_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net944),
    .D(net2300),
    .Q_N(_00172_),
    .Q(\i_core.cpu.i_core.i_shift.a[26] ));
 sg13g2_dfrbp_1 _10425_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net943),
    .D(net2378),
    .Q_N(_00170_),
    .Q(\i_core.cpu.i_core.i_shift.a[27] ));
 sg13g2_dfrbp_1 _10426_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net942),
    .D(_00370_),
    .Q_N(_00195_),
    .Q(\i_core.cpu.i_core.i_shift.a[30] ));
 sg13g2_dfrbp_1 _10427_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net941),
    .D(_00371_),
    .Q_N(_00197_),
    .Q(\i_core.cpu.i_core.i_shift.a[31] ));
 sg13g2_dfrbp_1 _10428_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net940),
    .D(net2439),
    .Q_N(_04299_),
    .Q(\i_core.cpu.instr_data[1][0] ));
 sg13g2_dfrbp_1 _10429_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net938),
    .D(net2342),
    .Q_N(_00100_),
    .Q(\i_core.cpu.instr_data[1][1] ));
 sg13g2_dfrbp_1 _10430_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net936),
    .D(net2159),
    .Q_N(_04298_),
    .Q(\i_core.cpu.instr_data[0][2] ));
 sg13g2_dfrbp_1 _10431_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net935),
    .D(net2113),
    .Q_N(_04297_),
    .Q(\i_core.cpu.instr_data[0][3] ));
 sg13g2_dfrbp_1 _10432_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net934),
    .D(net1932),
    .Q_N(_00103_),
    .Q(\i_core.cpu.instr_data[0][4] ));
 sg13g2_dfrbp_1 _10433_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net933),
    .D(net1942),
    .Q_N(_00107_),
    .Q(\i_core.cpu.instr_data[0][5] ));
 sg13g2_dfrbp_1 _10434_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net932),
    .D(net1913),
    .Q_N(_00111_),
    .Q(\i_core.cpu.instr_data[0][6] ));
 sg13g2_dfrbp_1 _10435_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net931),
    .D(net1940),
    .Q_N(_00127_),
    .Q(\i_core.cpu.instr_data[0][7] ));
 sg13g2_dfrbp_1 _10436_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net930),
    .D(net1934),
    .Q_N(_00131_),
    .Q(\i_core.cpu.instr_data[0][8] ));
 sg13g2_dfrbp_1 _10437_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net929),
    .D(net1949),
    .Q_N(_00135_),
    .Q(\i_core.cpu.instr_data[0][9] ));
 sg13g2_dfrbp_1 _10438_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net928),
    .D(net1962),
    .Q_N(_00139_),
    .Q(\i_core.cpu.instr_data[0][10] ));
 sg13g2_dfrbp_1 _10439_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net927),
    .D(net1900),
    .Q_N(_00147_),
    .Q(\i_core.cpu.instr_data[0][11] ));
 sg13g2_dfrbp_1 _10440_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net926),
    .D(net1911),
    .Q_N(_00143_),
    .Q(\i_core.cpu.instr_data[0][12] ));
 sg13g2_dfrbp_1 _10441_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net925),
    .D(net1951),
    .Q_N(_00115_),
    .Q(\i_core.cpu.instr_data[0][13] ));
 sg13g2_dfrbp_1 _10442_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net924),
    .D(net1923),
    .Q_N(_00119_),
    .Q(\i_core.cpu.instr_data[0][14] ));
 sg13g2_dfrbp_1 _10443_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net923),
    .D(net1955),
    .Q_N(_00123_),
    .Q(\i_core.cpu.instr_data[0][15] ));
 sg13g2_dfrbp_1 _10444_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net922),
    .D(net2319),
    .Q_N(_04296_),
    .Q(\i_core.cpu.instr_data[2][2] ));
 sg13g2_dfrbp_1 _10445_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net921),
    .D(net2350),
    .Q_N(_04295_),
    .Q(\i_core.cpu.instr_data[2][3] ));
 sg13g2_dfrbp_1 _10446_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net920),
    .D(net2013),
    .Q_N(_00105_),
    .Q(\i_core.cpu.instr_data[2][4] ));
 sg13g2_dfrbp_1 _10447_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net919),
    .D(net2109),
    .Q_N(_00109_),
    .Q(\i_core.cpu.instr_data[2][5] ));
 sg13g2_dfrbp_1 _10448_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net918),
    .D(net2022),
    .Q_N(_00113_),
    .Q(\i_core.cpu.instr_data[2][6] ));
 sg13g2_dfrbp_1 _10449_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net917),
    .D(net2050),
    .Q_N(_00129_),
    .Q(\i_core.cpu.instr_data[2][7] ));
 sg13g2_dfrbp_1 _10450_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net916),
    .D(net1868),
    .Q_N(_00133_),
    .Q(\i_core.cpu.instr_data[2][8] ));
 sg13g2_dfrbp_1 _10451_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net915),
    .D(net1856),
    .Q_N(_00137_),
    .Q(\i_core.cpu.instr_data[2][9] ));
 sg13g2_dfrbp_1 _10452_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net914),
    .D(net1850),
    .Q_N(_00141_),
    .Q(\i_core.cpu.instr_data[2][10] ));
 sg13g2_dfrbp_1 _10453_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net913),
    .D(net1870),
    .Q_N(_00149_),
    .Q(\i_core.cpu.instr_data[2][11] ));
 sg13g2_dfrbp_1 _10454_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net912),
    .D(net1846),
    .Q_N(_00145_),
    .Q(\i_core.cpu.instr_data[2][12] ));
 sg13g2_dfrbp_1 _10455_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net911),
    .D(net1829),
    .Q_N(_00117_),
    .Q(\i_core.cpu.instr_data[2][13] ));
 sg13g2_dfrbp_1 _10456_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net910),
    .D(net1877),
    .Q_N(_00121_),
    .Q(\i_core.cpu.instr_data[2][14] ));
 sg13g2_dfrbp_1 _10457_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net909),
    .D(net1844),
    .Q_N(_00125_),
    .Q(\i_core.cpu.instr_data[2][15] ));
 sg13g2_dfrbp_1 _10458_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net908),
    .D(net2373),
    .Q_N(_04294_),
    .Q(\i_core.cpu.instr_data[3][2] ));
 sg13g2_dfrbp_1 _10459_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net907),
    .D(net2289),
    .Q_N(_04293_),
    .Q(\i_core.cpu.instr_data[3][3] ));
 sg13g2_dfrbp_1 _10460_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net906),
    .D(net2074),
    .Q_N(_00106_),
    .Q(\i_core.cpu.instr_data[3][4] ));
 sg13g2_dfrbp_1 _10461_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net905),
    .D(net2018),
    .Q_N(_00110_),
    .Q(\i_core.cpu.instr_data[3][5] ));
 sg13g2_dfrbp_1 _10462_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net904),
    .D(net2080),
    .Q_N(_00114_),
    .Q(\i_core.cpu.instr_data[3][6] ));
 sg13g2_dfrbp_1 _10463_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net903),
    .D(net2020),
    .Q_N(_00130_),
    .Q(\i_core.cpu.instr_data[3][7] ));
 sg13g2_dfrbp_1 _10464_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net902),
    .D(net1864),
    .Q_N(_00134_),
    .Q(\i_core.cpu.instr_data[3][8] ));
 sg13g2_dfrbp_1 _10465_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net901),
    .D(net1866),
    .Q_N(_00138_),
    .Q(\i_core.cpu.instr_data[3][9] ));
 sg13g2_dfrbp_1 _10466_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net900),
    .D(net1854),
    .Q_N(_00142_),
    .Q(\i_core.cpu.instr_data[3][10] ));
 sg13g2_dfrbp_1 _10467_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net899),
    .D(net1858),
    .Q_N(_00150_),
    .Q(\i_core.cpu.instr_data[3][11] ));
 sg13g2_dfrbp_1 _10468_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net898),
    .D(net1886),
    .Q_N(_00146_),
    .Q(\i_core.cpu.instr_data[3][12] ));
 sg13g2_dfrbp_1 _10469_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net897),
    .D(net1834),
    .Q_N(_00118_),
    .Q(\i_core.cpu.instr_data[3][13] ));
 sg13g2_dfrbp_1 _10470_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net896),
    .D(net1840),
    .Q_N(_00122_),
    .Q(\i_core.cpu.instr_data[3][14] ));
 sg13g2_dfrbp_1 _10471_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net895),
    .D(net1884),
    .Q_N(_00126_),
    .Q(\i_core.cpu.instr_data[3][15] ));
 sg13g2_dfrbp_1 _10472_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net894),
    .D(net2002),
    .Q_N(_04292_),
    .Q(\i_spi.data[1] ));
 sg13g2_dfrbp_1 _10473_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net893),
    .D(net2040),
    .Q_N(_04291_),
    .Q(\i_spi.data[2] ));
 sg13g2_dfrbp_1 _10474_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net892),
    .D(net1998),
    .Q_N(_04290_),
    .Q(\i_spi.data[3] ));
 sg13g2_dfrbp_1 _10475_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net891),
    .D(net1953),
    .Q_N(_04289_),
    .Q(\i_spi.data[4] ));
 sg13g2_dfrbp_1 _10476_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net890),
    .D(_00420_),
    .Q_N(_04288_),
    .Q(\i_spi.data[5] ));
 sg13g2_dfrbp_1 _10477_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net889),
    .D(net1994),
    .Q_N(_04287_),
    .Q(\i_spi.data[6] ));
 sg13g2_dfrbp_1 _10478_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net888),
    .D(net1960),
    .Q_N(_04286_),
    .Q(\i_spi.data[7] ));
 sg13g2_dfrbp_1 _10479_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net887),
    .D(net2234),
    .Q_N(_04285_),
    .Q(\addr[0] ));
 sg13g2_dfrbp_1 _10480_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net886),
    .D(net2052),
    .Q_N(_04284_),
    .Q(\addr[1] ));
 sg13g2_dfrbp_1 _10481_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net885),
    .D(_00425_),
    .Q_N(_04283_),
    .Q(\addr[2] ));
 sg13g2_dfrbp_1 _10482_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net884),
    .D(_00426_),
    .Q_N(_04282_),
    .Q(\addr[3] ));
 sg13g2_dfrbp_1 _10483_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net883),
    .D(_00427_),
    .Q_N(_04281_),
    .Q(\addr[4] ));
 sg13g2_dfrbp_1 _10484_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net882),
    .D(_00428_),
    .Q_N(_04280_),
    .Q(\addr[5] ));
 sg13g2_dfrbp_1 _10485_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net881),
    .D(_00429_),
    .Q_N(_04279_),
    .Q(\addr[6] ));
 sg13g2_dfrbp_1 _10486_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net880),
    .D(_00430_),
    .Q_N(_04278_),
    .Q(\addr[7] ));
 sg13g2_dfrbp_1 _10487_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net879),
    .D(_00431_),
    .Q_N(_04277_),
    .Q(\addr[8] ));
 sg13g2_dfrbp_1 _10488_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net878),
    .D(_00432_),
    .Q_N(_04276_),
    .Q(\addr[9] ));
 sg13g2_dfrbp_1 _10489_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net877),
    .D(_00433_),
    .Q_N(_04275_),
    .Q(\addr[10] ));
 sg13g2_dfrbp_1 _10490_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net876),
    .D(_00434_),
    .Q_N(_04274_),
    .Q(\addr[11] ));
 sg13g2_dfrbp_1 _10491_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net875),
    .D(_00435_),
    .Q_N(_04273_),
    .Q(\addr[12] ));
 sg13g2_dfrbp_1 _10492_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net874),
    .D(_00436_),
    .Q_N(_04272_),
    .Q(\addr[13] ));
 sg13g2_dfrbp_1 _10493_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net873),
    .D(_00437_),
    .Q_N(_04271_),
    .Q(\addr[14] ));
 sg13g2_dfrbp_1 _10494_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net872),
    .D(net2231),
    .Q_N(_04270_),
    .Q(\addr[15] ));
 sg13g2_dfrbp_1 _10495_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net871),
    .D(_00439_),
    .Q_N(_04269_),
    .Q(\addr[16] ));
 sg13g2_dfrbp_1 _10496_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net870),
    .D(_00440_),
    .Q_N(_04268_),
    .Q(\addr[17] ));
 sg13g2_dfrbp_1 _10497_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net869),
    .D(_00441_),
    .Q_N(_04267_),
    .Q(\addr[18] ));
 sg13g2_dfrbp_1 _10498_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net868),
    .D(_00442_),
    .Q_N(_04266_),
    .Q(\addr[19] ));
 sg13g2_dfrbp_1 _10499_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net867),
    .D(_00443_),
    .Q_N(_04265_),
    .Q(\addr[20] ));
 sg13g2_dfrbp_1 _10500_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net866),
    .D(net2206),
    .Q_N(_04264_),
    .Q(\addr[21] ));
 sg13g2_dfrbp_1 _10501_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net865),
    .D(net2199),
    .Q_N(_04263_),
    .Q(\addr[22] ));
 sg13g2_dfrbp_1 _10502_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net864),
    .D(net2111),
    .Q_N(_00161_),
    .Q(\addr[23] ));
 sg13g2_dfrbp_1 _10503_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net863),
    .D(_00447_),
    .Q_N(_04262_),
    .Q(\addr[24] ));
 sg13g2_dfrbp_1 _10504_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net861),
    .D(_00448_),
    .Q_N(_04261_),
    .Q(\addr[25] ));
 sg13g2_dfrbp_1 _10505_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net859),
    .D(_00449_),
    .Q_N(_04260_),
    .Q(\addr[26] ));
 sg13g2_dfrbp_1 _10506_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net857),
    .D(_00450_),
    .Q_N(_04259_),
    .Q(\addr[27] ));
 sg13g2_dfrbp_1 _10507_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net855),
    .D(net2266),
    .Q_N(_04258_),
    .Q(\i_core.cpu.instr_data[1][2] ));
 sg13g2_dfrbp_1 _10508_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net854),
    .D(net2222),
    .Q_N(_04257_),
    .Q(\i_core.cpu.instr_data[1][3] ));
 sg13g2_dfrbp_1 _10509_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net853),
    .D(net2078),
    .Q_N(_00104_),
    .Q(\i_core.cpu.instr_data[1][4] ));
 sg13g2_dfrbp_1 _10510_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net852),
    .D(net2057),
    .Q_N(_00108_),
    .Q(\i_core.cpu.instr_data[1][5] ));
 sg13g2_dfrbp_1 _10511_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net851),
    .D(net2118),
    .Q_N(_00112_),
    .Q(\i_core.cpu.instr_data[1][6] ));
 sg13g2_dfrbp_1 _10512_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net850),
    .D(net2076),
    .Q_N(_00128_),
    .Q(\i_core.cpu.instr_data[1][7] ));
 sg13g2_dfrbp_1 _10513_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net849),
    .D(net1838),
    .Q_N(_00132_),
    .Q(\i_core.cpu.instr_data[1][8] ));
 sg13g2_dfrbp_1 _10514_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net848),
    .D(net1852),
    .Q_N(_00136_),
    .Q(\i_core.cpu.instr_data[1][9] ));
 sg13g2_dfrbp_1 _10515_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net847),
    .D(net1860),
    .Q_N(_00140_),
    .Q(\i_core.cpu.instr_data[1][10] ));
 sg13g2_dfrbp_1 _10516_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net846),
    .D(net1879),
    .Q_N(_00148_),
    .Q(\i_core.cpu.instr_data[1][11] ));
 sg13g2_dfrbp_1 _10517_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net845),
    .D(net1848),
    .Q_N(_00144_),
    .Q(\i_core.cpu.instr_data[1][12] ));
 sg13g2_dfrbp_1 _10518_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net844),
    .D(net1836),
    .Q_N(_00116_),
    .Q(\i_core.cpu.instr_data[1][13] ));
 sg13g2_dfrbp_1 _10519_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net843),
    .D(net1842),
    .Q_N(_00120_),
    .Q(\i_core.cpu.instr_data[1][14] ));
 sg13g2_dfrbp_1 _10520_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net842),
    .D(net1862),
    .Q_N(_00124_),
    .Q(\i_core.cpu.instr_data[1][15] ));
 sg13g2_dfrbp_1 _10521_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net840),
    .D(net2336),
    .Q_N(_04256_),
    .Q(\i_core.cpu.i_core.mepc[0] ));
 sg13g2_dfrbp_1 _10522_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net839),
    .D(net2347),
    .Q_N(_04255_),
    .Q(\i_core.cpu.i_core.mepc[1] ));
 sg13g2_dfrbp_1 _10523_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net838),
    .D(_00467_),
    .Q_N(_04254_),
    .Q(\i_core.cpu.i_core.mepc[2] ));
 sg13g2_dfrbp_1 _10524_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net837),
    .D(net2353),
    .Q_N(_04253_),
    .Q(\i_core.cpu.i_core.mepc[3] ));
 sg13g2_dfrbp_1 _10525_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net836),
    .D(net2229),
    .Q_N(_04252_),
    .Q(\i_core.cpu.i_core.mepc[4] ));
 sg13g2_dfrbp_1 _10526_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net835),
    .D(net2270),
    .Q_N(_04251_),
    .Q(\i_core.cpu.i_core.mepc[5] ));
 sg13g2_dfrbp_1 _10527_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net834),
    .D(net2356),
    .Q_N(_04250_),
    .Q(\i_core.cpu.i_core.mepc[6] ));
 sg13g2_dfrbp_1 _10528_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net833),
    .D(net2044),
    .Q_N(_04249_),
    .Q(\i_core.cpu.i_core.mepc[7] ));
 sg13g2_dfrbp_1 _10529_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net832),
    .D(net2152),
    .Q_N(_04248_),
    .Q(\i_core.cpu.i_core.mepc[8] ));
 sg13g2_dfrbp_1 _10530_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net831),
    .D(net2209),
    .Q_N(_04247_),
    .Q(\i_core.cpu.i_core.mepc[9] ));
 sg13g2_dfrbp_1 _10531_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net830),
    .D(net2261),
    .Q_N(_04246_),
    .Q(\i_core.cpu.i_core.mepc[10] ));
 sg13g2_dfrbp_1 _10532_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net829),
    .D(_00476_),
    .Q_N(_04245_),
    .Q(\i_core.cpu.i_core.mepc[11] ));
 sg13g2_dfrbp_1 _10533_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net828),
    .D(_00477_),
    .Q_N(_04244_),
    .Q(\i_core.cpu.i_core.mepc[12] ));
 sg13g2_dfrbp_1 _10534_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net827),
    .D(_00478_),
    .Q_N(_04243_),
    .Q(\i_core.cpu.i_core.mepc[13] ));
 sg13g2_dfrbp_1 _10535_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net826),
    .D(net2167),
    .Q_N(_04242_),
    .Q(\i_core.cpu.i_core.mepc[14] ));
 sg13g2_dfrbp_1 _10536_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net825),
    .D(_00480_),
    .Q_N(_04241_),
    .Q(\i_core.cpu.i_core.mepc[15] ));
 sg13g2_dfrbp_1 _10537_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net824),
    .D(net2174),
    .Q_N(_04240_),
    .Q(\i_core.cpu.i_core.mepc[16] ));
 sg13g2_dfrbp_1 _10538_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net823),
    .D(net2236),
    .Q_N(_04239_),
    .Q(\i_core.cpu.i_core.mepc[17] ));
 sg13g2_dfrbp_1 _10539_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net822),
    .D(_00483_),
    .Q_N(_04238_),
    .Q(\i_core.cpu.i_core.mepc[18] ));
 sg13g2_dfrbp_1 _10540_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net821),
    .D(net2127),
    .Q_N(_04237_),
    .Q(\i_core.cpu.i_core.mepc[19] ));
 sg13g2_dfrbp_1 _10541_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net820),
    .D(_00485_),
    .Q_N(_04236_),
    .Q(\i_core.cpu.i_core.i_shift.adjusted_shift_amt[0] ));
 sg13g2_dfrbp_1 _10542_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net819),
    .D(_00486_),
    .Q_N(_04235_),
    .Q(\i_core.cpu.i_core.i_shift.adjusted_shift_amt[1] ));
 sg13g2_dfrbp_1 _10543_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net818),
    .D(_00487_),
    .Q_N(_04234_),
    .Q(\i_core.cpu.i_core.i_shift.b[2] ));
 sg13g2_dfrbp_1 _10544_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net708),
    .D(_00488_),
    .Q_N(_04843_),
    .Q(\i_core.cpu.i_core.i_shift.b[3] ));
 sg13g2_dfrbp_1 _10545_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net709),
    .D(_00016_),
    .Q_N(_04844_),
    .Q(\i_core.cpu.i_core.multiplier.accum[0] ));
 sg13g2_dfrbp_1 _10546_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net710),
    .D(_00019_),
    .Q_N(_00200_),
    .Q(\i_core.cpu.i_core.multiplier.accum[1] ));
 sg13g2_dfrbp_1 _10547_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net711),
    .D(_00020_),
    .Q_N(_04845_),
    .Q(\i_core.cpu.i_core.multiplier.accum[2] ));
 sg13g2_dfrbp_1 _10548_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net712),
    .D(_00021_),
    .Q_N(_04846_),
    .Q(\i_core.cpu.i_core.multiplier.accum[3] ));
 sg13g2_dfrbp_1 _10549_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net713),
    .D(_00022_),
    .Q_N(_04847_),
    .Q(\i_core.cpu.i_core.multiplier.accum[4] ));
 sg13g2_dfrbp_1 _10550_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net714),
    .D(_00023_),
    .Q_N(_04848_),
    .Q(\i_core.cpu.i_core.multiplier.accum[5] ));
 sg13g2_dfrbp_1 _10551_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net715),
    .D(_00024_),
    .Q_N(_04849_),
    .Q(\i_core.cpu.i_core.multiplier.accum[6] ));
 sg13g2_dfrbp_1 _10552_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net716),
    .D(_00025_),
    .Q_N(_04850_),
    .Q(\i_core.cpu.i_core.multiplier.accum[7] ));
 sg13g2_dfrbp_1 _10553_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net717),
    .D(_00026_),
    .Q_N(_04851_),
    .Q(\i_core.cpu.i_core.multiplier.accum[8] ));
 sg13g2_dfrbp_1 _10554_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net718),
    .D(_00027_),
    .Q_N(_04852_),
    .Q(\i_core.cpu.i_core.multiplier.accum[9] ));
 sg13g2_dfrbp_1 _10555_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net723),
    .D(_00017_),
    .Q_N(_04853_),
    .Q(\i_core.cpu.i_core.multiplier.accum[10] ));
 sg13g2_dfrbp_1 _10556_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net817),
    .D(_00018_),
    .Q_N(_04233_),
    .Q(\i_core.cpu.i_core.multiplier.accum[11] ));
 sg13g2_dfrbp_1 _10557_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net816),
    .D(net2452),
    .Q_N(_04232_),
    .Q(\i_core.cpu.instr_data[0][0] ));
 sg13g2_dfrbp_1 _10558_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net814),
    .D(net2404),
    .Q_N(_00099_),
    .Q(\i_core.cpu.instr_data[0][1] ));
 sg13g2_dfrbp_1 _10559_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net812),
    .D(_00491_),
    .Q_N(_04231_),
    .Q(debug_register_data));
 sg13g2_dfrbp_1 _10560_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net841),
    .D(net2238),
    .Q_N(_04854_),
    .Q(\i_core.mem.data_stall ));
 sg13g2_dfrbp_1 _10561_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net811),
    .D(net2506),
    .Q_N(_00151_),
    .Q(\i_core.mem.qspi_write_done ));
 sg13g2_dfrbp_1 _10562_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net809),
    .D(_00493_),
    .Q_N(_04230_),
    .Q(\i_core.cpu.i_core.multiplier.accum[12] ));
 sg13g2_dfrbp_1 _10563_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net808),
    .D(_00494_),
    .Q_N(_04229_),
    .Q(\i_core.cpu.i_core.multiplier.accum[13] ));
 sg13g2_dfrbp_1 _10564_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net807),
    .D(_00495_),
    .Q_N(_04228_),
    .Q(\i_core.cpu.i_core.multiplier.accum[14] ));
 sg13g2_dfrbp_1 _10565_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net806),
    .D(_00496_),
    .Q_N(_04227_),
    .Q(\i_core.cpu.i_core.multiplier.accum[15] ));
 sg13g2_dfrbp_1 _10566_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net805),
    .D(_00497_),
    .Q_N(_00157_),
    .Q(\i_core.mem.qspi_data_byte_idx[0] ));
 sg13g2_dfrbp_1 _10567_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net803),
    .D(_00498_),
    .Q_N(_04226_),
    .Q(\i_core.mem.qspi_data_byte_idx[1] ));
 sg13g2_dfrbp_1 _10568_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net801),
    .D(_00499_),
    .Q_N(_04225_),
    .Q(\i_core.cpu.instr_data_in[0] ));
 sg13g2_dfrbp_1 _10569_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net800),
    .D(_00500_),
    .Q_N(_04224_),
    .Q(\i_core.cpu.instr_data_in[1] ));
 sg13g2_dfrbp_1 _10570_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net799),
    .D(net2627),
    .Q_N(_04223_),
    .Q(\i_core.cpu.instr_data_in[2] ));
 sg13g2_dfrbp_1 _10571_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net798),
    .D(_00502_),
    .Q_N(_04222_),
    .Q(\i_core.cpu.instr_data_in[3] ));
 sg13g2_dfrbp_1 _10572_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net797),
    .D(_00503_),
    .Q_N(_04221_),
    .Q(\i_core.cpu.instr_data_in[4] ));
 sg13g2_dfrbp_1 _10573_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net796),
    .D(net2291),
    .Q_N(_04220_),
    .Q(\i_core.cpu.instr_data_in[5] ));
 sg13g2_dfrbp_1 _10574_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net795),
    .D(net2412),
    .Q_N(_04219_),
    .Q(\i_core.cpu.instr_data_in[6] ));
 sg13g2_dfrbp_1 _10575_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net794),
    .D(net2463),
    .Q_N(_04218_),
    .Q(\i_core.cpu.instr_data_in[7] ));
 sg13g2_dfrbp_1 _10576_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net793),
    .D(net2086),
    .Q_N(_04217_),
    .Q(\i_core.mem.qspi_data_buf[8] ));
 sg13g2_dfrbp_1 _10577_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net792),
    .D(net2100),
    .Q_N(_04216_),
    .Q(\i_core.mem.qspi_data_buf[9] ));
 sg13g2_dfrbp_1 _10578_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net791),
    .D(_00509_),
    .Q_N(_04215_),
    .Q(\i_core.mem.qspi_data_buf[10] ));
 sg13g2_dfrbp_1 _10579_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net790),
    .D(_00510_),
    .Q_N(_04214_),
    .Q(\i_core.mem.qspi_data_buf[11] ));
 sg13g2_dfrbp_1 _10580_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net789),
    .D(_00511_),
    .Q_N(_04213_),
    .Q(\i_core.mem.qspi_data_buf[12] ));
 sg13g2_dfrbp_1 _10581_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net788),
    .D(_00512_),
    .Q_N(_04212_),
    .Q(\i_core.mem.qspi_data_buf[13] ));
 sg13g2_dfrbp_1 _10582_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net787),
    .D(net2054),
    .Q_N(_04211_),
    .Q(\i_core.mem.qspi_data_buf[14] ));
 sg13g2_dfrbp_1 _10583_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net786),
    .D(_00514_),
    .Q_N(_04210_),
    .Q(\i_core.mem.qspi_data_buf[15] ));
 sg13g2_dfrbp_1 _10584_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net785),
    .D(net1889),
    .Q_N(_04209_),
    .Q(\i_core.mem.data_from_read[16] ));
 sg13g2_dfrbp_1 _10585_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net784),
    .D(net1919),
    .Q_N(_04208_),
    .Q(\i_core.mem.data_from_read[17] ));
 sg13g2_dfrbp_1 _10586_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net783),
    .D(net1894),
    .Q_N(_04207_),
    .Q(\i_core.mem.data_from_read[18] ));
 sg13g2_dfrbp_1 _10587_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net782),
    .D(net1896),
    .Q_N(_04206_),
    .Q(\i_core.mem.data_from_read[19] ));
 sg13g2_dfrbp_1 _10588_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net781),
    .D(net1972),
    .Q_N(_04205_),
    .Q(\i_core.mem.data_from_read[20] ));
 sg13g2_dfrbp_1 _10589_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net780),
    .D(net1905),
    .Q_N(_04204_),
    .Q(\i_core.mem.data_from_read[21] ));
 sg13g2_dfrbp_1 _10590_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net779),
    .D(net1908),
    .Q_N(_04203_),
    .Q(\i_core.mem.data_from_read[22] ));
 sg13g2_dfrbp_1 _10591_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net778),
    .D(net1892),
    .Q_N(_04202_),
    .Q(\i_core.mem.data_from_read[23] ));
 sg13g2_dfrbp_1 _10592_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net777),
    .D(_00523_),
    .Q_N(_04201_),
    .Q(\i_core.mem.qspi_data_buf[24] ));
 sg13g2_dfrbp_1 _10593_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net776),
    .D(_00524_),
    .Q_N(_04200_),
    .Q(\i_core.mem.qspi_data_buf[25] ));
 sg13g2_dfrbp_1 _10594_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net775),
    .D(_00525_),
    .Q_N(_04199_),
    .Q(\i_core.mem.qspi_data_buf[26] ));
 sg13g2_dfrbp_1 _10595_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net774),
    .D(_00526_),
    .Q_N(_04198_),
    .Q(\i_core.mem.qspi_data_buf[27] ));
 sg13g2_dfrbp_1 _10596_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net773),
    .D(_00527_),
    .Q_N(_04197_),
    .Q(\i_core.mem.qspi_data_buf[28] ));
 sg13g2_dfrbp_1 _10597_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net772),
    .D(_00528_),
    .Q_N(_04196_),
    .Q(\i_core.mem.qspi_data_buf[29] ));
 sg13g2_dfrbp_1 _10598_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net771),
    .D(_00529_),
    .Q_N(_04195_),
    .Q(\i_core.mem.qspi_data_buf[30] ));
 sg13g2_dfrbp_1 _10599_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net770),
    .D(_00530_),
    .Q_N(_04194_),
    .Q(\i_core.mem.qspi_data_buf[31] ));
 sg13g2_dfrbp_1 _10600_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net769),
    .D(net2502),
    .Q_N(_04193_),
    .Q(\i_core.cpu.instr_fetch_started ));
 sg13g2_dfrbp_1 _10601_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net768),
    .D(_00532_),
    .Q_N(_00089_),
    .Q(\i_core.mem.instr_active ));
 sg13g2_dfrbp_1 _10602_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net766),
    .D(net2511),
    .Q_N(_00160_),
    .Q(\i_core.mem.q_ctrl.read_cycles_count[0] ));
 sg13g2_dfrbp_1 _10603_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net765),
    .D(_00534_),
    .Q_N(_04192_),
    .Q(\i_core.mem.q_ctrl.read_cycles_count[1] ));
 sg13g2_dfrbp_1 _10604_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net764),
    .D(_00535_),
    .Q_N(_04191_),
    .Q(\i_core.mem.q_ctrl.read_cycles_count[2] ));
 sg13g2_dfrbp_1 _10605_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net763),
    .D(_00536_),
    .Q_N(_04190_),
    .Q(\i_core.mem.q_ctrl.data_req ));
 sg13g2_dfrbp_1 _10606_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net762),
    .D(_00537_),
    .Q_N(_04189_),
    .Q(\i_core.mem.q_ctrl.nibbles_remaining[0] ));
 sg13g2_dfrbp_1 _10607_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net760),
    .D(_00538_),
    .Q_N(_04188_),
    .Q(\i_core.mem.q_ctrl.nibbles_remaining[1] ));
 sg13g2_dfrbp_1 _10608_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net758),
    .D(_00539_),
    .Q_N(_04187_),
    .Q(\i_core.mem.q_ctrl.nibbles_remaining[2] ));
 sg13g2_dfrbp_1 _10609_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net756),
    .D(_00540_),
    .Q_N(_00159_),
    .Q(\i_core.mem.q_ctrl.is_writing ));
 sg13g2_dfrbp_1 _10610_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net754),
    .D(_00541_),
    .Q_N(_04186_),
    .Q(\i_core.mem.q_ctrl.data_ready ));
 sg13g2_dfrbp_1 _10611_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net753),
    .D(_00542_),
    .Q_N(_00213_),
    .Q(\i_core.mem.q_ctrl.fsm_state[0] ));
 sg13g2_dfrbp_1 _10612_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net751),
    .D(_00543_),
    .Q_N(_04185_),
    .Q(\i_core.mem.q_ctrl.fsm_state[1] ));
 sg13g2_dfrbp_1 _10613_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net749),
    .D(_00544_),
    .Q_N(_00152_),
    .Q(\i_core.mem.q_ctrl.fsm_state[2] ));
 sg13g2_dfrbp_1 _10614_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net747),
    .D(_00545_),
    .Q_N(_04184_),
    .Q(\i_core.mem.q_ctrl.spi_ram_b_select ));
 sg13g2_dfrbp_1 _10615_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net745),
    .D(_00546_),
    .Q_N(_04183_),
    .Q(\i_core.mem.q_ctrl.spi_ram_a_select ));
 sg13g2_dfrbp_1 _10616_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net743),
    .D(net2541),
    .Q_N(_04182_),
    .Q(\i_core.mem.q_ctrl.spi_flash_select ));
 sg13g2_dfrbp_1 _10617_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net741),
    .D(_00548_),
    .Q_N(_00158_),
    .Q(\i_core.mem.q_ctrl.spi_clk_out ));
 sg13g2_dfrbp_1 _10618_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net739),
    .D(net2064),
    .Q_N(_04181_),
    .Q(\i_core.mem.q_ctrl.spi_data_oe[0] ));
 sg13g2_dfrbp_1 _10619_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net737),
    .D(_00550_),
    .Q_N(_00167_),
    .Q(\i_core.cpu.i_core.i_shift.a[28] ));
 sg13g2_dfrbp_1 _10620_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net735),
    .D(_00551_),
    .Q_N(_00193_),
    .Q(\i_core.cpu.i_core.i_shift.a[29] ));
 sg13g2_dfrbp_1 _10621_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net733),
    .D(_00552_),
    .Q_N(_04180_),
    .Q(\i_core.mem.q_ctrl.spi_in_buffer[0] ));
 sg13g2_dfrbp_1 _10622_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net732),
    .D(_00553_),
    .Q_N(_04179_),
    .Q(\i_core.mem.q_ctrl.spi_in_buffer[1] ));
 sg13g2_dfrbp_1 _10623_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net731),
    .D(_00554_),
    .Q_N(_04178_),
    .Q(\i_core.mem.q_ctrl.spi_in_buffer[2] ));
 sg13g2_dfrbp_1 _10624_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net730),
    .D(_00555_),
    .Q_N(_04177_),
    .Q(\i_core.mem.q_ctrl.spi_in_buffer[3] ));
 sg13g2_dfrbp_1 _10625_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net729),
    .D(net2031),
    .Q_N(_04176_),
    .Q(\i_core.mem.q_ctrl.spi_in_buffer[4] ));
 sg13g2_dfrbp_1 _10626_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net728),
    .D(net2000),
    .Q_N(_04175_),
    .Q(\i_core.mem.q_ctrl.spi_in_buffer[5] ));
 sg13g2_dfrbp_1 _10627_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net727),
    .D(net1958),
    .Q_N(_04174_),
    .Q(\i_core.mem.q_ctrl.spi_in_buffer[6] ));
 sg13g2_dfrbp_1 _10628_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net726),
    .D(net1996),
    .Q_N(_04173_),
    .Q(\i_core.mem.q_ctrl.spi_in_buffer[7] ));
 sg13g2_dfrbp_1 _10629_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net725),
    .D(_00560_),
    .Q_N(_00208_),
    .Q(\i_core.cpu.instr_data_in[8] ));
 sg13g2_dfrbp_1 _10630_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net724),
    .D(_00561_),
    .Q_N(_00209_),
    .Q(\i_core.cpu.instr_data_in[9] ));
 sg13g2_dfrbp_1 _10631_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net722),
    .D(_00562_),
    .Q_N(_00210_),
    .Q(\i_core.cpu.instr_data_in[10] ));
 sg13g2_dfrbp_1 _10632_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net721),
    .D(_00563_),
    .Q_N(_00211_),
    .Q(\i_core.cpu.instr_data_in[11] ));
 sg13g2_dfrbp_1 _10633_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net720),
    .D(net2470),
    .Q_N(_00205_),
    .Q(\i_core.cpu.instr_data_in[12] ));
 sg13g2_dfrbp_1 _10634_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net719),
    .D(net2375),
    .Q_N(_00206_),
    .Q(\i_core.cpu.instr_data_in[13] ));
 sg13g2_dfrbp_1 _10635_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net706),
    .D(_00566_),
    .Q_N(_00212_),
    .Q(\i_core.cpu.instr_data_in[14] ));
 sg13g2_dfrbp_1 _10636_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net705),
    .D(_00567_),
    .Q_N(_00207_),
    .Q(\i_core.cpu.instr_data_in[15] ));
 sg13g2_dfrbp_1 _10637_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net704),
    .D(_00568_),
    .Q_N(_04172_),
    .Q(\i_core.mem.q_ctrl.last_ram_b_sel ));
 sg13g2_dfrbp_1 _10638_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net703),
    .D(_00569_),
    .Q_N(_04171_),
    .Q(\i_core.mem.q_ctrl.last_ram_a_sel ));
 sg13g2_dfrbp_1 _10639_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net702),
    .D(_00570_),
    .Q_N(_04170_),
    .Q(\i_core.cpu.instr_fetch_stopped ));
 sg13g2_dfrbp_1 _10640_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net701),
    .D(net2499),
    .Q_N(_04169_),
    .Q(\i_core.cpu.instr_data[2][0] ));
 sg13g2_dfrbp_1 _10641_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net699),
    .D(net2308),
    .Q_N(_00101_),
    .Q(\i_core.cpu.instr_data[2][1] ));
 sg13g2_dfrbp_1 _10642_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net697),
    .D(_00573_),
    .Q_N(_04168_),
    .Q(\i_core.mem.q_ctrl.delay_cycles_cfg[0] ));
 sg13g2_dfrbp_1 _10643_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net696),
    .D(_00574_),
    .Q_N(_04167_),
    .Q(\i_core.mem.q_ctrl.delay_cycles_cfg[1] ));
 sg13g2_dfrbp_1 _10644_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net695),
    .D(_00575_),
    .Q_N(_04166_),
    .Q(\i_core.mem.q_ctrl.delay_cycles_cfg[2] ));
 sg13g2_dfrbp_1 _10645_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net694),
    .D(_00576_),
    .Q_N(_00087_),
    .Q(\i_core.cpu.instr_write_offset[1] ));
 sg13g2_dfrbp_1 _10646_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net693),
    .D(_00577_),
    .Q_N(_04165_),
    .Q(\i_core.cpu.instr_write_offset[2] ));
 sg13g2_dfrbp_1 _10647_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net692),
    .D(net2144),
    .Q_N(_04164_),
    .Q(\i_core.mem.q_ctrl.addr[1] ));
 sg13g2_dfrbp_1 _10648_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net690),
    .D(_00579_),
    .Q_N(_04163_),
    .Q(\i_core.mem.q_ctrl.addr[2] ));
 sg13g2_dfrbp_1 _10649_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net688),
    .D(_00580_),
    .Q_N(_04162_),
    .Q(\i_core.mem.q_ctrl.addr[3] ));
 sg13g2_dfrbp_1 _10650_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net686),
    .D(_00581_),
    .Q_N(_00097_),
    .Q(\i_core.cpu.pc[1] ));
 sg13g2_dfrbp_1 _10651_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net684),
    .D(_00582_),
    .Q_N(_00098_),
    .Q(\i_core.cpu.pc[2] ));
 sg13g2_dfrbp_1 _10652_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net682),
    .D(_00583_),
    .Q_N(_04161_),
    .Q(\i_core.cpu.instr_data_start[3] ));
 sg13g2_dfrbp_1 _10653_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net680),
    .D(_00584_),
    .Q_N(_00163_),
    .Q(\i_core.cpu.instr_data_start[4] ));
 sg13g2_dfrbp_1 _10654_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net678),
    .D(_00585_),
    .Q_N(_04160_),
    .Q(\i_core.cpu.instr_data_start[5] ));
 sg13g2_dfrbp_1 _10655_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net676),
    .D(_00586_),
    .Q_N(_04159_),
    .Q(\i_core.cpu.instr_data_start[6] ));
 sg13g2_dfrbp_1 _10656_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net674),
    .D(_00587_),
    .Q_N(_04158_),
    .Q(\i_core.cpu.instr_data_start[7] ));
 sg13g2_dfrbp_1 _10657_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net672),
    .D(net2652),
    .Q_N(_04157_),
    .Q(\i_core.cpu.instr_data_start[8] ));
 sg13g2_dfrbp_1 _10658_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net670),
    .D(_00589_),
    .Q_N(_04156_),
    .Q(\i_core.cpu.instr_data_start[9] ));
 sg13g2_dfrbp_1 _10659_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net668),
    .D(_00590_),
    .Q_N(_04155_),
    .Q(\i_core.cpu.instr_data_start[10] ));
 sg13g2_dfrbp_1 _10660_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net666),
    .D(_00591_),
    .Q_N(_00201_),
    .Q(\i_core.cpu.instr_data_start[11] ));
 sg13g2_dfrbp_1 _10661_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net664),
    .D(_00592_),
    .Q_N(_04154_),
    .Q(\i_core.cpu.instr_data_start[12] ));
 sg13g2_dfrbp_1 _10662_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net662),
    .D(_00593_),
    .Q_N(_04153_),
    .Q(\i_core.cpu.instr_data_start[13] ));
 sg13g2_dfrbp_1 _10663_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net660),
    .D(_00594_),
    .Q_N(_04152_),
    .Q(\i_core.cpu.instr_data_start[14] ));
 sg13g2_dfrbp_1 _10664_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net658),
    .D(_00595_),
    .Q_N(_04151_),
    .Q(\i_core.cpu.instr_data_start[15] ));
 sg13g2_dfrbp_1 _10665_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net656),
    .D(_00596_),
    .Q_N(_04150_),
    .Q(\i_core.cpu.instr_data_start[16] ));
 sg13g2_dfrbp_1 _10666_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net654),
    .D(_00597_),
    .Q_N(_04149_),
    .Q(\i_core.cpu.instr_data_start[17] ));
 sg13g2_dfrbp_1 _10667_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net652),
    .D(_00598_),
    .Q_N(_04148_),
    .Q(\i_core.cpu.instr_data_start[18] ));
 sg13g2_dfrbp_1 _10668_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net650),
    .D(_00599_),
    .Q_N(_00165_),
    .Q(\i_core.cpu.instr_data_start[19] ));
 sg13g2_dfrbp_1 _10669_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net648),
    .D(_00600_),
    .Q_N(_04147_),
    .Q(\i_core.cpu.instr_data_start[20] ));
 sg13g2_dfrbp_1 _10670_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net646),
    .D(_00601_),
    .Q_N(_04146_),
    .Q(\i_core.cpu.instr_data_start[21] ));
 sg13g2_dfrbp_1 _10671_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net644),
    .D(_00602_),
    .Q_N(_04145_),
    .Q(\i_core.cpu.instr_data_start[22] ));
 sg13g2_dfrbp_1 _10672_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net642),
    .D(_00603_),
    .Q_N(_00162_),
    .Q(\i_core.cpu.instr_data_start[23] ));
 sg13g2_dfrbp_1 _10673_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net640),
    .D(_00604_),
    .Q_N(_00088_),
    .Q(\i_core.cpu.instr_fetch_running ));
 sg13g2_dfrbp_1 _10674_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net638),
    .D(_00605_),
    .Q_N(_00090_),
    .Q(\i_core.cpu.was_early_branch ));
 sg13g2_dfrbp_1 _10675_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net636),
    .D(_00606_),
    .Q_N(_04144_),
    .Q(\i_core.cpu.data_write_n[0] ));
 sg13g2_dfrbp_1 _10676_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net634),
    .D(net2490),
    .Q_N(_04143_),
    .Q(\i_core.cpu.data_write_n[1] ));
 sg13g2_dfrbp_1 _10677_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net632),
    .D(net2492),
    .Q_N(_04142_),
    .Q(\i_core.cpu.data_read_n[0] ));
 sg13g2_dfrbp_1 _10678_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net968),
    .D(net2534),
    .Q_N(_04855_),
    .Q(\i_core.cpu.data_read_n[1] ));
 sg13g2_dfrbp_1 _10679_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net630),
    .D(net2427),
    .Q_N(_04141_),
    .Q(debug_data_continue));
 sg13g2_dfrbp_1 _10680_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net625),
    .D(_00610_),
    .Q_N(_00083_),
    .Q(\i_core.cpu.no_write_in_progress ));
 sg13g2_dfrbp_1 _10681_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net621),
    .D(net1921),
    .Q_N(_04140_),
    .Q(\i_core.cpu.load_started ));
 sg13g2_dfrbp_1 _10682_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net617),
    .D(_00612_),
    .Q_N(_04139_),
    .Q(\data_to_write[0] ));
 sg13g2_dfrbp_1 _10683_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net614),
    .D(_00613_),
    .Q_N(_04138_),
    .Q(\data_to_write[1] ));
 sg13g2_dfrbp_1 _10684_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net612),
    .D(_00614_),
    .Q_N(_04137_),
    .Q(\data_to_write[2] ));
 sg13g2_dfrbp_1 _10685_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net610),
    .D(_00615_),
    .Q_N(_04136_),
    .Q(\data_to_write[3] ));
 sg13g2_dfrbp_1 _10686_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net606),
    .D(_00616_),
    .Q_N(_04135_),
    .Q(\data_to_write[4] ));
 sg13g2_dfrbp_1 _10687_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net604),
    .D(_00617_),
    .Q_N(_04134_),
    .Q(\data_to_write[5] ));
 sg13g2_dfrbp_1 _10688_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net602),
    .D(_00618_),
    .Q_N(_04133_),
    .Q(\data_to_write[6] ));
 sg13g2_dfrbp_1 _10689_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net600),
    .D(_00619_),
    .Q_N(_00202_),
    .Q(\data_to_write[7] ));
 sg13g2_dfrbp_1 _10690_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net598),
    .D(_00620_),
    .Q_N(_04132_),
    .Q(\data_to_write[8] ));
 sg13g2_dfrbp_1 _10691_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net596),
    .D(_00621_),
    .Q_N(_04131_),
    .Q(\data_to_write[9] ));
 sg13g2_dfrbp_1 _10692_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net594),
    .D(_00622_),
    .Q_N(_04130_),
    .Q(\data_to_write[10] ));
 sg13g2_dfrbp_1 _10693_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net588),
    .D(_00623_),
    .Q_N(_04129_),
    .Q(\data_to_write[11] ));
 sg13g2_dfrbp_1 _10694_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net586),
    .D(_00624_),
    .Q_N(_04128_),
    .Q(\data_to_write[12] ));
 sg13g2_dfrbp_1 _10695_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net584),
    .D(_00625_),
    .Q_N(_04127_),
    .Q(\data_to_write[13] ));
 sg13g2_dfrbp_1 _10696_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net582),
    .D(_00626_),
    .Q_N(_04126_),
    .Q(\data_to_write[14] ));
 sg13g2_dfrbp_1 _10697_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net580),
    .D(_00627_),
    .Q_N(_04125_),
    .Q(\data_to_write[15] ));
 sg13g2_dfrbp_1 _10698_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net578),
    .D(_00628_),
    .Q_N(_04124_),
    .Q(\data_to_write[16] ));
 sg13g2_dfrbp_1 _10699_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net576),
    .D(_00629_),
    .Q_N(_04123_),
    .Q(\data_to_write[17] ));
 sg13g2_dfrbp_1 _10700_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net574),
    .D(_00630_),
    .Q_N(_04122_),
    .Q(\data_to_write[18] ));
 sg13g2_dfrbp_1 _10701_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net572),
    .D(_00631_),
    .Q_N(_04121_),
    .Q(\data_to_write[19] ));
 sg13g2_dfrbp_1 _10702_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net570),
    .D(_00632_),
    .Q_N(_04120_),
    .Q(\data_to_write[20] ));
 sg13g2_dfrbp_1 _10703_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net568),
    .D(_00633_),
    .Q_N(_04119_),
    .Q(\data_to_write[21] ));
 sg13g2_dfrbp_1 _10704_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net566),
    .D(_00634_),
    .Q_N(_04118_),
    .Q(\data_to_write[22] ));
 sg13g2_dfrbp_1 _10705_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net564),
    .D(_00635_),
    .Q_N(_04117_),
    .Q(\data_to_write[23] ));
 sg13g2_dfrbp_1 _10706_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net562),
    .D(_00636_),
    .Q_N(_04116_),
    .Q(\data_to_write[24] ));
 sg13g2_dfrbp_1 _10707_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net560),
    .D(_00637_),
    .Q_N(_04115_),
    .Q(\data_to_write[25] ));
 sg13g2_dfrbp_1 _10708_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net540),
    .D(_00638_),
    .Q_N(_04114_),
    .Q(\data_to_write[26] ));
 sg13g2_dfrbp_1 _10709_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net534),
    .D(_00639_),
    .Q_N(_04113_),
    .Q(\data_to_write[27] ));
 sg13g2_dfrbp_1 _10710_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net532),
    .D(_00640_),
    .Q_N(_04112_),
    .Q(\data_to_write[28] ));
 sg13g2_dfrbp_1 _10711_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net530),
    .D(_00641_),
    .Q_N(_04111_),
    .Q(\data_to_write[29] ));
 sg13g2_dfrbp_1 _10712_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net528),
    .D(_00642_),
    .Q_N(_04110_),
    .Q(\data_to_write[30] ));
 sg13g2_dfrbp_1 _10713_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net526),
    .D(_00643_),
    .Q_N(_04109_),
    .Q(\data_to_write[31] ));
 sg13g2_dfrbp_1 _10714_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net524),
    .D(_00644_),
    .Q_N(_00218_),
    .Q(\i_core.cpu.counter[2] ));
 sg13g2_dfrbp_1 _10715_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net522),
    .D(_00645_),
    .Q_N(_00092_),
    .Q(\i_core.cpu.counter[3] ));
 sg13g2_dfrbp_1 _10716_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net520),
    .D(_00646_),
    .Q_N(_00084_),
    .Q(\i_core.cpu.counter[4] ));
 sg13g2_dfrbp_1 _10717_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net499),
    .D(_00647_),
    .Q_N(_04108_),
    .Q(\i_core.cpu.data_ready_core ));
 sg13g2_dfrbp_1 _10718_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net494),
    .D(net2177),
    .Q_N(_04107_),
    .Q(\i_core.cpu.data_ready_latch ));
 sg13g2_dfrbp_1 _10719_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net492),
    .D(_00649_),
    .Q_N(_04106_),
    .Q(\i_core.cpu.is_load ));
 sg13g2_dfrbp_1 _10720_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net483),
    .D(_00650_),
    .Q_N(_04105_),
    .Q(\i_core.cpu.is_alu_imm ));
 sg13g2_dfrbp_1 _10721_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net479),
    .D(_00651_),
    .Q_N(_04104_),
    .Q(\i_core.cpu.is_auipc ));
 sg13g2_dfrbp_1 _10722_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net475),
    .D(_00652_),
    .Q_N(_04103_),
    .Q(\i_core.cpu.is_store ));
 sg13g2_dfrbp_1 _10723_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net471),
    .D(_00653_),
    .Q_N(_04102_),
    .Q(\i_core.cpu.is_alu_reg ));
 sg13g2_dfrbp_1 _10724_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net467),
    .D(_00654_),
    .Q_N(_04101_),
    .Q(\i_core.cpu.is_lui ));
 sg13g2_dfrbp_1 _10725_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net463),
    .D(_00655_),
    .Q_N(_04100_),
    .Q(\i_core.cpu.is_branch ));
 sg13g2_dfrbp_1 _10726_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net459),
    .D(_00656_),
    .Q_N(_04099_),
    .Q(\i_core.cpu.is_jalr ));
 sg13g2_dfrbp_1 _10727_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net455),
    .D(_00657_),
    .Q_N(_04098_),
    .Q(\i_core.cpu.is_jal ));
 sg13g2_dfrbp_1 _10728_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net451),
    .D(_00658_),
    .Q_N(_04097_),
    .Q(\i_core.cpu.is_system ));
 sg13g2_dfrbp_1 _10729_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net446),
    .D(_00659_),
    .Q_N(_04096_),
    .Q(\i_core.cpu.instr_len[1] ));
 sg13g2_dfrbp_1 _10730_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net439),
    .D(_00660_),
    .Q_N(_04095_),
    .Q(\i_core.cpu.instr_len[2] ));
 sg13g2_dfrbp_1 _10731_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net435),
    .D(_00661_),
    .Q_N(_04094_),
    .Q(\i_core.cpu.i_core.imm_lo[0] ));
 sg13g2_dfrbp_1 _10732_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net431),
    .D(_00662_),
    .Q_N(_04093_),
    .Q(\i_core.cpu.i_core.imm_lo[1] ));
 sg13g2_dfrbp_1 _10733_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net429),
    .D(_00663_),
    .Q_N(_04092_),
    .Q(\i_core.cpu.i_core.imm_lo[2] ));
 sg13g2_dfrbp_1 _10734_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net425),
    .D(_00664_),
    .Q_N(_04091_),
    .Q(\i_core.cpu.i_core.imm_lo[3] ));
 sg13g2_dfrbp_1 _10735_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net423),
    .D(_00665_),
    .Q_N(_04090_),
    .Q(\i_core.cpu.i_core.imm_lo[4] ));
 sg13g2_dfrbp_1 _10736_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net421),
    .D(_00666_),
    .Q_N(_04089_),
    .Q(\i_core.cpu.i_core.imm_lo[5] ));
 sg13g2_dfrbp_1 _10737_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net419),
    .D(_00667_),
    .Q_N(_04088_),
    .Q(\i_core.cpu.i_core.imm_lo[6] ));
 sg13g2_dfrbp_1 _10738_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net417),
    .D(_00668_),
    .Q_N(_04087_),
    .Q(\i_core.cpu.i_core.imm_lo[7] ));
 sg13g2_dfrbp_1 _10739_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net1035),
    .D(_00669_),
    .Q_N(_04086_),
    .Q(\i_core.cpu.i_core.imm_lo[8] ));
 sg13g2_dfrbp_1 _10740_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net1033),
    .D(_00670_),
    .Q_N(_04085_),
    .Q(\i_core.cpu.i_core.imm_lo[9] ));
 sg13g2_dfrbp_1 _10741_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net1031),
    .D(_00671_),
    .Q_N(_04084_),
    .Q(\i_core.cpu.i_core.imm_lo[10] ));
 sg13g2_dfrbp_1 _10742_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net1029),
    .D(_00672_),
    .Q_N(_04083_),
    .Q(\i_core.cpu.i_core.imm_lo[11] ));
 sg13g2_dfrbp_1 _10743_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net939),
    .D(_00673_),
    .Q_N(_04082_),
    .Q(\i_core.cpu.imm[12] ));
 sg13g2_dfrbp_1 _10744_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net937),
    .D(_00674_),
    .Q_N(_04081_),
    .Q(\i_core.cpu.imm[13] ));
 sg13g2_dfrbp_1 _10745_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net862),
    .D(_00675_),
    .Q_N(_04080_),
    .Q(\i_core.cpu.imm[14] ));
 sg13g2_dfrbp_1 _10746_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net860),
    .D(_00676_),
    .Q_N(_04079_),
    .Q(\i_core.cpu.imm[15] ));
 sg13g2_dfrbp_1 _10747_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net858),
    .D(_00677_),
    .Q_N(_04078_),
    .Q(\i_core.cpu.imm[16] ));
 sg13g2_dfrbp_1 _10748_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net856),
    .D(_00678_),
    .Q_N(_04077_),
    .Q(\i_core.cpu.imm[17] ));
 sg13g2_dfrbp_1 _10749_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net815),
    .D(_00679_),
    .Q_N(_04076_),
    .Q(\i_core.cpu.imm[18] ));
 sg13g2_dfrbp_1 _10750_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net813),
    .D(_00680_),
    .Q_N(_04075_),
    .Q(\i_core.cpu.imm[19] ));
 sg13g2_dfrbp_1 _10751_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net810),
    .D(_00681_),
    .Q_N(_04074_),
    .Q(\i_core.cpu.imm[20] ));
 sg13g2_dfrbp_1 _10752_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net804),
    .D(_00682_),
    .Q_N(_04073_),
    .Q(\i_core.cpu.imm[21] ));
 sg13g2_dfrbp_1 _10753_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net802),
    .D(_00683_),
    .Q_N(_04072_),
    .Q(\i_core.cpu.imm[22] ));
 sg13g2_dfrbp_1 _10754_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net767),
    .D(_00684_),
    .Q_N(_04071_),
    .Q(\i_core.cpu.imm[23] ));
 sg13g2_dfrbp_1 _10755_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net761),
    .D(_00685_),
    .Q_N(_04070_),
    .Q(\i_core.cpu.imm[24] ));
 sg13g2_dfrbp_1 _10756_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net759),
    .D(_00686_),
    .Q_N(_04069_),
    .Q(\i_core.cpu.imm[25] ));
 sg13g2_dfrbp_1 _10757_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net757),
    .D(_00687_),
    .Q_N(_04068_),
    .Q(\i_core.cpu.imm[26] ));
 sg13g2_dfrbp_1 _10758_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net755),
    .D(_00688_),
    .Q_N(_04067_),
    .Q(\i_core.cpu.imm[27] ));
 sg13g2_dfrbp_1 _10759_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net752),
    .D(_00689_),
    .Q_N(_04066_),
    .Q(\i_core.cpu.imm[28] ));
 sg13g2_dfrbp_1 _10760_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net750),
    .D(_00690_),
    .Q_N(_04065_),
    .Q(\i_core.cpu.imm[29] ));
 sg13g2_dfrbp_1 _10761_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net748),
    .D(_00691_),
    .Q_N(_04064_),
    .Q(\i_core.cpu.imm[30] ));
 sg13g2_dfrbp_1 _10762_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net746),
    .D(_00692_),
    .Q_N(_04063_),
    .Q(\i_core.cpu.imm[31] ));
 sg13g2_dfrbp_1 _10763_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net744),
    .D(_00693_),
    .Q_N(_04062_),
    .Q(\i_core.cpu.alu_op[0] ));
 sg13g2_dfrbp_1 _10764_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net742),
    .D(_00694_),
    .Q_N(_04061_),
    .Q(\i_core.cpu.alu_op[1] ));
 sg13g2_dfrbp_1 _10765_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net740),
    .D(_00695_),
    .Q_N(_00166_),
    .Q(\i_core.cpu.alu_op[2] ));
 sg13g2_dfrbp_1 _10766_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net738),
    .D(_00696_),
    .Q_N(_04060_),
    .Q(\i_core.cpu.alu_op[3] ));
 sg13g2_dfrbp_1 _10767_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net736),
    .D(_00697_),
    .Q_N(_04059_),
    .Q(\i_core.cpu.i_core.mem_op[0] ));
 sg13g2_dfrbp_1 _10768_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net734),
    .D(_00698_),
    .Q_N(_04058_),
    .Q(\i_core.cpu.i_core.mem_op[1] ));
 sg13g2_dfrbp_1 _10769_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net700),
    .D(_00699_),
    .Q_N(_04057_),
    .Q(\i_core.cpu.i_core.mem_op[2] ));
 sg13g2_dfrbp_1 _10770_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net698),
    .D(_00700_),
    .Q_N(_04056_),
    .Q(\i_core.cpu.i_core.i_registers.rs1[0] ));
 sg13g2_dfrbp_1 _10771_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net691),
    .D(_00701_),
    .Q_N(_04055_),
    .Q(\i_core.cpu.i_core.i_registers.rs1[1] ));
 sg13g2_dfrbp_1 _10772_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net689),
    .D(_00702_),
    .Q_N(_04054_),
    .Q(\i_core.cpu.i_core.i_registers.rs1[2] ));
 sg13g2_dfrbp_1 _10773_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net687),
    .D(_00703_),
    .Q_N(_04053_),
    .Q(\i_core.cpu.i_core.i_registers.rs1[3] ));
 sg13g2_dfrbp_1 _10774_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net685),
    .D(_00704_),
    .Q_N(_04052_),
    .Q(\i_core.cpu.i_core.i_registers.rs2[0] ));
 sg13g2_dfrbp_1 _10775_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net683),
    .D(_00705_),
    .Q_N(_04051_),
    .Q(\i_core.cpu.i_core.i_registers.rs2[1] ));
 sg13g2_dfrbp_1 _10776_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net681),
    .D(_00706_),
    .Q_N(_04050_),
    .Q(\i_core.cpu.i_core.i_registers.rs2[2] ));
 sg13g2_dfrbp_1 _10777_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net679),
    .D(_00707_),
    .Q_N(_04049_),
    .Q(\i_core.cpu.i_core.i_registers.rs2[3] ));
 sg13g2_dfrbp_1 _10778_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net677),
    .D(_00708_),
    .Q_N(_00214_),
    .Q(\i_core.cpu.additional_mem_ops[0] ));
 sg13g2_dfrbp_1 _10779_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net673),
    .D(net2321),
    .Q_N(_04048_),
    .Q(\i_core.cpu.additional_mem_ops[1] ));
 sg13g2_dfrbp_1 _10780_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net669),
    .D(_00710_),
    .Q_N(_04047_),
    .Q(\i_core.cpu.additional_mem_ops[2] ));
 sg13g2_dfrbp_1 _10781_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net665),
    .D(_00711_),
    .Q_N(_04046_),
    .Q(\i_core.cpu.mem_op_increment_reg ));
 sg13g2_dfrbp_1 _10782_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net661),
    .D(_00712_),
    .Q_N(_00086_),
    .Q(\i_core.cpu.i_core.is_interrupt ));
 sg13g2_dfrbp_1 _10783_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net657),
    .D(_00713_),
    .Q_N(_00096_),
    .Q(debug_instr_valid));
 sg13g2_dfrbp_1 _10784_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net653),
    .D(_00714_),
    .Q_N(_04045_),
    .Q(\i_core.mem.q_ctrl.addr[0] ));
 sg13g2_dfrbp_1 _10785_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net649),
    .D(_00715_),
    .Q_N(_04044_),
    .Q(\i_core.cpu.instr_write_offset[3] ));
 sg13g2_dfrbp_1 _10786_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net647),
    .D(_00716_),
    .Q_N(_04043_),
    .Q(\i_core.mem.q_ctrl.addr[4] ));
 sg13g2_dfrbp_1 _10787_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net645),
    .D(net1930),
    .Q_N(_04042_),
    .Q(\i_core.mem.q_ctrl.addr[5] ));
 sg13g2_dfrbp_1 _10788_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net643),
    .D(net2062),
    .Q_N(_04041_),
    .Q(\i_core.mem.q_ctrl.addr[6] ));
 sg13g2_dfrbp_1 _10789_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net641),
    .D(net2034),
    .Q_N(_04040_),
    .Q(\i_core.mem.q_ctrl.addr[7] ));
 sg13g2_dfrbp_1 _10790_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net639),
    .D(_00720_),
    .Q_N(_04039_),
    .Q(\i_core.mem.q_ctrl.addr[8] ));
 sg13g2_dfrbp_1 _10791_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net637),
    .D(_00721_),
    .Q_N(_04038_),
    .Q(\i_core.mem.q_ctrl.addr[9] ));
 sg13g2_dfrbp_1 _10792_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net635),
    .D(_00722_),
    .Q_N(_04037_),
    .Q(\i_core.mem.q_ctrl.addr[10] ));
 sg13g2_dfrbp_1 _10793_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net633),
    .D(net2163),
    .Q_N(_04036_),
    .Q(\i_core.mem.q_ctrl.addr[11] ));
 sg13g2_dfrbp_1 _10794_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net631),
    .D(_00724_),
    .Q_N(_04035_),
    .Q(\i_core.mem.q_ctrl.addr[12] ));
 sg13g2_dfrbp_1 _10795_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net627),
    .D(net2070),
    .Q_N(_04034_),
    .Q(\i_core.mem.q_ctrl.addr[13] ));
 sg13g2_dfrbp_1 _10796_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net623),
    .D(_00726_),
    .Q_N(_04033_),
    .Q(\i_core.mem.q_ctrl.addr[14] ));
 sg13g2_dfrbp_1 _10797_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net619),
    .D(net2116),
    .Q_N(_04032_),
    .Q(\i_core.mem.q_ctrl.addr[15] ));
 sg13g2_dfrbp_1 _10798_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net496),
    .D(net2171),
    .Q_N(_04031_),
    .Q(\i_core.mem.q_ctrl.addr[16] ));
 sg13g2_dfrbp_1 _10799_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net490),
    .D(net2072),
    .Q_N(_04030_),
    .Q(\i_core.mem.q_ctrl.addr[17] ));
 sg13g2_dfrbp_1 _10800_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net481),
    .D(_00730_),
    .Q_N(_04029_),
    .Q(\i_core.mem.q_ctrl.addr[18] ));
 sg13g2_dfrbp_1 _10801_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net477),
    .D(net1977),
    .Q_N(_04028_),
    .Q(\i_core.mem.q_ctrl.addr[19] ));
 sg13g2_dfrbp_1 _10802_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net473),
    .D(_00732_),
    .Q_N(_04027_),
    .Q(\i_core.mem.q_ctrl.addr[20] ));
 sg13g2_dfrbp_1 _10803_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net469),
    .D(_00733_),
    .Q_N(_04026_),
    .Q(\i_core.mem.q_ctrl.addr[21] ));
 sg13g2_dfrbp_1 _10804_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net465),
    .D(_00734_),
    .Q_N(_04025_),
    .Q(\i_core.mem.q_ctrl.addr[22] ));
 sg13g2_dfrbp_1 _10805_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net969),
    .D(net2180),
    .Q_N(_04856_),
    .Q(\i_core.mem.q_ctrl.addr[23] ));
 sg13g2_dfrbp_1 _10806_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net970),
    .D(net1615),
    .Q_N(_00164_),
    .Q(\i_core.cpu.i_core.i_instrret.data[0] ));
 sg13g2_dfrbp_1 _10807_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net971),
    .D(net1559),
    .Q_N(_00199_),
    .Q(\i_core.cpu.i_core.i_instrret.data[1] ));
 sg13g2_dfrbp_1 _10808_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net972),
    .D(net1553),
    .Q_N(_04857_),
    .Q(\i_core.cpu.i_core.i_instrret.data[2] ));
 sg13g2_dfrbp_1 _10809_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net973),
    .D(net1529),
    .Q_N(_04858_),
    .Q(\i_core.cpu.i_core.i_instrret.data[3] ));
 sg13g2_dfrbp_1 _10810_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net974),
    .D(net1607),
    .Q_N(_04859_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10811_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net975),
    .D(net1735),
    .Q_N(_04860_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10812_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net976),
    .D(net1638),
    .Q_N(_04861_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10813_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net977),
    .D(net1621),
    .Q_N(_04862_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10814_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net978),
    .D(net1736),
    .Q_N(_04863_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10815_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net979),
    .D(net1688),
    .Q_N(_04864_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10816_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net980),
    .D(net1555),
    .Q_N(_04865_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10817_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net981),
    .D(net1623),
    .Q_N(_04866_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10818_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net982),
    .D(net1648),
    .Q_N(_04867_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10819_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net983),
    .D(net1079),
    .Q_N(_04868_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10820_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net984),
    .D(net1738),
    .Q_N(_04869_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10821_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net985),
    .D(net1620),
    .Q_N(_04870_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10822_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net986),
    .D(net1072),
    .Q_N(_04871_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10823_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net987),
    .D(net1649),
    .Q_N(_04872_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10824_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net988),
    .D(net1686),
    .Q_N(_04873_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10825_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net989),
    .D(net1577),
    .Q_N(_04874_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10826_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net990),
    .D(net1616),
    .Q_N(_04875_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10827_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net991),
    .D(net1728),
    .Q_N(_04876_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10828_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net992),
    .D(net1109),
    .Q_N(_04877_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10829_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net993),
    .D(net1609),
    .Q_N(_04878_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10830_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net994),
    .D(net1674),
    .Q_N(_04879_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10831_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net995),
    .D(net1677),
    .Q_N(_04880_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10832_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net1001),
    .D(net1752),
    .Q_N(_04881_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10833_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net461),
    .D(net1673),
    .Q_N(_04024_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10834_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net457),
    .D(net2525),
    .Q_N(_04023_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10835_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net453),
    .D(_00737_),
    .Q_N(_04022_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10836_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net448),
    .D(_00738_),
    .Q_N(_04021_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10837_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net441),
    .D(_00739_),
    .Q_N(_04020_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[31].A ));
 sg13g2_dfrbp_1 _10838_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net1002),
    .D(net2423),
    .Q_N(_00217_),
    .Q(\i_core.cpu.i_core.i_instrret.cy ));
 sg13g2_dfrbp_1 _10839_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net1003),
    .D(net1789),
    .Q_N(_04882_),
    .Q(\i_core.cpu.i_core.cycle_count[0] ));
 sg13g2_dfrbp_1 _10840_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net1004),
    .D(net1819),
    .Q_N(_04883_),
    .Q(\i_core.cpu.i_core.cycle_count[1] ));
 sg13g2_dfrbp_1 _10841_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1005),
    .D(net1817),
    .Q_N(_04884_),
    .Q(\i_core.cpu.i_core.cycle_count[2] ));
 sg13g2_dfrbp_1 _10842_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net1006),
    .D(net1692),
    .Q_N(_04885_),
    .Q(\i_core.cpu.i_core.cycle_count[3] ));
 sg13g2_dfrbp_1 _10843_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net1007),
    .D(net1092),
    .Q_N(_04886_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[4].A ));
 sg13g2_dfrbp_1 _10844_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net1008),
    .D(net1678),
    .Q_N(_04887_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[5].A ));
 sg13g2_dfrbp_1 _10845_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net1009),
    .D(net1665),
    .Q_N(_04888_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[6].A ));
 sg13g2_dfrbp_1 _10846_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net1010),
    .D(net1566),
    .Q_N(_04889_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[7].A ));
 sg13g2_dfrbp_1 _10847_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1011),
    .D(net1625),
    .Q_N(_04890_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[8].A ));
 sg13g2_dfrbp_1 _10848_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net1012),
    .D(net1089),
    .Q_N(_04891_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[9].A ));
 sg13g2_dfrbp_1 _10849_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1013),
    .D(net1596),
    .Q_N(_04892_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[10].A ));
 sg13g2_dfrbp_1 _10850_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net1014),
    .D(net1479),
    .Q_N(_04893_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[11].A ));
 sg13g2_dfrbp_1 _10851_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1015),
    .D(net1669),
    .Q_N(_04894_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[12].A ));
 sg13g2_dfrbp_1 _10852_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1016),
    .D(net1612),
    .Q_N(_04895_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[13].A ));
 sg13g2_dfrbp_1 _10853_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1017),
    .D(net1707),
    .Q_N(_04896_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[14].A ));
 sg13g2_dfrbp_1 _10854_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net1018),
    .D(net1622),
    .Q_N(_04897_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[15].A ));
 sg13g2_dfrbp_1 _10855_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1019),
    .D(net1633),
    .Q_N(_04898_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[16].A ));
 sg13g2_dfrbp_1 _10856_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1020),
    .D(net1618),
    .Q_N(_04899_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[17].A ));
 sg13g2_dfrbp_1 _10857_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1021),
    .D(net1617),
    .Q_N(_04900_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[18].A ));
 sg13g2_dfrbp_1 _10858_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net1022),
    .D(net1574),
    .Q_N(_04901_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[19].A ));
 sg13g2_dfrbp_1 _10859_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1023),
    .D(net1614),
    .Q_N(_04902_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[20].A ));
 sg13g2_dfrbp_1 _10860_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1024),
    .D(net1580),
    .Q_N(_04903_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[21].A ));
 sg13g2_dfrbp_1 _10861_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1025),
    .D(net1611),
    .Q_N(_04904_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[22].A ));
 sg13g2_dfrbp_1 _10862_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net1026),
    .D(net1511),
    .Q_N(_04905_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[23].A ));
 sg13g2_dfrbp_1 _10863_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1027),
    .D(net1734),
    .Q_N(_04906_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[24].A ));
 sg13g2_dfrbp_1 _10864_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net1028),
    .D(net1570),
    .Q_N(_04907_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[25].A ));
 sg13g2_dfrbp_1 _10865_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net651),
    .D(net1528),
    .Q_N(_04908_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[26].A ));
 sg13g2_dfrbp_1 _10866_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net437),
    .D(net1626),
    .Q_N(_04019_),
    .Q(\i_core.cpu.i_core.i_cycles.i_regbuf[27].A ));
 sg13g2_dfrbp_1 _10867_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net675),
    .D(_00741_),
    .Q_N(_04018_),
    .Q(\i_core.cpu.i_core.i_shift.b[4] ));
 sg13g2_dfrbp_1 _10868_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net671),
    .D(_00742_),
    .Q_N(_04017_),
    .Q(\i_core.cpu.i_core.i_cycles.cy ));
 sg13g2_dfrbp_1 _10869_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net667),
    .D(net2215),
    .Q_N(_04016_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[28].A ));
 sg13g2_dfrbp_1 _10870_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net663),
    .D(net1831),
    .Q_N(_04015_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[29].A ));
 sg13g2_dfrbp_1 _10871_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net659),
    .D(_00745_),
    .Q_N(_04014_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[30].A ));
 sg13g2_dfrbp_1 _10872_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net655),
    .D(_00746_),
    .Q_N(_04013_),
    .Q(\i_core.cpu.i_core.i_instrret.i_regbuf[31].A ));
 sg13g2_tiehi _09850__14 (.L_HI(net14));
 sg13g2_tiehi _09851__15 (.L_HI(net15));
 sg13g2_tiehi _09852__16 (.L_HI(net16));
 sg13g2_tiehi _09853__17 (.L_HI(net17));
 sg13g2_tiehi _09854__18 (.L_HI(net18));
 sg13g2_tiehi _09855__19 (.L_HI(net19));
 sg13g2_tiehi _09856__20 (.L_HI(net20));
 sg13g2_tiehi _09857__21 (.L_HI(net21));
 sg13g2_tiehi _09858__22 (.L_HI(net22));
 sg13g2_tiehi _09859__23 (.L_HI(net23));
 sg13g2_tiehi _09860__24 (.L_HI(net24));
 sg13g2_tiehi _09861__25 (.L_HI(net25));
 sg13g2_tiehi _09862__26 (.L_HI(net26));
 sg13g2_tiehi _09863__27 (.L_HI(net27));
 sg13g2_tiehi _09864__28 (.L_HI(net28));
 sg13g2_tiehi _09865__29 (.L_HI(net29));
 sg13g2_tiehi _09866__30 (.L_HI(net30));
 sg13g2_tiehi _09867__31 (.L_HI(net31));
 sg13g2_tiehi _09868__32 (.L_HI(net32));
 sg13g2_tiehi _09869__33 (.L_HI(net33));
 sg13g2_tiehi _09870__34 (.L_HI(net34));
 sg13g2_tiehi _09871__35 (.L_HI(net35));
 sg13g2_tiehi _09872__36 (.L_HI(net36));
 sg13g2_tiehi _09873__37 (.L_HI(net37));
 sg13g2_tiehi _09874__38 (.L_HI(net38));
 sg13g2_tiehi _09875__39 (.L_HI(net39));
 sg13g2_tiehi _09876__40 (.L_HI(net40));
 sg13g2_tiehi _09877__41 (.L_HI(net41));
 sg13g2_tiehi _09878__42 (.L_HI(net42));
 sg13g2_tiehi _09879__43 (.L_HI(net43));
 sg13g2_tiehi _09880__44 (.L_HI(net44));
 sg13g2_tiehi _09881__45 (.L_HI(net45));
 sg13g2_tiehi _09882__46 (.L_HI(net46));
 sg13g2_tiehi _09883__47 (.L_HI(net47));
 sg13g2_tiehi _09884__48 (.L_HI(net48));
 sg13g2_tiehi _09885__49 (.L_HI(net49));
 sg13g2_tiehi _09886__50 (.L_HI(net50));
 sg13g2_tiehi _09887__51 (.L_HI(net51));
 sg13g2_tiehi _09888__52 (.L_HI(net52));
 sg13g2_tiehi _09889__53 (.L_HI(net53));
 sg13g2_tiehi _09890__54 (.L_HI(net54));
 sg13g2_tiehi _09891__55 (.L_HI(net55));
 sg13g2_tiehi _09892__56 (.L_HI(net56));
 sg13g2_tiehi _09893__57 (.L_HI(net57));
 sg13g2_tiehi _09894__58 (.L_HI(net58));
 sg13g2_tiehi _09895__59 (.L_HI(net59));
 sg13g2_tiehi _09896__60 (.L_HI(net60));
 sg13g2_tiehi _09897__61 (.L_HI(net61));
 sg13g2_tiehi _09898__62 (.L_HI(net62));
 sg13g2_tiehi _09899__63 (.L_HI(net63));
 sg13g2_tiehi _09900__64 (.L_HI(net64));
 sg13g2_tiehi _09901__65 (.L_HI(net65));
 sg13g2_tiehi _09902__66 (.L_HI(net66));
 sg13g2_tiehi _09903__67 (.L_HI(net67));
 sg13g2_tiehi _09904__68 (.L_HI(net68));
 sg13g2_tiehi _09905__69 (.L_HI(net69));
 sg13g2_tiehi _09906__70 (.L_HI(net70));
 sg13g2_tiehi _09907__71 (.L_HI(net71));
 sg13g2_tiehi _09908__72 (.L_HI(net72));
 sg13g2_tiehi _09909__73 (.L_HI(net73));
 sg13g2_tiehi _09910__74 (.L_HI(net74));
 sg13g2_tiehi _09911__75 (.L_HI(net75));
 sg13g2_tiehi _09912__76 (.L_HI(net76));
 sg13g2_tiehi _09913__77 (.L_HI(net77));
 sg13g2_tiehi _09914__78 (.L_HI(net78));
 sg13g2_tiehi _09915__79 (.L_HI(net79));
 sg13g2_tiehi _09916__80 (.L_HI(net80));
 sg13g2_tiehi _09917__81 (.L_HI(net81));
 sg13g2_tiehi _09918__82 (.L_HI(net82));
 sg13g2_tiehi _09919__83 (.L_HI(net83));
 sg13g2_tiehi _09920__84 (.L_HI(net84));
 sg13g2_tiehi _09921__85 (.L_HI(net85));
 sg13g2_tiehi _09922__86 (.L_HI(net86));
 sg13g2_tiehi _09923__87 (.L_HI(net87));
 sg13g2_tiehi _09924__88 (.L_HI(net88));
 sg13g2_tiehi _09925__89 (.L_HI(net89));
 sg13g2_tiehi _09926__90 (.L_HI(net90));
 sg13g2_tiehi _09927__91 (.L_HI(net91));
 sg13g2_tiehi _09928__92 (.L_HI(net92));
 sg13g2_tiehi _09929__93 (.L_HI(net93));
 sg13g2_tiehi _09930__94 (.L_HI(net94));
 sg13g2_tiehi _09931__95 (.L_HI(net95));
 sg13g2_tiehi _09932__96 (.L_HI(net96));
 sg13g2_tiehi _09933__97 (.L_HI(net97));
 sg13g2_tiehi _09934__98 (.L_HI(net98));
 sg13g2_tiehi _09935__99 (.L_HI(net99));
 sg13g2_tiehi _09936__100 (.L_HI(net100));
 sg13g2_tiehi _09937__101 (.L_HI(net101));
 sg13g2_tiehi _09938__102 (.L_HI(net102));
 sg13g2_tiehi _09939__103 (.L_HI(net103));
 sg13g2_tiehi _09940__104 (.L_HI(net104));
 sg13g2_tiehi _09941__105 (.L_HI(net105));
 sg13g2_tiehi _09942__106 (.L_HI(net106));
 sg13g2_tiehi _09943__107 (.L_HI(net107));
 sg13g2_tiehi _09944__108 (.L_HI(net108));
 sg13g2_tiehi _09945__109 (.L_HI(net109));
 sg13g2_tiehi _09946__110 (.L_HI(net110));
 sg13g2_tiehi _09947__111 (.L_HI(net111));
 sg13g2_tiehi _09948__112 (.L_HI(net112));
 sg13g2_tiehi _09949__113 (.L_HI(net113));
 sg13g2_tiehi _09950__114 (.L_HI(net114));
 sg13g2_tiehi _09951__115 (.L_HI(net115));
 sg13g2_tiehi _09952__116 (.L_HI(net116));
 sg13g2_tiehi _09953__117 (.L_HI(net117));
 sg13g2_tiehi _09954__118 (.L_HI(net118));
 sg13g2_tiehi _09955__119 (.L_HI(net119));
 sg13g2_tiehi _09956__120 (.L_HI(net120));
 sg13g2_tiehi _09957__121 (.L_HI(net121));
 sg13g2_tiehi _09958__122 (.L_HI(net122));
 sg13g2_tiehi _09959__123 (.L_HI(net123));
 sg13g2_tiehi _09960__124 (.L_HI(net124));
 sg13g2_tiehi _09961__125 (.L_HI(net125));
 sg13g2_tiehi _09962__126 (.L_HI(net126));
 sg13g2_tiehi _09963__127 (.L_HI(net127));
 sg13g2_tiehi _09964__128 (.L_HI(net128));
 sg13g2_tiehi _09965__129 (.L_HI(net129));
 sg13g2_tiehi _09966__130 (.L_HI(net130));
 sg13g2_tiehi _09967__131 (.L_HI(net131));
 sg13g2_tiehi _09968__132 (.L_HI(net132));
 sg13g2_tiehi _09969__133 (.L_HI(net133));
 sg13g2_tiehi _09970__134 (.L_HI(net134));
 sg13g2_tiehi _09971__135 (.L_HI(net135));
 sg13g2_tiehi _09972__136 (.L_HI(net136));
 sg13g2_tiehi _09973__137 (.L_HI(net137));
 sg13g2_tiehi _09974__138 (.L_HI(net138));
 sg13g2_tiehi _09975__139 (.L_HI(net139));
 sg13g2_tiehi _09976__140 (.L_HI(net140));
 sg13g2_tiehi _09977__141 (.L_HI(net141));
 sg13g2_tiehi _09978__142 (.L_HI(net142));
 sg13g2_tiehi _09979__143 (.L_HI(net143));
 sg13g2_tiehi _09980__144 (.L_HI(net144));
 sg13g2_tiehi _09981__145 (.L_HI(net145));
 sg13g2_tiehi _09982__146 (.L_HI(net146));
 sg13g2_tiehi _09983__147 (.L_HI(net147));
 sg13g2_tiehi _09984__148 (.L_HI(net148));
 sg13g2_tiehi _09985__149 (.L_HI(net149));
 sg13g2_tiehi _09986__150 (.L_HI(net150));
 sg13g2_tiehi _09987__151 (.L_HI(net151));
 sg13g2_tiehi _09988__152 (.L_HI(net152));
 sg13g2_tiehi _09989__153 (.L_HI(net153));
 sg13g2_tiehi _09990__154 (.L_HI(net154));
 sg13g2_tiehi _09991__155 (.L_HI(net155));
 sg13g2_tiehi _09992__156 (.L_HI(net156));
 sg13g2_tiehi _09993__157 (.L_HI(net157));
 sg13g2_tiehi _09994__158 (.L_HI(net158));
 sg13g2_tiehi _09995__159 (.L_HI(net159));
 sg13g2_tiehi _09996__160 (.L_HI(net160));
 sg13g2_tiehi _09997__161 (.L_HI(net161));
 sg13g2_tiehi _09998__162 (.L_HI(net162));
 sg13g2_tiehi _09999__163 (.L_HI(net163));
 sg13g2_tiehi _10000__164 (.L_HI(net164));
 sg13g2_tiehi _10001__165 (.L_HI(net165));
 sg13g2_tiehi _10002__166 (.L_HI(net166));
 sg13g2_tiehi _10003__167 (.L_HI(net167));
 sg13g2_tiehi _10004__168 (.L_HI(net168));
 sg13g2_tiehi _10005__169 (.L_HI(net169));
 sg13g2_tiehi _10006__170 (.L_HI(net170));
 sg13g2_tiehi _10007__171 (.L_HI(net171));
 sg13g2_tiehi _10008__172 (.L_HI(net172));
 sg13g2_tiehi _10009__173 (.L_HI(net173));
 sg13g2_tiehi _10010__174 (.L_HI(net174));
 sg13g2_tiehi _10011__175 (.L_HI(net175));
 sg13g2_tiehi _10012__176 (.L_HI(net176));
 sg13g2_tiehi _10013__177 (.L_HI(net177));
 sg13g2_tiehi _10014__178 (.L_HI(net178));
 sg13g2_tiehi _10015__179 (.L_HI(net179));
 sg13g2_tiehi _10016__180 (.L_HI(net180));
 sg13g2_tiehi _10017__181 (.L_HI(net181));
 sg13g2_tiehi _10018__182 (.L_HI(net182));
 sg13g2_tiehi _10019__183 (.L_HI(net183));
 sg13g2_tiehi _10020__184 (.L_HI(net184));
 sg13g2_tiehi _10021__185 (.L_HI(net185));
 sg13g2_tiehi _10022__186 (.L_HI(net186));
 sg13g2_tiehi _10023__187 (.L_HI(net187));
 sg13g2_tiehi _10024__188 (.L_HI(net188));
 sg13g2_tiehi _10025__189 (.L_HI(net189));
 sg13g2_tiehi _10026__190 (.L_HI(net190));
 sg13g2_tiehi _10027__191 (.L_HI(net191));
 sg13g2_tiehi _10028__192 (.L_HI(net192));
 sg13g2_tiehi _10029__193 (.L_HI(net193));
 sg13g2_tiehi _10030__194 (.L_HI(net194));
 sg13g2_tiehi _10031__195 (.L_HI(net195));
 sg13g2_tiehi _10032__196 (.L_HI(net196));
 sg13g2_tiehi _10033__197 (.L_HI(net197));
 sg13g2_tiehi _10034__198 (.L_HI(net198));
 sg13g2_tiehi _10035__199 (.L_HI(net199));
 sg13g2_tiehi _10036__200 (.L_HI(net200));
 sg13g2_tiehi _10037__201 (.L_HI(net201));
 sg13g2_tiehi _10038__202 (.L_HI(net202));
 sg13g2_tiehi _10039__203 (.L_HI(net203));
 sg13g2_tiehi _10040__204 (.L_HI(net204));
 sg13g2_tiehi _10041__205 (.L_HI(net205));
 sg13g2_tiehi _10042__206 (.L_HI(net206));
 sg13g2_tiehi _10043__207 (.L_HI(net207));
 sg13g2_tiehi _10044__208 (.L_HI(net208));
 sg13g2_tiehi _10045__209 (.L_HI(net209));
 sg13g2_tiehi _10046__210 (.L_HI(net210));
 sg13g2_tiehi _10047__211 (.L_HI(net211));
 sg13g2_tiehi _10048__212 (.L_HI(net212));
 sg13g2_tiehi _10049__213 (.L_HI(net213));
 sg13g2_tiehi _10050__214 (.L_HI(net214));
 sg13g2_tiehi _10051__215 (.L_HI(net215));
 sg13g2_tiehi _10052__216 (.L_HI(net216));
 sg13g2_tiehi _10053__217 (.L_HI(net217));
 sg13g2_tiehi _10054__218 (.L_HI(net218));
 sg13g2_tiehi _10055__219 (.L_HI(net219));
 sg13g2_tiehi _10056__220 (.L_HI(net220));
 sg13g2_tiehi _10057__221 (.L_HI(net221));
 sg13g2_tiehi _10058__222 (.L_HI(net222));
 sg13g2_tiehi _10059__223 (.L_HI(net223));
 sg13g2_tiehi _10060__224 (.L_HI(net224));
 sg13g2_tiehi _10061__225 (.L_HI(net225));
 sg13g2_tiehi _10062__226 (.L_HI(net226));
 sg13g2_tiehi _10063__227 (.L_HI(net227));
 sg13g2_tiehi _10064__228 (.L_HI(net228));
 sg13g2_tiehi _10065__229 (.L_HI(net229));
 sg13g2_tiehi _10066__230 (.L_HI(net230));
 sg13g2_tiehi _10067__231 (.L_HI(net231));
 sg13g2_tiehi _10068__232 (.L_HI(net232));
 sg13g2_tiehi _10069__233 (.L_HI(net233));
 sg13g2_tiehi _10070__234 (.L_HI(net234));
 sg13g2_tiehi _10071__235 (.L_HI(net235));
 sg13g2_tiehi _10072__236 (.L_HI(net236));
 sg13g2_tiehi _10073__237 (.L_HI(net237));
 sg13g2_tiehi _10074__238 (.L_HI(net238));
 sg13g2_tiehi _10075__239 (.L_HI(net239));
 sg13g2_tiehi _10076__240 (.L_HI(net240));
 sg13g2_tiehi _10077__241 (.L_HI(net241));
 sg13g2_tiehi _10078__242 (.L_HI(net242));
 sg13g2_tiehi _10079__243 (.L_HI(net243));
 sg13g2_tiehi _10080__244 (.L_HI(net244));
 sg13g2_tiehi _10081__245 (.L_HI(net245));
 sg13g2_tiehi _10082__246 (.L_HI(net246));
 sg13g2_tiehi _10083__247 (.L_HI(net247));
 sg13g2_tiehi _10084__248 (.L_HI(net248));
 sg13g2_tiehi _10085__249 (.L_HI(net249));
 sg13g2_tiehi _10086__250 (.L_HI(net250));
 sg13g2_tiehi _10087__251 (.L_HI(net251));
 sg13g2_tiehi _10088__252 (.L_HI(net252));
 sg13g2_tiehi _10089__253 (.L_HI(net253));
 sg13g2_tiehi _10090__254 (.L_HI(net254));
 sg13g2_tiehi _10091__255 (.L_HI(net255));
 sg13g2_tiehi _10092__256 (.L_HI(net256));
 sg13g2_tiehi _10093__257 (.L_HI(net257));
 sg13g2_tiehi _10094__258 (.L_HI(net258));
 sg13g2_tiehi _10095__259 (.L_HI(net259));
 sg13g2_tiehi _10096__260 (.L_HI(net260));
 sg13g2_tiehi _10097__261 (.L_HI(net261));
 sg13g2_tiehi _10098__262 (.L_HI(net262));
 sg13g2_tiehi _10099__263 (.L_HI(net263));
 sg13g2_tiehi _10100__264 (.L_HI(net264));
 sg13g2_tiehi _10101__265 (.L_HI(net265));
 sg13g2_tiehi _10102__266 (.L_HI(net266));
 sg13g2_tiehi _10103__267 (.L_HI(net267));
 sg13g2_tiehi _10104__268 (.L_HI(net268));
 sg13g2_tiehi _10105__269 (.L_HI(net269));
 sg13g2_tiehi _10106__270 (.L_HI(net270));
 sg13g2_tiehi _10107__271 (.L_HI(net271));
 sg13g2_tiehi _10108__272 (.L_HI(net272));
 sg13g2_tiehi _10109__273 (.L_HI(net273));
 sg13g2_tiehi _10110__274 (.L_HI(net274));
 sg13g2_tiehi _10111__275 (.L_HI(net275));
 sg13g2_tiehi _10112__276 (.L_HI(net276));
 sg13g2_tiehi _10113__277 (.L_HI(net277));
 sg13g2_tiehi _10114__278 (.L_HI(net278));
 sg13g2_tiehi _10115__279 (.L_HI(net279));
 sg13g2_tiehi _10116__280 (.L_HI(net280));
 sg13g2_tiehi _10117__281 (.L_HI(net281));
 sg13g2_tiehi _10118__282 (.L_HI(net282));
 sg13g2_tiehi _10119__283 (.L_HI(net283));
 sg13g2_tiehi _10120__284 (.L_HI(net284));
 sg13g2_tiehi _10121__285 (.L_HI(net285));
 sg13g2_tiehi _10122__286 (.L_HI(net286));
 sg13g2_tiehi _10123__287 (.L_HI(net287));
 sg13g2_tiehi _10124__288 (.L_HI(net288));
 sg13g2_tiehi _10125__289 (.L_HI(net289));
 sg13g2_tiehi _10126__290 (.L_HI(net290));
 sg13g2_tiehi _10127__291 (.L_HI(net291));
 sg13g2_tiehi _10128__292 (.L_HI(net292));
 sg13g2_tiehi _10129__293 (.L_HI(net293));
 sg13g2_tiehi _10130__294 (.L_HI(net294));
 sg13g2_tiehi _10131__295 (.L_HI(net295));
 sg13g2_tiehi _10132__296 (.L_HI(net296));
 sg13g2_tiehi _10133__297 (.L_HI(net297));
 sg13g2_tiehi _10134__298 (.L_HI(net298));
 sg13g2_tiehi _10135__299 (.L_HI(net299));
 sg13g2_tiehi _10136__300 (.L_HI(net300));
 sg13g2_tiehi _10137__301 (.L_HI(net301));
 sg13g2_tiehi _10138__302 (.L_HI(net302));
 sg13g2_tiehi _10139__303 (.L_HI(net303));
 sg13g2_tiehi _10140__304 (.L_HI(net304));
 sg13g2_tiehi _10141__305 (.L_HI(net305));
 sg13g2_tiehi _10142__306 (.L_HI(net306));
 sg13g2_tiehi _10143__307 (.L_HI(net307));
 sg13g2_tiehi _10144__308 (.L_HI(net308));
 sg13g2_tiehi _10145__309 (.L_HI(net309));
 sg13g2_tiehi _10146__310 (.L_HI(net310));
 sg13g2_tiehi _10147__311 (.L_HI(net311));
 sg13g2_tiehi _10148__312 (.L_HI(net312));
 sg13g2_tiehi _10149__313 (.L_HI(net313));
 sg13g2_tiehi _10150__314 (.L_HI(net314));
 sg13g2_tiehi _10151__315 (.L_HI(net315));
 sg13g2_tiehi _10152__316 (.L_HI(net316));
 sg13g2_tiehi _10153__317 (.L_HI(net317));
 sg13g2_tiehi _10154__318 (.L_HI(net318));
 sg13g2_tiehi _10155__319 (.L_HI(net319));
 sg13g2_tiehi _10156__320 (.L_HI(net320));
 sg13g2_tiehi _10157__321 (.L_HI(net321));
 sg13g2_tiehi _10158__322 (.L_HI(net322));
 sg13g2_tiehi _10159__323 (.L_HI(net323));
 sg13g2_tiehi _10160__324 (.L_HI(net324));
 sg13g2_tiehi _10161__325 (.L_HI(net325));
 sg13g2_tiehi _10162__326 (.L_HI(net326));
 sg13g2_tiehi _10163__327 (.L_HI(net327));
 sg13g2_tiehi _10164__328 (.L_HI(net328));
 sg13g2_tiehi _10165__329 (.L_HI(net329));
 sg13g2_tiehi _10166__330 (.L_HI(net330));
 sg13g2_tiehi _10167__331 (.L_HI(net331));
 sg13g2_tiehi _10168__332 (.L_HI(net332));
 sg13g2_tiehi _10169__333 (.L_HI(net333));
 sg13g2_tiehi _10170__334 (.L_HI(net334));
 sg13g2_tiehi _10171__335 (.L_HI(net335));
 sg13g2_tiehi _10172__336 (.L_HI(net336));
 sg13g2_tiehi _10173__337 (.L_HI(net337));
 sg13g2_tiehi _10174__338 (.L_HI(net338));
 sg13g2_tiehi _10175__339 (.L_HI(net339));
 sg13g2_tiehi _10176__340 (.L_HI(net340));
 sg13g2_tiehi _10177__341 (.L_HI(net341));
 sg13g2_tiehi _10178__342 (.L_HI(net342));
 sg13g2_tiehi _10179__343 (.L_HI(net343));
 sg13g2_tiehi _10180__344 (.L_HI(net344));
 sg13g2_tiehi _10181__345 (.L_HI(net345));
 sg13g2_tiehi _10182__346 (.L_HI(net346));
 sg13g2_tiehi _10183__347 (.L_HI(net347));
 sg13g2_tiehi _10184__348 (.L_HI(net348));
 sg13g2_tiehi _10185__349 (.L_HI(net349));
 sg13g2_tiehi _10186__350 (.L_HI(net350));
 sg13g2_tiehi _10187__351 (.L_HI(net351));
 sg13g2_tiehi _10188__352 (.L_HI(net352));
 sg13g2_tiehi _10189__353 (.L_HI(net353));
 sg13g2_tiehi _10190__354 (.L_HI(net354));
 sg13g2_tiehi _10191__355 (.L_HI(net355));
 sg13g2_tiehi _10192__356 (.L_HI(net356));
 sg13g2_tiehi _10193__357 (.L_HI(net357));
 sg13g2_tiehi _10194__358 (.L_HI(net358));
 sg13g2_tiehi _10195__359 (.L_HI(net359));
 sg13g2_tiehi _10196__360 (.L_HI(net360));
 sg13g2_tiehi _10197__361 (.L_HI(net361));
 sg13g2_tiehi _10198__362 (.L_HI(net362));
 sg13g2_tiehi _10199__363 (.L_HI(net363));
 sg13g2_tiehi _10200__364 (.L_HI(net364));
 sg13g2_tiehi _10201__365 (.L_HI(net365));
 sg13g2_tiehi _10202__366 (.L_HI(net366));
 sg13g2_tiehi _10203__367 (.L_HI(net367));
 sg13g2_tiehi _10204__368 (.L_HI(net368));
 sg13g2_tiehi _10205__369 (.L_HI(net369));
 sg13g2_tiehi _10206__370 (.L_HI(net370));
 sg13g2_tiehi _10207__371 (.L_HI(net371));
 sg13g2_tiehi _10208__372 (.L_HI(net372));
 sg13g2_tiehi _10209__373 (.L_HI(net373));
 sg13g2_tiehi _10210__374 (.L_HI(net374));
 sg13g2_tiehi _10211__375 (.L_HI(net375));
 sg13g2_tiehi _10212__376 (.L_HI(net376));
 sg13g2_tiehi _10213__377 (.L_HI(net377));
 sg13g2_tiehi _10214__378 (.L_HI(net378));
 sg13g2_tiehi _10215__379 (.L_HI(net379));
 sg13g2_tiehi _10216__380 (.L_HI(net380));
 sg13g2_tiehi _10217__381 (.L_HI(net381));
 sg13g2_tiehi _10218__382 (.L_HI(net382));
 sg13g2_tiehi _10219__383 (.L_HI(net383));
 sg13g2_tiehi _10220__384 (.L_HI(net384));
 sg13g2_tiehi _10221__385 (.L_HI(net385));
 sg13g2_tiehi _10222__386 (.L_HI(net386));
 sg13g2_tiehi _10223__387 (.L_HI(net387));
 sg13g2_tiehi _10224__388 (.L_HI(net388));
 sg13g2_tiehi _10225__389 (.L_HI(net389));
 sg13g2_tiehi _10226__390 (.L_HI(net390));
 sg13g2_tiehi _10227__391 (.L_HI(net391));
 sg13g2_tiehi _10228__392 (.L_HI(net392));
 sg13g2_tiehi _10229__393 (.L_HI(net393));
 sg13g2_tiehi _10230__394 (.L_HI(net394));
 sg13g2_tiehi _10231__395 (.L_HI(net395));
 sg13g2_tiehi _10232__396 (.L_HI(net396));
 sg13g2_tiehi _10233__397 (.L_HI(net397));
 sg13g2_tiehi _10234__398 (.L_HI(net398));
 sg13g2_tiehi _10235__399 (.L_HI(net399));
 sg13g2_tiehi _10236__400 (.L_HI(net400));
 sg13g2_tiehi _10237__401 (.L_HI(net401));
 sg13g2_tiehi _10238__402 (.L_HI(net402));
 sg13g2_tiehi _10239__403 (.L_HI(net403));
 sg13g2_tiehi _10240__404 (.L_HI(net404));
 sg13g2_tiehi _10241__405 (.L_HI(net405));
 sg13g2_tiehi _10242__406 (.L_HI(net406));
 sg13g2_tiehi _10243__407 (.L_HI(net407));
 sg13g2_tiehi _10244__408 (.L_HI(net408));
 sg13g2_tiehi _10245__409 (.L_HI(net409));
 sg13g2_tiehi _10246__410 (.L_HI(net410));
 sg13g2_tiehi _10247__411 (.L_HI(net411));
 sg13g2_tiehi _10248__412 (.L_HI(net412));
 sg13g2_tiehi _10249__413 (.L_HI(net413));
 sg13g2_tiehi _10250__414 (.L_HI(net414));
 sg13g2_tiehi _10251__415 (.L_HI(net415));
 sg13g2_tiehi _10370__416 (.L_HI(net416));
 sg13g2_tiehi _10738__417 (.L_HI(net417));
 sg13g2_tiehi _10369__418 (.L_HI(net418));
 sg13g2_tiehi _10737__419 (.L_HI(net419));
 sg13g2_tiehi _10368__420 (.L_HI(net420));
 sg13g2_tiehi _10736__421 (.L_HI(net421));
 sg13g2_tiehi _10367__422 (.L_HI(net422));
 sg13g2_tiehi _10735__423 (.L_HI(net423));
 sg13g2_tiehi _10366__424 (.L_HI(net424));
 sg13g2_tiehi _10734__425 (.L_HI(net425));
 sg13g2_tiehi _10365__426 (.L_HI(net426));
 sg13g2_tiehi _10252__427 (.L_HI(net427));
 sg13g2_tiehi _10364__428 (.L_HI(net428));
 sg13g2_tiehi _10733__429 (.L_HI(net429));
 sg13g2_tiehi _10363__430 (.L_HI(net430));
 sg13g2_tiehi _10732__431 (.L_HI(net431));
 sg13g2_tiehi _10362__432 (.L_HI(net432));
 sg13g2_tiehi _10361__433 (.L_HI(net433));
 sg13g2_tiehi _10360__434 (.L_HI(net434));
 sg13g2_tiehi _10731__435 (.L_HI(net435));
 sg13g2_tiehi _10359__436 (.L_HI(net436));
 sg13g2_tiehi _10866__437 (.L_HI(net437));
 sg13g2_tiehi _10358__438 (.L_HI(net438));
 sg13g2_tiehi _10730__439 (.L_HI(net439));
 sg13g2_tiehi _10357__440 (.L_HI(net440));
 sg13g2_tiehi _10837__441 (.L_HI(net441));
 sg13g2_tiehi _10264__442 (.L_HI(net442));
 sg13g2_tiehi _10279__443 (.L_HI(net443));
 sg13g2_tiehi _10356__444 (.L_HI(net444));
 sg13g2_tiehi _10355__445 (.L_HI(net445));
 sg13g2_tiehi _10729__446 (.L_HI(net446));
 sg13g2_tiehi _10354__447 (.L_HI(net447));
 sg13g2_tiehi _10836__448 (.L_HI(net448));
 sg13g2_tiehi _10353__449 (.L_HI(net449));
 sg13g2_tiehi _10352__450 (.L_HI(net450));
 sg13g2_tiehi _10728__451 (.L_HI(net451));
 sg13g2_tiehi _10351__452 (.L_HI(net452));
 sg13g2_tiehi _10835__453 (.L_HI(net453));
 sg13g2_tiehi _10350__454 (.L_HI(net454));
 sg13g2_tiehi _10727__455 (.L_HI(net455));
 sg13g2_tiehi _10349__456 (.L_HI(net456));
 sg13g2_tiehi _10834__457 (.L_HI(net457));
 sg13g2_tiehi _10348__458 (.L_HI(net458));
 sg13g2_tiehi _10726__459 (.L_HI(net459));
 sg13g2_tiehi _10347__460 (.L_HI(net460));
 sg13g2_tiehi _10833__461 (.L_HI(net461));
 sg13g2_tiehi _10346__462 (.L_HI(net462));
 sg13g2_tiehi _10725__463 (.L_HI(net463));
 sg13g2_tiehi _10345__464 (.L_HI(net464));
 sg13g2_tiehi _10804__465 (.L_HI(net465));
 sg13g2_tiehi _10344__466 (.L_HI(net466));
 sg13g2_tiehi _10724__467 (.L_HI(net467));
 sg13g2_tiehi _10343__468 (.L_HI(net468));
 sg13g2_tiehi _10803__469 (.L_HI(net469));
 sg13g2_tiehi _10342__470 (.L_HI(net470));
 sg13g2_tiehi _10723__471 (.L_HI(net471));
 sg13g2_tiehi _10341__472 (.L_HI(net472));
 sg13g2_tiehi _10802__473 (.L_HI(net473));
 sg13g2_tiehi _10340__474 (.L_HI(net474));
 sg13g2_tiehi _10722__475 (.L_HI(net475));
 sg13g2_tiehi _10339__476 (.L_HI(net476));
 sg13g2_tiehi _10801__477 (.L_HI(net477));
 sg13g2_tiehi _10338__478 (.L_HI(net478));
 sg13g2_tiehi _10721__479 (.L_HI(net479));
 sg13g2_tiehi _10337__480 (.L_HI(net480));
 sg13g2_tiehi _10800__481 (.L_HI(net481));
 sg13g2_tiehi _10336__482 (.L_HI(net482));
 sg13g2_tiehi _10720__483 (.L_HI(net483));
 sg13g2_tiehi _10335__484 (.L_HI(net484));
 sg13g2_tiehi _10334__485 (.L_HI(net485));
 sg13g2_tiehi _10333__486 (.L_HI(net486));
 sg13g2_tiehi _10332__487 (.L_HI(net487));
 sg13g2_tiehi _10331__488 (.L_HI(net488));
 sg13g2_tiehi _10330__489 (.L_HI(net489));
 sg13g2_tiehi _10799__490 (.L_HI(net490));
 sg13g2_tiehi _10329__491 (.L_HI(net491));
 sg13g2_tiehi _10719__492 (.L_HI(net492));
 sg13g2_tiehi _10328__493 (.L_HI(net493));
 sg13g2_tiehi _10718__494 (.L_HI(net494));
 sg13g2_tiehi _10327__495 (.L_HI(net495));
 sg13g2_tiehi _10798__496 (.L_HI(net496));
 sg13g2_tiehi _10326__497 (.L_HI(net497));
 sg13g2_tiehi _10325__498 (.L_HI(net498));
 sg13g2_tiehi _10717__499 (.L_HI(net499));
 sg13g2_tiehi _10324__500 (.L_HI(net500));
 sg13g2_tiehi _10323__501 (.L_HI(net501));
 sg13g2_tiehi _10322__502 (.L_HI(net502));
 sg13g2_tiehi _10321__503 (.L_HI(net503));
 sg13g2_tiehi _10320__504 (.L_HI(net504));
 sg13g2_tiehi _10319__505 (.L_HI(net505));
 sg13g2_tiehi _10318__506 (.L_HI(net506));
 sg13g2_tiehi _10317__507 (.L_HI(net507));
 sg13g2_tiehi _10316__508 (.L_HI(net508));
 sg13g2_tiehi _10315__509 (.L_HI(net509));
 sg13g2_tiehi _10314__510 (.L_HI(net510));
 sg13g2_tiehi _10313__511 (.L_HI(net511));
 sg13g2_tiehi _10312__512 (.L_HI(net512));
 sg13g2_tiehi _10311__513 (.L_HI(net513));
 sg13g2_tiehi _10310__514 (.L_HI(net514));
 sg13g2_tiehi _10309__515 (.L_HI(net515));
 sg13g2_tiehi _10308__516 (.L_HI(net516));
 sg13g2_tiehi _10307__517 (.L_HI(net517));
 sg13g2_tiehi _10306__518 (.L_HI(net518));
 sg13g2_tiehi _10305__519 (.L_HI(net519));
 sg13g2_tiehi _10716__520 (.L_HI(net520));
 sg13g2_tiehi _10304__521 (.L_HI(net521));
 sg13g2_tiehi _10715__522 (.L_HI(net522));
 sg13g2_tiehi _10303__523 (.L_HI(net523));
 sg13g2_tiehi _10714__524 (.L_HI(net524));
 sg13g2_tiehi _10302__525 (.L_HI(net525));
 sg13g2_tiehi _10713__526 (.L_HI(net526));
 sg13g2_tiehi _10301__527 (.L_HI(net527));
 sg13g2_tiehi _10712__528 (.L_HI(net528));
 sg13g2_tiehi _10300__529 (.L_HI(net529));
 sg13g2_tiehi _10711__530 (.L_HI(net530));
 sg13g2_tiehi _10299__531 (.L_HI(net531));
 sg13g2_tiehi _10710__532 (.L_HI(net532));
 sg13g2_tiehi _10298__533 (.L_HI(net533));
 sg13g2_tiehi _10709__534 (.L_HI(net534));
 sg13g2_tiehi _10297__535 (.L_HI(net535));
 sg13g2_tiehi _10280__536 (.L_HI(net536));
 sg13g2_tiehi _10373__537 (.L_HI(net537));
 sg13g2_tiehi _10374__538 (.L_HI(net538));
 sg13g2_tiehi _10375__539 (.L_HI(net539));
 sg13g2_tiehi _10708__540 (.L_HI(net540));
 sg13g2_tiehi _10376__541 (.L_HI(net541));
 sg13g2_tiehi _10378__542 (.L_HI(net542));
 sg13g2_tiehi _10379__543 (.L_HI(net543));
 sg13g2_tiehi _10380__544 (.L_HI(net544));
 sg13g2_tiehi _10381__545 (.L_HI(net545));
 sg13g2_tiehi _10382__546 (.L_HI(net546));
 sg13g2_tiehi _10383__547 (.L_HI(net547));
 sg13g2_tiehi _10384__548 (.L_HI(net548));
 sg13g2_tiehi _10385__549 (.L_HI(net549));
 sg13g2_tiehi _10386__550 (.L_HI(net550));
 sg13g2_tiehi _10387__551 (.L_HI(net551));
 sg13g2_tiehi _10388__552 (.L_HI(net552));
 sg13g2_tiehi _10389__553 (.L_HI(net553));
 sg13g2_tiehi _10390__554 (.L_HI(net554));
 sg13g2_tiehi _10391__555 (.L_HI(net555));
 sg13g2_tiehi _10392__556 (.L_HI(net556));
 sg13g2_tiehi _10393__557 (.L_HI(net557));
 sg13g2_tiehi _10394__558 (.L_HI(net558));
 sg13g2_tiehi _10296__559 (.L_HI(net559));
 sg13g2_tiehi _10707__560 (.L_HI(net560));
 sg13g2_tiehi _10295__561 (.L_HI(net561));
 sg13g2_tiehi _10706__562 (.L_HI(net562));
 sg13g2_tiehi _10294__563 (.L_HI(net563));
 sg13g2_tiehi _10705__564 (.L_HI(net564));
 sg13g2_tiehi _10293__565 (.L_HI(net565));
 sg13g2_tiehi _10704__566 (.L_HI(net566));
 sg13g2_tiehi _10292__567 (.L_HI(net567));
 sg13g2_tiehi _10703__568 (.L_HI(net568));
 sg13g2_tiehi _10291__569 (.L_HI(net569));
 sg13g2_tiehi _10702__570 (.L_HI(net570));
 sg13g2_tiehi _10290__571 (.L_HI(net571));
 sg13g2_tiehi _10701__572 (.L_HI(net572));
 sg13g2_tiehi _10289__573 (.L_HI(net573));
 sg13g2_tiehi _10700__574 (.L_HI(net574));
 sg13g2_tiehi _10288__575 (.L_HI(net575));
 sg13g2_tiehi _10699__576 (.L_HI(net576));
 sg13g2_tiehi _10287__577 (.L_HI(net577));
 sg13g2_tiehi _10698__578 (.L_HI(net578));
 sg13g2_tiehi _10286__579 (.L_HI(net579));
 sg13g2_tiehi _10697__580 (.L_HI(net580));
 sg13g2_tiehi _10285__581 (.L_HI(net581));
 sg13g2_tiehi _10696__582 (.L_HI(net582));
 sg13g2_tiehi _10284__583 (.L_HI(net583));
 sg13g2_tiehi _10695__584 (.L_HI(net584));
 sg13g2_tiehi _10283__585 (.L_HI(net585));
 sg13g2_tiehi _10694__586 (.L_HI(net586));
 sg13g2_tiehi _10282__587 (.L_HI(net587));
 sg13g2_tiehi _10693__588 (.L_HI(net588));
 sg13g2_tiehi _10281__589 (.L_HI(net589));
 sg13g2_tiehi _10278__590 (.L_HI(net590));
 sg13g2_tiehi _10277__591 (.L_HI(net591));
 sg13g2_tiehi _10276__592 (.L_HI(net592));
 sg13g2_tiehi _10275__593 (.L_HI(net593));
 sg13g2_tiehi _10692__594 (.L_HI(net594));
 sg13g2_tiehi _10274__595 (.L_HI(net595));
 sg13g2_tiehi _10691__596 (.L_HI(net596));
 sg13g2_tiehi _10273__597 (.L_HI(net597));
 sg13g2_tiehi _10690__598 (.L_HI(net598));
 sg13g2_tiehi _10272__599 (.L_HI(net599));
 sg13g2_tiehi _10689__600 (.L_HI(net600));
 sg13g2_tiehi _10271__601 (.L_HI(net601));
 sg13g2_tiehi _10688__602 (.L_HI(net602));
 sg13g2_tiehi _10270__603 (.L_HI(net603));
 sg13g2_tiehi _10687__604 (.L_HI(net604));
 sg13g2_tiehi _10269__605 (.L_HI(net605));
 sg13g2_tiehi _10686__606 (.L_HI(net606));
 sg13g2_tiehi _10268__607 (.L_HI(net607));
 sg13g2_tiehi _10267__608 (.L_HI(net608));
 sg13g2_tiehi _10266__609 (.L_HI(net609));
 sg13g2_tiehi _10685__610 (.L_HI(net610));
 sg13g2_tiehi _10265__611 (.L_HI(net611));
 sg13g2_tiehi _10684__612 (.L_HI(net612));
 sg13g2_tiehi _10263__613 (.L_HI(net613));
 sg13g2_tiehi _10683__614 (.L_HI(net614));
 sg13g2_tiehi _10262__615 (.L_HI(net615));
 sg13g2_tiehi _10261__616 (.L_HI(net616));
 sg13g2_tiehi _10682__617 (.L_HI(net617));
 sg13g2_tiehi _10260__618 (.L_HI(net618));
 sg13g2_tiehi _10797__619 (.L_HI(net619));
 sg13g2_tiehi _10259__620 (.L_HI(net620));
 sg13g2_tiehi _10681__621 (.L_HI(net621));
 sg13g2_tiehi _10258__622 (.L_HI(net622));
 sg13g2_tiehi _10796__623 (.L_HI(net623));
 sg13g2_tiehi _10257__624 (.L_HI(net624));
 sg13g2_tiehi _10680__625 (.L_HI(net625));
 sg13g2_tiehi _10256__626 (.L_HI(net626));
 sg13g2_tiehi _10795__627 (.L_HI(net627));
 sg13g2_tiehi _10255__628 (.L_HI(net628));
 sg13g2_tiehi _10254__629 (.L_HI(net629));
 sg13g2_tiehi _10679__630 (.L_HI(net630));
 sg13g2_tiehi _10794__631 (.L_HI(net631));
 sg13g2_tiehi _10677__632 (.L_HI(net632));
 sg13g2_tiehi _10793__633 (.L_HI(net633));
 sg13g2_tiehi _10676__634 (.L_HI(net634));
 sg13g2_tiehi _10792__635 (.L_HI(net635));
 sg13g2_tiehi _10675__636 (.L_HI(net636));
 sg13g2_tiehi _10791__637 (.L_HI(net637));
 sg13g2_tiehi _10674__638 (.L_HI(net638));
 sg13g2_tiehi _10790__639 (.L_HI(net639));
 sg13g2_tiehi _10673__640 (.L_HI(net640));
 sg13g2_tiehi _10789__641 (.L_HI(net641));
 sg13g2_tiehi _10672__642 (.L_HI(net642));
 sg13g2_tiehi _10788__643 (.L_HI(net643));
 sg13g2_tiehi _10671__644 (.L_HI(net644));
 sg13g2_tiehi _10787__645 (.L_HI(net645));
 sg13g2_tiehi _10670__646 (.L_HI(net646));
 sg13g2_tiehi _10786__647 (.L_HI(net647));
 sg13g2_tiehi _10669__648 (.L_HI(net648));
 sg13g2_tiehi _10785__649 (.L_HI(net649));
 sg13g2_tiehi _10668__650 (.L_HI(net650));
 sg13g2_tiehi _10865__651 (.L_HI(net651));
 sg13g2_tiehi _10667__652 (.L_HI(net652));
 sg13g2_tiehi _10784__653 (.L_HI(net653));
 sg13g2_tiehi _10666__654 (.L_HI(net654));
 sg13g2_tiehi _10872__655 (.L_HI(net655));
 sg13g2_tiehi _10665__656 (.L_HI(net656));
 sg13g2_tiehi _10783__657 (.L_HI(net657));
 sg13g2_tiehi _10664__658 (.L_HI(net658));
 sg13g2_tiehi _10871__659 (.L_HI(net659));
 sg13g2_tiehi _10663__660 (.L_HI(net660));
 sg13g2_tiehi _10782__661 (.L_HI(net661));
 sg13g2_tiehi _10662__662 (.L_HI(net662));
 sg13g2_tiehi _10870__663 (.L_HI(net663));
 sg13g2_tiehi _10661__664 (.L_HI(net664));
 sg13g2_tiehi _10781__665 (.L_HI(net665));
 sg13g2_tiehi _10660__666 (.L_HI(net666));
 sg13g2_tiehi _10869__667 (.L_HI(net667));
 sg13g2_tiehi _10659__668 (.L_HI(net668));
 sg13g2_tiehi _10780__669 (.L_HI(net669));
 sg13g2_tiehi _10658__670 (.L_HI(net670));
 sg13g2_tiehi _10868__671 (.L_HI(net671));
 sg13g2_tiehi _10657__672 (.L_HI(net672));
 sg13g2_tiehi _10779__673 (.L_HI(net673));
 sg13g2_tiehi _10656__674 (.L_HI(net674));
 sg13g2_tiehi _10867__675 (.L_HI(net675));
 sg13g2_tiehi _10655__676 (.L_HI(net676));
 sg13g2_tiehi _10778__677 (.L_HI(net677));
 sg13g2_tiehi _10654__678 (.L_HI(net678));
 sg13g2_tiehi _10777__679 (.L_HI(net679));
 sg13g2_tiehi _10653__680 (.L_HI(net680));
 sg13g2_tiehi _10776__681 (.L_HI(net681));
 sg13g2_tiehi _10652__682 (.L_HI(net682));
 sg13g2_tiehi _10775__683 (.L_HI(net683));
 sg13g2_tiehi _10651__684 (.L_HI(net684));
 sg13g2_tiehi _10774__685 (.L_HI(net685));
 sg13g2_tiehi _10650__686 (.L_HI(net686));
 sg13g2_tiehi _10773__687 (.L_HI(net687));
 sg13g2_tiehi _10649__688 (.L_HI(net688));
 sg13g2_tiehi _10772__689 (.L_HI(net689));
 sg13g2_tiehi _10648__690 (.L_HI(net690));
 sg13g2_tiehi _10771__691 (.L_HI(net691));
 sg13g2_tiehi _10647__692 (.L_HI(net692));
 sg13g2_tiehi _10646__693 (.L_HI(net693));
 sg13g2_tiehi _10645__694 (.L_HI(net694));
 sg13g2_tiehi _10644__695 (.L_HI(net695));
 sg13g2_tiehi _10643__696 (.L_HI(net696));
 sg13g2_tiehi _10642__697 (.L_HI(net697));
 sg13g2_tiehi _10770__698 (.L_HI(net698));
 sg13g2_tiehi _10641__699 (.L_HI(net699));
 sg13g2_tiehi _10769__700 (.L_HI(net700));
 sg13g2_tiehi _10640__701 (.L_HI(net701));
 sg13g2_tiehi _10639__702 (.L_HI(net702));
 sg13g2_tiehi _10638__703 (.L_HI(net703));
 sg13g2_tiehi _10637__704 (.L_HI(net704));
 sg13g2_tiehi _10636__705 (.L_HI(net705));
 sg13g2_tiehi _10635__706 (.L_HI(net706));
 sg13g2_tiehi _10395__707 (.L_HI(net707));
 sg13g2_tiehi _10544__708 (.L_HI(net708));
 sg13g2_tiehi _10545__709 (.L_HI(net709));
 sg13g2_tiehi _10546__710 (.L_HI(net710));
 sg13g2_tiehi _10547__711 (.L_HI(net711));
 sg13g2_tiehi _10548__712 (.L_HI(net712));
 sg13g2_tiehi _10549__713 (.L_HI(net713));
 sg13g2_tiehi _10550__714 (.L_HI(net714));
 sg13g2_tiehi _10551__715 (.L_HI(net715));
 sg13g2_tiehi _10552__716 (.L_HI(net716));
 sg13g2_tiehi _10553__717 (.L_HI(net717));
 sg13g2_tiehi _10554__718 (.L_HI(net718));
 sg13g2_tiehi _10634__719 (.L_HI(net719));
 sg13g2_tiehi _10633__720 (.L_HI(net720));
 sg13g2_tiehi _10632__721 (.L_HI(net721));
 sg13g2_tiehi _10631__722 (.L_HI(net722));
 sg13g2_tiehi _10555__723 (.L_HI(net723));
 sg13g2_tiehi _10630__724 (.L_HI(net724));
 sg13g2_tiehi _10629__725 (.L_HI(net725));
 sg13g2_tiehi _10628__726 (.L_HI(net726));
 sg13g2_tiehi _10627__727 (.L_HI(net727));
 sg13g2_tiehi _10626__728 (.L_HI(net728));
 sg13g2_tiehi _10625__729 (.L_HI(net729));
 sg13g2_tiehi _10624__730 (.L_HI(net730));
 sg13g2_tiehi _10623__731 (.L_HI(net731));
 sg13g2_tiehi _10622__732 (.L_HI(net732));
 sg13g2_tiehi _10621__733 (.L_HI(net733));
 sg13g2_tiehi _10768__734 (.L_HI(net734));
 sg13g2_tiehi _10620__735 (.L_HI(net735));
 sg13g2_tiehi _10767__736 (.L_HI(net736));
 sg13g2_tiehi _10619__737 (.L_HI(net737));
 sg13g2_tiehi _10766__738 (.L_HI(net738));
 sg13g2_tiehi _10618__739 (.L_HI(net739));
 sg13g2_tiehi _10765__740 (.L_HI(net740));
 sg13g2_tiehi _10617__741 (.L_HI(net741));
 sg13g2_tiehi _10764__742 (.L_HI(net742));
 sg13g2_tiehi _10616__743 (.L_HI(net743));
 sg13g2_tiehi _10763__744 (.L_HI(net744));
 sg13g2_tiehi _10615__745 (.L_HI(net745));
 sg13g2_tiehi _10762__746 (.L_HI(net746));
 sg13g2_tiehi _10614__747 (.L_HI(net747));
 sg13g2_tiehi _10761__748 (.L_HI(net748));
 sg13g2_tiehi _10613__749 (.L_HI(net749));
 sg13g2_tiehi _10760__750 (.L_HI(net750));
 sg13g2_tiehi _10612__751 (.L_HI(net751));
 sg13g2_tiehi _10759__752 (.L_HI(net752));
 sg13g2_tiehi _10611__753 (.L_HI(net753));
 sg13g2_tiehi _10610__754 (.L_HI(net754));
 sg13g2_tiehi _10758__755 (.L_HI(net755));
 sg13g2_tiehi _10609__756 (.L_HI(net756));
 sg13g2_tiehi _10757__757 (.L_HI(net757));
 sg13g2_tiehi _10608__758 (.L_HI(net758));
 sg13g2_tiehi _10756__759 (.L_HI(net759));
 sg13g2_tiehi _10607__760 (.L_HI(net760));
 sg13g2_tiehi _10755__761 (.L_HI(net761));
 sg13g2_tiehi _10606__762 (.L_HI(net762));
 sg13g2_tiehi _10605__763 (.L_HI(net763));
 sg13g2_tiehi _10604__764 (.L_HI(net764));
 sg13g2_tiehi _10603__765 (.L_HI(net765));
 sg13g2_tiehi _10602__766 (.L_HI(net766));
 sg13g2_tiehi _10754__767 (.L_HI(net767));
 sg13g2_tiehi _10601__768 (.L_HI(net768));
 sg13g2_tiehi _10600__769 (.L_HI(net769));
 sg13g2_tiehi _10599__770 (.L_HI(net770));
 sg13g2_tiehi _10598__771 (.L_HI(net771));
 sg13g2_tiehi _10597__772 (.L_HI(net772));
 sg13g2_tiehi _10596__773 (.L_HI(net773));
 sg13g2_tiehi _10595__774 (.L_HI(net774));
 sg13g2_tiehi _10594__775 (.L_HI(net775));
 sg13g2_tiehi _10593__776 (.L_HI(net776));
 sg13g2_tiehi _10592__777 (.L_HI(net777));
 sg13g2_tiehi _10591__778 (.L_HI(net778));
 sg13g2_tiehi _10590__779 (.L_HI(net779));
 sg13g2_tiehi _10589__780 (.L_HI(net780));
 sg13g2_tiehi _10588__781 (.L_HI(net781));
 sg13g2_tiehi _10587__782 (.L_HI(net782));
 sg13g2_tiehi _10586__783 (.L_HI(net783));
 sg13g2_tiehi _10585__784 (.L_HI(net784));
 sg13g2_tiehi _10584__785 (.L_HI(net785));
 sg13g2_tiehi _10583__786 (.L_HI(net786));
 sg13g2_tiehi _10582__787 (.L_HI(net787));
 sg13g2_tiehi _10581__788 (.L_HI(net788));
 sg13g2_tiehi _10580__789 (.L_HI(net789));
 sg13g2_tiehi _10579__790 (.L_HI(net790));
 sg13g2_tiehi _10578__791 (.L_HI(net791));
 sg13g2_tiehi _10577__792 (.L_HI(net792));
 sg13g2_tiehi _10576__793 (.L_HI(net793));
 sg13g2_tiehi _10575__794 (.L_HI(net794));
 sg13g2_tiehi _10574__795 (.L_HI(net795));
 sg13g2_tiehi _10573__796 (.L_HI(net796));
 sg13g2_tiehi _10572__797 (.L_HI(net797));
 sg13g2_tiehi _10571__798 (.L_HI(net798));
 sg13g2_tiehi _10570__799 (.L_HI(net799));
 sg13g2_tiehi _10569__800 (.L_HI(net800));
 sg13g2_tiehi _10568__801 (.L_HI(net801));
 sg13g2_tiehi _10753__802 (.L_HI(net802));
 sg13g2_tiehi _10567__803 (.L_HI(net803));
 sg13g2_tiehi _10752__804 (.L_HI(net804));
 sg13g2_tiehi _10566__805 (.L_HI(net805));
 sg13g2_tiehi _10565__806 (.L_HI(net806));
 sg13g2_tiehi _10564__807 (.L_HI(net807));
 sg13g2_tiehi _10563__808 (.L_HI(net808));
 sg13g2_tiehi _10562__809 (.L_HI(net809));
 sg13g2_tiehi _10751__810 (.L_HI(net810));
 sg13g2_tiehi _10561__811 (.L_HI(net811));
 sg13g2_tiehi _10559__812 (.L_HI(net812));
 sg13g2_tiehi _10750__813 (.L_HI(net813));
 sg13g2_tiehi _10558__814 (.L_HI(net814));
 sg13g2_tiehi _10749__815 (.L_HI(net815));
 sg13g2_tiehi _10557__816 (.L_HI(net816));
 sg13g2_tiehi _10556__817 (.L_HI(net817));
 sg13g2_tiehi _10543__818 (.L_HI(net818));
 sg13g2_tiehi _10542__819 (.L_HI(net819));
 sg13g2_tiehi _10541__820 (.L_HI(net820));
 sg13g2_tiehi _10540__821 (.L_HI(net821));
 sg13g2_tiehi _10539__822 (.L_HI(net822));
 sg13g2_tiehi _10538__823 (.L_HI(net823));
 sg13g2_tiehi _10537__824 (.L_HI(net824));
 sg13g2_tiehi _10536__825 (.L_HI(net825));
 sg13g2_tiehi _10535__826 (.L_HI(net826));
 sg13g2_tiehi _10534__827 (.L_HI(net827));
 sg13g2_tiehi _10533__828 (.L_HI(net828));
 sg13g2_tiehi _10532__829 (.L_HI(net829));
 sg13g2_tiehi _10531__830 (.L_HI(net830));
 sg13g2_tiehi _10530__831 (.L_HI(net831));
 sg13g2_tiehi _10529__832 (.L_HI(net832));
 sg13g2_tiehi _10528__833 (.L_HI(net833));
 sg13g2_tiehi _10527__834 (.L_HI(net834));
 sg13g2_tiehi _10526__835 (.L_HI(net835));
 sg13g2_tiehi _10525__836 (.L_HI(net836));
 sg13g2_tiehi _10524__837 (.L_HI(net837));
 sg13g2_tiehi _10523__838 (.L_HI(net838));
 sg13g2_tiehi _10522__839 (.L_HI(net839));
 sg13g2_tiehi _10521__840 (.L_HI(net840));
 sg13g2_tiehi _10560__841 (.L_HI(net841));
 sg13g2_tiehi _10520__842 (.L_HI(net842));
 sg13g2_tiehi _10519__843 (.L_HI(net843));
 sg13g2_tiehi _10518__844 (.L_HI(net844));
 sg13g2_tiehi _10517__845 (.L_HI(net845));
 sg13g2_tiehi _10516__846 (.L_HI(net846));
 sg13g2_tiehi _10515__847 (.L_HI(net847));
 sg13g2_tiehi _10514__848 (.L_HI(net848));
 sg13g2_tiehi _10513__849 (.L_HI(net849));
 sg13g2_tiehi _10512__850 (.L_HI(net850));
 sg13g2_tiehi _10511__851 (.L_HI(net851));
 sg13g2_tiehi _10510__852 (.L_HI(net852));
 sg13g2_tiehi _10509__853 (.L_HI(net853));
 sg13g2_tiehi _10508__854 (.L_HI(net854));
 sg13g2_tiehi _10507__855 (.L_HI(net855));
 sg13g2_tiehi _10748__856 (.L_HI(net856));
 sg13g2_tiehi _10506__857 (.L_HI(net857));
 sg13g2_tiehi _10747__858 (.L_HI(net858));
 sg13g2_tiehi _10505__859 (.L_HI(net859));
 sg13g2_tiehi _10746__860 (.L_HI(net860));
 sg13g2_tiehi _10504__861 (.L_HI(net861));
 sg13g2_tiehi _10745__862 (.L_HI(net862));
 sg13g2_tiehi _10503__863 (.L_HI(net863));
 sg13g2_tiehi _10502__864 (.L_HI(net864));
 sg13g2_tiehi _10501__865 (.L_HI(net865));
 sg13g2_tiehi _10500__866 (.L_HI(net866));
 sg13g2_tiehi _10499__867 (.L_HI(net867));
 sg13g2_tiehi _10498__868 (.L_HI(net868));
 sg13g2_tiehi _10497__869 (.L_HI(net869));
 sg13g2_tiehi _10496__870 (.L_HI(net870));
 sg13g2_tiehi _10495__871 (.L_HI(net871));
 sg13g2_tiehi _10494__872 (.L_HI(net872));
 sg13g2_tiehi _10493__873 (.L_HI(net873));
 sg13g2_tiehi _10492__874 (.L_HI(net874));
 sg13g2_tiehi _10491__875 (.L_HI(net875));
 sg13g2_tiehi _10490__876 (.L_HI(net876));
 sg13g2_tiehi _10489__877 (.L_HI(net877));
 sg13g2_tiehi _10488__878 (.L_HI(net878));
 sg13g2_tiehi _10487__879 (.L_HI(net879));
 sg13g2_tiehi _10486__880 (.L_HI(net880));
 sg13g2_tiehi _10485__881 (.L_HI(net881));
 sg13g2_tiehi _10484__882 (.L_HI(net882));
 sg13g2_tiehi _10483__883 (.L_HI(net883));
 sg13g2_tiehi _10482__884 (.L_HI(net884));
 sg13g2_tiehi _10481__885 (.L_HI(net885));
 sg13g2_tiehi _10480__886 (.L_HI(net886));
 sg13g2_tiehi _10479__887 (.L_HI(net887));
 sg13g2_tiehi _10478__888 (.L_HI(net888));
 sg13g2_tiehi _10477__889 (.L_HI(net889));
 sg13g2_tiehi _10476__890 (.L_HI(net890));
 sg13g2_tiehi _10475__891 (.L_HI(net891));
 sg13g2_tiehi _10474__892 (.L_HI(net892));
 sg13g2_tiehi _10473__893 (.L_HI(net893));
 sg13g2_tiehi _10472__894 (.L_HI(net894));
 sg13g2_tiehi _10471__895 (.L_HI(net895));
 sg13g2_tiehi _10470__896 (.L_HI(net896));
 sg13g2_tiehi _10469__897 (.L_HI(net897));
 sg13g2_tiehi _10468__898 (.L_HI(net898));
 sg13g2_tiehi _10467__899 (.L_HI(net899));
 sg13g2_tiehi _10466__900 (.L_HI(net900));
 sg13g2_tiehi _10465__901 (.L_HI(net901));
 sg13g2_tiehi _10464__902 (.L_HI(net902));
 sg13g2_tiehi _10463__903 (.L_HI(net903));
 sg13g2_tiehi _10462__904 (.L_HI(net904));
 sg13g2_tiehi _10461__905 (.L_HI(net905));
 sg13g2_tiehi _10460__906 (.L_HI(net906));
 sg13g2_tiehi _10459__907 (.L_HI(net907));
 sg13g2_tiehi _10458__908 (.L_HI(net908));
 sg13g2_tiehi _10457__909 (.L_HI(net909));
 sg13g2_tiehi _10456__910 (.L_HI(net910));
 sg13g2_tiehi _10455__911 (.L_HI(net911));
 sg13g2_tiehi _10454__912 (.L_HI(net912));
 sg13g2_tiehi _10453__913 (.L_HI(net913));
 sg13g2_tiehi _10452__914 (.L_HI(net914));
 sg13g2_tiehi _10451__915 (.L_HI(net915));
 sg13g2_tiehi _10450__916 (.L_HI(net916));
 sg13g2_tiehi _10449__917 (.L_HI(net917));
 sg13g2_tiehi _10448__918 (.L_HI(net918));
 sg13g2_tiehi _10447__919 (.L_HI(net919));
 sg13g2_tiehi _10446__920 (.L_HI(net920));
 sg13g2_tiehi _10445__921 (.L_HI(net921));
 sg13g2_tiehi _10444__922 (.L_HI(net922));
 sg13g2_tiehi _10443__923 (.L_HI(net923));
 sg13g2_tiehi _10442__924 (.L_HI(net924));
 sg13g2_tiehi _10441__925 (.L_HI(net925));
 sg13g2_tiehi _10440__926 (.L_HI(net926));
 sg13g2_tiehi _10439__927 (.L_HI(net927));
 sg13g2_tiehi _10438__928 (.L_HI(net928));
 sg13g2_tiehi _10437__929 (.L_HI(net929));
 sg13g2_tiehi _10436__930 (.L_HI(net930));
 sg13g2_tiehi _10435__931 (.L_HI(net931));
 sg13g2_tiehi _10434__932 (.L_HI(net932));
 sg13g2_tiehi _10433__933 (.L_HI(net933));
 sg13g2_tiehi _10432__934 (.L_HI(net934));
 sg13g2_tiehi _10431__935 (.L_HI(net935));
 sg13g2_tiehi _10430__936 (.L_HI(net936));
 sg13g2_tiehi _10744__937 (.L_HI(net937));
 sg13g2_tiehi _10429__938 (.L_HI(net938));
 sg13g2_tiehi _10743__939 (.L_HI(net939));
 sg13g2_tiehi _10428__940 (.L_HI(net940));
 sg13g2_tiehi _10427__941 (.L_HI(net941));
 sg13g2_tiehi _10426__942 (.L_HI(net942));
 sg13g2_tiehi _10425__943 (.L_HI(net943));
 sg13g2_tiehi _10424__944 (.L_HI(net944));
 sg13g2_tiehi _10423__945 (.L_HI(net945));
 sg13g2_tiehi _10422__946 (.L_HI(net946));
 sg13g2_tiehi _10421__947 (.L_HI(net947));
 sg13g2_tiehi _10420__948 (.L_HI(net948));
 sg13g2_tiehi _10419__949 (.L_HI(net949));
 sg13g2_tiehi _10418__950 (.L_HI(net950));
 sg13g2_tiehi _10417__951 (.L_HI(net951));
 sg13g2_tiehi _10416__952 (.L_HI(net952));
 sg13g2_tiehi _10415__953 (.L_HI(net953));
 sg13g2_tiehi _10414__954 (.L_HI(net954));
 sg13g2_tiehi _10413__955 (.L_HI(net955));
 sg13g2_tiehi _10412__956 (.L_HI(net956));
 sg13g2_tiehi _10411__957 (.L_HI(net957));
 sg13g2_tiehi _10410__958 (.L_HI(net958));
 sg13g2_tiehi _10409__959 (.L_HI(net959));
 sg13g2_tiehi _10408__960 (.L_HI(net960));
 sg13g2_tiehi _10407__961 (.L_HI(net961));
 sg13g2_tiehi _10406__962 (.L_HI(net962));
 sg13g2_tiehi _10405__963 (.L_HI(net963));
 sg13g2_tiehi _10404__964 (.L_HI(net964));
 sg13g2_tiehi _10403__965 (.L_HI(net965));
 sg13g2_tiehi _10402__966 (.L_HI(net966));
 sg13g2_tiehi _10401__967 (.L_HI(net967));
 sg13g2_tiehi _10678__968 (.L_HI(net968));
 sg13g2_tiehi _10805__969 (.L_HI(net969));
 sg13g2_tiehi _10806__970 (.L_HI(net970));
 sg13g2_tiehi _10807__971 (.L_HI(net971));
 sg13g2_tiehi _10808__972 (.L_HI(net972));
 sg13g2_tiehi _10809__973 (.L_HI(net973));
 sg13g2_tiehi _10810__974 (.L_HI(net974));
 sg13g2_tiehi _10811__975 (.L_HI(net975));
 sg13g2_tiehi _10812__976 (.L_HI(net976));
 sg13g2_tiehi _10813__977 (.L_HI(net977));
 sg13g2_tiehi _10814__978 (.L_HI(net978));
 sg13g2_tiehi _10815__979 (.L_HI(net979));
 sg13g2_tiehi _10816__980 (.L_HI(net980));
 sg13g2_tiehi _10817__981 (.L_HI(net981));
 sg13g2_tiehi _10818__982 (.L_HI(net982));
 sg13g2_tiehi _10819__983 (.L_HI(net983));
 sg13g2_tiehi _10820__984 (.L_HI(net984));
 sg13g2_tiehi _10821__985 (.L_HI(net985));
 sg13g2_tiehi _10822__986 (.L_HI(net986));
 sg13g2_tiehi _10823__987 (.L_HI(net987));
 sg13g2_tiehi _10824__988 (.L_HI(net988));
 sg13g2_tiehi _10825__989 (.L_HI(net989));
 sg13g2_tiehi _10826__990 (.L_HI(net990));
 sg13g2_tiehi _10827__991 (.L_HI(net991));
 sg13g2_tiehi _10828__992 (.L_HI(net992));
 sg13g2_tiehi _10829__993 (.L_HI(net993));
 sg13g2_tiehi _10830__994 (.L_HI(net994));
 sg13g2_tiehi _10831__995 (.L_HI(net995));
 sg13g2_tiehi _10400__996 (.L_HI(net996));
 sg13g2_tiehi _10399__997 (.L_HI(net997));
 sg13g2_tiehi _10398__998 (.L_HI(net998));
 sg13g2_tiehi _10397__999 (.L_HI(net999));
 sg13g2_tiehi _10396__1000 (.L_HI(net1000));
 sg13g2_tiehi _10832__1001 (.L_HI(net1001));
 sg13g2_tiehi _10838__1002 (.L_HI(net1002));
 sg13g2_tiehi _10839__1003 (.L_HI(net1003));
 sg13g2_tiehi _10840__1004 (.L_HI(net1004));
 sg13g2_tiehi _10841__1005 (.L_HI(net1005));
 sg13g2_tiehi _10842__1006 (.L_HI(net1006));
 sg13g2_tiehi _10843__1007 (.L_HI(net1007));
 sg13g2_tiehi _10844__1008 (.L_HI(net1008));
 sg13g2_tiehi _10845__1009 (.L_HI(net1009));
 sg13g2_tiehi _10846__1010 (.L_HI(net1010));
 sg13g2_tiehi _10847__1011 (.L_HI(net1011));
 sg13g2_tiehi _10848__1012 (.L_HI(net1012));
 sg13g2_tiehi _10849__1013 (.L_HI(net1013));
 sg13g2_tiehi _10850__1014 (.L_HI(net1014));
 sg13g2_tiehi _10851__1015 (.L_HI(net1015));
 sg13g2_tiehi _10852__1016 (.L_HI(net1016));
 sg13g2_tiehi _10853__1017 (.L_HI(net1017));
 sg13g2_tiehi _10854__1018 (.L_HI(net1018));
 sg13g2_tiehi _10855__1019 (.L_HI(net1019));
 sg13g2_tiehi _10856__1020 (.L_HI(net1020));
 sg13g2_tiehi _10857__1021 (.L_HI(net1021));
 sg13g2_tiehi _10858__1022 (.L_HI(net1022));
 sg13g2_tiehi _10859__1023 (.L_HI(net1023));
 sg13g2_tiehi _10860__1024 (.L_HI(net1024));
 sg13g2_tiehi _10861__1025 (.L_HI(net1025));
 sg13g2_tiehi _10862__1026 (.L_HI(net1026));
 sg13g2_tiehi _10863__1027 (.L_HI(net1027));
 sg13g2_tiehi _10864__1028 (.L_HI(net1028));
 sg13g2_tiehi _10742__1029 (.L_HI(net1029));
 sg13g2_tiehi _10377__1030 (.L_HI(net1030));
 sg13g2_tiehi _10741__1031 (.L_HI(net1031));
 sg13g2_tiehi _10372__1032 (.L_HI(net1032));
 sg13g2_tiehi _10740__1033 (.L_HI(net1033));
 sg13g2_tiehi _10371__1034 (.L_HI(net1034));
 sg13g2_tiehi _10739__1035 (.L_HI(net1035));
 sg13g2_tiehi _10253__1036 (.L_HI(net1036));
 sg13g2_tiehi _09837__1037 (.L_HI(net1037));
 sg13g2_tiehi _09838__1038 (.L_HI(net1038));
 sg13g2_tiehi _09839__1039 (.L_HI(net1039));
 sg13g2_tiehi _09840__1040 (.L_HI(net1040));
 sg13g2_tiehi _09841__1041 (.L_HI(net1041));
 sg13g2_tiehi _09842__1042 (.L_HI(net1042));
 sg13g2_tiehi _09843__1043 (.L_HI(net1043));
 sg13g2_tiehi _09844__1044 (.L_HI(net1044));
 sg13g2_tiehi _09845__1045 (.L_HI(net1045));
 sg13g2_tiehi _09846__1046 (.L_HI(net1046));
 sg13g2_tiehi _09847__1047 (.L_HI(net1047));
 sg13g2_tiehi _09848__1048 (.L_HI(net1048));
 sg13g2_inv_1 _06071__1 (.Y(net1049),
    .A(clknet_1_0__leaf_clk));
 sg13g2_buf_2 _11909_ (.A(net1),
    .X(uio_oe[0]));
 sg13g2_buf_2 _11910_ (.A(uio_oe[5]),
    .X(uio_oe[1]));
 sg13g2_buf_2 _11911_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_2 _11912_ (.A(net1),
    .X(uio_oe[3]));
 sg13g2_buf_2 _11913_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_2 _11914_ (.A(net1),
    .X(uio_oe[6]));
 sg13g2_buf_2 _11915_ (.A(net1),
    .X(uio_oe[7]));
 sg13g2_buf_2 _11916_ (.A(\i_core.mem.q_ctrl.spi_flash_select ),
    .X(uio_out[0]));
 sg13g2_buf_2 _11917_ (.A(\i_core.mem.q_ctrl.spi_clk_out ),
    .X(uio_out[3]));
 sg13g2_buf_2 _11918_ (.A(\i_core.mem.q_ctrl.spi_ram_a_select ),
    .X(uio_out[6]));
 sg13g2_buf_2 _11919_ (.A(\i_core.mem.q_ctrl.spi_ram_b_select ),
    .X(uio_out[7]));
 sg13g2_buf_4 fanout1110 (.X(net1110),
    .A(net1111));
 sg13g2_buf_4 fanout1111 (.X(net1111),
    .A(\debug_rd[3] ));
 sg13g2_buf_2 fanout1112 (.A(_03056_),
    .X(net1112));
 sg13g2_buf_4 fanout1113 (.X(net1113),
    .A(net1114));
 sg13g2_buf_4 fanout1114 (.X(net1114),
    .A(_03221_));
 sg13g2_buf_2 fanout1115 (.A(net1119),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(net1119),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(net1118),
    .X(net1117));
 sg13g2_buf_4 fanout1118 (.X(net1118),
    .A(net1119));
 sg13g2_buf_2 fanout1119 (.A(_03220_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(net1122),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_03218_),
    .X(net1122));
 sg13g2_buf_4 fanout1123 (.X(net1123),
    .A(net1124));
 sg13g2_buf_2 fanout1124 (.A(_02992_),
    .X(net1124));
 sg13g2_buf_4 fanout1125 (.X(net1125),
    .A(_02944_));
 sg13g2_buf_4 fanout1126 (.X(net1126),
    .A(\debug_rd[2] ));
 sg13g2_buf_4 fanout1127 (.X(net1127),
    .A(\debug_rd[2] ));
 sg13g2_buf_4 fanout1128 (.X(net1128),
    .A(net1129));
 sg13g2_buf_4 fanout1129 (.X(net1129),
    .A(net1130));
 sg13g2_buf_4 fanout1130 (.X(net1130),
    .A(_02584_));
 sg13g2_buf_4 fanout1131 (.X(net1131),
    .A(net1132));
 sg13g2_buf_4 fanout1132 (.X(net1132),
    .A(\debug_rd[1] ));
 sg13g2_buf_2 fanout1133 (.A(net1134),
    .X(net1133));
 sg13g2_buf_4 fanout1134 (.X(net1134),
    .A(net1135));
 sg13g2_buf_4 fanout1135 (.X(net1135),
    .A(net1136));
 sg13g2_buf_2 fanout1136 (.A(_03575_),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(net1138),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(net1144),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(net1144),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(net1141),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(net1144),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(net1144),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(net1144),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(_03574_),
    .X(net1144));
 sg13g2_buf_4 fanout1145 (.X(net1145),
    .A(net1146));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(net1147));
 sg13g2_buf_4 fanout1147 (.X(net1147),
    .A(_02746_));
 sg13g2_buf_2 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_4 fanout1149 (.X(net1149),
    .A(net1151));
 sg13g2_buf_2 fanout1150 (.A(net1151),
    .X(net1150));
 sg13g2_buf_2 fanout1151 (.A(_02737_),
    .X(net1151));
 sg13g2_buf_2 fanout1152 (.A(net1153),
    .X(net1152));
 sg13g2_buf_2 fanout1153 (.A(_02733_),
    .X(net1153));
 sg13g2_buf_4 fanout1154 (.X(net1154),
    .A(_02733_));
 sg13g2_buf_2 fanout1155 (.A(_02391_),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(_03500_),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(_03500_),
    .X(net1157));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(_03499_));
 sg13g2_buf_1 fanout1159 (.A(_03499_),
    .X(net1159));
 sg13g2_buf_4 fanout1160 (.X(net1160),
    .A(net1162));
 sg13g2_buf_4 fanout1161 (.X(net1161),
    .A(_03241_));
 sg13g2_buf_2 fanout1162 (.A(_03241_),
    .X(net1162));
 sg13g2_buf_2 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(_03240_),
    .X(net1164));
 sg13g2_buf_4 fanout1165 (.X(net1165),
    .A(net1166));
 sg13g2_buf_2 fanout1166 (.A(\debug_rd[0] ),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(net1169),
    .X(net1167));
 sg13g2_buf_4 fanout1168 (.X(net1168),
    .A(net1169));
 sg13g2_buf_2 fanout1169 (.A(net1170),
    .X(net1169));
 sg13g2_buf_2 fanout1170 (.A(_02578_),
    .X(net1170));
 sg13g2_buf_4 fanout1171 (.X(net1171),
    .A(_01833_));
 sg13g2_buf_4 fanout1172 (.X(net1172),
    .A(net1174));
 sg13g2_buf_4 fanout1173 (.X(net1173),
    .A(_01832_));
 sg13g2_buf_2 fanout1174 (.A(_01832_),
    .X(net1174));
 sg13g2_buf_2 fanout1175 (.A(_03745_),
    .X(net1175));
 sg13g2_buf_4 fanout1176 (.X(net1176),
    .A(net1178));
 sg13g2_buf_1 fanout1177 (.A(net1178),
    .X(net1177));
 sg13g2_buf_4 fanout1178 (.X(net1178),
    .A(_01739_));
 sg13g2_buf_2 fanout1179 (.A(net1181),
    .X(net1179));
 sg13g2_buf_4 fanout1180 (.X(net1180),
    .A(net1181));
 sg13g2_buf_4 fanout1181 (.X(net1181),
    .A(_01738_));
 sg13g2_buf_2 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_2 fanout1183 (.A(_02764_),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(_02416_),
    .X(net1184));
 sg13g2_buf_4 fanout1185 (.X(net1185),
    .A(_01776_));
 sg13g2_buf_2 fanout1186 (.A(net1187),
    .X(net1186));
 sg13g2_buf_4 fanout1187 (.X(net1187),
    .A(_01775_));
 sg13g2_buf_4 fanout1188 (.X(net1188),
    .A(net1189));
 sg13g2_buf_4 fanout1189 (.X(net1189),
    .A(_01773_));
 sg13g2_buf_2 fanout1190 (.A(_01433_),
    .X(net1190));
 sg13g2_buf_2 fanout1191 (.A(_03526_),
    .X(net1191));
 sg13g2_buf_2 fanout1192 (.A(net1193),
    .X(net1192));
 sg13g2_buf_4 fanout1193 (.X(net1193),
    .A(_03525_));
 sg13g2_buf_2 fanout1194 (.A(net1199),
    .X(net1194));
 sg13g2_buf_2 fanout1195 (.A(net1196),
    .X(net1195));
 sg13g2_buf_4 fanout1196 (.X(net1196),
    .A(net1199));
 sg13g2_buf_4 fanout1197 (.X(net1197),
    .A(net1198));
 sg13g2_buf_2 fanout1198 (.A(net1199),
    .X(net1198));
 sg13g2_buf_2 fanout1199 (.A(_01754_),
    .X(net1199));
 sg13g2_buf_2 fanout1200 (.A(net1201),
    .X(net1200));
 sg13g2_buf_4 fanout1201 (.X(net1201),
    .A(_01753_));
 sg13g2_buf_2 fanout1202 (.A(_01429_),
    .X(net1202));
 sg13g2_buf_2 fanout1203 (.A(net1205),
    .X(net1203));
 sg13g2_buf_1 fanout1204 (.A(net1205),
    .X(net1204));
 sg13g2_buf_2 fanout1205 (.A(_02587_),
    .X(net1205));
 sg13g2_buf_2 fanout1206 (.A(net1208),
    .X(net1206));
 sg13g2_buf_1 fanout1207 (.A(net1208),
    .X(net1207));
 sg13g2_buf_2 fanout1208 (.A(_02444_),
    .X(net1208));
 sg13g2_buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_4 fanout1210 (.X(net1210),
    .A(_02050_));
 sg13g2_buf_2 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_4 fanout1212 (.X(net1212),
    .A(_02033_));
 sg13g2_buf_4 fanout1213 (.X(net1213),
    .A(_01827_));
 sg13g2_buf_2 fanout1214 (.A(_01827_),
    .X(net1214));
 sg13g2_buf_4 fanout1215 (.X(net1215),
    .A(_01751_));
 sg13g2_buf_2 fanout1216 (.A(net1217),
    .X(net1216));
 sg13g2_buf_4 fanout1217 (.X(net1217),
    .A(_01581_));
 sg13g2_buf_2 fanout1218 (.A(_03132_),
    .X(net1218));
 sg13g2_buf_2 fanout1219 (.A(_03132_),
    .X(net1219));
 sg13g2_buf_2 fanout1220 (.A(net1223),
    .X(net1220));
 sg13g2_buf_2 fanout1221 (.A(net1222),
    .X(net1221));
 sg13g2_buf_2 fanout1222 (.A(net1223),
    .X(net1222));
 sg13g2_buf_1 fanout1223 (.A(_02786_),
    .X(net1223));
 sg13g2_buf_2 fanout1224 (.A(net1227),
    .X(net1224));
 sg13g2_buf_2 fanout1225 (.A(net1226),
    .X(net1225));
 sg13g2_buf_2 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_buf_2 fanout1227 (.A(_02786_),
    .X(net1227));
 sg13g2_buf_2 fanout1228 (.A(_02528_),
    .X(net1228));
 sg13g2_buf_2 fanout1229 (.A(_02479_),
    .X(net1229));
 sg13g2_buf_2 fanout1230 (.A(net1231),
    .X(net1230));
 sg13g2_buf_2 fanout1231 (.A(_01893_),
    .X(net1231));
 sg13g2_buf_2 fanout1232 (.A(net1233),
    .X(net1232));
 sg13g2_buf_2 fanout1233 (.A(_01649_),
    .X(net1233));
 sg13g2_buf_2 fanout1234 (.A(_01493_),
    .X(net1234));
 sg13g2_buf_2 fanout1235 (.A(_01474_),
    .X(net1235));
 sg13g2_buf_2 fanout1236 (.A(_01458_),
    .X(net1236));
 sg13g2_buf_2 fanout1237 (.A(net1238),
    .X(net1237));
 sg13g2_buf_2 fanout1238 (.A(_01419_),
    .X(net1238));
 sg13g2_buf_2 fanout1239 (.A(net1240),
    .X(net1239));
 sg13g2_buf_4 fanout1240 (.X(net1240),
    .A(net1243));
 sg13g2_buf_4 fanout1241 (.X(net1241),
    .A(net1243));
 sg13g2_buf_1 fanout1242 (.A(net1243),
    .X(net1242));
 sg13g2_buf_2 fanout1243 (.A(_03579_),
    .X(net1243));
 sg13g2_buf_4 fanout1244 (.X(net1244),
    .A(_03578_));
 sg13g2_buf_2 fanout1245 (.A(_03578_),
    .X(net1245));
 sg13g2_buf_4 fanout1246 (.X(net1246),
    .A(_03501_));
 sg13g2_buf_4 fanout1247 (.X(net1247),
    .A(_02069_));
 sg13g2_buf_4 fanout1248 (.X(net1248),
    .A(_01829_));
 sg13g2_buf_4 fanout1249 (.X(net1249),
    .A(_01821_));
 sg13g2_buf_4 fanout1250 (.X(net1250),
    .A(_01795_));
 sg13g2_buf_2 fanout1251 (.A(_01795_),
    .X(net1251));
 sg13g2_buf_4 fanout1252 (.X(net1252),
    .A(_01792_));
 sg13g2_buf_2 fanout1253 (.A(_01788_),
    .X(net1253));
 sg13g2_buf_4 fanout1254 (.X(net1254),
    .A(_01788_));
 sg13g2_buf_2 fanout1255 (.A(net1256),
    .X(net1255));
 sg13g2_buf_4 fanout1256 (.X(net1256),
    .A(_01787_));
 sg13g2_buf_4 fanout1257 (.X(net1257),
    .A(_01781_));
 sg13g2_buf_2 fanout1258 (.A(_03126_),
    .X(net1258));
 sg13g2_buf_2 fanout1259 (.A(_03121_),
    .X(net1259));
 sg13g2_buf_1 fanout1260 (.A(_03121_),
    .X(net1260));
 sg13g2_buf_2 fanout1261 (.A(net1263),
    .X(net1261));
 sg13g2_buf_1 fanout1262 (.A(net1263),
    .X(net1262));
 sg13g2_buf_4 fanout1263 (.X(net1263),
    .A(_03108_));
 sg13g2_buf_4 fanout1264 (.X(net1264),
    .A(net1265));
 sg13g2_buf_4 fanout1265 (.X(net1265),
    .A(net1266));
 sg13g2_buf_4 fanout1266 (.X(net1266),
    .A(_02717_));
 sg13g2_buf_4 fanout1267 (.X(net1267),
    .A(_02717_));
 sg13g2_buf_4 fanout1268 (.X(net1268),
    .A(net1270));
 sg13g2_buf_2 fanout1269 (.A(net1270),
    .X(net1269));
 sg13g2_buf_4 fanout1270 (.X(net1270),
    .A(net1273));
 sg13g2_buf_4 fanout1271 (.X(net1271),
    .A(net1272));
 sg13g2_buf_2 fanout1272 (.A(net1273),
    .X(net1272));
 sg13g2_buf_4 fanout1273 (.X(net1273),
    .A(_01742_));
 sg13g2_buf_4 fanout1274 (.X(net1274),
    .A(net1276));
 sg13g2_buf_4 fanout1275 (.X(net1275),
    .A(net1276));
 sg13g2_buf_4 fanout1276 (.X(net1276),
    .A(_01732_));
 sg13g2_buf_2 fanout1277 (.A(_01327_),
    .X(net1277));
 sg13g2_buf_4 fanout1278 (.X(net1278),
    .A(net1279));
 sg13g2_buf_2 fanout1279 (.A(_01132_),
    .X(net1279));
 sg13g2_buf_2 fanout1280 (.A(_03136_),
    .X(net1280));
 sg13g2_buf_2 fanout1281 (.A(_03136_),
    .X(net1281));
 sg13g2_buf_2 fanout1282 (.A(net1283),
    .X(net1282));
 sg13g2_buf_1 fanout1283 (.A(net1284),
    .X(net1283));
 sg13g2_buf_1 fanout1284 (.A(_02955_),
    .X(net1284));
 sg13g2_buf_2 fanout1285 (.A(net1286),
    .X(net1285));
 sg13g2_buf_1 fanout1286 (.A(net1287),
    .X(net1286));
 sg13g2_buf_2 fanout1287 (.A(_02947_),
    .X(net1287));
 sg13g2_buf_4 fanout1288 (.X(net1288),
    .A(_01838_));
 sg13g2_buf_8 fanout1289 (.A(net1291),
    .X(net1289));
 sg13g2_buf_4 fanout1290 (.X(net1290),
    .A(net1291));
 sg13g2_buf_4 fanout1291 (.X(net1291),
    .A(_01745_));
 sg13g2_buf_4 fanout1292 (.X(net1292),
    .A(net1293));
 sg13g2_buf_2 fanout1293 (.A(_01744_),
    .X(net1293));
 sg13g2_buf_4 fanout1294 (.X(net1294),
    .A(_01744_));
 sg13g2_buf_2 fanout1295 (.A(net1296),
    .X(net1295));
 sg13g2_buf_1 fanout1296 (.A(net1300),
    .X(net1296));
 sg13g2_buf_2 fanout1297 (.A(net1300),
    .X(net1297));
 sg13g2_buf_2 fanout1298 (.A(net1299),
    .X(net1298));
 sg13g2_buf_2 fanout1299 (.A(net1300),
    .X(net1299));
 sg13g2_buf_4 fanout1300 (.X(net1300),
    .A(_01733_));
 sg13g2_buf_2 fanout1301 (.A(net1302),
    .X(net1301));
 sg13g2_buf_2 fanout1302 (.A(net1303),
    .X(net1302));
 sg13g2_buf_1 fanout1303 (.A(_01305_),
    .X(net1303));
 sg13g2_buf_2 fanout1304 (.A(_01304_),
    .X(net1304));
 sg13g2_buf_2 fanout1305 (.A(_01304_),
    .X(net1305));
 sg13g2_buf_2 fanout1306 (.A(net1307),
    .X(net1306));
 sg13g2_buf_2 fanout1307 (.A(_01165_),
    .X(net1307));
 sg13g2_buf_4 fanout1308 (.X(net1308),
    .A(net1309));
 sg13g2_buf_2 fanout1309 (.A(_01160_),
    .X(net1309));
 sg13g2_buf_4 fanout1310 (.X(net1310),
    .A(_01159_));
 sg13g2_buf_4 fanout1311 (.X(net1311),
    .A(net1312));
 sg13g2_buf_4 fanout1312 (.X(net1312),
    .A(_01133_));
 sg13g2_buf_2 fanout1313 (.A(net1316),
    .X(net1313));
 sg13g2_buf_4 fanout1314 (.X(net1314),
    .A(net1316));
 sg13g2_buf_2 fanout1315 (.A(net1316),
    .X(net1315));
 sg13g2_buf_2 fanout1316 (.A(net1318),
    .X(net1316));
 sg13g2_buf_2 fanout1317 (.A(net1318),
    .X(net1317));
 sg13g2_buf_2 fanout1318 (.A(_00818_),
    .X(net1318));
 sg13g2_buf_4 fanout1319 (.X(net1319),
    .A(_00154_));
 sg13g2_buf_4 fanout1320 (.X(net1320),
    .A(net1322));
 sg13g2_buf_4 fanout1321 (.X(net1321),
    .A(net1322));
 sg13g2_buf_2 fanout1322 (.A(net1327),
    .X(net1322));
 sg13g2_buf_2 fanout1323 (.A(net1324),
    .X(net1323));
 sg13g2_buf_1 fanout1324 (.A(net1327),
    .X(net1324));
 sg13g2_buf_4 fanout1325 (.X(net1325),
    .A(net1327));
 sg13g2_buf_2 fanout1326 (.A(net1327),
    .X(net1326));
 sg13g2_buf_2 fanout1327 (.A(\i_core.mem.q_ctrl.rstn ),
    .X(net1327));
 sg13g2_buf_4 fanout1328 (.X(net1328),
    .A(_03135_));
 sg13g2_buf_2 fanout1329 (.A(_03135_),
    .X(net1329));
 sg13g2_buf_2 fanout1330 (.A(_03134_),
    .X(net1330));
 sg13g2_buf_2 fanout1331 (.A(net1332),
    .X(net1331));
 sg13g2_buf_2 fanout1332 (.A(_02972_),
    .X(net1332));
 sg13g2_buf_2 fanout1333 (.A(_02024_),
    .X(net1333));
 sg13g2_buf_1 fanout1334 (.A(_02024_),
    .X(net1334));
 sg13g2_buf_4 fanout1335 (.X(net1335),
    .A(_01185_));
 sg13g2_buf_4 fanout1336 (.X(net1336),
    .A(_01173_));
 sg13g2_buf_2 fanout1337 (.A(_00949_),
    .X(net1337));
 sg13g2_buf_2 fanout1338 (.A(_00939_),
    .X(net1338));
 sg13g2_buf_2 fanout1339 (.A(_00938_),
    .X(net1339));
 sg13g2_buf_2 fanout1340 (.A(_00935_),
    .X(net1340));
 sg13g2_buf_2 fanout1341 (.A(_00934_),
    .X(net1341));
 sg13g2_buf_1 fanout1342 (.A(_00934_),
    .X(net1342));
 sg13g2_buf_2 fanout1343 (.A(net1345),
    .X(net1343));
 sg13g2_buf_4 fanout1344 (.X(net1344),
    .A(net1345));
 sg13g2_buf_4 fanout1345 (.X(net1345),
    .A(_00931_));
 sg13g2_buf_4 fanout1346 (.X(net1346),
    .A(net1349));
 sg13g2_buf_2 fanout1347 (.A(net1348),
    .X(net1347));
 sg13g2_buf_2 fanout1348 (.A(net1349),
    .X(net1348));
 sg13g2_buf_2 fanout1349 (.A(_00930_),
    .X(net1349));
 sg13g2_buf_4 fanout1350 (.X(net1350),
    .A(net1351));
 sg13g2_buf_4 fanout1351 (.X(net1351),
    .A(net1352));
 sg13g2_buf_2 fanout1352 (.A(net1353),
    .X(net1352));
 sg13g2_buf_2 fanout1353 (.A(_00908_),
    .X(net1353));
 sg13g2_buf_4 fanout1354 (.X(net1354),
    .A(_00907_));
 sg13g2_buf_2 fanout1355 (.A(_00893_),
    .X(net1355));
 sg13g2_buf_2 fanout1356 (.A(_00891_),
    .X(net1356));
 sg13g2_buf_4 fanout1357 (.X(net1357),
    .A(net1359));
 sg13g2_buf_4 fanout1358 (.X(net1358),
    .A(net1359));
 sg13g2_buf_4 fanout1359 (.X(net1359),
    .A(_00881_));
 sg13g2_buf_4 fanout1360 (.X(net1360),
    .A(_00879_));
 sg13g2_buf_2 fanout1361 (.A(net1362),
    .X(net1361));
 sg13g2_buf_4 fanout1362 (.X(net1362),
    .A(_00879_));
 sg13g2_buf_2 fanout1363 (.A(net1365),
    .X(net1363));
 sg13g2_buf_2 fanout1364 (.A(net1365),
    .X(net1364));
 sg13g2_buf_4 fanout1365 (.X(net1365),
    .A(_00876_));
 sg13g2_buf_4 fanout1366 (.X(net1366),
    .A(net1367));
 sg13g2_buf_2 fanout1367 (.A(_00874_),
    .X(net1367));
 sg13g2_buf_2 fanout1368 (.A(_00874_),
    .X(net1368));
 sg13g2_buf_2 fanout1369 (.A(net1370),
    .X(net1369));
 sg13g2_buf_1 fanout1370 (.A(_00829_),
    .X(net1370));
 sg13g2_buf_2 fanout1371 (.A(net1372),
    .X(net1371));
 sg13g2_buf_2 fanout1372 (.A(net1373),
    .X(net1372));
 sg13g2_buf_2 fanout1373 (.A(_00829_),
    .X(net1373));
 sg13g2_buf_4 fanout1374 (.X(net1374),
    .A(_00791_));
 sg13g2_buf_4 fanout1375 (.X(net1375),
    .A(_00790_));
 sg13g2_buf_2 fanout1376 (.A(_00790_),
    .X(net1376));
 sg13g2_buf_2 fanout1377 (.A(net1378),
    .X(net1377));
 sg13g2_buf_4 fanout1378 (.X(net1378),
    .A(net1379));
 sg13g2_buf_4 fanout1379 (.X(net1379),
    .A(_00788_));
 sg13g2_buf_2 fanout1380 (.A(net1382),
    .X(net1380));
 sg13g2_buf_4 fanout1381 (.X(net1381),
    .A(net1382));
 sg13g2_buf_4 fanout1382 (.X(net1382),
    .A(_00786_));
 sg13g2_buf_2 fanout1383 (.A(net1384),
    .X(net1383));
 sg13g2_buf_2 fanout1384 (.A(net1387),
    .X(net1384));
 sg13g2_buf_4 fanout1385 (.X(net1385),
    .A(net1387));
 sg13g2_buf_2 fanout1386 (.A(net1387),
    .X(net1386));
 sg13g2_buf_2 fanout1387 (.A(_00783_),
    .X(net1387));
 sg13g2_buf_2 fanout1388 (.A(net1389),
    .X(net1388));
 sg13g2_buf_2 fanout1389 (.A(_00755_),
    .X(net1389));
 sg13g2_buf_2 fanout1390 (.A(net1392),
    .X(net1390));
 sg13g2_buf_1 fanout1391 (.A(net1392),
    .X(net1391));
 sg13g2_buf_2 fanout1392 (.A(net1393),
    .X(net1392));
 sg13g2_buf_2 fanout1393 (.A(debug_instr_valid),
    .X(net1393));
 sg13g2_buf_4 fanout1394 (.X(net1394),
    .A(net2681));
 sg13g2_buf_4 fanout1395 (.X(net1395),
    .A(net1401));
 sg13g2_buf_4 fanout1396 (.X(net1396),
    .A(net1400));
 sg13g2_buf_1 fanout1397 (.A(net1400),
    .X(net1397));
 sg13g2_buf_8 fanout1398 (.A(net1400),
    .X(net1398));
 sg13g2_buf_2 fanout1399 (.A(net1400),
    .X(net1399));
 sg13g2_buf_2 fanout1400 (.A(net1401),
    .X(net1400));
 sg13g2_buf_2 fanout1401 (.A(\i_core.cpu.alu_op[2] ),
    .X(net1401));
 sg13g2_buf_4 fanout1402 (.X(net1402),
    .A(\i_core.cpu.alu_op[1] ));
 sg13g2_buf_2 fanout1403 (.A(\i_core.cpu.alu_op[1] ),
    .X(net1403));
 sg13g2_buf_4 fanout1404 (.X(net1404),
    .A(net1405));
 sg13g2_buf_2 fanout1405 (.A(net1407),
    .X(net1405));
 sg13g2_buf_2 fanout1406 (.A(net1407),
    .X(net1406));
 sg13g2_buf_2 fanout1407 (.A(\i_core.cpu.counter[4] ),
    .X(net1407));
 sg13g2_buf_2 fanout1408 (.A(net1409),
    .X(net1408));
 sg13g2_buf_2 fanout1409 (.A(net1410),
    .X(net1409));
 sg13g2_buf_4 fanout1410 (.X(net1410),
    .A(\i_core.cpu.counter[3] ));
 sg13g2_buf_4 fanout1411 (.X(net1411),
    .A(net1412));
 sg13g2_buf_2 fanout1412 (.A(net1415),
    .X(net1412));
 sg13g2_buf_2 fanout1413 (.A(net1414),
    .X(net1413));
 sg13g2_buf_4 fanout1414 (.X(net1414),
    .A(net1415));
 sg13g2_buf_4 fanout1415 (.X(net1415),
    .A(net1416));
 sg13g2_buf_8 fanout1416 (.A(\i_core.cpu.counter[2] ),
    .X(net1416));
 sg13g2_buf_2 fanout1417 (.A(net1419),
    .X(net1417));
 sg13g2_buf_2 fanout1418 (.A(net1419),
    .X(net1418));
 sg13g2_buf_1 fanout1419 (.A(net2671),
    .X(net1419));
 sg13g2_buf_2 fanout1420 (.A(net1421),
    .X(net1420));
 sg13g2_buf_2 fanout1421 (.A(net1422),
    .X(net1421));
 sg13g2_buf_2 fanout1422 (.A(\i_core.cpu.was_early_branch ),
    .X(net1422));
 sg13g2_buf_2 fanout1423 (.A(net2670),
    .X(net1423));
 sg13g2_buf_2 fanout1424 (.A(net2664),
    .X(net1424));
 sg13g2_buf_2 fanout1425 (.A(net2494),
    .X(net1425));
 sg13g2_buf_2 fanout1426 (.A(\i_core.cpu.instr_data_start[14] ),
    .X(net1426));
 sg13g2_buf_4 fanout1427 (.X(net1427),
    .A(\i_core.cpu.instr_data_start[7] ));
 sg13g2_buf_2 fanout1428 (.A(net2631),
    .X(net1428));
 sg13g2_buf_2 fanout1429 (.A(_00152_),
    .X(net1429));
 sg13g2_buf_2 fanout1430 (.A(\i_core.mem.q_ctrl.fsm_state[2] ),
    .X(net1430));
 sg13g2_buf_4 fanout1431 (.X(net1431),
    .A(net2663));
 sg13g2_buf_2 fanout1432 (.A(net1433),
    .X(net1432));
 sg13g2_buf_1 fanout1433 (.A(net1435),
    .X(net1433));
 sg13g2_buf_2 fanout1434 (.A(net1435),
    .X(net1434));
 sg13g2_buf_1 fanout1435 (.A(\i_core.mem.q_ctrl.is_writing ),
    .X(net1435));
 sg13g2_buf_2 fanout1436 (.A(net2672),
    .X(net1436));
 sg13g2_buf_4 fanout1437 (.X(net1437),
    .A(\i_core.mem.qspi_data_byte_idx[0] ));
 sg13g2_buf_2 fanout1438 (.A(\i_core.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .X(net1438));
 sg13g2_buf_2 fanout1439 (.A(net1440),
    .X(net1439));
 sg13g2_buf_2 fanout1440 (.A(net1441),
    .X(net1440));
 sg13g2_buf_1 fanout1441 (.A(\i_core.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .X(net1441));
 sg13g2_buf_2 fanout1442 (.A(net1444),
    .X(net1442));
 sg13g2_buf_1 fanout1443 (.A(net1444),
    .X(net1443));
 sg13g2_buf_1 fanout1444 (.A(net2673),
    .X(net1444));
 sg13g2_buf_2 fanout1445 (.A(net1446),
    .X(net1445));
 sg13g2_buf_1 fanout1446 (.A(net1447),
    .X(net1446));
 sg13g2_buf_2 fanout1447 (.A(\i_core.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .X(net1447));
 sg13g2_buf_2 fanout1448 (.A(net1449),
    .X(net1448));
 sg13g2_buf_4 fanout1449 (.X(net1449),
    .A(\i_core.cpu.i_core.i_shift.adjusted_shift_amt[0] ));
 sg13g2_buf_2 fanout1450 (.A(\addr[4] ),
    .X(net1450));
 sg13g2_buf_2 fanout1451 (.A(net1452),
    .X(net1451));
 sg13g2_buf_1 fanout1452 (.A(net2587),
    .X(net1452));
 sg13g2_buf_2 fanout1453 (.A(net1456),
    .X(net1453));
 sg13g2_buf_2 fanout1454 (.A(net1456),
    .X(net1454));
 sg13g2_buf_2 fanout1455 (.A(net1456),
    .X(net1455));
 sg13g2_buf_2 fanout1456 (.A(\i_spi.busy ),
    .X(net1456));
 sg13g2_buf_4 fanout1457 (.X(net1457),
    .A(net1458));
 sg13g2_buf_4 fanout1458 (.X(net1458),
    .A(net2426));
 sg13g2_buf_2 fanout1459 (.A(net1460),
    .X(net1459));
 sg13g2_buf_2 fanout1460 (.A(net1461),
    .X(net1460));
 sg13g2_buf_4 fanout1461 (.X(net1461),
    .A(net2442));
 sg13g2_buf_4 fanout1462 (.X(net1462),
    .A(net2443));
 sg13g2_buf_2 fanout1463 (.A(net1464),
    .X(net1463));
 sg13g2_buf_4 fanout1464 (.X(net1464),
    .A(net2443));
 sg13g2_buf_4 fanout1465 (.X(net1465),
    .A(net1467));
 sg13g2_buf_2 fanout1466 (.A(net1467),
    .X(net1466));
 sg13g2_buf_2 fanout1467 (.A(net2480),
    .X(net1467));
 sg13g2_buf_2 fanout1468 (.A(net5),
    .X(net1468));
 sg13g2_buf_2 fanout1469 (.A(net1470),
    .X(net1469));
 sg13g2_buf_2 fanout1470 (.A(ui_in[3]),
    .X(net1470));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_4 input9 (.X(net9),
    .A(uio_in[1]));
 sg13g2_buf_4 input10 (.X(net10),
    .A(uio_in[2]));
 sg13g2_buf_4 input11 (.X(net11),
    .A(uio_in[4]));
 sg13g2_buf_2 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_tiehi _09849__13 (.L_HI(net13));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_leaf_0_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_1_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_2_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_3_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_4_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_5_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_6_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_7_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_8_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_9_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_10_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_11_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_12_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_13_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_14_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_15_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_16_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_17_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_18_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_19_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_20_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_21_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_22_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_23_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_24_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_25_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_26_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_27_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_28_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_29_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_30_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_31_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_32_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_33_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_34_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_35_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_36_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_37_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_38_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_39_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_40_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_41_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_42_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_43_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_43_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_44_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_44_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_45_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_45_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_46_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_46_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_47_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_47_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_48_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_48_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_49_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_49_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_50_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_50_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_51_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_51_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_52_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_52_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_53_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_53_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_54_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_54_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_55_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_55_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_56_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_56_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_57_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_57_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_58_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_58_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_59_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_59_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_60_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_60_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_61_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_61_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_62_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_62_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_63_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_63_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_64_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_64_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_65_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_65_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_66_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_66_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_67_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_67_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_68_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_68_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_69_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_69_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_70_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_70_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_71_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_71_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_72_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_72_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_73_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_73_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_74_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_74_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_75_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_75_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_76_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_76_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_77_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_77_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_78_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_78_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_79_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_79_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_80_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_80_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_81_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_81_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_82_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_82_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_83_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_83_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_84_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_84_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_85_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_85_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_86_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_86_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_87_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_87_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_88_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_88_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_89_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_89_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_90_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_90_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_91_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_91_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_92_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_92_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_93_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_93_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_94_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_94_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_95_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_95_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_96_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_96_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_97_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_97_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_98_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_98_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_99_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_99_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_100_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_100_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_101_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_101_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_102_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_102_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_103_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_103_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_104_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_104_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_105_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_105_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_106_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_106_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_107_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_107_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_108_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_108_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_109_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_109_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_110_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_110_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_111_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_111_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_112_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_112_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_113_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_113_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_114_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_114_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_115_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_115_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_116_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_116_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_117_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_117_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_118_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_118_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_119_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_119_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_120_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_120_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_121_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_121_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_122_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_122_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_123_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_123_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_124_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_124_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_125_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_125_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_126_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_126_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_128_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_128_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_129_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_129_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_130_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_130_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_131_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_131_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_132_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_132_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_133_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_133_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_134_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_134_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_135_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_135_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_136_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_136_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_137_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_137_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_138_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_138_clk_regs));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_1 clkload0 (.A(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkload1 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkload2 (.A(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkload3 (.A(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkload4 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkload5 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkload6 (.A(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkload7 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkload8 (.A(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkload9 (.A(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkload10 (.A(clknet_5_29__leaf_clk_regs));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_0_clk_regs));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_138_clk_regs));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_9_clk_regs));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_126_clk_regs));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_13_clk_regs));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_16_clk_regs));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_15_clk_regs));
 sg13g2_inv_8 clkload18 (.A(clknet_leaf_73_clk_regs));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_123_clk_regs));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_19_clk_regs));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_20_clk_regs));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_21_clk_regs));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_28_clk_regs));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_35_clk_regs));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_49_clk_regs));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_38_clk_regs));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_122_clk_regs));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_97_clk_regs));
 sg13g2_inv_2 clkload29 (.A(clknet_leaf_72_clk_regs));
 sg13g2_inv_4 clkload30 (.A(clknet_leaf_119_clk_regs));
 sg13g2_inv_4 clkload31 (.A(clknet_leaf_53_clk_regs));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_54_clk_regs));
 sg13g2_inv_2 clkload33 (.A(clknet_leaf_59_clk_regs));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_76_clk_regs));
 sg13g2_inv_2 clkload35 (.A(clknet_leaf_61_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(delaynet_1_clk));
 sg13g2_buf_2 delaybuf_1_clk (.A(delaynet_1_clk),
    .X(delaynet_2_clk));
 sg13g2_buf_2 delaybuf_2_clk (.A(delaynet_2_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold2 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold3 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold4 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[20].A ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[17].A ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold33 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold37 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[13].A ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold43 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[8].A ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold45 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold47 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold51 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold57 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[26].A ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold61 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold64 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold67 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold69 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[15].A ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold71 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold73 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold77 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold79 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold83 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold85 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold90 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold92 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold94 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold100 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[27].A ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold102 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold104 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold105 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold107 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold115 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold117 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[30].A ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[7].A ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold121 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold136 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold137 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold142 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[6].A ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[14].A ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[5].A ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold150 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold152 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[11].A ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[29].A ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[23].A ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[23].A ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[25].A ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold172 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold180 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold184 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[14].A ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold189 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold190 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold193 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold196 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold197 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[8].A ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold198 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[27].A ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold201 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[26].A ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold202 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[17].A ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold203 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[24].A ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold205 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[4].A ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[24].A ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[22].A ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold208 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[21].A ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold209 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold210 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[19].A ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[11].A ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold212 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[19].A ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[15].A ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold214 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[12].A ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold216 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[31].A ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold218 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold221 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[20].A ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold224 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold225 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold226 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold227 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[10].A ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold229 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold231 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold233 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold236 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[16].A ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold239 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[21].A ),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold240 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold241 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold242 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold243 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold245 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold247 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold249 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold251 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold253 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[10].A ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold256 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold257 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold258 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold259 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[16].A ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold260 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold262 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold263 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[31].A ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold264 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[28].A ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold266 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold267 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[29].A ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold268 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[9].A ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold269 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold270 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold271 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold272 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold273 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold274 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold275 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[22].A ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold277 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[13].A ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold279 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold280 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold281 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[7].A ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold283 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold284 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold285 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold287 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold288 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold289 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold290 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold291 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold293 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold294 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold295 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold296 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold297 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[18].A ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold298 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold299 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold300 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold301 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold302 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold303 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold304 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold305 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold306 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold307 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold308 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold309 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold310 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold311 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold312 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold313 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold314 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold315 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold316 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold317 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[15].A ),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold318 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[25].A ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold319 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold320 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold321 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold322 (.A(\i_core.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold323 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold324 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[28].A ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold325 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[9].A ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold326 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[12].A ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold327 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold328 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[18].A ),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold329 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold330 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold331 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold332 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold333 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold334 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold335 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold336 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold337 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold338 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold339 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold340 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[23].A ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold341 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold342 (.A(\i_core.cpu.i_core.i_instrret.i_regbuf[30].A ),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold343 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold344 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold345 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[16].A ),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold346 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold347 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold348 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[20].A ),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold349 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold350 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold351 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold352 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold353 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold354 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[30].A ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold355 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold356 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[18].A ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold357 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold358 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold359 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold360 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[28].A ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold361 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[22].A ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold362 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold363 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[17].A ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold364 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold365 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold366 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold367 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold368 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold369 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold370 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold371 (.A(\i_core.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold372 (.A(\i_core.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold373 (.A(\i_core.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold374 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold375 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold376 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold377 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[21].A ),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold378 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold379 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[4].A ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold380 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[8].A ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold381 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[14].A ),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold382 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[29].A ),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold383 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold384 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[19].A ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold385 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold386 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold387 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[13].A ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold388 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold389 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold390 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold391 (.A(\i_core.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold392 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold393 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold394 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold395 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold396 (.A(\i_core.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold397 (.A(\i_core.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold398 (.A(\i_core.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold399 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold400 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[9].A ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold401 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[31].A ),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold402 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[11].A ),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold403 (.A(\i_core.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold404 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[10].A ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold405 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold406 (.A(_00220_),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold407 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[6].A ),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold408 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[12].A ),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold409 (.A(\i_core.cpu.i_core.i_cycles.i_regbuf[5].A ),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold410 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold411 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold412 (.A(\i_core.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold413 (.A(\i_core.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold414 (.A(\i_core.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[4].A ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold415 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[5].A ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold416 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[6].A ),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold417 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[7].A ),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold418 (.A(\i_core.cpu.instr_data[2][13] ),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold419 (.A(_00399_),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold420 (.A(\i_core.cpu.i_core.i_instrret.data[1] ),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold421 (.A(_00744_),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold422 (.A(\i_uart_rx.rxd_reg[1] ),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold423 (.A(\i_core.cpu.instr_data[3][13] ),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold424 (.A(_00413_),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold425 (.A(\i_core.cpu.instr_data[1][13] ),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold426 (.A(_00462_),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold427 (.A(\i_core.cpu.instr_data[1][8] ),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold428 (.A(_00457_),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold429 (.A(\i_core.cpu.instr_data[3][14] ),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold430 (.A(_00414_),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold431 (.A(\i_core.cpu.instr_data[1][14] ),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold432 (.A(_00463_),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold433 (.A(\i_core.cpu.instr_data[2][15] ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold434 (.A(_00401_),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold435 (.A(\i_core.cpu.instr_data[2][12] ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold436 (.A(_00398_),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold437 (.A(\i_core.cpu.instr_data[1][12] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold438 (.A(_00461_),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold439 (.A(\i_core.cpu.instr_data[2][10] ),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold440 (.A(_00396_),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold441 (.A(\i_core.cpu.instr_data[1][9] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold442 (.A(_00458_),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold443 (.A(\i_core.cpu.instr_data[3][10] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold444 (.A(_00410_),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold445 (.A(\i_core.cpu.instr_data[2][9] ),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold446 (.A(_00395_),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold447 (.A(\i_core.cpu.instr_data[3][11] ),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold448 (.A(_00411_),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold449 (.A(\i_core.cpu.instr_data[1][10] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold450 (.A(_00459_),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold451 (.A(\i_core.cpu.instr_data[1][15] ),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold452 (.A(_00464_),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold453 (.A(\i_core.cpu.instr_data[3][8] ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold454 (.A(_00408_),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold455 (.A(\i_core.cpu.instr_data[3][9] ),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold456 (.A(_00409_),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold457 (.A(\i_core.cpu.instr_data[2][8] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold458 (.A(_00394_),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold459 (.A(\i_core.cpu.instr_data[2][11] ),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold460 (.A(_00397_),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold461 (.A(_00219_),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold462 (.A(_02616_),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold463 (.A(_00310_),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold464 (.A(\i_core.mem.q_ctrl.addr[0] ),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold465 (.A(_03880_),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold466 (.A(\i_core.cpu.instr_data[2][14] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold467 (.A(_00400_),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold468 (.A(\i_core.cpu.instr_data[1][11] ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold469 (.A(_00460_),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold470 (.A(\data_to_write[29] ),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold471 (.A(\i_debug_uart_tx.cycle_counter[4] ),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold472 (.A(_02625_),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold473 (.A(\i_core.cpu.instr_data[3][15] ),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold474 (.A(_00415_),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold475 (.A(\i_core.cpu.instr_data[3][12] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold476 (.A(_00412_),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold477 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[24].A ),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold478 (.A(\i_core.mem.data_from_read[16] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold479 (.A(_00515_),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold480 (.A(\data_to_write[30] ),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold481 (.A(\i_core.mem.data_from_read[23] ),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold482 (.A(_00522_),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold483 (.A(\i_core.mem.data_from_read[18] ),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold484 (.A(_00517_),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold485 (.A(\i_core.mem.data_from_read[19] ),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold486 (.A(_00518_),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold487 (.A(\data_to_write[26] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold488 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[27].A ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold489 (.A(\i_core.cpu.instr_data[0][11] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold490 (.A(_00383_),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold491 (.A(\data_to_write[10] ),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold492 (.A(\data_to_write[27] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold493 (.A(\data_to_write[28] ),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold494 (.A(\i_core.mem.data_from_read[21] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold495 (.A(_00520_),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold496 (.A(\i_core.mem.q_ctrl.spi_ram_b_select ),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold497 (.A(\i_core.mem.data_from_read[22] ),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold498 (.A(_00521_),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold499 (.A(\data_to_write[31] ),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold500 (.A(\i_core.cpu.instr_data[0][12] ),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold501 (.A(_00384_),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold502 (.A(\i_core.cpu.instr_data[0][6] ),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold503 (.A(_00378_),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold504 (.A(\i_uart_tx.data_to_send[7] ),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold505 (.A(_00256_),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold506 (.A(\i_spi.bits_remaining[1] ),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold507 (.A(_02668_),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold508 (.A(\i_core.mem.data_from_read[17] ),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold509 (.A(_00516_),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold510 (.A(\i_core.cpu.load_started ),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold511 (.A(_00611_),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold512 (.A(\i_core.cpu.instr_data[0][14] ),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold513 (.A(_00386_),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold514 (.A(\data_to_write[11] ),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold515 (.A(_00215_),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold516 (.A(_00244_),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold517 (.A(\data_to_write[19] ),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold518 (.A(_03479_),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold519 (.A(\i_core.mem.q_ctrl.addr[5] ),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold520 (.A(_00717_),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold521 (.A(\i_core.cpu.instr_data[0][4] ),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold522 (.A(_00376_),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold523 (.A(\i_core.cpu.instr_data[0][8] ),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold524 (.A(_00380_),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold525 (.A(\i_debug_uart_tx.data_to_send[7] ),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold526 (.A(_00309_),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold527 (.A(\i_core.mem.q_ctrl.spi_ram_a_select ),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold528 (.A(\data_to_write[24] ),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold529 (.A(\i_core.cpu.instr_data[0][7] ),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold530 (.A(_00379_),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold531 (.A(\i_core.cpu.instr_data[0][5] ),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold532 (.A(_00377_),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold533 (.A(_00222_),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold534 (.A(_02348_),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold535 (.A(_00232_),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold536 (.A(\i_core.cpu.instr_data[3][1] ),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold537 (.A(_00301_),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold538 (.A(\i_core.cpu.instr_data[0][9] ),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold539 (.A(_00381_),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold540 (.A(\i_core.cpu.instr_data[0][13] ),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold541 (.A(_00385_),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold542 (.A(\i_spi.data[4] ),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold543 (.A(_00419_),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold544 (.A(\i_core.cpu.instr_data[0][15] ),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold545 (.A(_00387_),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold546 (.A(\i_core.cpu.imm[31] ),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold547 (.A(\i_core.mem.q_ctrl.spi_in_buffer[2] ),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold548 (.A(_00558_),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold549 (.A(\i_spi.data[7] ),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold550 (.A(_00422_),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold551 (.A(\i_core.cpu.instr_data[0][10] ),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold552 (.A(_00382_),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold553 (.A(\i_core.mem.qspi_data_buf[24] ),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold554 (.A(_02983_),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold555 (.A(\i_spi.read_latency ),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold556 (.A(\i_core.cpu.i_core.mcause[3] ),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold557 (.A(_00229_),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold558 (.A(\i_uart_tx.cycle_counter[1] ),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold559 (.A(_02482_),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold560 (.A(_00258_),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold561 (.A(\i_core.mem.data_from_read[20] ),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold562 (.A(_00519_),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold563 (.A(\i_core.cpu.imm[26] ),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold564 (.A(\data_to_write[17] ),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold565 (.A(_03477_),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold566 (.A(\i_core.mem.q_ctrl.addr[19] ),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold567 (.A(_00731_),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold568 (.A(\i_spi.bits_remaining[0] ),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold569 (.A(_00323_),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold570 (.A(_00221_),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold571 (.A(_02481_),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold572 (.A(\i_core.mem.qspi_data_buf[31] ),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold573 (.A(_02990_),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold574 (.A(\i_core.mem.qspi_data_buf[27] ),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold575 (.A(_02986_),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold576 (.A(\gpio_out[4] ),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold577 (.A(_00004_),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold578 (.A(\gpio_out[7] ),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold579 (.A(_00007_),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold580 (.A(\data_to_write[16] ),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold581 (.A(_03476_),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold582 (.A(\i_core.cpu.imm[28] ),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold583 (.A(\i_spi.data[6] ),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold584 (.A(_00421_),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold585 (.A(\i_core.mem.q_ctrl.spi_in_buffer[7] ),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold586 (.A(_00559_),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold587 (.A(\i_spi.data[3] ),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold588 (.A(_00418_),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold589 (.A(\i_core.mem.q_ctrl.spi_in_buffer[5] ),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold590 (.A(_00557_),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold591 (.A(\i_spi.data[1] ),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold592 (.A(_00416_),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold593 (.A(\i_core.mem.qspi_data_buf[15] ),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold594 (.A(\gpio_out[1] ),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold595 (.A(\i_spi.data[5] ),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold596 (.A(\i_core.mem.qspi_data_buf[29] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold597 (.A(\i_core.cpu.i_core.time_hi[2] ),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold598 (.A(_02351_),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold599 (.A(_00234_),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold600 (.A(\gpio_out[2] ),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold601 (.A(_00002_),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold602 (.A(\i_core.cpu.instr_data[2][4] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold603 (.A(_00390_),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold604 (.A(\gpio_out[3] ),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold605 (.A(_00003_),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold606 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[25].A ),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold607 (.A(\i_core.cpu.instr_data[3][5] ),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold608 (.A(_00405_),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold609 (.A(\i_core.cpu.instr_data[3][7] ),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold610 (.A(_00407_),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold611 (.A(\i_core.cpu.instr_data[2][6] ),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold612 (.A(_00392_),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold613 (.A(\i_uart_rx.rxd_reg[0] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold614 (.A(_00291_),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold615 (.A(\i_core.mem.qspi_data_buf[28] ),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold616 (.A(\i_uart_rx.bit_sample ),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold617 (.A(_00279_),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold618 (.A(\i_core.cpu.imm[27] ),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold619 (.A(\i_core.cpu.i_core.i_registers.reg_access[7][0] ),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold620 (.A(\i_core.mem.q_ctrl.spi_in_buffer[4] ),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold621 (.A(_00556_),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold622 (.A(\i_core.cpu.imm[25] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold623 (.A(\i_core.mem.q_ctrl.addr[3] ),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold624 (.A(_00719_),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold625 (.A(\i_core.mem.q_ctrl.addr[4] ),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold626 (.A(_03885_),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold627 (.A(\data_to_write[18] ),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold628 (.A(_03478_),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold629 (.A(\i_spi.data[2] ),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold630 (.A(_00417_),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold631 (.A(\i_core.cpu.i_core.i_registers.reg_access[15][2] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold632 (.A(\i_spi.clock_divider[1] ),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold633 (.A(\i_core.cpu.i_core.mepc[11] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold634 (.A(_00472_),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold635 (.A(\i_core.cpu.instr_data[3][0] ),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold636 (.A(_00300_),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold637 (.A(\i_core.mem.qspi_data_buf[26] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold638 (.A(_02985_),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold639 (.A(\i_core.cpu.instr_data[2][7] ),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold640 (.A(_00393_),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold641 (.A(\addr[1] ),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold642 (.A(_00424_),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold643 (.A(\i_core.mem.qspi_data_buf[14] ),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold644 (.A(_00513_),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold645 (.A(\i_core.mem.qspi_data_buf[13] ),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold646 (.A(\i_core.cpu.instr_data[1][5] ),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold647 (.A(_00454_),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold648 (.A(\i_core.mem.qspi_data_buf[12] ),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold649 (.A(\i_core.mem.qspi_data_buf[30] ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold650 (.A(_02989_),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold651 (.A(\i_core.mem.q_ctrl.addr[6] ),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold652 (.A(_00718_),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold653 (.A(\i_core.mem.q_ctrl.spi_data_oe[0] ),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold654 (.A(_00549_),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold655 (.A(\i_core.cpu.imm[24] ),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold656 (.A(\gpio_out[6] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold657 (.A(_00006_),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold658 (.A(\i_core.mem.q_ctrl.addr[13] ),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold659 (.A(_03938_),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold660 (.A(_00725_),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold661 (.A(\i_core.mem.q_ctrl.addr[17] ),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold662 (.A(_00729_),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold663 (.A(\i_core.cpu.instr_data[3][4] ),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold664 (.A(_00404_),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold665 (.A(\i_core.cpu.instr_data[1][7] ),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold666 (.A(_00456_),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold667 (.A(\i_core.cpu.instr_data[1][4] ),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold668 (.A(_00453_),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold669 (.A(\i_core.cpu.instr_data[3][6] ),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold670 (.A(_00406_),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold671 (.A(\i_core.mem.qspi_data_buf[10] ),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold672 (.A(\i_core.mem.q_ctrl.addr[9] ),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold673 (.A(_03916_),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold674 (.A(\i_core.cpu.i_core.i_registers.reg_access[10][0] ),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold675 (.A(\i_core.mem.qspi_data_buf[8] ),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold676 (.A(_00507_),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold677 (.A(\data_to_write[25] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold678 (.A(\i_core.mem.q_ctrl.addr[2] ),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold679 (.A(_03228_),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold680 (.A(\i_core.mem.q_ctrl.spi_in_buffer[0] ),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold681 (.A(_03122_),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold682 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[26].A ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold683 (.A(\i_core.mem.q_ctrl.delay_cycles_cfg[0] ),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold684 (.A(\i_uart_rx.cycle_counter[1] ),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold685 (.A(_02529_),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold686 (.A(_00281_),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold687 (.A(\i_core.cpu.imm[30] ),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold688 (.A(\addr[3] ),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold689 (.A(\i_core.mem.qspi_data_buf[9] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold690 (.A(_00508_),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold691 (.A(\gpio_out[5] ),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold692 (.A(_00005_),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold693 (.A(\i_uart_tx.cycle_counter[7] ),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold694 (.A(_02493_),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold695 (.A(_00264_),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold696 (.A(\i_core.mem.q_ctrl.addr[10] ),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold697 (.A(_03922_),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold698 (.A(\i_core.cpu.instr_data[2][5] ),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold699 (.A(_00391_),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold700 (.A(\addr[23] ),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold701 (.A(_00446_),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold702 (.A(\i_core.cpu.instr_data[0][3] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold703 (.A(_00375_),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold704 (.A(\i_core.mem.q_ctrl.addr[15] ),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold705 (.A(_03949_),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold706 (.A(_00727_),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold707 (.A(\i_core.cpu.instr_data[1][6] ),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold708 (.A(_00455_),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold709 (.A(\i_core.mem.q_ctrl.addr[14] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold710 (.A(_03944_),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold711 (.A(\i_core.mem.qspi_data_buf[25] ),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold712 (.A(_02984_),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold713 (.A(\i_core.mem.q_ctrl.stop_txn_reg ),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold714 (.A(\i_core.mem.qspi_data_buf[11] ),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold715 (.A(\i_core.cpu.imm[29] ),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold716 (.A(\i_core.cpu.i_core.mepc[19] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold717 (.A(_00484_),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold718 (.A(\i_core.cpu.i_core.time_hi[1] ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold719 (.A(_00233_),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold720 (.A(\i_core.cpu.i_core.last_interrupt_req[0] ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold721 (.A(_00235_),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold722 (.A(\data_to_write[13] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold723 (.A(\data_to_write[12] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold724 (.A(\i_spi.spi_select ),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold725 (.A(_00329_),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold726 (.A(\addr[6] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold727 (.A(\i_core.mem.q_ctrl.spi_in_buffer[3] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold728 (.A(_03124_),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold729 (.A(\i_core.cpu.i_core.is_interrupt ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold730 (.A(\addr[18] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold731 (.A(\i_core.mem.q_ctrl.addr[8] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold732 (.A(_03910_),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold733 (.A(\i_core.mem.q_ctrl.addr[1] ),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold734 (.A(_00578_),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold735 (.A(\i_core.cpu.i_core.i_shift.a[21] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold736 (.A(_00359_),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold737 (.A(\i_core.cpu.i_core.last_interrupt_req[1] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold738 (.A(_00236_),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold739 (.A(\i_core.cpu.i_core.i_shift.a[18] ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold740 (.A(_00360_),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold741 (.A(\i_core.cpu.i_core.mepc[12] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold742 (.A(_00473_),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold743 (.A(\addr[7] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold744 (.A(\i_spi.clock_count[0] ),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold745 (.A(\i_spi.spi_dc ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold746 (.A(_00328_),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold747 (.A(\i_core.mem.q_ctrl.delay_cycles_cfg[1] ),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold748 (.A(\i_core.cpu.instr_data[0][2] ),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold749 (.A(_00374_),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold750 (.A(\gpio_out[0] ),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold751 (.A(\i_core.mem.q_ctrl.addr[11] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold752 (.A(_03927_),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold753 (.A(_00723_),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold754 (.A(\i_uart_rx.recieved_data[0] ),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold755 (.A(_00272_),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold756 (.A(\i_core.cpu.i_core.mepc[18] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold757 (.A(_00479_),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold758 (.A(\i_core.cpu.i_core.mie[19] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold759 (.A(_00337_),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold760 (.A(\i_core.mem.q_ctrl.addr[16] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold761 (.A(_00728_),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold762 (.A(\addr[20] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold763 (.A(\i_core.cpu.i_core.mepc[16] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold764 (.A(_00481_),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold765 (.A(\data_to_write[23] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold766 (.A(\i_core.cpu.data_ready_latch ),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold767 (.A(_00648_),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold768 (.A(\i_core.cpu.i_core.i_shift.a[25] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold769 (.A(\i_core.mem.q_ctrl.addr[23] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold770 (.A(_00735_),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold771 (.A(\data_to_write[22] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold772 (.A(\i_core.mem.q_ctrl.addr[18] ),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold773 (.A(\data_to_write[14] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold774 (.A(\data_to_write[21] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold775 (.A(\i_core.cpu.i_core.i_registers.reg_access[15][3] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold776 (.A(\addr[14] ),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold777 (.A(\i_core.mem.q_ctrl.spi_in_buffer[1] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold778 (.A(\data_to_write[15] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold779 (.A(\i_core.cpu.i_core.load_done ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold780 (.A(_00224_),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold781 (.A(\data_to_write[20] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold782 (.A(\i_core.cpu.i_core.i_registers.reg_access[7][1] ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold783 (.A(\gpio_out_sel[2] ),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold784 (.A(_00010_),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold785 (.A(\gpio_out_sel[3] ),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold786 (.A(_00011_),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold787 (.A(\i_core.cpu.i_core.i_registers.reg_access[15][1] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold788 (.A(\addr[22] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold789 (.A(_00445_),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold790 (.A(\i_core.cpu.additional_mem_ops[2] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold791 (.A(\i_spi.end_txn_reg ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold792 (.A(_00299_),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold793 (.A(_00160_),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold794 (.A(_03120_),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold795 (.A(\addr[21] ),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold796 (.A(_00444_),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold797 (.A(\i_core.cpu.i_core.i_registers.reg_access[2][1] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold798 (.A(\i_core.cpu.i_core.mepc[13] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold799 (.A(_00474_),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold800 (.A(\i_core.cpu.is_auipc ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold801 (.A(\i_spi.bits_remaining[2] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold802 (.A(_02670_),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold803 (.A(_00217_),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold804 (.A(_04004_),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold805 (.A(_00743_),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold806 (.A(\i_core.cpu.i_core.i_shift.a[17] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold807 (.A(_00355_),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold808 (.A(\i_core.cpu.i_core.i_registers.reg_access[2][3] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold809 (.A(\i_uart_tx.cycle_counter[2] ),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold810 (.A(_02484_),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold811 (.A(\i_core.cpu.instr_data[1][3] ),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold812 (.A(_00452_),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold813 (.A(\i_debug_uart_tx.cycle_counter[1] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold814 (.A(_02619_),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold815 (.A(_00311_),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold816 (.A(\i_uart_rx.recieved_data[5] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold817 (.A(_00276_),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold818 (.A(\i_core.cpu.i_core.mepc[8] ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold819 (.A(_00469_),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold820 (.A(\addr[15] ),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold821 (.A(_00438_),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold822 (.A(\gpio_out_sel[1] ),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold823 (.A(\addr[0] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold824 (.A(_00423_),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold825 (.A(\i_core.cpu.i_core.mepc[17] ),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold826 (.A(_00482_),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold827 (.A(debug_data_continue),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold828 (.A(_00492_),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold829 (.A(\i_core.cpu.i_core.i_registers.reg_access[13][0] ),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold830 (.A(\i_core.mem.q_ctrl.addr[12] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold831 (.A(_03933_),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold832 (.A(\i_core.cpu.i_core.i_registers.reg_access[13][1] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold833 (.A(\i_core.cpu.i_core.i_registers.reg_access[1][3] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold834 (.A(\addr[17] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold835 (.A(\i_core.cpu.i_core.i_registers.reg_access[7][3] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold836 (.A(\gpio_out_sel[4] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold837 (.A(_00012_),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold838 (.A(\i_uart_rx.recieved_data[2] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold839 (.A(_00273_),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold840 (.A(\i_core.cpu.i_core.i_shift.a[29] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold841 (.A(\i_core.cpu.i_core.mepc[15] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold842 (.A(\i_uart_rx.recieved_data[6] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold843 (.A(\gpio_out_sel[5] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold844 (.A(_00013_),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold845 (.A(\i_core.cpu.i_core.i_shift.a[14] ),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold846 (.A(\addr[16] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold847 (.A(\i_core.cpu.i_core.i_registers.reg_access[1][2] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold848 (.A(\gpio_out_sel[0] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold849 (.A(\i_core.cpu.i_core.mepc[22] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold850 (.A(\i_core.cpu.i_core.mepc[14] ),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold851 (.A(_00475_),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold852 (.A(\i_core.cpu.is_jal ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold853 (.A(\i_uart_rx.recieved_data[3] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold854 (.A(\i_uart_rx.recieved_data[7] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold855 (.A(\i_core.cpu.instr_data[1][2] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold856 (.A(_00451_),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold857 (.A(\addr[13] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold858 (.A(\i_core.cpu.i_core.i_shift.b[3] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold859 (.A(\i_core.cpu.i_core.mepc[9] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold860 (.A(_00470_),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold861 (.A(\i_core.cpu.i_core.i_shift.a[22] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold862 (.A(_00364_),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold863 (.A(\i_core.cpu.i_core.i_shift.a[23] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold864 (.A(_00365_),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold865 (.A(\i_core.cpu.i_core.i_registers.reg_access[8][2] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold866 (.A(\i_uart_tx.cycle_counter[9] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold867 (.A(_02497_),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold868 (.A(\i_core.cpu.i_core.i_shift.a[20] ),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold869 (.A(_00362_),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold870 (.A(\i_core.cpu.i_core.i_registers.reg_access[2][2] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold871 (.A(\i_uart_rx.cycle_counter[4] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold872 (.A(_02534_),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold873 (.A(\i_core.cpu.i_core.mie[17] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold874 (.A(_00339_),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold875 (.A(\i_core.cpu.i_core.is_double_fault_r ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold876 (.A(_00231_),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold877 (.A(\i_core.cpu.i_core.mem_op[2] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold878 (.A(\i_core.cpu.instr_data[3][3] ),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold879 (.A(_00403_),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold880 (.A(\i_core.cpu.instr_data_in[13] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold881 (.A(_00504_),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold882 (.A(\i_debug_uart_tx.fsm_state[2] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold883 (.A(_00317_),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold884 (.A(\i_core.cpu.i_core.i_registers.reg_access[7][2] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold885 (.A(\i_core.cpu.i_core.i_registers.reg_access[2][0] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold886 (.A(\i_core.cpu.i_core.i_registers.reg_access[14][1] ),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold887 (.A(\i_core.cpu.i_core.mepc[21] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold888 (.A(\i_core.cpu.i_core.i_registers.reg_access[14][0] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold889 (.A(\i_core.cpu.i_core.i_shift.a[26] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold890 (.A(_00368_),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold891 (.A(\i_core.cpu.i_core.i_shift.a[28] ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold892 (.A(\addr[12] ),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold893 (.A(\i_uart_rx.cycle_counter[8] ),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold894 (.A(_02542_),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold895 (.A(\i_core.mem.q_ctrl.addr[22] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold896 (.A(\i_core.cpu.i_core.i_registers.reg_access[8][1] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold897 (.A(\i_core.cpu.instr_data[2][1] ),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold898 (.A(_00572_),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold899 (.A(\i_uart_rx.recieved_data[4] ),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold900 (.A(\gpio_out_sel[6] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold901 (.A(_00014_),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold902 (.A(\i_core.cpu.i_core.i_registers.reg_access[10][1] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold903 (.A(\i_core.cpu.i_core.mie[18] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold904 (.A(\i_spi.clock_divider[0] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold905 (.A(\i_spi.bits_remaining[3] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold906 (.A(_02672_),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold907 (.A(_00326_),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold908 (.A(\i_core.cpu.instr_data[2][2] ),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold909 (.A(_00388_),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold910 (.A(\i_core.cpu.additional_mem_ops[1] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold911 (.A(_00709_),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold912 (.A(\i_core.cpu.i_core.i_registers.reg_access[8][0] ),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold913 (.A(\i_uart_rx.cycle_counter[3] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold914 (.A(_02532_),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold915 (.A(\i_core.cpu.i_core.i_shift.a[16] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold916 (.A(\i_core.cpu.i_core.mie[16] ),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold917 (.A(\i_core.mem.q_ctrl.last_ram_b_sel ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold918 (.A(_03102_),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold919 (.A(\i_uart_tx.cycle_counter[3] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold920 (.A(\i_core.cpu.i_core.i_registers.reg_access[1][0] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold921 (.A(\addr[25] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold922 (.A(\i_uart_rx.cycle_counter[2] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold923 (.A(_02530_),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold924 (.A(\i_uart_tx.cycle_counter[4] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold925 (.A(\i_core.cpu.i_core.mepc[4] ),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold926 (.A(_00465_),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold927 (.A(\i_core.cpu.i_core.i_shift.a[19] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold928 (.A(\i_core.cpu.i_core.mip[16] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold929 (.A(_00336_),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold930 (.A(\i_core.cpu.i_core.i_registers.reg_access[14][3] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold931 (.A(\i_core.cpu.instr_data[1][1] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold932 (.A(_00373_),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold933 (.A(\i_uart_tx.cycle_counter[8] ),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold934 (.A(_02495_),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold935 (.A(\i_uart_tx.cycle_counter[5] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold936 (.A(\i_core.cpu.i_core.mepc[5] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold937 (.A(_00466_),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold938 (.A(_00161_),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold939 (.A(\i_core.cpu.instr_data[2][3] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold940 (.A(_00389_),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold941 (.A(\i_core.cpu.i_core.i_shift.a[12] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold942 (.A(\i_core.cpu.i_core.mepc[7] ),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold943 (.A(_00468_),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold944 (.A(\i_core.mem.q_ctrl.addr[20] ),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold945 (.A(\i_core.cpu.i_core.mepc[6] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold946 (.A(_00471_),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold947 (.A(\i_uart_rx.cycle_counter[6] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold948 (.A(_02538_),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold949 (.A(\i_uart_tx.cycle_counter[6] ),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold950 (.A(\i_core.cpu.i_core.i_registers.reg_access[10][3] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold951 (.A(\i_core.cpu.i_core.mstatus_mpie ),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold952 (.A(_02383_),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold953 (.A(_00241_),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold954 (.A(\i_core.cpu.i_core.mepc[2] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold955 (.A(\i_uart_tx.fsm_state[2] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold956 (.A(_02511_),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold957 (.A(_00270_),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold958 (.A(\i_core.mem.q_ctrl.addr[21] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold959 (.A(\i_uart_rx.cycle_counter[5] ),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold960 (.A(\i_core.cpu.instr_data_in[11] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold961 (.A(\i_core.cpu.i_core.i_registers.reg_access[13][3] ),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold962 (.A(\i_core.cpu.instr_data[3][2] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold963 (.A(_00402_),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold964 (.A(\i_core.cpu.instr_data_in[9] ),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold965 (.A(_00565_),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold966 (.A(\i_core.mem.q_ctrl.spi_clk_out ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold967 (.A(\i_core.cpu.i_core.i_shift.a[27] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold968 (.A(_00369_),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold969 (.A(\i_uart_rx.cycle_counter[9] ),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold970 (.A(\i_core.cpu.i_core.i_registers.reg_access[12][1] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold971 (.A(\i_core.cpu.instr_len[1] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold972 (.A(\addr[19] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold973 (.A(\i_core.cpu.i_core.mcause[1] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold974 (.A(_00228_),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold975 (.A(\i_core.cpu.i_core.i_registers.reg_access[6][3] ),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold976 (.A(\i_uart_tx.data_to_send[0] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold977 (.A(_00341_),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold978 (.A(\addr[9] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold979 (.A(\i_uart_rx.cycle_counter[7] ),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold980 (.A(\i_core.cpu.i_core.i_registers.reg_access[9][1] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold981 (.A(\addr[11] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold982 (.A(\i_core.cpu.no_write_in_progress ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold983 (.A(_00159_),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold984 (.A(_03079_),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold985 (.A(\i_debug_uart_tx.fsm_state[3] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold986 (.A(_02641_),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold987 (.A(\i_uart_tx.fsm_state[1] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold988 (.A(\i_debug_uart_tx.data_to_send[0] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold989 (.A(_02681_),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold990 (.A(_00331_),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold991 (.A(\i_core.cpu.data_ready_core ),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold992 (.A(\i_core.cpu.i_core.i_registers.reg_access[1][1] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold993 (.A(\i_core.cpu.instr_data[0][1] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold994 (.A(_00490_),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold995 (.A(\addr[27] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold996 (.A(_02863_),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold997 (.A(_00214_),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold998 (.A(_03861_),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold999 (.A(\i_core.cpu.i_core.i_shift.a[15] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\i_core.cpu.i_core.mepc[23] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\i_core.cpu.instr_data_in[6] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold1002 (.A(_00505_),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\i_core.cpu.i_core.cycle_count[3] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold1004 (.A(_02346_),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\addr[24] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\i_core.cpu.i_core.mcause[4] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\i_core.cpu.instr_data_in[1] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\i_core.cpu.i_core.cycle[0] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold1009 (.A(_02326_),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\i_core.cpu.i_core.mip[17] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold1011 (.A(_00335_),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\i_core.cpu.i_core.i_instrret.data[3] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold1013 (.A(_00740_),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold1014 (.A(_00086_),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\i_core.cpu.i_core.i_registers.reg_access[6][1] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold1016 (.A(_00153_),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold1017 (.A(_00028_),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\i_core.cpu.imm[12] ),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\addr[10] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\addr[26] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold1021 (.A(_02862_),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\i_spi.data[0] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\i_core.mem.q_ctrl.nibbles_remaining[2] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\addr[8] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\i_core.cpu.instr_data_start[7] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\i_core.cpu.i_core.i_registers.reg_access[10][2] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\i_core.cpu.i_core.i_registers.reg_access[14][2] ),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\i_core.cpu.instr_data[1][0] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold1029 (.A(_00372_),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\i_core.cpu.i_core.mstatus_mte ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold1031 (.A(_00243_),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\i_core.cpu.i_core.i_cycles.rstn ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold1033 (.A(net1467),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\addr[5] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\i_core.cpu.i_core.i_registers.reg_access[12][3] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\i_core.cpu.i_core.i_registers.reg_access[12][0] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\i_debug_uart_tx.cycle_counter[2] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold1038 (.A(_02623_),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\addr[4] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\i_core.cpu.i_core.i_registers.rs1[1] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\i_core.cpu.instr_data[0][0] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold1042 (.A(_00489_),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\i_core.cpu.i_core.i_registers.reg_access[15][0] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\i_core.cpu.i_core.i_registers.reg_access[8][3] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\i_core.cpu.i_core.i_registers.reg_access[9][2] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\i_core.cpu.instr_data_start[14] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\i_core.cpu.i_core.i_registers.reg_access[9][3] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\data_to_write[8] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\i_core.cpu.imm[15] ),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\i_core.cpu.mem_op_increment_reg ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\data_to_write[9] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\i_core.cpu.instr_data_in[15] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold1053 (.A(_00506_),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\i_core.mem.instr_active ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold1055 (.A(_02991_),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\i_core.cpu.imm[23] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\i_core.cpu.i_core.i_shift.a[1] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold1058 (.A(_00343_),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\i_core.cpu.instr_data_in[12] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold1060 (.A(_00564_),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\data_to_write[7] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\i_uart_rx.fsm_state[0] ),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold1063 (.A(_00293_),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\i_core.cpu.i_core.i_shift.a[3] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold1065 (.A(_00345_),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\i_core.cpu.i_core.i_shift.a[24] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\i_core.cpu.instr_data_start[9] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\i_core.cpu.i_core.i_shift.b[4] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\i_core.cpu.i_core.i_registers.reg_access[12][2] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\i_core.cpu.i_core.i_cycles.rstn ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\i_uart_tx.cycle_counter[10] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\i_core.cpu.i_core.i_registers.rs1[0] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\i_core.cpu.instr_data_in[8] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\i_spi.clock_count[1] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold1075 (.A(_00321_),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\i_core.cpu.is_alu_reg ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\i_core.cpu.i_core.cycle_count[2] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold1078 (.A(_04002_),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\i_core.cpu.data_write_n[1] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold1080 (.A(_00607_),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\i_core.cpu.data_read_n[0] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold1082 (.A(_00608_),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\i_core.cpu.instr_len[2] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\i_core.cpu.instr_data_start[15] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\i_core.cpu.i_core.i_registers.reg_access[11][1] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\i_debug_uart_tx.fsm_state[1] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold1087 (.A(_02634_),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\i_core.cpu.instr_data[2][0] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold1089 (.A(_00571_),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\i_core.cpu.imm[19] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold1091 (.A(_00151_),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold1092 (.A(_00531_),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold1093 (.A(_00218_),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\i_core.cpu.imm[16] ),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\i_core.mem.q_ctrl.data_req ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold1096 (.A(_00082_),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\i_core.cpu.i_core.i_registers.reg_access[6][0] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\i_core.cpu.i_core.i_registers.reg_access[9][0] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\i_core.cpu.i_core.i_registers.rs1[2] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\i_core.mem.q_ctrl.read_cycles_count[0] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold1101 (.A(_00533_),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\i_uart_rx.fsm_state[2] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold1103 (.A(_02569_),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold1104 (.A(_00295_),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\i_core.cpu.instr_data_start[23] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\i_core.cpu.imm[22] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\i_core.cpu.imm[17] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\i_uart_tx.fsm_state[3] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold1109 (.A(_00271_),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\i_core.cpu.imm[13] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\i_core.cpu.i_core.i_registers.rs2[1] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\i_core.cpu.instr_data_start[17] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\i_core.cpu.i_core.cycle_count[0] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold1114 (.A(_03999_),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold1115 (.A(_00736_),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\i_core.cpu.imm[20] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\i_core.cpu.i_core.i_shift.a[2] ),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold1118 (.A(_00344_),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\i_core.cpu.i_core.imm_lo[0] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\i_core.cpu.i_core.i_registers.reg_access[13][2] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\i_uart_rx.cycle_counter[10] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\i_core.cpu.data_write_n[0] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\i_core.cpu.data_read_n[1] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold1124 (.A(_00609_),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\i_debug_uart_tx.cycle_counter[3] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold1126 (.A(_02624_),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold1127 (.A(_00157_),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold1128 (.A(_02939_),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\i_core.cpu.i_core.i_registers.reg_access[6][2] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\i_core.mem.q_ctrl.spi_flash_select ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold1131 (.A(_00547_),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\i_core.cpu.i_core.i_shift.a[30] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\i_core.cpu.i_core.i_shift.a[0] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold1134 (.A(_00342_),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\i_debug_uart_tx.fsm_state[0] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold1136 (.A(_02632_),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\i_core.cpu.instr_data_in[0] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\i_core.cpu.i_core.i_registers.reg_access[11][2] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\i_uart_tx.fsm_state[0] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\i_core.cpu.i_core.i_registers.rs1[3] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\i_core.mem.q_ctrl.delay_cycles_cfg[2] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\i_core.cpu.instr_data_in[4] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\i_core.cpu.imm[14] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\i_core.mem.q_ctrl.nibbles_remaining[1] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\i_core.cpu.instr_data_start[5] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\i_core.cpu.i_core.mepc[20] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\i_core.cpu.i_core.i_registers.reg_access[11][3] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\i_core.cpu.i_core.mstatus_mte ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold1149 (.A(_00242_),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\i_core.cpu.i_core.imm_lo[4] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\i_core.cpu.i_core.i_registers.reg_access[11][0] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\i_spi.spi_clk_out ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\i_core.cpu.i_core.imm_lo[7] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\i_core.cpu.instr_data_in[3] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\i_debug_uart_tx.data_to_send[6] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold1156 (.A(_00308_),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\i_core.cpu.i_core.i_registers.reg_access[5][3] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\i_core.cpu.is_lui ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\i_uart_rx.fsm_state[3] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold1160 (.A(_00296_),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\i_core.cpu.i_core.i_instrret.data[2] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold1162 (.A(_04011_),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\i_core.mem.q_ctrl.read_cycles_count[2] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\i_core.cpu.i_core.i_registers.reg_access[5][0] ),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\i_uart_rx.fsm_state[1] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\i_core.cpu.i_core.i_shift.b[2] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\i_debug_uart_tx.data_to_send[1] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\i_core.cpu.instr_data_start[4] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\i_core.cpu.instr_data_start[12] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\i_core.cpu.imm[18] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\i_uart_tx.data_to_send[2] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold1172 (.A(_02460_),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\i_core.cpu.i_core.load_top_bit ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\i_core.cpu.i_core.i_registers.reg_access[5][1] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\i_core.cpu.i_core.i_registers.rs2[3] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\i_core.cpu.i_core.imm_lo[6] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\addr[2] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\i_core.cpu.i_core.mem_op[1] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\i_debug_uart_tx.data_to_send[2] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\i_core.cpu.i_core.i_registers.reg_access[5][2] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\i_core.cpu.is_system ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\i_uart_tx.data_to_send[1] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\i_core.cpu.i_core.imm_lo[1] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\i_core.cpu.imm[21] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\i_core.cpu.i_core.i_registers.rs2[2] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\i_debug_uart_tx.data_to_send[4] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_02603_),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold1188 (.A(_00305_),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\i_core.cpu.instr_data_start[19] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\i_debug_uart_tx.data_to_send[5] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold1191 (.A(_00307_),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\i_uart_tx.data_to_send[6] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold1193 (.A(_00255_),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\i_core.cpu.i_core.imm_lo[2] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\i_core.cpu.i_core.mcause[0] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\i_core.cpu.i_core.i_registers.rs2[0] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\i_uart_tx.data_to_send[4] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold1198 (.A(_02466_),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold1199 (.A(_00252_),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\i_uart_tx.data_to_send[5] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold1201 (.A(_00254_),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\i_core.cpu.i_core.i_shift.a[11] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\i_core.mem.q_ctrl.nibbles_remaining[0] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\i_core.cpu.i_core.imm_lo[3] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\i_core.cpu.i_core.i_shift.a[10] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\i_core.cpu.i_core.i_shift.a[8] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold1207 (.A(_00158_),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\i_core.cpu.is_store ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\i_core.cpu.i_core.cycle_count[1] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold1210 (.A(debug_register_data),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\i_core.cpu.instr_data_start[13] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\data_to_write[4] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\i_debug_uart_tx.data_to_send[3] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold1214 (.A(_00304_),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\i_core.cpu.i_core.imm_lo[5] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\i_core.cpu.instr_data_in[2] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold1217 (.A(_00501_),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\i_core.cpu.is_alu_imm ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\i_core.cpu.i_core.i_shift.a[6] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\i_core.cpu.instr_data_in[10] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\i_core.cpu.instr_data_start[3] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\i_core.cpu.i_core.i_shift.a[13] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold1223 (.A(_00351_),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\i_uart_tx.data_to_send[3] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\i_core.cpu.i_core.i_registers.rd[2] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\i_core.cpu.i_core.i_shift.a[7] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\i_core.cpu.i_core.imm_lo[11] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\i_core.cpu.pc[1] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\i_core.cpu.i_core.i_registers.rd[1] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\i_core.cpu.instr_fetch_running ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold1231 (.A(_03430_),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold1232 (.A(_00087_),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\i_core.cpu.i_core.imm_lo[9] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\i_core.cpu.pc[2] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\i_core.cpu.i_core.i_registers.rd[3] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\i_core.cpu.i_core.i_shift.a[5] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold1237 (.A(_00347_),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\i_core.cpu.instr_data_start[11] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\i_core.cpu.i_core.i_shift.a[4] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\i_core.cpu.instr_data_start[22] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\i_core.cpu.instr_data_start[8] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold1242 (.A(_00588_),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\i_core.cpu.i_core.imm_lo[8] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\i_core.mem.qspi_data_byte_idx[1] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\i_core.cpu.i_core.i_shift.a[31] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\i_core.cpu.instr_data_start[6] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\i_core.cpu.instr_data_start[21] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\i_core.cpu.i_core.imm_lo[10] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\i_core.cpu.instr_data_in[14] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\i_core.cpu.is_jalr ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\gpio_out_sel[7] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\i_core.cpu.instr_data_start[10] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\i_core.mem.q_ctrl.fsm_state[1] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\i_core.cpu.instr_data_start[16] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\i_core.cpu.i_core.mem_op[0] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\i_core.cpu.alu_op[3] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\i_core.cpu.is_branch ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\i_core.mem.q_ctrl.last_ram_a_sel ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold1259 (.A(_03077_),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\i_core.cpu.instr_data_start[20] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\i_core.cpu.was_early_branch ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\i_core.mem.q_ctrl.read_cycles_count[1] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\i_core.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\data_to_write[3] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\i_core.cpu.alu_op[0] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\i_core.cpu.is_load ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\i_core.mem.instr_active ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\data_to_write[2] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\i_core.mem.q_ctrl.fsm_state[0] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\i_uart_rx.fsm_state[0] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\i_core.cpu.alu_op[2] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\data_to_write[5] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\i_core.cpu.alu_op[0] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\data_to_write[2] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\i_core.mem.q_ctrl.spi_clk_out ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\i_core.cpu.i_core.mepc[20] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\i_core.mem.q_ctrl.spi_clk_out ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\data_to_write[2] ),
    .X(net2688));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_6 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_7 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_8 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_9 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_10 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_11 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_12 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_13 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_14 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_15 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_16 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_17 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_18 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_19 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_20 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_21 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_22 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_23 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_24 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_25 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_26 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_27 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_28 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_29 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_30 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_31 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_32 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_33 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_34 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_35 (.A(clknet_0_clk_regs));
 sg13g2_antennanp ANTENNA_36 (.A(clk));
 sg13g2_antennanp ANTENNA_37 (.A(clk));
 sg13g2_antennanp ANTENNA_38 (.A(\i_core.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[27].A ));
 sg13g2_antennanp ANTENNA_39 (.A(clk));
 sg13g2_antennanp ANTENNA_40 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_fill_1 FILLER_0_268 ();
 sg13g2_fill_2 FILLER_0_279 ();
 sg13g2_fill_1 FILLER_0_337 ();
 sg13g2_fill_1 FILLER_0_375 ();
 sg13g2_fill_2 FILLER_0_389 ();
 sg13g2_fill_1 FILLER_0_391 ();
 sg13g2_fill_2 FILLER_0_396 ();
 sg13g2_fill_1 FILLER_0_398 ();
 sg13g2_decap_4 FILLER_0_438 ();
 sg13g2_decap_4 FILLER_0_542 ();
 sg13g2_decap_8 FILLER_0_550 ();
 sg13g2_fill_1 FILLER_0_557 ();
 sg13g2_decap_8 FILLER_0_562 ();
 sg13g2_decap_8 FILLER_0_569 ();
 sg13g2_decap_8 FILLER_0_576 ();
 sg13g2_decap_8 FILLER_0_583 ();
 sg13g2_decap_8 FILLER_0_590 ();
 sg13g2_decap_8 FILLER_0_597 ();
 sg13g2_decap_8 FILLER_0_604 ();
 sg13g2_decap_8 FILLER_0_611 ();
 sg13g2_decap_8 FILLER_0_618 ();
 sg13g2_decap_8 FILLER_0_625 ();
 sg13g2_decap_8 FILLER_0_632 ();
 sg13g2_decap_8 FILLER_0_639 ();
 sg13g2_decap_8 FILLER_0_646 ();
 sg13g2_decap_8 FILLER_0_653 ();
 sg13g2_decap_8 FILLER_0_660 ();
 sg13g2_decap_8 FILLER_0_667 ();
 sg13g2_decap_8 FILLER_0_674 ();
 sg13g2_decap_8 FILLER_0_681 ();
 sg13g2_decap_8 FILLER_0_688 ();
 sg13g2_decap_8 FILLER_0_695 ();
 sg13g2_decap_8 FILLER_0_702 ();
 sg13g2_decap_8 FILLER_0_709 ();
 sg13g2_decap_8 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_723 ();
 sg13g2_decap_8 FILLER_0_730 ();
 sg13g2_decap_8 FILLER_0_737 ();
 sg13g2_decap_8 FILLER_0_744 ();
 sg13g2_decap_8 FILLER_0_751 ();
 sg13g2_decap_8 FILLER_0_758 ();
 sg13g2_decap_8 FILLER_0_765 ();
 sg13g2_decap_8 FILLER_0_772 ();
 sg13g2_decap_8 FILLER_0_779 ();
 sg13g2_decap_8 FILLER_0_786 ();
 sg13g2_decap_4 FILLER_0_793 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_4 FILLER_0_808 ();
 sg13g2_fill_1 FILLER_0_812 ();
 sg13g2_decap_4 FILLER_0_826 ();
 sg13g2_fill_2 FILLER_0_830 ();
 sg13g2_fill_1 FILLER_0_940 ();
 sg13g2_decap_8 FILLER_0_958 ();
 sg13g2_decap_8 FILLER_0_965 ();
 sg13g2_decap_8 FILLER_0_972 ();
 sg13g2_decap_8 FILLER_0_979 ();
 sg13g2_decap_8 FILLER_0_986 ();
 sg13g2_decap_8 FILLER_0_993 ();
 sg13g2_decap_8 FILLER_0_1000 ();
 sg13g2_decap_8 FILLER_0_1007 ();
 sg13g2_decap_8 FILLER_0_1014 ();
 sg13g2_decap_8 FILLER_0_1021 ();
 sg13g2_decap_8 FILLER_0_1028 ();
 sg13g2_decap_8 FILLER_0_1035 ();
 sg13g2_decap_8 FILLER_0_1042 ();
 sg13g2_decap_8 FILLER_0_1049 ();
 sg13g2_decap_8 FILLER_0_1056 ();
 sg13g2_decap_8 FILLER_0_1063 ();
 sg13g2_decap_8 FILLER_0_1070 ();
 sg13g2_decap_8 FILLER_0_1077 ();
 sg13g2_decap_8 FILLER_0_1084 ();
 sg13g2_decap_8 FILLER_0_1091 ();
 sg13g2_decap_8 FILLER_0_1098 ();
 sg13g2_decap_8 FILLER_0_1105 ();
 sg13g2_decap_8 FILLER_0_1112 ();
 sg13g2_decap_8 FILLER_0_1119 ();
 sg13g2_decap_8 FILLER_0_1126 ();
 sg13g2_decap_8 FILLER_0_1133 ();
 sg13g2_decap_8 FILLER_0_1140 ();
 sg13g2_decap_8 FILLER_0_1147 ();
 sg13g2_decap_8 FILLER_0_1154 ();
 sg13g2_decap_8 FILLER_0_1161 ();
 sg13g2_decap_8 FILLER_0_1168 ();
 sg13g2_decap_8 FILLER_0_1175 ();
 sg13g2_decap_8 FILLER_0_1182 ();
 sg13g2_decap_8 FILLER_0_1189 ();
 sg13g2_decap_8 FILLER_0_1196 ();
 sg13g2_decap_8 FILLER_0_1203 ();
 sg13g2_decap_8 FILLER_0_1210 ();
 sg13g2_decap_8 FILLER_0_1217 ();
 sg13g2_decap_8 FILLER_0_1224 ();
 sg13g2_decap_8 FILLER_0_1231 ();
 sg13g2_decap_8 FILLER_0_1238 ();
 sg13g2_decap_8 FILLER_0_1245 ();
 sg13g2_decap_8 FILLER_0_1252 ();
 sg13g2_decap_8 FILLER_0_1259 ();
 sg13g2_decap_8 FILLER_0_1266 ();
 sg13g2_decap_8 FILLER_0_1273 ();
 sg13g2_decap_8 FILLER_0_1280 ();
 sg13g2_decap_8 FILLER_0_1287 ();
 sg13g2_decap_8 FILLER_0_1294 ();
 sg13g2_decap_8 FILLER_0_1301 ();
 sg13g2_decap_8 FILLER_0_1308 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_fill_2 FILLER_1_175 ();
 sg13g2_fill_1 FILLER_1_177 ();
 sg13g2_fill_2 FILLER_1_243 ();
 sg13g2_fill_1 FILLER_1_245 ();
 sg13g2_fill_2 FILLER_1_324 ();
 sg13g2_fill_1 FILLER_1_352 ();
 sg13g2_fill_2 FILLER_1_379 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_fill_1 FILLER_1_409 ();
 sg13g2_fill_2 FILLER_1_475 ();
 sg13g2_decap_4 FILLER_1_499 ();
 sg13g2_fill_1 FILLER_1_512 ();
 sg13g2_decap_8 FILLER_1_577 ();
 sg13g2_decap_4 FILLER_1_584 ();
 sg13g2_decap_8 FILLER_1_592 ();
 sg13g2_decap_8 FILLER_1_599 ();
 sg13g2_decap_8 FILLER_1_610 ();
 sg13g2_decap_8 FILLER_1_617 ();
 sg13g2_decap_8 FILLER_1_624 ();
 sg13g2_decap_8 FILLER_1_631 ();
 sg13g2_decap_4 FILLER_1_638 ();
 sg13g2_decap_8 FILLER_1_646 ();
 sg13g2_decap_8 FILLER_1_653 ();
 sg13g2_decap_8 FILLER_1_660 ();
 sg13g2_decap_4 FILLER_1_667 ();
 sg13g2_decap_8 FILLER_1_675 ();
 sg13g2_decap_8 FILLER_1_682 ();
 sg13g2_decap_8 FILLER_1_689 ();
 sg13g2_decap_8 FILLER_1_696 ();
 sg13g2_decap_8 FILLER_1_703 ();
 sg13g2_decap_8 FILLER_1_710 ();
 sg13g2_decap_8 FILLER_1_717 ();
 sg13g2_decap_8 FILLER_1_724 ();
 sg13g2_decap_8 FILLER_1_731 ();
 sg13g2_decap_4 FILLER_1_738 ();
 sg13g2_fill_1 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_747 ();
 sg13g2_decap_8 FILLER_1_754 ();
 sg13g2_decap_8 FILLER_1_761 ();
 sg13g2_decap_8 FILLER_1_768 ();
 sg13g2_decap_8 FILLER_1_775 ();
 sg13g2_decap_4 FILLER_1_782 ();
 sg13g2_fill_1 FILLER_1_786 ();
 sg13g2_fill_1 FILLER_1_857 ();
 sg13g2_fill_1 FILLER_1_913 ();
 sg13g2_fill_2 FILLER_1_939 ();
 sg13g2_fill_2 FILLER_1_967 ();
 sg13g2_decap_8 FILLER_1_995 ();
 sg13g2_decap_8 FILLER_1_1002 ();
 sg13g2_decap_8 FILLER_1_1009 ();
 sg13g2_decap_8 FILLER_1_1016 ();
 sg13g2_decap_8 FILLER_1_1023 ();
 sg13g2_decap_8 FILLER_1_1030 ();
 sg13g2_decap_8 FILLER_1_1037 ();
 sg13g2_decap_8 FILLER_1_1044 ();
 sg13g2_decap_8 FILLER_1_1051 ();
 sg13g2_decap_8 FILLER_1_1058 ();
 sg13g2_decap_8 FILLER_1_1065 ();
 sg13g2_decap_8 FILLER_1_1072 ();
 sg13g2_decap_8 FILLER_1_1079 ();
 sg13g2_decap_8 FILLER_1_1086 ();
 sg13g2_decap_8 FILLER_1_1093 ();
 sg13g2_decap_8 FILLER_1_1100 ();
 sg13g2_decap_8 FILLER_1_1107 ();
 sg13g2_decap_8 FILLER_1_1114 ();
 sg13g2_decap_8 FILLER_1_1121 ();
 sg13g2_decap_8 FILLER_1_1128 ();
 sg13g2_decap_8 FILLER_1_1135 ();
 sg13g2_decap_8 FILLER_1_1142 ();
 sg13g2_decap_8 FILLER_1_1149 ();
 sg13g2_decap_8 FILLER_1_1156 ();
 sg13g2_decap_8 FILLER_1_1163 ();
 sg13g2_decap_8 FILLER_1_1170 ();
 sg13g2_decap_8 FILLER_1_1177 ();
 sg13g2_decap_8 FILLER_1_1184 ();
 sg13g2_decap_8 FILLER_1_1191 ();
 sg13g2_decap_8 FILLER_1_1198 ();
 sg13g2_decap_8 FILLER_1_1205 ();
 sg13g2_decap_8 FILLER_1_1212 ();
 sg13g2_decap_8 FILLER_1_1219 ();
 sg13g2_decap_8 FILLER_1_1226 ();
 sg13g2_decap_8 FILLER_1_1233 ();
 sg13g2_decap_8 FILLER_1_1240 ();
 sg13g2_decap_8 FILLER_1_1247 ();
 sg13g2_decap_8 FILLER_1_1254 ();
 sg13g2_decap_8 FILLER_1_1261 ();
 sg13g2_decap_8 FILLER_1_1268 ();
 sg13g2_decap_8 FILLER_1_1275 ();
 sg13g2_decap_8 FILLER_1_1282 ();
 sg13g2_decap_8 FILLER_1_1289 ();
 sg13g2_decap_8 FILLER_1_1296 ();
 sg13g2_decap_8 FILLER_1_1303 ();
 sg13g2_decap_4 FILLER_1_1310 ();
 sg13g2_fill_1 FILLER_1_1314 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_fill_2 FILLER_2_214 ();
 sg13g2_fill_2 FILLER_2_240 ();
 sg13g2_fill_1 FILLER_2_242 ();
 sg13g2_fill_2 FILLER_2_298 ();
 sg13g2_fill_1 FILLER_2_300 ();
 sg13g2_fill_2 FILLER_2_340 ();
 sg13g2_fill_1 FILLER_2_355 ();
 sg13g2_fill_2 FILLER_2_409 ();
 sg13g2_fill_1 FILLER_2_411 ();
 sg13g2_fill_2 FILLER_2_425 ();
 sg13g2_fill_2 FILLER_2_453 ();
 sg13g2_fill_1 FILLER_2_455 ();
 sg13g2_fill_2 FILLER_2_526 ();
 sg13g2_fill_1 FILLER_2_528 ();
 sg13g2_fill_1 FILLER_2_612 ();
 sg13g2_fill_1 FILLER_2_648 ();
 sg13g2_decap_4 FILLER_2_688 ();
 sg13g2_fill_1 FILLER_2_692 ();
 sg13g2_decap_8 FILLER_2_706 ();
 sg13g2_decap_8 FILLER_2_713 ();
 sg13g2_decap_8 FILLER_2_720 ();
 sg13g2_fill_1 FILLER_2_727 ();
 sg13g2_fill_2 FILLER_2_758 ();
 sg13g2_decap_8 FILLER_2_769 ();
 sg13g2_decap_4 FILLER_2_776 ();
 sg13g2_fill_2 FILLER_2_784 ();
 sg13g2_fill_2 FILLER_2_842 ();
 sg13g2_fill_1 FILLER_2_844 ();
 sg13g2_fill_1 FILLER_2_901 ();
 sg13g2_fill_2 FILLER_2_919 ();
 sg13g2_fill_1 FILLER_2_926 ();
 sg13g2_decap_8 FILLER_2_979 ();
 sg13g2_decap_8 FILLER_2_995 ();
 sg13g2_decap_8 FILLER_2_1002 ();
 sg13g2_decap_8 FILLER_2_1009 ();
 sg13g2_decap_8 FILLER_2_1016 ();
 sg13g2_decap_8 FILLER_2_1023 ();
 sg13g2_decap_8 FILLER_2_1030 ();
 sg13g2_decap_8 FILLER_2_1037 ();
 sg13g2_decap_8 FILLER_2_1044 ();
 sg13g2_decap_8 FILLER_2_1051 ();
 sg13g2_decap_8 FILLER_2_1058 ();
 sg13g2_decap_8 FILLER_2_1065 ();
 sg13g2_decap_8 FILLER_2_1072 ();
 sg13g2_decap_8 FILLER_2_1079 ();
 sg13g2_decap_8 FILLER_2_1086 ();
 sg13g2_decap_8 FILLER_2_1093 ();
 sg13g2_decap_8 FILLER_2_1100 ();
 sg13g2_decap_8 FILLER_2_1107 ();
 sg13g2_decap_8 FILLER_2_1114 ();
 sg13g2_decap_8 FILLER_2_1121 ();
 sg13g2_decap_8 FILLER_2_1128 ();
 sg13g2_decap_8 FILLER_2_1135 ();
 sg13g2_decap_8 FILLER_2_1142 ();
 sg13g2_decap_8 FILLER_2_1149 ();
 sg13g2_decap_8 FILLER_2_1156 ();
 sg13g2_decap_8 FILLER_2_1163 ();
 sg13g2_decap_8 FILLER_2_1170 ();
 sg13g2_decap_8 FILLER_2_1177 ();
 sg13g2_decap_8 FILLER_2_1184 ();
 sg13g2_decap_8 FILLER_2_1191 ();
 sg13g2_decap_8 FILLER_2_1198 ();
 sg13g2_decap_8 FILLER_2_1205 ();
 sg13g2_decap_8 FILLER_2_1212 ();
 sg13g2_decap_8 FILLER_2_1219 ();
 sg13g2_decap_8 FILLER_2_1226 ();
 sg13g2_decap_8 FILLER_2_1233 ();
 sg13g2_decap_8 FILLER_2_1240 ();
 sg13g2_decap_8 FILLER_2_1247 ();
 sg13g2_decap_8 FILLER_2_1254 ();
 sg13g2_decap_8 FILLER_2_1261 ();
 sg13g2_decap_8 FILLER_2_1268 ();
 sg13g2_decap_8 FILLER_2_1275 ();
 sg13g2_decap_8 FILLER_2_1282 ();
 sg13g2_decap_8 FILLER_2_1289 ();
 sg13g2_decap_8 FILLER_2_1296 ();
 sg13g2_decap_8 FILLER_2_1303 ();
 sg13g2_decap_4 FILLER_2_1310 ();
 sg13g2_fill_1 FILLER_2_1314 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_4 FILLER_3_140 ();
 sg13g2_fill_2 FILLER_3_144 ();
 sg13g2_decap_4 FILLER_3_150 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_fill_1 FILLER_3_168 ();
 sg13g2_fill_2 FILLER_3_193 ();
 sg13g2_fill_1 FILLER_3_275 ();
 sg13g2_fill_2 FILLER_3_287 ();
 sg13g2_fill_1 FILLER_3_307 ();
 sg13g2_fill_2 FILLER_3_358 ();
 sg13g2_fill_2 FILLER_3_379 ();
 sg13g2_fill_2 FILLER_3_472 ();
 sg13g2_fill_1 FILLER_3_474 ();
 sg13g2_decap_8 FILLER_3_487 ();
 sg13g2_fill_2 FILLER_3_494 ();
 sg13g2_fill_1 FILLER_3_496 ();
 sg13g2_decap_8 FILLER_3_501 ();
 sg13g2_fill_1 FILLER_3_534 ();
 sg13g2_fill_2 FILLER_3_587 ();
 sg13g2_fill_1 FILLER_3_589 ();
 sg13g2_fill_1 FILLER_3_594 ();
 sg13g2_fill_1 FILLER_3_630 ();
 sg13g2_fill_1 FILLER_3_666 ();
 sg13g2_fill_2 FILLER_3_810 ();
 sg13g2_fill_2 FILLER_3_878 ();
 sg13g2_decap_8 FILLER_3_997 ();
 sg13g2_decap_8 FILLER_3_1004 ();
 sg13g2_decap_8 FILLER_3_1011 ();
 sg13g2_decap_8 FILLER_3_1018 ();
 sg13g2_decap_8 FILLER_3_1025 ();
 sg13g2_decap_8 FILLER_3_1032 ();
 sg13g2_decap_8 FILLER_3_1039 ();
 sg13g2_decap_8 FILLER_3_1046 ();
 sg13g2_decap_8 FILLER_3_1053 ();
 sg13g2_decap_8 FILLER_3_1060 ();
 sg13g2_decap_8 FILLER_3_1067 ();
 sg13g2_decap_8 FILLER_3_1074 ();
 sg13g2_decap_8 FILLER_3_1081 ();
 sg13g2_decap_8 FILLER_3_1088 ();
 sg13g2_decap_8 FILLER_3_1095 ();
 sg13g2_decap_8 FILLER_3_1102 ();
 sg13g2_decap_8 FILLER_3_1109 ();
 sg13g2_decap_8 FILLER_3_1116 ();
 sg13g2_decap_8 FILLER_3_1123 ();
 sg13g2_decap_8 FILLER_3_1130 ();
 sg13g2_decap_8 FILLER_3_1137 ();
 sg13g2_decap_8 FILLER_3_1144 ();
 sg13g2_decap_8 FILLER_3_1151 ();
 sg13g2_decap_8 FILLER_3_1158 ();
 sg13g2_decap_8 FILLER_3_1165 ();
 sg13g2_decap_8 FILLER_3_1172 ();
 sg13g2_decap_8 FILLER_3_1179 ();
 sg13g2_decap_8 FILLER_3_1186 ();
 sg13g2_decap_8 FILLER_3_1193 ();
 sg13g2_decap_8 FILLER_3_1200 ();
 sg13g2_decap_8 FILLER_3_1207 ();
 sg13g2_decap_8 FILLER_3_1214 ();
 sg13g2_decap_8 FILLER_3_1221 ();
 sg13g2_decap_8 FILLER_3_1228 ();
 sg13g2_decap_8 FILLER_3_1235 ();
 sg13g2_decap_8 FILLER_3_1242 ();
 sg13g2_decap_8 FILLER_3_1249 ();
 sg13g2_decap_8 FILLER_3_1256 ();
 sg13g2_decap_8 FILLER_3_1263 ();
 sg13g2_decap_8 FILLER_3_1270 ();
 sg13g2_decap_8 FILLER_3_1277 ();
 sg13g2_decap_8 FILLER_3_1284 ();
 sg13g2_decap_8 FILLER_3_1291 ();
 sg13g2_decap_8 FILLER_3_1298 ();
 sg13g2_decap_8 FILLER_3_1305 ();
 sg13g2_fill_2 FILLER_3_1312 ();
 sg13g2_fill_1 FILLER_3_1314 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_4 FILLER_4_133 ();
 sg13g2_fill_1 FILLER_4_137 ();
 sg13g2_fill_2 FILLER_4_152 ();
 sg13g2_fill_1 FILLER_4_154 ();
 sg13g2_fill_2 FILLER_4_455 ();
 sg13g2_fill_2 FILLER_4_492 ();
 sg13g2_fill_1 FILLER_4_494 ();
 sg13g2_fill_2 FILLER_4_521 ();
 sg13g2_fill_1 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_605 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_fill_2 FILLER_4_675 ();
 sg13g2_fill_1 FILLER_4_677 ();
 sg13g2_decap_4 FILLER_4_730 ();
 sg13g2_fill_1 FILLER_4_734 ();
 sg13g2_fill_2 FILLER_4_762 ();
 sg13g2_fill_1 FILLER_4_764 ();
 sg13g2_decap_4 FILLER_4_821 ();
 sg13g2_fill_1 FILLER_4_825 ();
 sg13g2_fill_2 FILLER_4_896 ();
 sg13g2_decap_8 FILLER_4_1002 ();
 sg13g2_decap_8 FILLER_4_1009 ();
 sg13g2_decap_8 FILLER_4_1016 ();
 sg13g2_decap_8 FILLER_4_1023 ();
 sg13g2_decap_8 FILLER_4_1030 ();
 sg13g2_decap_8 FILLER_4_1037 ();
 sg13g2_decap_8 FILLER_4_1044 ();
 sg13g2_decap_8 FILLER_4_1051 ();
 sg13g2_decap_8 FILLER_4_1058 ();
 sg13g2_decap_8 FILLER_4_1065 ();
 sg13g2_decap_8 FILLER_4_1072 ();
 sg13g2_decap_8 FILLER_4_1079 ();
 sg13g2_decap_8 FILLER_4_1086 ();
 sg13g2_decap_8 FILLER_4_1093 ();
 sg13g2_decap_8 FILLER_4_1100 ();
 sg13g2_decap_8 FILLER_4_1107 ();
 sg13g2_decap_8 FILLER_4_1114 ();
 sg13g2_decap_8 FILLER_4_1121 ();
 sg13g2_decap_8 FILLER_4_1128 ();
 sg13g2_decap_8 FILLER_4_1135 ();
 sg13g2_decap_8 FILLER_4_1142 ();
 sg13g2_decap_8 FILLER_4_1149 ();
 sg13g2_decap_8 FILLER_4_1156 ();
 sg13g2_decap_8 FILLER_4_1163 ();
 sg13g2_decap_8 FILLER_4_1170 ();
 sg13g2_decap_8 FILLER_4_1177 ();
 sg13g2_decap_8 FILLER_4_1184 ();
 sg13g2_decap_8 FILLER_4_1191 ();
 sg13g2_decap_8 FILLER_4_1198 ();
 sg13g2_decap_8 FILLER_4_1205 ();
 sg13g2_decap_8 FILLER_4_1212 ();
 sg13g2_decap_8 FILLER_4_1219 ();
 sg13g2_decap_8 FILLER_4_1226 ();
 sg13g2_decap_8 FILLER_4_1233 ();
 sg13g2_decap_8 FILLER_4_1240 ();
 sg13g2_decap_8 FILLER_4_1247 ();
 sg13g2_decap_8 FILLER_4_1254 ();
 sg13g2_decap_8 FILLER_4_1261 ();
 sg13g2_decap_8 FILLER_4_1268 ();
 sg13g2_decap_8 FILLER_4_1275 ();
 sg13g2_decap_8 FILLER_4_1282 ();
 sg13g2_decap_8 FILLER_4_1289 ();
 sg13g2_decap_8 FILLER_4_1296 ();
 sg13g2_decap_8 FILLER_4_1303 ();
 sg13g2_decap_4 FILLER_4_1310 ();
 sg13g2_fill_1 FILLER_4_1314 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_165 ();
 sg13g2_fill_2 FILLER_5_239 ();
 sg13g2_fill_2 FILLER_5_251 ();
 sg13g2_fill_1 FILLER_5_253 ();
 sg13g2_fill_2 FILLER_5_307 ();
 sg13g2_fill_1 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_4 FILLER_5_392 ();
 sg13g2_fill_1 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_421 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_fill_1 FILLER_5_430 ();
 sg13g2_decap_8 FILLER_5_435 ();
 sg13g2_fill_1 FILLER_5_442 ();
 sg13g2_fill_2 FILLER_5_647 ();
 sg13g2_fill_2 FILLER_5_693 ();
 sg13g2_fill_2 FILLER_5_791 ();
 sg13g2_fill_1 FILLER_5_793 ();
 sg13g2_fill_2 FILLER_5_803 ();
 sg13g2_fill_2 FILLER_5_836 ();
 sg13g2_fill_1 FILLER_5_838 ();
 sg13g2_decap_8 FILLER_5_908 ();
 sg13g2_fill_1 FILLER_5_915 ();
 sg13g2_fill_2 FILLER_5_991 ();
 sg13g2_decap_8 FILLER_5_1010 ();
 sg13g2_decap_8 FILLER_5_1017 ();
 sg13g2_decap_8 FILLER_5_1024 ();
 sg13g2_decap_8 FILLER_5_1031 ();
 sg13g2_decap_8 FILLER_5_1038 ();
 sg13g2_decap_8 FILLER_5_1045 ();
 sg13g2_decap_8 FILLER_5_1052 ();
 sg13g2_decap_8 FILLER_5_1059 ();
 sg13g2_decap_8 FILLER_5_1066 ();
 sg13g2_decap_8 FILLER_5_1073 ();
 sg13g2_decap_8 FILLER_5_1080 ();
 sg13g2_decap_8 FILLER_5_1087 ();
 sg13g2_decap_8 FILLER_5_1094 ();
 sg13g2_decap_8 FILLER_5_1101 ();
 sg13g2_decap_8 FILLER_5_1108 ();
 sg13g2_decap_8 FILLER_5_1115 ();
 sg13g2_decap_8 FILLER_5_1122 ();
 sg13g2_decap_8 FILLER_5_1129 ();
 sg13g2_decap_8 FILLER_5_1136 ();
 sg13g2_decap_8 FILLER_5_1143 ();
 sg13g2_decap_8 FILLER_5_1150 ();
 sg13g2_decap_8 FILLER_5_1157 ();
 sg13g2_decap_8 FILLER_5_1164 ();
 sg13g2_decap_8 FILLER_5_1171 ();
 sg13g2_decap_8 FILLER_5_1178 ();
 sg13g2_decap_8 FILLER_5_1185 ();
 sg13g2_decap_8 FILLER_5_1192 ();
 sg13g2_decap_8 FILLER_5_1199 ();
 sg13g2_decap_8 FILLER_5_1206 ();
 sg13g2_decap_8 FILLER_5_1213 ();
 sg13g2_decap_8 FILLER_5_1220 ();
 sg13g2_decap_8 FILLER_5_1227 ();
 sg13g2_decap_8 FILLER_5_1234 ();
 sg13g2_decap_8 FILLER_5_1241 ();
 sg13g2_decap_8 FILLER_5_1248 ();
 sg13g2_decap_8 FILLER_5_1255 ();
 sg13g2_decap_8 FILLER_5_1262 ();
 sg13g2_decap_8 FILLER_5_1269 ();
 sg13g2_decap_8 FILLER_5_1276 ();
 sg13g2_decap_8 FILLER_5_1283 ();
 sg13g2_decap_8 FILLER_5_1290 ();
 sg13g2_decap_8 FILLER_5_1297 ();
 sg13g2_decap_8 FILLER_5_1304 ();
 sg13g2_decap_4 FILLER_5_1311 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_fill_2 FILLER_6_119 ();
 sg13g2_fill_1 FILLER_6_294 ();
 sg13g2_fill_2 FILLER_6_384 ();
 sg13g2_fill_2 FILLER_6_412 ();
 sg13g2_fill_1 FILLER_6_414 ();
 sg13g2_fill_2 FILLER_6_419 ();
 sg13g2_fill_1 FILLER_6_421 ();
 sg13g2_decap_8 FILLER_6_433 ();
 sg13g2_fill_2 FILLER_6_448 ();
 sg13g2_fill_1 FILLER_6_480 ();
 sg13g2_decap_4 FILLER_6_487 ();
 sg13g2_fill_1 FILLER_6_491 ();
 sg13g2_fill_2 FILLER_6_501 ();
 sg13g2_fill_1 FILLER_6_503 ();
 sg13g2_decap_4 FILLER_6_508 ();
 sg13g2_fill_2 FILLER_6_512 ();
 sg13g2_fill_1 FILLER_6_527 ();
 sg13g2_fill_2 FILLER_6_536 ();
 sg13g2_fill_1 FILLER_6_538 ();
 sg13g2_fill_2 FILLER_6_557 ();
 sg13g2_fill_2 FILLER_6_598 ();
 sg13g2_fill_1 FILLER_6_661 ();
 sg13g2_fill_2 FILLER_6_671 ();
 sg13g2_fill_2 FILLER_6_704 ();
 sg13g2_fill_1 FILLER_6_706 ();
 sg13g2_fill_2 FILLER_6_741 ();
 sg13g2_fill_1 FILLER_6_743 ();
 sg13g2_fill_2 FILLER_6_848 ();
 sg13g2_fill_2 FILLER_6_868 ();
 sg13g2_fill_1 FILLER_6_870 ();
 sg13g2_fill_1 FILLER_6_902 ();
 sg13g2_decap_8 FILLER_6_1007 ();
 sg13g2_decap_8 FILLER_6_1014 ();
 sg13g2_decap_8 FILLER_6_1021 ();
 sg13g2_decap_8 FILLER_6_1028 ();
 sg13g2_decap_8 FILLER_6_1035 ();
 sg13g2_decap_8 FILLER_6_1042 ();
 sg13g2_decap_8 FILLER_6_1049 ();
 sg13g2_decap_8 FILLER_6_1056 ();
 sg13g2_decap_8 FILLER_6_1063 ();
 sg13g2_decap_8 FILLER_6_1070 ();
 sg13g2_decap_8 FILLER_6_1077 ();
 sg13g2_decap_8 FILLER_6_1084 ();
 sg13g2_decap_8 FILLER_6_1091 ();
 sg13g2_decap_8 FILLER_6_1098 ();
 sg13g2_decap_8 FILLER_6_1105 ();
 sg13g2_decap_8 FILLER_6_1112 ();
 sg13g2_decap_8 FILLER_6_1119 ();
 sg13g2_decap_8 FILLER_6_1126 ();
 sg13g2_decap_8 FILLER_6_1133 ();
 sg13g2_decap_8 FILLER_6_1140 ();
 sg13g2_decap_8 FILLER_6_1147 ();
 sg13g2_decap_8 FILLER_6_1154 ();
 sg13g2_decap_8 FILLER_6_1161 ();
 sg13g2_decap_8 FILLER_6_1168 ();
 sg13g2_decap_8 FILLER_6_1175 ();
 sg13g2_decap_8 FILLER_6_1182 ();
 sg13g2_decap_8 FILLER_6_1189 ();
 sg13g2_decap_8 FILLER_6_1196 ();
 sg13g2_decap_8 FILLER_6_1203 ();
 sg13g2_decap_8 FILLER_6_1210 ();
 sg13g2_decap_8 FILLER_6_1217 ();
 sg13g2_decap_8 FILLER_6_1224 ();
 sg13g2_decap_8 FILLER_6_1231 ();
 sg13g2_decap_8 FILLER_6_1238 ();
 sg13g2_decap_8 FILLER_6_1245 ();
 sg13g2_decap_8 FILLER_6_1252 ();
 sg13g2_decap_8 FILLER_6_1259 ();
 sg13g2_decap_8 FILLER_6_1266 ();
 sg13g2_decap_8 FILLER_6_1273 ();
 sg13g2_decap_8 FILLER_6_1280 ();
 sg13g2_decap_8 FILLER_6_1287 ();
 sg13g2_decap_8 FILLER_6_1294 ();
 sg13g2_decap_8 FILLER_6_1301 ();
 sg13g2_decap_8 FILLER_6_1308 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_147 ();
 sg13g2_fill_2 FILLER_7_163 ();
 sg13g2_fill_1 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_199 ();
 sg13g2_fill_2 FILLER_7_230 ();
 sg13g2_fill_1 FILLER_7_232 ();
 sg13g2_fill_2 FILLER_7_247 ();
 sg13g2_fill_1 FILLER_7_258 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_288 ();
 sg13g2_fill_2 FILLER_7_294 ();
 sg13g2_fill_1 FILLER_7_301 ();
 sg13g2_fill_2 FILLER_7_324 ();
 sg13g2_fill_2 FILLER_7_339 ();
 sg13g2_fill_1 FILLER_7_341 ();
 sg13g2_fill_1 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_4 FILLER_7_394 ();
 sg13g2_fill_2 FILLER_7_410 ();
 sg13g2_fill_1 FILLER_7_412 ();
 sg13g2_fill_1 FILLER_7_418 ();
 sg13g2_decap_4 FILLER_7_431 ();
 sg13g2_fill_2 FILLER_7_451 ();
 sg13g2_fill_2 FILLER_7_480 ();
 sg13g2_fill_1 FILLER_7_491 ();
 sg13g2_fill_2 FILLER_7_510 ();
 sg13g2_fill_1 FILLER_7_512 ();
 sg13g2_fill_2 FILLER_7_547 ();
 sg13g2_decap_8 FILLER_7_557 ();
 sg13g2_decap_4 FILLER_7_573 ();
 sg13g2_fill_2 FILLER_7_638 ();
 sg13g2_fill_1 FILLER_7_683 ();
 sg13g2_fill_2 FILLER_7_701 ();
 sg13g2_fill_1 FILLER_7_703 ();
 sg13g2_fill_2 FILLER_7_716 ();
 sg13g2_fill_1 FILLER_7_718 ();
 sg13g2_fill_1 FILLER_7_750 ();
 sg13g2_fill_1 FILLER_7_849 ();
 sg13g2_fill_2 FILLER_7_876 ();
 sg13g2_fill_1 FILLER_7_878 ();
 sg13g2_decap_8 FILLER_7_897 ();
 sg13g2_fill_1 FILLER_7_904 ();
 sg13g2_decap_8 FILLER_7_1005 ();
 sg13g2_decap_8 FILLER_7_1012 ();
 sg13g2_decap_8 FILLER_7_1019 ();
 sg13g2_decap_8 FILLER_7_1026 ();
 sg13g2_decap_8 FILLER_7_1033 ();
 sg13g2_decap_8 FILLER_7_1040 ();
 sg13g2_decap_8 FILLER_7_1047 ();
 sg13g2_decap_8 FILLER_7_1054 ();
 sg13g2_decap_8 FILLER_7_1061 ();
 sg13g2_decap_8 FILLER_7_1068 ();
 sg13g2_decap_8 FILLER_7_1075 ();
 sg13g2_decap_8 FILLER_7_1082 ();
 sg13g2_decap_8 FILLER_7_1089 ();
 sg13g2_decap_8 FILLER_7_1096 ();
 sg13g2_decap_8 FILLER_7_1103 ();
 sg13g2_decap_8 FILLER_7_1110 ();
 sg13g2_decap_8 FILLER_7_1117 ();
 sg13g2_decap_8 FILLER_7_1124 ();
 sg13g2_decap_8 FILLER_7_1131 ();
 sg13g2_decap_8 FILLER_7_1138 ();
 sg13g2_decap_8 FILLER_7_1145 ();
 sg13g2_decap_8 FILLER_7_1152 ();
 sg13g2_decap_8 FILLER_7_1159 ();
 sg13g2_decap_8 FILLER_7_1166 ();
 sg13g2_decap_8 FILLER_7_1173 ();
 sg13g2_decap_8 FILLER_7_1180 ();
 sg13g2_decap_8 FILLER_7_1187 ();
 sg13g2_decap_8 FILLER_7_1194 ();
 sg13g2_decap_8 FILLER_7_1201 ();
 sg13g2_decap_8 FILLER_7_1208 ();
 sg13g2_decap_8 FILLER_7_1215 ();
 sg13g2_decap_8 FILLER_7_1222 ();
 sg13g2_decap_8 FILLER_7_1229 ();
 sg13g2_decap_8 FILLER_7_1236 ();
 sg13g2_decap_8 FILLER_7_1243 ();
 sg13g2_decap_8 FILLER_7_1250 ();
 sg13g2_decap_8 FILLER_7_1257 ();
 sg13g2_decap_8 FILLER_7_1264 ();
 sg13g2_decap_8 FILLER_7_1271 ();
 sg13g2_decap_8 FILLER_7_1278 ();
 sg13g2_decap_8 FILLER_7_1285 ();
 sg13g2_decap_8 FILLER_7_1292 ();
 sg13g2_decap_8 FILLER_7_1299 ();
 sg13g2_decap_8 FILLER_7_1306 ();
 sg13g2_fill_2 FILLER_7_1313 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_fill_1 FILLER_8_112 ();
 sg13g2_fill_1 FILLER_8_144 ();
 sg13g2_fill_1 FILLER_8_226 ();
 sg13g2_fill_2 FILLER_8_274 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_fill_2 FILLER_8_330 ();
 sg13g2_fill_1 FILLER_8_332 ();
 sg13g2_fill_2 FILLER_8_352 ();
 sg13g2_fill_1 FILLER_8_367 ();
 sg13g2_fill_1 FILLER_8_373 ();
 sg13g2_decap_4 FILLER_8_389 ();
 sg13g2_fill_2 FILLER_8_393 ();
 sg13g2_decap_4 FILLER_8_426 ();
 sg13g2_fill_2 FILLER_8_453 ();
 sg13g2_fill_1 FILLER_8_455 ();
 sg13g2_fill_2 FILLER_8_495 ();
 sg13g2_fill_1 FILLER_8_497 ();
 sg13g2_fill_2 FILLER_8_513 ();
 sg13g2_fill_1 FILLER_8_515 ();
 sg13g2_fill_2 FILLER_8_524 ();
 sg13g2_fill_2 FILLER_8_540 ();
 sg13g2_fill_1 FILLER_8_542 ();
 sg13g2_fill_1 FILLER_8_593 ();
 sg13g2_fill_1 FILLER_8_602 ();
 sg13g2_fill_1 FILLER_8_612 ();
 sg13g2_fill_2 FILLER_8_652 ();
 sg13g2_fill_1 FILLER_8_723 ();
 sg13g2_fill_2 FILLER_8_733 ();
 sg13g2_fill_1 FILLER_8_770 ();
 sg13g2_fill_2 FILLER_8_808 ();
 sg13g2_fill_1 FILLER_8_810 ();
 sg13g2_fill_2 FILLER_8_821 ();
 sg13g2_fill_1 FILLER_8_823 ();
 sg13g2_fill_2 FILLER_8_850 ();
 sg13g2_fill_1 FILLER_8_878 ();
 sg13g2_fill_1 FILLER_8_923 ();
 sg13g2_fill_2 FILLER_8_936 ();
 sg13g2_fill_1 FILLER_8_938 ();
 sg13g2_decap_8 FILLER_8_1009 ();
 sg13g2_decap_8 FILLER_8_1016 ();
 sg13g2_decap_8 FILLER_8_1023 ();
 sg13g2_decap_8 FILLER_8_1030 ();
 sg13g2_decap_8 FILLER_8_1037 ();
 sg13g2_decap_8 FILLER_8_1044 ();
 sg13g2_decap_8 FILLER_8_1051 ();
 sg13g2_decap_8 FILLER_8_1058 ();
 sg13g2_decap_8 FILLER_8_1065 ();
 sg13g2_decap_8 FILLER_8_1072 ();
 sg13g2_decap_8 FILLER_8_1079 ();
 sg13g2_decap_8 FILLER_8_1086 ();
 sg13g2_decap_8 FILLER_8_1093 ();
 sg13g2_decap_8 FILLER_8_1100 ();
 sg13g2_decap_8 FILLER_8_1107 ();
 sg13g2_decap_8 FILLER_8_1114 ();
 sg13g2_decap_8 FILLER_8_1121 ();
 sg13g2_decap_8 FILLER_8_1128 ();
 sg13g2_decap_8 FILLER_8_1135 ();
 sg13g2_decap_8 FILLER_8_1142 ();
 sg13g2_decap_8 FILLER_8_1149 ();
 sg13g2_decap_8 FILLER_8_1156 ();
 sg13g2_decap_8 FILLER_8_1163 ();
 sg13g2_decap_8 FILLER_8_1170 ();
 sg13g2_decap_8 FILLER_8_1177 ();
 sg13g2_decap_8 FILLER_8_1184 ();
 sg13g2_decap_8 FILLER_8_1191 ();
 sg13g2_decap_8 FILLER_8_1198 ();
 sg13g2_decap_8 FILLER_8_1205 ();
 sg13g2_decap_8 FILLER_8_1212 ();
 sg13g2_decap_8 FILLER_8_1219 ();
 sg13g2_decap_8 FILLER_8_1226 ();
 sg13g2_decap_8 FILLER_8_1233 ();
 sg13g2_decap_8 FILLER_8_1240 ();
 sg13g2_decap_8 FILLER_8_1247 ();
 sg13g2_decap_8 FILLER_8_1254 ();
 sg13g2_decap_8 FILLER_8_1261 ();
 sg13g2_decap_8 FILLER_8_1268 ();
 sg13g2_decap_8 FILLER_8_1275 ();
 sg13g2_decap_8 FILLER_8_1282 ();
 sg13g2_decap_8 FILLER_8_1289 ();
 sg13g2_decap_8 FILLER_8_1296 ();
 sg13g2_decap_8 FILLER_8_1303 ();
 sg13g2_decap_4 FILLER_8_1310 ();
 sg13g2_fill_1 FILLER_8_1314 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_4 FILLER_9_112 ();
 sg13g2_fill_2 FILLER_9_116 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_221 ();
 sg13g2_fill_2 FILLER_9_232 ();
 sg13g2_fill_2 FILLER_9_290 ();
 sg13g2_fill_1 FILLER_9_306 ();
 sg13g2_fill_2 FILLER_9_370 ();
 sg13g2_fill_1 FILLER_9_372 ();
 sg13g2_fill_2 FILLER_9_384 ();
 sg13g2_fill_1 FILLER_9_386 ();
 sg13g2_fill_2 FILLER_9_394 ();
 sg13g2_fill_1 FILLER_9_396 ();
 sg13g2_fill_1 FILLER_9_419 ();
 sg13g2_fill_2 FILLER_9_450 ();
 sg13g2_fill_1 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_458 ();
 sg13g2_decap_8 FILLER_9_465 ();
 sg13g2_fill_2 FILLER_9_472 ();
 sg13g2_fill_1 FILLER_9_474 ();
 sg13g2_decap_4 FILLER_9_485 ();
 sg13g2_fill_1 FILLER_9_489 ();
 sg13g2_decap_4 FILLER_9_519 ();
 sg13g2_decap_4 FILLER_9_554 ();
 sg13g2_decap_8 FILLER_9_562 ();
 sg13g2_fill_2 FILLER_9_569 ();
 sg13g2_fill_1 FILLER_9_571 ();
 sg13g2_fill_2 FILLER_9_633 ();
 sg13g2_fill_2 FILLER_9_692 ();
 sg13g2_fill_1 FILLER_9_694 ();
 sg13g2_fill_2 FILLER_9_760 ();
 sg13g2_fill_2 FILLER_9_766 ();
 sg13g2_fill_1 FILLER_9_768 ();
 sg13g2_fill_1 FILLER_9_851 ();
 sg13g2_fill_2 FILLER_9_861 ();
 sg13g2_fill_1 FILLER_9_871 ();
 sg13g2_fill_1 FILLER_9_881 ();
 sg13g2_fill_1 FILLER_9_887 ();
 sg13g2_fill_1 FILLER_9_897 ();
 sg13g2_fill_2 FILLER_9_907 ();
 sg13g2_fill_1 FILLER_9_999 ();
 sg13g2_decap_4 FILLER_9_1021 ();
 sg13g2_fill_1 FILLER_9_1025 ();
 sg13g2_decap_8 FILLER_9_1035 ();
 sg13g2_decap_8 FILLER_9_1042 ();
 sg13g2_fill_2 FILLER_9_1049 ();
 sg13g2_fill_1 FILLER_9_1051 ();
 sg13g2_decap_8 FILLER_9_1056 ();
 sg13g2_decap_8 FILLER_9_1063 ();
 sg13g2_decap_8 FILLER_9_1070 ();
 sg13g2_decap_8 FILLER_9_1077 ();
 sg13g2_decap_8 FILLER_9_1084 ();
 sg13g2_decap_8 FILLER_9_1091 ();
 sg13g2_decap_8 FILLER_9_1098 ();
 sg13g2_decap_8 FILLER_9_1105 ();
 sg13g2_decap_8 FILLER_9_1112 ();
 sg13g2_decap_8 FILLER_9_1119 ();
 sg13g2_decap_8 FILLER_9_1126 ();
 sg13g2_decap_8 FILLER_9_1133 ();
 sg13g2_decap_8 FILLER_9_1140 ();
 sg13g2_decap_8 FILLER_9_1147 ();
 sg13g2_decap_8 FILLER_9_1154 ();
 sg13g2_decap_8 FILLER_9_1161 ();
 sg13g2_decap_8 FILLER_9_1168 ();
 sg13g2_decap_8 FILLER_9_1175 ();
 sg13g2_decap_8 FILLER_9_1182 ();
 sg13g2_decap_8 FILLER_9_1189 ();
 sg13g2_decap_8 FILLER_9_1196 ();
 sg13g2_decap_8 FILLER_9_1203 ();
 sg13g2_decap_8 FILLER_9_1210 ();
 sg13g2_decap_8 FILLER_9_1217 ();
 sg13g2_decap_8 FILLER_9_1224 ();
 sg13g2_decap_8 FILLER_9_1231 ();
 sg13g2_decap_8 FILLER_9_1238 ();
 sg13g2_decap_8 FILLER_9_1245 ();
 sg13g2_decap_8 FILLER_9_1252 ();
 sg13g2_decap_8 FILLER_9_1259 ();
 sg13g2_decap_8 FILLER_9_1266 ();
 sg13g2_decap_8 FILLER_9_1273 ();
 sg13g2_decap_8 FILLER_9_1280 ();
 sg13g2_decap_8 FILLER_9_1287 ();
 sg13g2_decap_8 FILLER_9_1294 ();
 sg13g2_decap_8 FILLER_9_1301 ();
 sg13g2_decap_8 FILLER_9_1308 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_fill_2 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_160 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_fill_2 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_202 ();
 sg13g2_fill_1 FILLER_10_217 ();
 sg13g2_fill_2 FILLER_10_283 ();
 sg13g2_fill_2 FILLER_10_312 ();
 sg13g2_fill_1 FILLER_10_314 ();
 sg13g2_fill_2 FILLER_10_323 ();
 sg13g2_fill_2 FILLER_10_334 ();
 sg13g2_fill_1 FILLER_10_336 ();
 sg13g2_fill_2 FILLER_10_401 ();
 sg13g2_fill_2 FILLER_10_419 ();
 sg13g2_fill_1 FILLER_10_421 ();
 sg13g2_fill_1 FILLER_10_449 ();
 sg13g2_fill_1 FILLER_10_476 ();
 sg13g2_fill_1 FILLER_10_549 ();
 sg13g2_fill_2 FILLER_10_563 ();
 sg13g2_fill_1 FILLER_10_565 ();
 sg13g2_fill_2 FILLER_10_584 ();
 sg13g2_fill_2 FILLER_10_596 ();
 sg13g2_fill_1 FILLER_10_598 ();
 sg13g2_fill_2 FILLER_10_616 ();
 sg13g2_fill_1 FILLER_10_618 ();
 sg13g2_fill_2 FILLER_10_627 ();
 sg13g2_fill_1 FILLER_10_629 ();
 sg13g2_fill_2 FILLER_10_639 ();
 sg13g2_fill_2 FILLER_10_659 ();
 sg13g2_fill_2 FILLER_10_687 ();
 sg13g2_fill_1 FILLER_10_693 ();
 sg13g2_fill_1 FILLER_10_720 ();
 sg13g2_decap_4 FILLER_10_759 ();
 sg13g2_fill_1 FILLER_10_763 ();
 sg13g2_fill_1 FILLER_10_845 ();
 sg13g2_fill_1 FILLER_10_942 ();
 sg13g2_fill_2 FILLER_10_1056 ();
 sg13g2_fill_1 FILLER_10_1058 ();
 sg13g2_decap_8 FILLER_10_1068 ();
 sg13g2_decap_8 FILLER_10_1075 ();
 sg13g2_decap_8 FILLER_10_1082 ();
 sg13g2_decap_8 FILLER_10_1089 ();
 sg13g2_decap_8 FILLER_10_1096 ();
 sg13g2_decap_8 FILLER_10_1103 ();
 sg13g2_decap_8 FILLER_10_1110 ();
 sg13g2_decap_8 FILLER_10_1117 ();
 sg13g2_decap_8 FILLER_10_1124 ();
 sg13g2_decap_8 FILLER_10_1131 ();
 sg13g2_decap_8 FILLER_10_1138 ();
 sg13g2_decap_8 FILLER_10_1145 ();
 sg13g2_decap_8 FILLER_10_1152 ();
 sg13g2_decap_8 FILLER_10_1159 ();
 sg13g2_decap_8 FILLER_10_1166 ();
 sg13g2_decap_8 FILLER_10_1173 ();
 sg13g2_decap_8 FILLER_10_1180 ();
 sg13g2_decap_8 FILLER_10_1187 ();
 sg13g2_decap_8 FILLER_10_1194 ();
 sg13g2_decap_8 FILLER_10_1201 ();
 sg13g2_decap_8 FILLER_10_1208 ();
 sg13g2_decap_8 FILLER_10_1215 ();
 sg13g2_decap_8 FILLER_10_1222 ();
 sg13g2_decap_8 FILLER_10_1229 ();
 sg13g2_decap_8 FILLER_10_1236 ();
 sg13g2_decap_8 FILLER_10_1243 ();
 sg13g2_decap_8 FILLER_10_1250 ();
 sg13g2_decap_8 FILLER_10_1257 ();
 sg13g2_decap_8 FILLER_10_1264 ();
 sg13g2_decap_8 FILLER_10_1271 ();
 sg13g2_decap_8 FILLER_10_1278 ();
 sg13g2_decap_8 FILLER_10_1285 ();
 sg13g2_decap_8 FILLER_10_1292 ();
 sg13g2_decap_8 FILLER_10_1299 ();
 sg13g2_decap_8 FILLER_10_1306 ();
 sg13g2_fill_2 FILLER_10_1313 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_fill_2 FILLER_11_187 ();
 sg13g2_fill_1 FILLER_11_205 ();
 sg13g2_fill_1 FILLER_11_241 ();
 sg13g2_fill_2 FILLER_11_268 ();
 sg13g2_fill_2 FILLER_11_336 ();
 sg13g2_fill_1 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_4 FILLER_11_368 ();
 sg13g2_fill_1 FILLER_11_372 ();
 sg13g2_fill_2 FILLER_11_379 ();
 sg13g2_fill_1 FILLER_11_381 ();
 sg13g2_fill_2 FILLER_11_387 ();
 sg13g2_fill_1 FILLER_11_389 ();
 sg13g2_fill_2 FILLER_11_399 ();
 sg13g2_fill_1 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_427 ();
 sg13g2_decap_4 FILLER_11_434 ();
 sg13g2_fill_2 FILLER_11_461 ();
 sg13g2_fill_1 FILLER_11_463 ();
 sg13g2_fill_1 FILLER_11_475 ();
 sg13g2_fill_2 FILLER_11_498 ();
 sg13g2_fill_1 FILLER_11_500 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_fill_1 FILLER_11_518 ();
 sg13g2_fill_1 FILLER_11_571 ();
 sg13g2_fill_1 FILLER_11_592 ();
 sg13g2_fill_2 FILLER_11_654 ();
 sg13g2_fill_1 FILLER_11_704 ();
 sg13g2_fill_1 FILLER_11_709 ();
 sg13g2_fill_2 FILLER_11_802 ();
 sg13g2_fill_1 FILLER_11_804 ();
 sg13g2_fill_1 FILLER_11_815 ();
 sg13g2_fill_2 FILLER_11_846 ();
 sg13g2_fill_1 FILLER_11_865 ();
 sg13g2_fill_1 FILLER_11_884 ();
 sg13g2_fill_2 FILLER_11_911 ();
 sg13g2_fill_1 FILLER_11_913 ();
 sg13g2_fill_1 FILLER_11_940 ();
 sg13g2_fill_1 FILLER_11_1002 ();
 sg13g2_fill_1 FILLER_11_1016 ();
 sg13g2_decap_8 FILLER_11_1069 ();
 sg13g2_decap_8 FILLER_11_1076 ();
 sg13g2_decap_8 FILLER_11_1083 ();
 sg13g2_decap_8 FILLER_11_1090 ();
 sg13g2_decap_8 FILLER_11_1097 ();
 sg13g2_decap_8 FILLER_11_1104 ();
 sg13g2_decap_8 FILLER_11_1111 ();
 sg13g2_decap_8 FILLER_11_1118 ();
 sg13g2_decap_8 FILLER_11_1125 ();
 sg13g2_decap_8 FILLER_11_1132 ();
 sg13g2_decap_8 FILLER_11_1139 ();
 sg13g2_decap_8 FILLER_11_1146 ();
 sg13g2_decap_8 FILLER_11_1153 ();
 sg13g2_decap_8 FILLER_11_1160 ();
 sg13g2_decap_8 FILLER_11_1167 ();
 sg13g2_decap_8 FILLER_11_1174 ();
 sg13g2_decap_8 FILLER_11_1181 ();
 sg13g2_decap_8 FILLER_11_1188 ();
 sg13g2_decap_8 FILLER_11_1195 ();
 sg13g2_decap_8 FILLER_11_1202 ();
 sg13g2_decap_8 FILLER_11_1209 ();
 sg13g2_decap_8 FILLER_11_1216 ();
 sg13g2_decap_8 FILLER_11_1223 ();
 sg13g2_decap_8 FILLER_11_1230 ();
 sg13g2_decap_8 FILLER_11_1237 ();
 sg13g2_decap_8 FILLER_11_1244 ();
 sg13g2_decap_8 FILLER_11_1251 ();
 sg13g2_decap_8 FILLER_11_1258 ();
 sg13g2_decap_8 FILLER_11_1265 ();
 sg13g2_decap_8 FILLER_11_1272 ();
 sg13g2_decap_8 FILLER_11_1279 ();
 sg13g2_decap_8 FILLER_11_1286 ();
 sg13g2_decap_8 FILLER_11_1293 ();
 sg13g2_decap_8 FILLER_11_1300 ();
 sg13g2_decap_8 FILLER_11_1307 ();
 sg13g2_fill_1 FILLER_11_1314 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_4 FILLER_12_105 ();
 sg13g2_fill_2 FILLER_12_109 ();
 sg13g2_fill_2 FILLER_12_150 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_fill_2 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_169 ();
 sg13g2_fill_1 FILLER_12_197 ();
 sg13g2_fill_2 FILLER_12_224 ();
 sg13g2_fill_2 FILLER_12_240 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_fill_1 FILLER_12_291 ();
 sg13g2_fill_2 FILLER_12_301 ();
 sg13g2_fill_1 FILLER_12_338 ();
 sg13g2_fill_2 FILLER_12_374 ();
 sg13g2_fill_2 FILLER_12_382 ();
 sg13g2_fill_1 FILLER_12_384 ();
 sg13g2_fill_2 FILLER_12_398 ();
 sg13g2_fill_1 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_416 ();
 sg13g2_fill_2 FILLER_12_422 ();
 sg13g2_fill_1 FILLER_12_424 ();
 sg13g2_fill_2 FILLER_12_458 ();
 sg13g2_fill_1 FILLER_12_473 ();
 sg13g2_fill_2 FILLER_12_483 ();
 sg13g2_decap_4 FILLER_12_505 ();
 sg13g2_fill_2 FILLER_12_517 ();
 sg13g2_fill_1 FILLER_12_519 ();
 sg13g2_decap_4 FILLER_12_525 ();
 sg13g2_fill_2 FILLER_12_529 ();
 sg13g2_fill_2 FILLER_12_544 ();
 sg13g2_fill_1 FILLER_12_555 ();
 sg13g2_fill_1 FILLER_12_586 ();
 sg13g2_fill_1 FILLER_12_631 ();
 sg13g2_decap_4 FILLER_12_684 ();
 sg13g2_fill_2 FILLER_12_688 ();
 sg13g2_fill_1 FILLER_12_725 ();
 sg13g2_fill_2 FILLER_12_743 ();
 sg13g2_fill_1 FILLER_12_745 ();
 sg13g2_fill_1 FILLER_12_785 ();
 sg13g2_fill_1 FILLER_12_812 ();
 sg13g2_fill_1 FILLER_12_823 ();
 sg13g2_fill_1 FILLER_12_904 ();
 sg13g2_fill_2 FILLER_12_910 ();
 sg13g2_fill_1 FILLER_12_912 ();
 sg13g2_fill_1 FILLER_12_922 ();
 sg13g2_fill_2 FILLER_12_949 ();
 sg13g2_fill_2 FILLER_12_1050 ();
 sg13g2_decap_8 FILLER_12_1069 ();
 sg13g2_decap_8 FILLER_12_1076 ();
 sg13g2_decap_8 FILLER_12_1083 ();
 sg13g2_decap_8 FILLER_12_1090 ();
 sg13g2_decap_8 FILLER_12_1097 ();
 sg13g2_decap_8 FILLER_12_1104 ();
 sg13g2_decap_8 FILLER_12_1111 ();
 sg13g2_decap_8 FILLER_12_1118 ();
 sg13g2_decap_8 FILLER_12_1125 ();
 sg13g2_decap_8 FILLER_12_1132 ();
 sg13g2_decap_8 FILLER_12_1139 ();
 sg13g2_decap_8 FILLER_12_1146 ();
 sg13g2_decap_8 FILLER_12_1153 ();
 sg13g2_decap_8 FILLER_12_1160 ();
 sg13g2_decap_8 FILLER_12_1167 ();
 sg13g2_decap_8 FILLER_12_1174 ();
 sg13g2_decap_8 FILLER_12_1181 ();
 sg13g2_decap_8 FILLER_12_1188 ();
 sg13g2_decap_8 FILLER_12_1195 ();
 sg13g2_decap_8 FILLER_12_1202 ();
 sg13g2_decap_8 FILLER_12_1209 ();
 sg13g2_decap_8 FILLER_12_1216 ();
 sg13g2_decap_8 FILLER_12_1223 ();
 sg13g2_decap_8 FILLER_12_1230 ();
 sg13g2_decap_8 FILLER_12_1237 ();
 sg13g2_decap_8 FILLER_12_1244 ();
 sg13g2_decap_8 FILLER_12_1251 ();
 sg13g2_decap_8 FILLER_12_1258 ();
 sg13g2_decap_8 FILLER_12_1265 ();
 sg13g2_decap_8 FILLER_12_1272 ();
 sg13g2_decap_8 FILLER_12_1279 ();
 sg13g2_decap_8 FILLER_12_1286 ();
 sg13g2_decap_8 FILLER_12_1293 ();
 sg13g2_decap_8 FILLER_12_1300 ();
 sg13g2_decap_8 FILLER_12_1307 ();
 sg13g2_fill_1 FILLER_12_1314 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_218 ();
 sg13g2_fill_2 FILLER_13_267 ();
 sg13g2_fill_1 FILLER_13_269 ();
 sg13g2_fill_1 FILLER_13_331 ();
 sg13g2_fill_2 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_342 ();
 sg13g2_decap_4 FILLER_13_355 ();
 sg13g2_decap_4 FILLER_13_391 ();
 sg13g2_fill_1 FILLER_13_395 ();
 sg13g2_fill_2 FILLER_13_418 ();
 sg13g2_fill_1 FILLER_13_430 ();
 sg13g2_fill_2 FILLER_13_447 ();
 sg13g2_fill_2 FILLER_13_459 ();
 sg13g2_fill_1 FILLER_13_461 ();
 sg13g2_fill_2 FILLER_13_468 ();
 sg13g2_fill_1 FILLER_13_470 ();
 sg13g2_decap_4 FILLER_13_493 ();
 sg13g2_fill_2 FILLER_13_497 ();
 sg13g2_fill_2 FILLER_13_564 ();
 sg13g2_fill_2 FILLER_13_579 ();
 sg13g2_fill_1 FILLER_13_614 ();
 sg13g2_fill_2 FILLER_13_641 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_fill_1 FILLER_13_707 ();
 sg13g2_fill_2 FILLER_13_800 ();
 sg13g2_fill_1 FILLER_13_802 ();
 sg13g2_decap_8 FILLER_13_850 ();
 sg13g2_fill_2 FILLER_13_857 ();
 sg13g2_fill_2 FILLER_13_983 ();
 sg13g2_fill_1 FILLER_13_985 ();
 sg13g2_fill_1 FILLER_13_1015 ();
 sg13g2_fill_1 FILLER_13_1020 ();
 sg13g2_decap_8 FILLER_13_1063 ();
 sg13g2_decap_8 FILLER_13_1070 ();
 sg13g2_decap_8 FILLER_13_1077 ();
 sg13g2_decap_8 FILLER_13_1084 ();
 sg13g2_decap_8 FILLER_13_1091 ();
 sg13g2_decap_8 FILLER_13_1098 ();
 sg13g2_decap_8 FILLER_13_1105 ();
 sg13g2_decap_8 FILLER_13_1112 ();
 sg13g2_decap_8 FILLER_13_1119 ();
 sg13g2_decap_8 FILLER_13_1126 ();
 sg13g2_decap_8 FILLER_13_1133 ();
 sg13g2_decap_8 FILLER_13_1140 ();
 sg13g2_decap_8 FILLER_13_1147 ();
 sg13g2_decap_8 FILLER_13_1154 ();
 sg13g2_decap_8 FILLER_13_1161 ();
 sg13g2_decap_8 FILLER_13_1168 ();
 sg13g2_decap_8 FILLER_13_1175 ();
 sg13g2_decap_8 FILLER_13_1182 ();
 sg13g2_decap_8 FILLER_13_1189 ();
 sg13g2_decap_8 FILLER_13_1196 ();
 sg13g2_decap_8 FILLER_13_1203 ();
 sg13g2_decap_8 FILLER_13_1210 ();
 sg13g2_decap_8 FILLER_13_1217 ();
 sg13g2_decap_8 FILLER_13_1224 ();
 sg13g2_decap_8 FILLER_13_1231 ();
 sg13g2_decap_8 FILLER_13_1238 ();
 sg13g2_decap_8 FILLER_13_1245 ();
 sg13g2_decap_8 FILLER_13_1252 ();
 sg13g2_decap_8 FILLER_13_1259 ();
 sg13g2_decap_8 FILLER_13_1266 ();
 sg13g2_decap_8 FILLER_13_1273 ();
 sg13g2_decap_8 FILLER_13_1280 ();
 sg13g2_decap_8 FILLER_13_1287 ();
 sg13g2_decap_8 FILLER_13_1294 ();
 sg13g2_decap_8 FILLER_13_1301 ();
 sg13g2_decap_8 FILLER_13_1308 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_170 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_fill_2 FILLER_14_211 ();
 sg13g2_fill_1 FILLER_14_213 ();
 sg13g2_fill_1 FILLER_14_227 ();
 sg13g2_fill_2 FILLER_14_250 ();
 sg13g2_fill_1 FILLER_14_252 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_322 ();
 sg13g2_fill_2 FILLER_14_328 ();
 sg13g2_fill_1 FILLER_14_330 ();
 sg13g2_decap_4 FILLER_14_336 ();
 sg13g2_fill_1 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_351 ();
 sg13g2_fill_1 FILLER_14_358 ();
 sg13g2_fill_2 FILLER_14_364 ();
 sg13g2_fill_2 FILLER_14_436 ();
 sg13g2_fill_2 FILLER_14_448 ();
 sg13g2_fill_1 FILLER_14_450 ();
 sg13g2_fill_2 FILLER_14_455 ();
 sg13g2_fill_1 FILLER_14_457 ();
 sg13g2_decap_4 FILLER_14_470 ();
 sg13g2_fill_2 FILLER_14_474 ();
 sg13g2_decap_4 FILLER_14_481 ();
 sg13g2_fill_1 FILLER_14_485 ();
 sg13g2_decap_4 FILLER_14_494 ();
 sg13g2_decap_8 FILLER_14_505 ();
 sg13g2_decap_4 FILLER_14_512 ();
 sg13g2_fill_1 FILLER_14_578 ();
 sg13g2_fill_1 FILLER_14_592 ();
 sg13g2_fill_2 FILLER_14_607 ();
 sg13g2_decap_4 FILLER_14_696 ();
 sg13g2_fill_1 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_705 ();
 sg13g2_fill_1 FILLER_14_726 ();
 sg13g2_fill_2 FILLER_14_811 ();
 sg13g2_fill_1 FILLER_14_813 ();
 sg13g2_fill_2 FILLER_14_828 ();
 sg13g2_decap_4 FILLER_14_1068 ();
 sg13g2_fill_2 FILLER_14_1077 ();
 sg13g2_fill_1 FILLER_14_1079 ();
 sg13g2_decap_8 FILLER_14_1084 ();
 sg13g2_decap_8 FILLER_14_1091 ();
 sg13g2_decap_8 FILLER_14_1098 ();
 sg13g2_decap_8 FILLER_14_1105 ();
 sg13g2_decap_8 FILLER_14_1112 ();
 sg13g2_decap_8 FILLER_14_1119 ();
 sg13g2_decap_8 FILLER_14_1126 ();
 sg13g2_decap_8 FILLER_14_1133 ();
 sg13g2_decap_8 FILLER_14_1140 ();
 sg13g2_decap_8 FILLER_14_1147 ();
 sg13g2_decap_8 FILLER_14_1154 ();
 sg13g2_decap_8 FILLER_14_1161 ();
 sg13g2_decap_8 FILLER_14_1168 ();
 sg13g2_decap_8 FILLER_14_1175 ();
 sg13g2_decap_8 FILLER_14_1182 ();
 sg13g2_decap_8 FILLER_14_1189 ();
 sg13g2_decap_8 FILLER_14_1196 ();
 sg13g2_decap_8 FILLER_14_1203 ();
 sg13g2_decap_8 FILLER_14_1210 ();
 sg13g2_decap_8 FILLER_14_1217 ();
 sg13g2_decap_8 FILLER_14_1224 ();
 sg13g2_decap_8 FILLER_14_1231 ();
 sg13g2_decap_8 FILLER_14_1238 ();
 sg13g2_decap_8 FILLER_14_1245 ();
 sg13g2_decap_8 FILLER_14_1252 ();
 sg13g2_decap_8 FILLER_14_1259 ();
 sg13g2_decap_8 FILLER_14_1266 ();
 sg13g2_decap_8 FILLER_14_1273 ();
 sg13g2_decap_8 FILLER_14_1280 ();
 sg13g2_decap_8 FILLER_14_1287 ();
 sg13g2_decap_8 FILLER_14_1294 ();
 sg13g2_decap_8 FILLER_14_1301 ();
 sg13g2_decap_8 FILLER_14_1308 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_4 FILLER_15_98 ();
 sg13g2_fill_2 FILLER_15_102 ();
 sg13g2_fill_2 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_2 FILLER_15_182 ();
 sg13g2_fill_1 FILLER_15_184 ();
 sg13g2_fill_2 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_fill_2 FILLER_15_328 ();
 sg13g2_decap_4 FILLER_15_357 ();
 sg13g2_fill_2 FILLER_15_361 ();
 sg13g2_fill_1 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_4 FILLER_15_410 ();
 sg13g2_fill_1 FILLER_15_414 ();
 sg13g2_fill_2 FILLER_15_431 ();
 sg13g2_fill_2 FILLER_15_442 ();
 sg13g2_fill_2 FILLER_15_450 ();
 sg13g2_fill_1 FILLER_15_452 ();
 sg13g2_fill_2 FILLER_15_475 ();
 sg13g2_fill_1 FILLER_15_477 ();
 sg13g2_decap_4 FILLER_15_503 ();
 sg13g2_fill_1 FILLER_15_507 ();
 sg13g2_fill_1 FILLER_15_631 ();
 sg13g2_decap_4 FILLER_15_658 ();
 sg13g2_fill_1 FILLER_15_662 ();
 sg13g2_fill_2 FILLER_15_671 ();
 sg13g2_fill_2 FILLER_15_682 ();
 sg13g2_decap_4 FILLER_15_688 ();
 sg13g2_fill_2 FILLER_15_692 ();
 sg13g2_fill_2 FILLER_15_803 ();
 sg13g2_decap_8 FILLER_15_845 ();
 sg13g2_decap_4 FILLER_15_852 ();
 sg13g2_decap_8 FILLER_15_869 ();
 sg13g2_fill_2 FILLER_15_923 ();
 sg13g2_fill_1 FILLER_15_925 ();
 sg13g2_fill_1 FILLER_15_987 ();
 sg13g2_decap_8 FILLER_15_1101 ();
 sg13g2_decap_8 FILLER_15_1108 ();
 sg13g2_decap_8 FILLER_15_1115 ();
 sg13g2_decap_8 FILLER_15_1122 ();
 sg13g2_decap_8 FILLER_15_1129 ();
 sg13g2_decap_8 FILLER_15_1136 ();
 sg13g2_decap_8 FILLER_15_1143 ();
 sg13g2_decap_8 FILLER_15_1150 ();
 sg13g2_decap_8 FILLER_15_1157 ();
 sg13g2_decap_8 FILLER_15_1164 ();
 sg13g2_decap_8 FILLER_15_1171 ();
 sg13g2_decap_8 FILLER_15_1178 ();
 sg13g2_decap_8 FILLER_15_1185 ();
 sg13g2_decap_8 FILLER_15_1192 ();
 sg13g2_decap_8 FILLER_15_1199 ();
 sg13g2_decap_8 FILLER_15_1206 ();
 sg13g2_decap_8 FILLER_15_1213 ();
 sg13g2_decap_8 FILLER_15_1220 ();
 sg13g2_decap_8 FILLER_15_1227 ();
 sg13g2_decap_8 FILLER_15_1234 ();
 sg13g2_decap_8 FILLER_15_1241 ();
 sg13g2_decap_8 FILLER_15_1248 ();
 sg13g2_decap_8 FILLER_15_1255 ();
 sg13g2_decap_8 FILLER_15_1262 ();
 sg13g2_decap_8 FILLER_15_1269 ();
 sg13g2_decap_8 FILLER_15_1276 ();
 sg13g2_decap_8 FILLER_15_1283 ();
 sg13g2_decap_8 FILLER_15_1290 ();
 sg13g2_decap_8 FILLER_15_1297 ();
 sg13g2_decap_8 FILLER_15_1304 ();
 sg13g2_decap_4 FILLER_15_1311 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_147 ();
 sg13g2_fill_1 FILLER_16_196 ();
 sg13g2_fill_2 FILLER_16_215 ();
 sg13g2_fill_1 FILLER_16_243 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_decap_4 FILLER_16_328 ();
 sg13g2_fill_2 FILLER_16_344 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_16_415 ();
 sg13g2_fill_1 FILLER_16_419 ();
 sg13g2_fill_2 FILLER_16_434 ();
 sg13g2_fill_2 FILLER_16_453 ();
 sg13g2_decap_4 FILLER_16_476 ();
 sg13g2_fill_2 FILLER_16_480 ();
 sg13g2_fill_2 FILLER_16_487 ();
 sg13g2_fill_2 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_513 ();
 sg13g2_fill_2 FILLER_16_520 ();
 sg13g2_fill_2 FILLER_16_527 ();
 sg13g2_fill_1 FILLER_16_533 ();
 sg13g2_fill_1 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_712 ();
 sg13g2_fill_1 FILLER_16_719 ();
 sg13g2_decap_4 FILLER_16_737 ();
 sg13g2_fill_2 FILLER_16_741 ();
 sg13g2_fill_2 FILLER_16_779 ();
 sg13g2_fill_1 FILLER_16_781 ();
 sg13g2_fill_1 FILLER_16_820 ();
 sg13g2_decap_8 FILLER_16_834 ();
 sg13g2_decap_4 FILLER_16_841 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_fill_2 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_936 ();
 sg13g2_fill_1 FILLER_16_938 ();
 sg13g2_fill_2 FILLER_16_970 ();
 sg13g2_fill_2 FILLER_16_1033 ();
 sg13g2_fill_1 FILLER_16_1061 ();
 sg13g2_fill_1 FILLER_16_1074 ();
 sg13g2_decap_8 FILLER_16_1123 ();
 sg13g2_decap_8 FILLER_16_1130 ();
 sg13g2_decap_8 FILLER_16_1137 ();
 sg13g2_decap_8 FILLER_16_1144 ();
 sg13g2_decap_8 FILLER_16_1151 ();
 sg13g2_decap_8 FILLER_16_1158 ();
 sg13g2_decap_8 FILLER_16_1165 ();
 sg13g2_decap_8 FILLER_16_1172 ();
 sg13g2_decap_8 FILLER_16_1179 ();
 sg13g2_decap_8 FILLER_16_1186 ();
 sg13g2_decap_8 FILLER_16_1193 ();
 sg13g2_decap_8 FILLER_16_1200 ();
 sg13g2_decap_8 FILLER_16_1207 ();
 sg13g2_decap_8 FILLER_16_1214 ();
 sg13g2_decap_8 FILLER_16_1221 ();
 sg13g2_decap_8 FILLER_16_1228 ();
 sg13g2_decap_8 FILLER_16_1235 ();
 sg13g2_decap_8 FILLER_16_1242 ();
 sg13g2_decap_8 FILLER_16_1249 ();
 sg13g2_decap_8 FILLER_16_1256 ();
 sg13g2_decap_8 FILLER_16_1263 ();
 sg13g2_decap_8 FILLER_16_1270 ();
 sg13g2_decap_8 FILLER_16_1277 ();
 sg13g2_decap_8 FILLER_16_1284 ();
 sg13g2_decap_8 FILLER_16_1291 ();
 sg13g2_decap_8 FILLER_16_1298 ();
 sg13g2_decap_8 FILLER_16_1305 ();
 sg13g2_fill_2 FILLER_16_1312 ();
 sg13g2_fill_1 FILLER_16_1314 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_179 ();
 sg13g2_fill_1 FILLER_17_186 ();
 sg13g2_fill_2 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_258 ();
 sg13g2_fill_1 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_275 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_fill_2 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_4 FILLER_17_355 ();
 sg13g2_fill_1 FILLER_17_365 ();
 sg13g2_fill_2 FILLER_17_388 ();
 sg13g2_fill_2 FILLER_17_405 ();
 sg13g2_fill_1 FILLER_17_417 ();
 sg13g2_fill_1 FILLER_17_422 ();
 sg13g2_decap_4 FILLER_17_433 ();
 sg13g2_decap_4 FILLER_17_453 ();
 sg13g2_fill_2 FILLER_17_457 ();
 sg13g2_fill_2 FILLER_17_468 ();
 sg13g2_fill_1 FILLER_17_470 ();
 sg13g2_decap_8 FILLER_17_475 ();
 sg13g2_fill_1 FILLER_17_612 ();
 sg13g2_fill_2 FILLER_17_622 ();
 sg13g2_fill_1 FILLER_17_624 ();
 sg13g2_decap_8 FILLER_17_657 ();
 sg13g2_decap_4 FILLER_17_664 ();
 sg13g2_fill_1 FILLER_17_677 ();
 sg13g2_fill_2 FILLER_17_765 ();
 sg13g2_fill_1 FILLER_17_767 ();
 sg13g2_fill_2 FILLER_17_787 ();
 sg13g2_fill_1 FILLER_17_789 ();
 sg13g2_fill_2 FILLER_17_904 ();
 sg13g2_fill_1 FILLER_17_906 ();
 sg13g2_fill_2 FILLER_17_916 ();
 sg13g2_fill_1 FILLER_17_918 ();
 sg13g2_fill_2 FILLER_17_959 ();
 sg13g2_fill_2 FILLER_17_995 ();
 sg13g2_fill_1 FILLER_17_997 ();
 sg13g2_fill_1 FILLER_17_1011 ();
 sg13g2_fill_1 FILLER_17_1015 ();
 sg13g2_fill_1 FILLER_17_1086 ();
 sg13g2_decap_8 FILLER_17_1104 ();
 sg13g2_decap_8 FILLER_17_1111 ();
 sg13g2_decap_8 FILLER_17_1118 ();
 sg13g2_decap_8 FILLER_17_1125 ();
 sg13g2_decap_8 FILLER_17_1132 ();
 sg13g2_decap_8 FILLER_17_1139 ();
 sg13g2_decap_8 FILLER_17_1146 ();
 sg13g2_decap_8 FILLER_17_1153 ();
 sg13g2_decap_8 FILLER_17_1160 ();
 sg13g2_decap_8 FILLER_17_1167 ();
 sg13g2_decap_8 FILLER_17_1174 ();
 sg13g2_decap_8 FILLER_17_1181 ();
 sg13g2_decap_8 FILLER_17_1188 ();
 sg13g2_decap_8 FILLER_17_1195 ();
 sg13g2_decap_8 FILLER_17_1202 ();
 sg13g2_decap_8 FILLER_17_1209 ();
 sg13g2_decap_8 FILLER_17_1216 ();
 sg13g2_decap_8 FILLER_17_1223 ();
 sg13g2_decap_8 FILLER_17_1230 ();
 sg13g2_decap_8 FILLER_17_1237 ();
 sg13g2_decap_8 FILLER_17_1244 ();
 sg13g2_decap_8 FILLER_17_1251 ();
 sg13g2_decap_8 FILLER_17_1258 ();
 sg13g2_decap_8 FILLER_17_1265 ();
 sg13g2_decap_8 FILLER_17_1272 ();
 sg13g2_decap_8 FILLER_17_1279 ();
 sg13g2_decap_8 FILLER_17_1286 ();
 sg13g2_decap_8 FILLER_17_1293 ();
 sg13g2_decap_8 FILLER_17_1300 ();
 sg13g2_decap_8 FILLER_17_1307 ();
 sg13g2_fill_1 FILLER_17_1314 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_fill_2 FILLER_18_98 ();
 sg13g2_decap_4 FILLER_18_113 ();
 sg13g2_fill_2 FILLER_18_117 ();
 sg13g2_fill_1 FILLER_18_122 ();
 sg13g2_fill_2 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_135 ();
 sg13g2_fill_2 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_190 ();
 sg13g2_fill_2 FILLER_18_205 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_fill_2 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_337 ();
 sg13g2_fill_2 FILLER_18_355 ();
 sg13g2_fill_1 FILLER_18_357 ();
 sg13g2_fill_2 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_fill_2 FILLER_18_389 ();
 sg13g2_fill_1 FILLER_18_391 ();
 sg13g2_fill_1 FILLER_18_402 ();
 sg13g2_fill_2 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_431 ();
 sg13g2_decap_4 FILLER_18_445 ();
 sg13g2_fill_2 FILLER_18_449 ();
 sg13g2_fill_2 FILLER_18_466 ();
 sg13g2_fill_2 FILLER_18_487 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_fill_2 FILLER_18_525 ();
 sg13g2_fill_1 FILLER_18_527 ();
 sg13g2_decap_4 FILLER_18_556 ();
 sg13g2_fill_2 FILLER_18_560 ();
 sg13g2_fill_1 FILLER_18_590 ();
 sg13g2_fill_2 FILLER_18_601 ();
 sg13g2_fill_1 FILLER_18_603 ();
 sg13g2_decap_8 FILLER_18_695 ();
 sg13g2_fill_2 FILLER_18_702 ();
 sg13g2_decap_8 FILLER_18_717 ();
 sg13g2_fill_2 FILLER_18_724 ();
 sg13g2_fill_2 FILLER_18_739 ();
 sg13g2_fill_2 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_fill_2 FILLER_18_850 ();
 sg13g2_fill_1 FILLER_18_852 ();
 sg13g2_fill_2 FILLER_18_857 ();
 sg13g2_fill_1 FILLER_18_877 ();
 sg13g2_fill_2 FILLER_18_901 ();
 sg13g2_fill_1 FILLER_18_903 ();
 sg13g2_fill_2 FILLER_18_982 ();
 sg13g2_fill_2 FILLER_18_1006 ();
 sg13g2_fill_1 FILLER_18_1008 ();
 sg13g2_fill_2 FILLER_18_1057 ();
 sg13g2_decap_8 FILLER_18_1102 ();
 sg13g2_decap_8 FILLER_18_1109 ();
 sg13g2_decap_8 FILLER_18_1116 ();
 sg13g2_decap_8 FILLER_18_1123 ();
 sg13g2_decap_8 FILLER_18_1130 ();
 sg13g2_decap_8 FILLER_18_1137 ();
 sg13g2_decap_8 FILLER_18_1144 ();
 sg13g2_decap_8 FILLER_18_1151 ();
 sg13g2_decap_8 FILLER_18_1158 ();
 sg13g2_decap_8 FILLER_18_1165 ();
 sg13g2_decap_8 FILLER_18_1172 ();
 sg13g2_decap_8 FILLER_18_1179 ();
 sg13g2_decap_8 FILLER_18_1186 ();
 sg13g2_decap_8 FILLER_18_1193 ();
 sg13g2_decap_8 FILLER_18_1200 ();
 sg13g2_decap_8 FILLER_18_1207 ();
 sg13g2_decap_8 FILLER_18_1214 ();
 sg13g2_decap_8 FILLER_18_1221 ();
 sg13g2_decap_8 FILLER_18_1228 ();
 sg13g2_decap_8 FILLER_18_1235 ();
 sg13g2_decap_8 FILLER_18_1242 ();
 sg13g2_decap_8 FILLER_18_1249 ();
 sg13g2_decap_8 FILLER_18_1256 ();
 sg13g2_decap_8 FILLER_18_1263 ();
 sg13g2_decap_8 FILLER_18_1270 ();
 sg13g2_decap_8 FILLER_18_1277 ();
 sg13g2_decap_8 FILLER_18_1284 ();
 sg13g2_decap_8 FILLER_18_1291 ();
 sg13g2_decap_8 FILLER_18_1298 ();
 sg13g2_decap_8 FILLER_18_1305 ();
 sg13g2_fill_2 FILLER_18_1312 ();
 sg13g2_fill_1 FILLER_18_1314 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_4 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_88 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_decap_4 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_4 FILLER_19_363 ();
 sg13g2_fill_1 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_4 FILLER_19_409 ();
 sg13g2_fill_1 FILLER_19_413 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_1 FILLER_19_428 ();
 sg13g2_fill_1 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_443 ();
 sg13g2_fill_1 FILLER_19_467 ();
 sg13g2_fill_2 FILLER_19_485 ();
 sg13g2_decap_4 FILLER_19_499 ();
 sg13g2_fill_2 FILLER_19_503 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_fill_1 FILLER_19_525 ();
 sg13g2_decap_4 FILLER_19_552 ();
 sg13g2_fill_2 FILLER_19_575 ();
 sg13g2_fill_1 FILLER_19_595 ();
 sg13g2_fill_1 FILLER_19_626 ();
 sg13g2_fill_1 FILLER_19_644 ();
 sg13g2_decap_4 FILLER_19_664 ();
 sg13g2_fill_1 FILLER_19_668 ();
 sg13g2_fill_1 FILLER_19_687 ();
 sg13g2_decap_8 FILLER_19_741 ();
 sg13g2_fill_1 FILLER_19_748 ();
 sg13g2_fill_2 FILLER_19_760 ();
 sg13g2_fill_1 FILLER_19_762 ();
 sg13g2_fill_1 FILLER_19_768 ();
 sg13g2_fill_2 FILLER_19_783 ();
 sg13g2_fill_1 FILLER_19_959 ();
 sg13g2_decap_8 FILLER_19_1107 ();
 sg13g2_decap_8 FILLER_19_1114 ();
 sg13g2_decap_8 FILLER_19_1121 ();
 sg13g2_decap_8 FILLER_19_1128 ();
 sg13g2_decap_8 FILLER_19_1135 ();
 sg13g2_decap_8 FILLER_19_1142 ();
 sg13g2_decap_8 FILLER_19_1149 ();
 sg13g2_decap_8 FILLER_19_1156 ();
 sg13g2_decap_8 FILLER_19_1163 ();
 sg13g2_decap_8 FILLER_19_1170 ();
 sg13g2_decap_8 FILLER_19_1177 ();
 sg13g2_decap_8 FILLER_19_1184 ();
 sg13g2_decap_8 FILLER_19_1191 ();
 sg13g2_decap_8 FILLER_19_1198 ();
 sg13g2_decap_8 FILLER_19_1205 ();
 sg13g2_decap_8 FILLER_19_1212 ();
 sg13g2_decap_8 FILLER_19_1219 ();
 sg13g2_decap_8 FILLER_19_1226 ();
 sg13g2_decap_8 FILLER_19_1233 ();
 sg13g2_decap_8 FILLER_19_1240 ();
 sg13g2_decap_8 FILLER_19_1247 ();
 sg13g2_decap_8 FILLER_19_1254 ();
 sg13g2_decap_8 FILLER_19_1261 ();
 sg13g2_decap_8 FILLER_19_1268 ();
 sg13g2_decap_8 FILLER_19_1275 ();
 sg13g2_decap_8 FILLER_19_1282 ();
 sg13g2_decap_8 FILLER_19_1289 ();
 sg13g2_decap_8 FILLER_19_1296 ();
 sg13g2_decap_8 FILLER_19_1303 ();
 sg13g2_decap_4 FILLER_19_1310 ();
 sg13g2_fill_1 FILLER_19_1314 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_4 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_127 ();
 sg13g2_fill_2 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_244 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_decap_8 FILLER_20_330 ();
 sg13g2_fill_1 FILLER_20_337 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_20_387 ();
 sg13g2_fill_1 FILLER_20_397 ();
 sg13g2_fill_2 FILLER_20_403 ();
 sg13g2_fill_1 FILLER_20_405 ();
 sg13g2_fill_2 FILLER_20_411 ();
 sg13g2_fill_1 FILLER_20_413 ();
 sg13g2_fill_1 FILLER_20_420 ();
 sg13g2_decap_4 FILLER_20_446 ();
 sg13g2_decap_4 FILLER_20_466 ();
 sg13g2_decap_4 FILLER_20_483 ();
 sg13g2_fill_1 FILLER_20_494 ();
 sg13g2_fill_1 FILLER_20_526 ();
 sg13g2_fill_2 FILLER_20_537 ();
 sg13g2_fill_1 FILLER_20_548 ();
 sg13g2_fill_2 FILLER_20_613 ();
 sg13g2_decap_4 FILLER_20_641 ();
 sg13g2_decap_8 FILLER_20_649 ();
 sg13g2_decap_8 FILLER_20_656 ();
 sg13g2_fill_1 FILLER_20_663 ();
 sg13g2_decap_4 FILLER_20_704 ();
 sg13g2_fill_2 FILLER_20_708 ();
 sg13g2_fill_1 FILLER_20_783 ();
 sg13g2_fill_2 FILLER_20_816 ();
 sg13g2_fill_1 FILLER_20_818 ();
 sg13g2_fill_2 FILLER_20_823 ();
 sg13g2_decap_8 FILLER_20_838 ();
 sg13g2_decap_8 FILLER_20_845 ();
 sg13g2_decap_4 FILLER_20_856 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_fill_2 FILLER_20_888 ();
 sg13g2_fill_2 FILLER_20_951 ();
 sg13g2_fill_1 FILLER_20_953 ();
 sg13g2_fill_1 FILLER_20_972 ();
 sg13g2_fill_2 FILLER_20_1061 ();
 sg13g2_fill_1 FILLER_20_1063 ();
 sg13g2_fill_2 FILLER_20_1082 ();
 sg13g2_fill_1 FILLER_20_1084 ();
 sg13g2_decap_8 FILLER_20_1124 ();
 sg13g2_decap_8 FILLER_20_1131 ();
 sg13g2_decap_8 FILLER_20_1138 ();
 sg13g2_decap_8 FILLER_20_1145 ();
 sg13g2_decap_8 FILLER_20_1152 ();
 sg13g2_decap_8 FILLER_20_1159 ();
 sg13g2_decap_8 FILLER_20_1166 ();
 sg13g2_decap_8 FILLER_20_1173 ();
 sg13g2_decap_8 FILLER_20_1180 ();
 sg13g2_decap_8 FILLER_20_1187 ();
 sg13g2_decap_8 FILLER_20_1194 ();
 sg13g2_decap_8 FILLER_20_1201 ();
 sg13g2_decap_8 FILLER_20_1208 ();
 sg13g2_decap_8 FILLER_20_1215 ();
 sg13g2_decap_8 FILLER_20_1222 ();
 sg13g2_decap_8 FILLER_20_1229 ();
 sg13g2_decap_8 FILLER_20_1236 ();
 sg13g2_decap_8 FILLER_20_1243 ();
 sg13g2_decap_8 FILLER_20_1250 ();
 sg13g2_decap_8 FILLER_20_1257 ();
 sg13g2_decap_8 FILLER_20_1264 ();
 sg13g2_decap_8 FILLER_20_1271 ();
 sg13g2_decap_8 FILLER_20_1278 ();
 sg13g2_decap_8 FILLER_20_1285 ();
 sg13g2_decap_8 FILLER_20_1292 ();
 sg13g2_decap_8 FILLER_20_1299 ();
 sg13g2_decap_8 FILLER_20_1306 ();
 sg13g2_fill_2 FILLER_20_1313 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_4 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_74 ();
 sg13g2_fill_1 FILLER_21_117 ();
 sg13g2_fill_2 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_decap_4 FILLER_21_340 ();
 sg13g2_fill_1 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_fill_2 FILLER_21_389 ();
 sg13g2_fill_1 FILLER_21_401 ();
 sg13g2_fill_2 FILLER_21_411 ();
 sg13g2_fill_1 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_419 ();
 sg13g2_fill_2 FILLER_21_426 ();
 sg13g2_decap_8 FILLER_21_445 ();
 sg13g2_fill_1 FILLER_21_452 ();
 sg13g2_fill_2 FILLER_21_473 ();
 sg13g2_fill_1 FILLER_21_475 ();
 sg13g2_decap_4 FILLER_21_521 ();
 sg13g2_fill_2 FILLER_21_525 ();
 sg13g2_fill_2 FILLER_21_558 ();
 sg13g2_decap_4 FILLER_21_564 ();
 sg13g2_fill_2 FILLER_21_629 ();
 sg13g2_fill_1 FILLER_21_631 ();
 sg13g2_fill_2 FILLER_21_636 ();
 sg13g2_fill_1 FILLER_21_638 ();
 sg13g2_fill_2 FILLER_21_728 ();
 sg13g2_fill_2 FILLER_21_745 ();
 sg13g2_fill_2 FILLER_21_751 ();
 sg13g2_decap_8 FILLER_21_761 ();
 sg13g2_fill_2 FILLER_21_768 ();
 sg13g2_decap_8 FILLER_21_787 ();
 sg13g2_decap_4 FILLER_21_794 ();
 sg13g2_fill_2 FILLER_21_798 ();
 sg13g2_decap_4 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_fill_2 FILLER_21_837 ();
 sg13g2_fill_1 FILLER_21_839 ();
 sg13g2_fill_1 FILLER_21_927 ();
 sg13g2_decap_8 FILLER_21_1136 ();
 sg13g2_decap_8 FILLER_21_1143 ();
 sg13g2_decap_8 FILLER_21_1150 ();
 sg13g2_decap_8 FILLER_21_1157 ();
 sg13g2_decap_8 FILLER_21_1164 ();
 sg13g2_decap_8 FILLER_21_1171 ();
 sg13g2_decap_8 FILLER_21_1178 ();
 sg13g2_decap_8 FILLER_21_1185 ();
 sg13g2_decap_8 FILLER_21_1192 ();
 sg13g2_decap_8 FILLER_21_1199 ();
 sg13g2_decap_8 FILLER_21_1206 ();
 sg13g2_decap_8 FILLER_21_1213 ();
 sg13g2_decap_8 FILLER_21_1220 ();
 sg13g2_decap_8 FILLER_21_1227 ();
 sg13g2_decap_8 FILLER_21_1234 ();
 sg13g2_decap_8 FILLER_21_1241 ();
 sg13g2_decap_8 FILLER_21_1248 ();
 sg13g2_decap_8 FILLER_21_1255 ();
 sg13g2_decap_8 FILLER_21_1262 ();
 sg13g2_decap_8 FILLER_21_1269 ();
 sg13g2_decap_8 FILLER_21_1276 ();
 sg13g2_decap_8 FILLER_21_1283 ();
 sg13g2_decap_8 FILLER_21_1290 ();
 sg13g2_decap_8 FILLER_21_1297 ();
 sg13g2_decap_8 FILLER_21_1304 ();
 sg13g2_decap_4 FILLER_21_1311 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_fill_2 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_65 ();
 sg13g2_fill_2 FILLER_22_92 ();
 sg13g2_decap_4 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_170 ();
 sg13g2_fill_1 FILLER_22_180 ();
 sg13g2_fill_2 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_232 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_364 ();
 sg13g2_fill_2 FILLER_22_377 ();
 sg13g2_fill_2 FILLER_22_384 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_decap_4 FILLER_22_430 ();
 sg13g2_fill_2 FILLER_22_450 ();
 sg13g2_fill_1 FILLER_22_452 ();
 sg13g2_fill_2 FILLER_22_457 ();
 sg13g2_fill_1 FILLER_22_473 ();
 sg13g2_fill_2 FILLER_22_500 ();
 sg13g2_decap_8 FILLER_22_524 ();
 sg13g2_fill_2 FILLER_22_531 ();
 sg13g2_fill_1 FILLER_22_533 ();
 sg13g2_fill_1 FILLER_22_544 ();
 sg13g2_fill_1 FILLER_22_558 ();
 sg13g2_fill_2 FILLER_22_565 ();
 sg13g2_fill_1 FILLER_22_567 ();
 sg13g2_fill_2 FILLER_22_647 ();
 sg13g2_fill_1 FILLER_22_649 ();
 sg13g2_fill_1 FILLER_22_707 ();
 sg13g2_fill_2 FILLER_22_756 ();
 sg13g2_fill_2 FILLER_22_779 ();
 sg13g2_fill_1 FILLER_22_793 ();
 sg13g2_fill_2 FILLER_22_861 ();
 sg13g2_fill_1 FILLER_22_863 ();
 sg13g2_fill_2 FILLER_22_894 ();
 sg13g2_fill_2 FILLER_22_952 ();
 sg13g2_fill_2 FILLER_22_963 ();
 sg13g2_fill_2 FILLER_22_983 ();
 sg13g2_fill_1 FILLER_22_985 ();
 sg13g2_fill_2 FILLER_22_1094 ();
 sg13g2_decap_8 FILLER_22_1131 ();
 sg13g2_decap_8 FILLER_22_1138 ();
 sg13g2_decap_8 FILLER_22_1145 ();
 sg13g2_decap_8 FILLER_22_1152 ();
 sg13g2_decap_8 FILLER_22_1159 ();
 sg13g2_decap_8 FILLER_22_1166 ();
 sg13g2_decap_8 FILLER_22_1173 ();
 sg13g2_decap_8 FILLER_22_1180 ();
 sg13g2_decap_8 FILLER_22_1187 ();
 sg13g2_decap_8 FILLER_22_1194 ();
 sg13g2_decap_8 FILLER_22_1201 ();
 sg13g2_decap_8 FILLER_22_1208 ();
 sg13g2_decap_8 FILLER_22_1215 ();
 sg13g2_decap_8 FILLER_22_1222 ();
 sg13g2_decap_8 FILLER_22_1229 ();
 sg13g2_decap_8 FILLER_22_1236 ();
 sg13g2_decap_8 FILLER_22_1243 ();
 sg13g2_decap_8 FILLER_22_1250 ();
 sg13g2_decap_8 FILLER_22_1257 ();
 sg13g2_decap_8 FILLER_22_1264 ();
 sg13g2_decap_8 FILLER_22_1271 ();
 sg13g2_decap_8 FILLER_22_1278 ();
 sg13g2_decap_8 FILLER_22_1285 ();
 sg13g2_decap_8 FILLER_22_1292 ();
 sg13g2_decap_8 FILLER_22_1299 ();
 sg13g2_decap_8 FILLER_22_1306 ();
 sg13g2_fill_2 FILLER_22_1313 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_fill_2 FILLER_23_198 ();
 sg13g2_fill_2 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_fill_1 FILLER_23_389 ();
 sg13g2_decap_4 FILLER_23_400 ();
 sg13g2_decap_8 FILLER_23_418 ();
 sg13g2_fill_2 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_437 ();
 sg13g2_decap_8 FILLER_23_478 ();
 sg13g2_decap_8 FILLER_23_489 ();
 sg13g2_fill_1 FILLER_23_496 ();
 sg13g2_fill_2 FILLER_23_507 ();
 sg13g2_fill_1 FILLER_23_518 ();
 sg13g2_fill_1 FILLER_23_541 ();
 sg13g2_decap_8 FILLER_23_554 ();
 sg13g2_fill_2 FILLER_23_561 ();
 sg13g2_fill_2 FILLER_23_578 ();
 sg13g2_fill_1 FILLER_23_586 ();
 sg13g2_fill_1 FILLER_23_642 ();
 sg13g2_fill_1 FILLER_23_676 ();
 sg13g2_fill_1 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_736 ();
 sg13g2_decap_4 FILLER_23_769 ();
 sg13g2_fill_2 FILLER_23_773 ();
 sg13g2_decap_8 FILLER_23_778 ();
 sg13g2_decap_4 FILLER_23_785 ();
 sg13g2_decap_4 FILLER_23_807 ();
 sg13g2_decap_8 FILLER_23_815 ();
 sg13g2_fill_1 FILLER_23_822 ();
 sg13g2_decap_8 FILLER_23_832 ();
 sg13g2_fill_1 FILLER_23_875 ();
 sg13g2_fill_2 FILLER_23_1036 ();
 sg13g2_fill_1 FILLER_23_1038 ();
 sg13g2_fill_2 FILLER_23_1062 ();
 sg13g2_fill_1 FILLER_23_1064 ();
 sg13g2_decap_8 FILLER_23_1117 ();
 sg13g2_decap_8 FILLER_23_1124 ();
 sg13g2_decap_8 FILLER_23_1131 ();
 sg13g2_decap_8 FILLER_23_1138 ();
 sg13g2_decap_8 FILLER_23_1145 ();
 sg13g2_decap_8 FILLER_23_1152 ();
 sg13g2_decap_8 FILLER_23_1159 ();
 sg13g2_decap_8 FILLER_23_1166 ();
 sg13g2_decap_8 FILLER_23_1173 ();
 sg13g2_decap_8 FILLER_23_1180 ();
 sg13g2_decap_8 FILLER_23_1187 ();
 sg13g2_decap_8 FILLER_23_1194 ();
 sg13g2_decap_8 FILLER_23_1201 ();
 sg13g2_decap_8 FILLER_23_1208 ();
 sg13g2_decap_8 FILLER_23_1215 ();
 sg13g2_decap_8 FILLER_23_1222 ();
 sg13g2_decap_8 FILLER_23_1229 ();
 sg13g2_decap_8 FILLER_23_1236 ();
 sg13g2_decap_8 FILLER_23_1243 ();
 sg13g2_decap_8 FILLER_23_1250 ();
 sg13g2_decap_8 FILLER_23_1257 ();
 sg13g2_decap_8 FILLER_23_1264 ();
 sg13g2_decap_8 FILLER_23_1271 ();
 sg13g2_decap_8 FILLER_23_1278 ();
 sg13g2_decap_8 FILLER_23_1285 ();
 sg13g2_decap_8 FILLER_23_1292 ();
 sg13g2_decap_8 FILLER_23_1299 ();
 sg13g2_decap_8 FILLER_23_1306 ();
 sg13g2_fill_2 FILLER_23_1313 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_51 ();
 sg13g2_decap_4 FILLER_24_115 ();
 sg13g2_fill_2 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_fill_2 FILLER_24_309 ();
 sg13g2_decap_4 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_380 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_fill_1 FILLER_24_409 ();
 sg13g2_fill_2 FILLER_24_464 ();
 sg13g2_fill_1 FILLER_24_488 ();
 sg13g2_decap_8 FILLER_24_498 ();
 sg13g2_decap_4 FILLER_24_505 ();
 sg13g2_fill_1 FILLER_24_509 ();
 sg13g2_fill_1 FILLER_24_541 ();
 sg13g2_fill_2 FILLER_24_546 ();
 sg13g2_fill_2 FILLER_24_566 ();
 sg13g2_fill_2 FILLER_24_587 ();
 sg13g2_fill_1 FILLER_24_622 ();
 sg13g2_decap_8 FILLER_24_649 ();
 sg13g2_decap_8 FILLER_24_656 ();
 sg13g2_fill_2 FILLER_24_663 ();
 sg13g2_fill_1 FILLER_24_665 ();
 sg13g2_fill_1 FILLER_24_702 ();
 sg13g2_decap_4 FILLER_24_716 ();
 sg13g2_fill_1 FILLER_24_733 ();
 sg13g2_decap_4 FILLER_24_769 ();
 sg13g2_fill_1 FILLER_24_773 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_4 FILLER_24_791 ();
 sg13g2_fill_2 FILLER_24_795 ();
 sg13g2_decap_4 FILLER_24_807 ();
 sg13g2_fill_2 FILLER_24_811 ();
 sg13g2_fill_1 FILLER_24_817 ();
 sg13g2_decap_8 FILLER_24_828 ();
 sg13g2_fill_1 FILLER_24_835 ();
 sg13g2_decap_8 FILLER_24_841 ();
 sg13g2_fill_1 FILLER_24_848 ();
 sg13g2_fill_2 FILLER_24_853 ();
 sg13g2_fill_2 FILLER_24_864 ();
 sg13g2_fill_1 FILLER_24_866 ();
 sg13g2_decap_4 FILLER_24_912 ();
 sg13g2_fill_2 FILLER_24_916 ();
 sg13g2_fill_2 FILLER_24_922 ();
 sg13g2_fill_2 FILLER_24_928 ();
 sg13g2_fill_1 FILLER_24_951 ();
 sg13g2_decap_8 FILLER_24_1121 ();
 sg13g2_decap_8 FILLER_24_1128 ();
 sg13g2_decap_8 FILLER_24_1135 ();
 sg13g2_decap_8 FILLER_24_1142 ();
 sg13g2_decap_8 FILLER_24_1149 ();
 sg13g2_decap_8 FILLER_24_1156 ();
 sg13g2_decap_8 FILLER_24_1163 ();
 sg13g2_decap_8 FILLER_24_1170 ();
 sg13g2_decap_8 FILLER_24_1177 ();
 sg13g2_decap_8 FILLER_24_1184 ();
 sg13g2_decap_8 FILLER_24_1191 ();
 sg13g2_decap_8 FILLER_24_1198 ();
 sg13g2_decap_8 FILLER_24_1205 ();
 sg13g2_decap_8 FILLER_24_1212 ();
 sg13g2_decap_8 FILLER_24_1219 ();
 sg13g2_decap_8 FILLER_24_1226 ();
 sg13g2_decap_8 FILLER_24_1233 ();
 sg13g2_decap_8 FILLER_24_1240 ();
 sg13g2_decap_8 FILLER_24_1247 ();
 sg13g2_decap_8 FILLER_24_1254 ();
 sg13g2_decap_8 FILLER_24_1261 ();
 sg13g2_decap_8 FILLER_24_1268 ();
 sg13g2_decap_8 FILLER_24_1275 ();
 sg13g2_decap_8 FILLER_24_1282 ();
 sg13g2_decap_8 FILLER_24_1289 ();
 sg13g2_decap_8 FILLER_24_1296 ();
 sg13g2_decap_8 FILLER_24_1303 ();
 sg13g2_decap_4 FILLER_24_1310 ();
 sg13g2_fill_1 FILLER_24_1314 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_4 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_85 ();
 sg13g2_decap_4 FILLER_25_92 ();
 sg13g2_fill_2 FILLER_25_96 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_fill_2 FILLER_25_291 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_decap_4 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_fill_2 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_4 FILLER_25_420 ();
 sg13g2_fill_2 FILLER_25_424 ();
 sg13g2_decap_4 FILLER_25_430 ();
 sg13g2_fill_2 FILLER_25_434 ();
 sg13g2_fill_2 FILLER_25_453 ();
 sg13g2_fill_1 FILLER_25_455 ();
 sg13g2_decap_4 FILLER_25_512 ();
 sg13g2_decap_8 FILLER_25_526 ();
 sg13g2_decap_4 FILLER_25_533 ();
 sg13g2_fill_1 FILLER_25_537 ();
 sg13g2_fill_2 FILLER_25_541 ();
 sg13g2_fill_1 FILLER_25_543 ();
 sg13g2_fill_1 FILLER_25_563 ();
 sg13g2_fill_1 FILLER_25_578 ();
 sg13g2_fill_2 FILLER_25_592 ();
 sg13g2_fill_1 FILLER_25_594 ();
 sg13g2_fill_2 FILLER_25_613 ();
 sg13g2_fill_1 FILLER_25_615 ();
 sg13g2_decap_8 FILLER_25_668 ();
 sg13g2_fill_1 FILLER_25_675 ();
 sg13g2_decap_4 FILLER_25_712 ();
 sg13g2_fill_1 FILLER_25_716 ();
 sg13g2_fill_2 FILLER_25_758 ();
 sg13g2_fill_1 FILLER_25_772 ();
 sg13g2_fill_1 FILLER_25_797 ();
 sg13g2_fill_2 FILLER_25_806 ();
 sg13g2_fill_1 FILLER_25_819 ();
 sg13g2_fill_2 FILLER_25_826 ();
 sg13g2_decap_4 FILLER_25_854 ();
 sg13g2_fill_2 FILLER_25_858 ();
 sg13g2_fill_2 FILLER_25_878 ();
 sg13g2_fill_2 FILLER_25_1044 ();
 sg13g2_fill_2 FILLER_25_1072 ();
 sg13g2_decap_8 FILLER_25_1129 ();
 sg13g2_decap_8 FILLER_25_1136 ();
 sg13g2_decap_8 FILLER_25_1143 ();
 sg13g2_decap_8 FILLER_25_1150 ();
 sg13g2_decap_8 FILLER_25_1157 ();
 sg13g2_decap_8 FILLER_25_1164 ();
 sg13g2_decap_8 FILLER_25_1171 ();
 sg13g2_decap_8 FILLER_25_1178 ();
 sg13g2_decap_8 FILLER_25_1185 ();
 sg13g2_decap_8 FILLER_25_1192 ();
 sg13g2_decap_8 FILLER_25_1199 ();
 sg13g2_decap_8 FILLER_25_1206 ();
 sg13g2_decap_8 FILLER_25_1213 ();
 sg13g2_decap_8 FILLER_25_1220 ();
 sg13g2_decap_8 FILLER_25_1227 ();
 sg13g2_decap_8 FILLER_25_1234 ();
 sg13g2_decap_8 FILLER_25_1241 ();
 sg13g2_decap_8 FILLER_25_1248 ();
 sg13g2_decap_8 FILLER_25_1255 ();
 sg13g2_decap_8 FILLER_25_1262 ();
 sg13g2_decap_8 FILLER_25_1269 ();
 sg13g2_decap_8 FILLER_25_1276 ();
 sg13g2_decap_8 FILLER_25_1283 ();
 sg13g2_decap_8 FILLER_25_1290 ();
 sg13g2_decap_8 FILLER_25_1297 ();
 sg13g2_decap_8 FILLER_25_1304 ();
 sg13g2_decap_4 FILLER_25_1311 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_4 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_53 ();
 sg13g2_fill_1 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_107 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_fill_2 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_350 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_fill_2 FILLER_26_383 ();
 sg13g2_fill_1 FILLER_26_385 ();
 sg13g2_fill_2 FILLER_26_391 ();
 sg13g2_fill_1 FILLER_26_464 ();
 sg13g2_fill_2 FILLER_26_483 ();
 sg13g2_fill_1 FILLER_26_560 ();
 sg13g2_fill_2 FILLER_26_588 ();
 sg13g2_fill_1 FILLER_26_590 ();
 sg13g2_decap_4 FILLER_26_683 ();
 sg13g2_fill_2 FILLER_26_687 ();
 sg13g2_fill_2 FILLER_26_694 ();
 sg13g2_fill_2 FILLER_26_714 ();
 sg13g2_fill_2 FILLER_26_745 ();
 sg13g2_fill_1 FILLER_26_752 ();
 sg13g2_decap_4 FILLER_26_773 ();
 sg13g2_fill_1 FILLER_26_777 ();
 sg13g2_fill_2 FILLER_26_788 ();
 sg13g2_fill_1 FILLER_26_790 ();
 sg13g2_fill_1 FILLER_26_801 ();
 sg13g2_fill_2 FILLER_26_807 ();
 sg13g2_fill_1 FILLER_26_809 ();
 sg13g2_decap_4 FILLER_26_848 ();
 sg13g2_fill_1 FILLER_26_852 ();
 sg13g2_decap_8 FILLER_26_889 ();
 sg13g2_decap_4 FILLER_26_896 ();
 sg13g2_fill_2 FILLER_26_939 ();
 sg13g2_fill_2 FILLER_26_985 ();
 sg13g2_fill_1 FILLER_26_1026 ();
 sg13g2_fill_1 FILLER_26_1058 ();
 sg13g2_fill_1 FILLER_26_1072 ();
 sg13g2_decap_8 FILLER_26_1128 ();
 sg13g2_decap_8 FILLER_26_1135 ();
 sg13g2_decap_8 FILLER_26_1142 ();
 sg13g2_decap_8 FILLER_26_1149 ();
 sg13g2_decap_8 FILLER_26_1156 ();
 sg13g2_decap_8 FILLER_26_1163 ();
 sg13g2_decap_8 FILLER_26_1170 ();
 sg13g2_decap_8 FILLER_26_1177 ();
 sg13g2_decap_8 FILLER_26_1184 ();
 sg13g2_decap_8 FILLER_26_1191 ();
 sg13g2_decap_8 FILLER_26_1198 ();
 sg13g2_decap_8 FILLER_26_1205 ();
 sg13g2_decap_8 FILLER_26_1212 ();
 sg13g2_decap_8 FILLER_26_1219 ();
 sg13g2_decap_8 FILLER_26_1226 ();
 sg13g2_decap_8 FILLER_26_1233 ();
 sg13g2_decap_8 FILLER_26_1240 ();
 sg13g2_decap_8 FILLER_26_1247 ();
 sg13g2_decap_8 FILLER_26_1254 ();
 sg13g2_decap_8 FILLER_26_1261 ();
 sg13g2_decap_8 FILLER_26_1268 ();
 sg13g2_decap_8 FILLER_26_1275 ();
 sg13g2_decap_8 FILLER_26_1282 ();
 sg13g2_decap_8 FILLER_26_1289 ();
 sg13g2_decap_8 FILLER_26_1296 ();
 sg13g2_decap_8 FILLER_26_1303 ();
 sg13g2_decap_4 FILLER_26_1310 ();
 sg13g2_fill_1 FILLER_26_1314 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_177 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_fill_2 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_296 ();
 sg13g2_decap_4 FILLER_27_307 ();
 sg13g2_fill_2 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_decap_4 FILLER_27_324 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_fill_2 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_388 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_fill_2 FILLER_27_404 ();
 sg13g2_fill_2 FILLER_27_411 ();
 sg13g2_fill_1 FILLER_27_413 ();
 sg13g2_fill_2 FILLER_27_430 ();
 sg13g2_decap_4 FILLER_27_441 ();
 sg13g2_fill_2 FILLER_27_445 ();
 sg13g2_fill_2 FILLER_27_514 ();
 sg13g2_fill_1 FILLER_27_530 ();
 sg13g2_decap_8 FILLER_27_535 ();
 sg13g2_decap_4 FILLER_27_542 ();
 sg13g2_fill_1 FILLER_27_581 ();
 sg13g2_fill_1 FILLER_27_594 ();
 sg13g2_fill_1 FILLER_27_647 ();
 sg13g2_decap_4 FILLER_27_693 ();
 sg13g2_fill_1 FILLER_27_774 ();
 sg13g2_fill_2 FILLER_27_796 ();
 sg13g2_fill_2 FILLER_27_804 ();
 sg13g2_fill_1 FILLER_27_816 ();
 sg13g2_fill_2 FILLER_27_823 ();
 sg13g2_fill_2 FILLER_27_837 ();
 sg13g2_fill_2 FILLER_27_849 ();
 sg13g2_fill_1 FILLER_27_851 ();
 sg13g2_fill_2 FILLER_27_882 ();
 sg13g2_decap_8 FILLER_27_903 ();
 sg13g2_fill_2 FILLER_27_910 ();
 sg13g2_fill_1 FILLER_27_912 ();
 sg13g2_fill_2 FILLER_27_922 ();
 sg13g2_fill_2 FILLER_27_968 ();
 sg13g2_fill_1 FILLER_27_1026 ();
 sg13g2_decap_8 FILLER_27_1131 ();
 sg13g2_decap_8 FILLER_27_1138 ();
 sg13g2_decap_8 FILLER_27_1145 ();
 sg13g2_decap_8 FILLER_27_1152 ();
 sg13g2_decap_8 FILLER_27_1159 ();
 sg13g2_decap_8 FILLER_27_1166 ();
 sg13g2_decap_8 FILLER_27_1173 ();
 sg13g2_decap_8 FILLER_27_1180 ();
 sg13g2_decap_8 FILLER_27_1187 ();
 sg13g2_decap_8 FILLER_27_1194 ();
 sg13g2_decap_8 FILLER_27_1201 ();
 sg13g2_decap_8 FILLER_27_1208 ();
 sg13g2_decap_8 FILLER_27_1215 ();
 sg13g2_decap_8 FILLER_27_1222 ();
 sg13g2_decap_8 FILLER_27_1229 ();
 sg13g2_decap_8 FILLER_27_1236 ();
 sg13g2_decap_8 FILLER_27_1243 ();
 sg13g2_decap_8 FILLER_27_1250 ();
 sg13g2_decap_8 FILLER_27_1257 ();
 sg13g2_decap_8 FILLER_27_1264 ();
 sg13g2_decap_8 FILLER_27_1271 ();
 sg13g2_decap_8 FILLER_27_1278 ();
 sg13g2_decap_8 FILLER_27_1285 ();
 sg13g2_decap_8 FILLER_27_1292 ();
 sg13g2_decap_8 FILLER_27_1299 ();
 sg13g2_decap_8 FILLER_27_1306 ();
 sg13g2_fill_2 FILLER_27_1313 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_37 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_fill_2 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_370 ();
 sg13g2_fill_1 FILLER_28_460 ();
 sg13g2_fill_2 FILLER_28_470 ();
 sg13g2_fill_1 FILLER_28_472 ();
 sg13g2_fill_2 FILLER_28_477 ();
 sg13g2_fill_1 FILLER_28_479 ();
 sg13g2_fill_1 FILLER_28_516 ();
 sg13g2_fill_2 FILLER_28_543 ();
 sg13g2_decap_8 FILLER_28_550 ();
 sg13g2_fill_2 FILLER_28_557 ();
 sg13g2_fill_1 FILLER_28_559 ();
 sg13g2_decap_8 FILLER_28_564 ();
 sg13g2_fill_2 FILLER_28_576 ();
 sg13g2_fill_1 FILLER_28_598 ();
 sg13g2_fill_2 FILLER_28_635 ();
 sg13g2_fill_1 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_696 ();
 sg13g2_decap_4 FILLER_28_703 ();
 sg13g2_fill_1 FILLER_28_707 ();
 sg13g2_decap_4 FILLER_28_712 ();
 sg13g2_fill_1 FILLER_28_716 ();
 sg13g2_fill_2 FILLER_28_730 ();
 sg13g2_fill_1 FILLER_28_732 ();
 sg13g2_fill_2 FILLER_28_742 ();
 sg13g2_fill_1 FILLER_28_744 ();
 sg13g2_fill_1 FILLER_28_755 ();
 sg13g2_fill_1 FILLER_28_761 ();
 sg13g2_decap_8 FILLER_28_767 ();
 sg13g2_fill_2 FILLER_28_774 ();
 sg13g2_fill_1 FILLER_28_782 ();
 sg13g2_fill_2 FILLER_28_789 ();
 sg13g2_fill_2 FILLER_28_812 ();
 sg13g2_fill_2 FILLER_28_819 ();
 sg13g2_fill_1 FILLER_28_821 ();
 sg13g2_fill_2 FILLER_28_854 ();
 sg13g2_fill_1 FILLER_28_879 ();
 sg13g2_fill_1 FILLER_28_958 ();
 sg13g2_fill_2 FILLER_28_985 ();
 sg13g2_fill_1 FILLER_28_987 ();
 sg13g2_fill_1 FILLER_28_1112 ();
 sg13g2_decap_8 FILLER_28_1130 ();
 sg13g2_decap_8 FILLER_28_1137 ();
 sg13g2_decap_8 FILLER_28_1144 ();
 sg13g2_decap_8 FILLER_28_1151 ();
 sg13g2_decap_8 FILLER_28_1158 ();
 sg13g2_decap_8 FILLER_28_1165 ();
 sg13g2_decap_8 FILLER_28_1172 ();
 sg13g2_decap_8 FILLER_28_1179 ();
 sg13g2_decap_8 FILLER_28_1186 ();
 sg13g2_decap_8 FILLER_28_1193 ();
 sg13g2_decap_8 FILLER_28_1200 ();
 sg13g2_decap_8 FILLER_28_1207 ();
 sg13g2_decap_8 FILLER_28_1214 ();
 sg13g2_decap_8 FILLER_28_1221 ();
 sg13g2_decap_8 FILLER_28_1228 ();
 sg13g2_decap_8 FILLER_28_1235 ();
 sg13g2_decap_8 FILLER_28_1242 ();
 sg13g2_decap_8 FILLER_28_1249 ();
 sg13g2_decap_8 FILLER_28_1256 ();
 sg13g2_decap_8 FILLER_28_1263 ();
 sg13g2_decap_8 FILLER_28_1270 ();
 sg13g2_decap_8 FILLER_28_1277 ();
 sg13g2_decap_8 FILLER_28_1284 ();
 sg13g2_decap_8 FILLER_28_1291 ();
 sg13g2_decap_8 FILLER_28_1298 ();
 sg13g2_decap_8 FILLER_28_1305 ();
 sg13g2_fill_2 FILLER_28_1312 ();
 sg13g2_fill_1 FILLER_28_1314 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_74 ();
 sg13g2_decap_4 FILLER_29_102 ();
 sg13g2_fill_2 FILLER_29_106 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_fill_2 FILLER_29_156 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_180 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_301 ();
 sg13g2_decap_4 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_361 ();
 sg13g2_decap_4 FILLER_29_368 ();
 sg13g2_decap_4 FILLER_29_377 ();
 sg13g2_fill_1 FILLER_29_381 ();
 sg13g2_fill_2 FILLER_29_391 ();
 sg13g2_fill_1 FILLER_29_393 ();
 sg13g2_fill_1 FILLER_29_398 ();
 sg13g2_fill_2 FILLER_29_425 ();
 sg13g2_fill_1 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_432 ();
 sg13g2_decap_4 FILLER_29_478 ();
 sg13g2_decap_8 FILLER_29_492 ();
 sg13g2_decap_4 FILLER_29_516 ();
 sg13g2_fill_1 FILLER_29_520 ();
 sg13g2_fill_2 FILLER_29_524 ();
 sg13g2_fill_1 FILLER_29_526 ();
 sg13g2_fill_2 FILLER_29_571 ();
 sg13g2_fill_1 FILLER_29_573 ();
 sg13g2_fill_2 FILLER_29_591 ();
 sg13g2_fill_2 FILLER_29_612 ();
 sg13g2_decap_4 FILLER_29_677 ();
 sg13g2_fill_2 FILLER_29_689 ();
 sg13g2_decap_4 FILLER_29_717 ();
 sg13g2_fill_2 FILLER_29_721 ();
 sg13g2_decap_4 FILLER_29_750 ();
 sg13g2_decap_4 FILLER_29_776 ();
 sg13g2_fill_1 FILLER_29_780 ();
 sg13g2_fill_1 FILLER_29_786 ();
 sg13g2_decap_4 FILLER_29_791 ();
 sg13g2_fill_2 FILLER_29_795 ();
 sg13g2_fill_1 FILLER_29_802 ();
 sg13g2_decap_4 FILLER_29_829 ();
 sg13g2_decap_8 FILLER_29_859 ();
 sg13g2_decap_4 FILLER_29_866 ();
 sg13g2_fill_2 FILLER_29_893 ();
 sg13g2_fill_1 FILLER_29_895 ();
 sg13g2_decap_4 FILLER_29_909 ();
 sg13g2_fill_1 FILLER_29_913 ();
 sg13g2_fill_2 FILLER_29_918 ();
 sg13g2_fill_1 FILLER_29_920 ();
 sg13g2_fill_2 FILLER_29_930 ();
 sg13g2_fill_1 FILLER_29_949 ();
 sg13g2_fill_1 FILLER_29_980 ();
 sg13g2_fill_1 FILLER_29_1016 ();
 sg13g2_fill_2 FILLER_29_1078 ();
 sg13g2_fill_1 FILLER_29_1089 ();
 sg13g2_decap_8 FILLER_29_1133 ();
 sg13g2_decap_8 FILLER_29_1140 ();
 sg13g2_decap_8 FILLER_29_1147 ();
 sg13g2_decap_8 FILLER_29_1154 ();
 sg13g2_decap_8 FILLER_29_1161 ();
 sg13g2_decap_8 FILLER_29_1168 ();
 sg13g2_decap_8 FILLER_29_1175 ();
 sg13g2_decap_8 FILLER_29_1182 ();
 sg13g2_decap_8 FILLER_29_1189 ();
 sg13g2_decap_8 FILLER_29_1196 ();
 sg13g2_decap_8 FILLER_29_1203 ();
 sg13g2_decap_8 FILLER_29_1210 ();
 sg13g2_decap_8 FILLER_29_1217 ();
 sg13g2_decap_8 FILLER_29_1224 ();
 sg13g2_decap_8 FILLER_29_1231 ();
 sg13g2_decap_8 FILLER_29_1238 ();
 sg13g2_decap_8 FILLER_29_1245 ();
 sg13g2_decap_8 FILLER_29_1252 ();
 sg13g2_decap_8 FILLER_29_1259 ();
 sg13g2_decap_8 FILLER_29_1266 ();
 sg13g2_decap_8 FILLER_29_1273 ();
 sg13g2_decap_8 FILLER_29_1280 ();
 sg13g2_decap_8 FILLER_29_1287 ();
 sg13g2_decap_8 FILLER_29_1294 ();
 sg13g2_decap_8 FILLER_29_1301 ();
 sg13g2_decap_8 FILLER_29_1308 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_73 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_fill_2 FILLER_30_132 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_309 ();
 sg13g2_fill_1 FILLER_30_394 ();
 sg13g2_fill_2 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_406 ();
 sg13g2_fill_2 FILLER_30_442 ();
 sg13g2_fill_1 FILLER_30_444 ();
 sg13g2_fill_2 FILLER_30_449 ();
 sg13g2_fill_1 FILLER_30_459 ();
 sg13g2_fill_2 FILLER_30_529 ();
 sg13g2_fill_1 FILLER_30_531 ();
 sg13g2_fill_1 FILLER_30_536 ();
 sg13g2_fill_1 FILLER_30_555 ();
 sg13g2_fill_2 FILLER_30_562 ();
 sg13g2_fill_1 FILLER_30_564 ();
 sg13g2_fill_1 FILLER_30_570 ();
 sg13g2_fill_2 FILLER_30_575 ();
 sg13g2_fill_2 FILLER_30_582 ();
 sg13g2_fill_1 FILLER_30_596 ();
 sg13g2_fill_1 FILLER_30_605 ();
 sg13g2_fill_2 FILLER_30_621 ();
 sg13g2_fill_1 FILLER_30_680 ();
 sg13g2_fill_2 FILLER_30_687 ();
 sg13g2_fill_1 FILLER_30_689 ();
 sg13g2_fill_2 FILLER_30_699 ();
 sg13g2_fill_1 FILLER_30_701 ();
 sg13g2_fill_2 FILLER_30_706 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_fill_1 FILLER_30_735 ();
 sg13g2_decap_4 FILLER_30_741 ();
 sg13g2_fill_2 FILLER_30_745 ();
 sg13g2_fill_2 FILLER_30_790 ();
 sg13g2_fill_1 FILLER_30_792 ();
 sg13g2_fill_2 FILLER_30_809 ();
 sg13g2_fill_1 FILLER_30_811 ();
 sg13g2_fill_2 FILLER_30_829 ();
 sg13g2_fill_1 FILLER_30_831 ();
 sg13g2_fill_2 FILLER_30_858 ();
 sg13g2_fill_1 FILLER_30_860 ();
 sg13g2_decap_4 FILLER_30_891 ();
 sg13g2_fill_2 FILLER_30_956 ();
 sg13g2_fill_1 FILLER_30_1010 ();
 sg13g2_fill_1 FILLER_30_1037 ();
 sg13g2_fill_1 FILLER_30_1120 ();
 sg13g2_decap_8 FILLER_30_1130 ();
 sg13g2_decap_8 FILLER_30_1137 ();
 sg13g2_decap_8 FILLER_30_1144 ();
 sg13g2_decap_8 FILLER_30_1151 ();
 sg13g2_decap_8 FILLER_30_1158 ();
 sg13g2_decap_8 FILLER_30_1165 ();
 sg13g2_decap_8 FILLER_30_1172 ();
 sg13g2_decap_8 FILLER_30_1179 ();
 sg13g2_decap_8 FILLER_30_1186 ();
 sg13g2_decap_8 FILLER_30_1193 ();
 sg13g2_decap_8 FILLER_30_1200 ();
 sg13g2_decap_8 FILLER_30_1207 ();
 sg13g2_decap_8 FILLER_30_1214 ();
 sg13g2_decap_8 FILLER_30_1221 ();
 sg13g2_decap_8 FILLER_30_1228 ();
 sg13g2_decap_8 FILLER_30_1235 ();
 sg13g2_decap_8 FILLER_30_1242 ();
 sg13g2_decap_8 FILLER_30_1249 ();
 sg13g2_decap_8 FILLER_30_1256 ();
 sg13g2_decap_8 FILLER_30_1263 ();
 sg13g2_decap_8 FILLER_30_1270 ();
 sg13g2_decap_8 FILLER_30_1277 ();
 sg13g2_decap_8 FILLER_30_1284 ();
 sg13g2_decap_8 FILLER_30_1291 ();
 sg13g2_decap_8 FILLER_30_1298 ();
 sg13g2_decap_8 FILLER_30_1305 ();
 sg13g2_fill_2 FILLER_30_1312 ();
 sg13g2_fill_1 FILLER_30_1314 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_107 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_fill_1 FILLER_31_242 ();
 sg13g2_decap_8 FILLER_31_256 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_decap_4 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_decap_4 FILLER_31_367 ();
 sg13g2_fill_2 FILLER_31_419 ();
 sg13g2_fill_1 FILLER_31_421 ();
 sg13g2_decap_4 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_435 ();
 sg13g2_decap_4 FILLER_31_442 ();
 sg13g2_fill_1 FILLER_31_446 ();
 sg13g2_fill_2 FILLER_31_461 ();
 sg13g2_decap_4 FILLER_31_476 ();
 sg13g2_fill_1 FILLER_31_480 ();
 sg13g2_decap_8 FILLER_31_494 ();
 sg13g2_decap_4 FILLER_31_501 ();
 sg13g2_fill_2 FILLER_31_505 ();
 sg13g2_fill_2 FILLER_31_515 ();
 sg13g2_decap_8 FILLER_31_522 ();
 sg13g2_fill_1 FILLER_31_529 ();
 sg13g2_fill_2 FILLER_31_534 ();
 sg13g2_fill_1 FILLER_31_536 ();
 sg13g2_decap_8 FILLER_31_560 ();
 sg13g2_fill_1 FILLER_31_567 ();
 sg13g2_fill_1 FILLER_31_576 ();
 sg13g2_decap_8 FILLER_31_580 ();
 sg13g2_decap_8 FILLER_31_587 ();
 sg13g2_fill_2 FILLER_31_594 ();
 sg13g2_fill_1 FILLER_31_608 ();
 sg13g2_decap_4 FILLER_31_644 ();
 sg13g2_fill_1 FILLER_31_657 ();
 sg13g2_fill_2 FILLER_31_671 ();
 sg13g2_fill_2 FILLER_31_684 ();
 sg13g2_fill_1 FILLER_31_686 ();
 sg13g2_decap_4 FILLER_31_739 ();
 sg13g2_fill_2 FILLER_31_743 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_fill_1 FILLER_31_767 ();
 sg13g2_fill_1 FILLER_31_773 ();
 sg13g2_fill_2 FILLER_31_783 ();
 sg13g2_fill_1 FILLER_31_785 ();
 sg13g2_decap_8 FILLER_31_796 ();
 sg13g2_fill_2 FILLER_31_803 ();
 sg13g2_fill_1 FILLER_31_805 ();
 sg13g2_decap_4 FILLER_31_816 ();
 sg13g2_fill_1 FILLER_31_820 ();
 sg13g2_decap_4 FILLER_31_830 ();
 sg13g2_fill_2 FILLER_31_834 ();
 sg13g2_fill_2 FILLER_31_857 ();
 sg13g2_fill_2 FILLER_31_869 ();
 sg13g2_fill_2 FILLER_31_920 ();
 sg13g2_fill_1 FILLER_31_1023 ();
 sg13g2_fill_2 FILLER_31_1067 ();
 sg13g2_fill_1 FILLER_31_1069 ();
 sg13g2_decap_8 FILLER_31_1122 ();
 sg13g2_decap_8 FILLER_31_1129 ();
 sg13g2_decap_8 FILLER_31_1136 ();
 sg13g2_decap_8 FILLER_31_1143 ();
 sg13g2_decap_8 FILLER_31_1150 ();
 sg13g2_decap_8 FILLER_31_1157 ();
 sg13g2_decap_8 FILLER_31_1164 ();
 sg13g2_decap_8 FILLER_31_1171 ();
 sg13g2_decap_8 FILLER_31_1178 ();
 sg13g2_decap_8 FILLER_31_1185 ();
 sg13g2_decap_8 FILLER_31_1192 ();
 sg13g2_decap_8 FILLER_31_1199 ();
 sg13g2_decap_8 FILLER_31_1206 ();
 sg13g2_decap_8 FILLER_31_1213 ();
 sg13g2_decap_8 FILLER_31_1220 ();
 sg13g2_decap_8 FILLER_31_1227 ();
 sg13g2_decap_8 FILLER_31_1234 ();
 sg13g2_decap_8 FILLER_31_1241 ();
 sg13g2_decap_8 FILLER_31_1248 ();
 sg13g2_decap_8 FILLER_31_1255 ();
 sg13g2_decap_8 FILLER_31_1262 ();
 sg13g2_decap_8 FILLER_31_1269 ();
 sg13g2_decap_8 FILLER_31_1276 ();
 sg13g2_decap_8 FILLER_31_1283 ();
 sg13g2_decap_8 FILLER_31_1290 ();
 sg13g2_decap_8 FILLER_31_1297 ();
 sg13g2_decap_8 FILLER_31_1304 ();
 sg13g2_decap_4 FILLER_31_1311 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_22 ();
 sg13g2_fill_2 FILLER_32_29 ();
 sg13g2_fill_1 FILLER_32_31 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_fill_1 FILLER_32_90 ();
 sg13g2_fill_2 FILLER_32_112 ();
 sg13g2_fill_1 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_173 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_4 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_decap_4 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_fill_2 FILLER_32_321 ();
 sg13g2_decap_4 FILLER_32_339 ();
 sg13g2_fill_1 FILLER_32_343 ();
 sg13g2_decap_4 FILLER_32_365 ();
 sg13g2_fill_2 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_379 ();
 sg13g2_decap_4 FILLER_32_416 ();
 sg13g2_fill_2 FILLER_32_420 ();
 sg13g2_fill_2 FILLER_32_439 ();
 sg13g2_decap_4 FILLER_32_469 ();
 sg13g2_fill_2 FILLER_32_473 ();
 sg13g2_fill_2 FILLER_32_493 ();
 sg13g2_fill_1 FILLER_32_508 ();
 sg13g2_fill_2 FILLER_32_574 ();
 sg13g2_fill_1 FILLER_32_585 ();
 sg13g2_fill_2 FILLER_32_602 ();
 sg13g2_fill_2 FILLER_32_617 ();
 sg13g2_fill_1 FILLER_32_619 ();
 sg13g2_fill_2 FILLER_32_632 ();
 sg13g2_fill_1 FILLER_32_649 ();
 sg13g2_decap_4 FILLER_32_676 ();
 sg13g2_decap_8 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_701 ();
 sg13g2_decap_8 FILLER_32_708 ();
 sg13g2_decap_4 FILLER_32_715 ();
 sg13g2_fill_2 FILLER_32_719 ();
 sg13g2_decap_8 FILLER_32_725 ();
 sg13g2_fill_1 FILLER_32_732 ();
 sg13g2_fill_1 FILLER_32_766 ();
 sg13g2_fill_2 FILLER_32_780 ();
 sg13g2_fill_1 FILLER_32_782 ();
 sg13g2_fill_1 FILLER_32_789 ();
 sg13g2_fill_2 FILLER_32_798 ();
 sg13g2_fill_1 FILLER_32_800 ();
 sg13g2_fill_2 FILLER_32_837 ();
 sg13g2_fill_1 FILLER_32_839 ();
 sg13g2_decap_4 FILLER_32_844 ();
 sg13g2_fill_1 FILLER_32_848 ();
 sg13g2_fill_2 FILLER_32_905 ();
 sg13g2_decap_4 FILLER_32_968 ();
 sg13g2_decap_4 FILLER_32_984 ();
 sg13g2_fill_2 FILLER_32_1006 ();
 sg13g2_fill_1 FILLER_32_1008 ();
 sg13g2_fill_1 FILLER_32_1100 ();
 sg13g2_decap_8 FILLER_32_1136 ();
 sg13g2_decap_8 FILLER_32_1143 ();
 sg13g2_decap_8 FILLER_32_1150 ();
 sg13g2_decap_8 FILLER_32_1157 ();
 sg13g2_decap_8 FILLER_32_1164 ();
 sg13g2_decap_8 FILLER_32_1171 ();
 sg13g2_decap_8 FILLER_32_1178 ();
 sg13g2_decap_8 FILLER_32_1185 ();
 sg13g2_decap_8 FILLER_32_1192 ();
 sg13g2_decap_8 FILLER_32_1199 ();
 sg13g2_decap_8 FILLER_32_1206 ();
 sg13g2_decap_8 FILLER_32_1213 ();
 sg13g2_decap_8 FILLER_32_1220 ();
 sg13g2_decap_8 FILLER_32_1227 ();
 sg13g2_decap_8 FILLER_32_1234 ();
 sg13g2_decap_8 FILLER_32_1241 ();
 sg13g2_decap_8 FILLER_32_1248 ();
 sg13g2_decap_8 FILLER_32_1255 ();
 sg13g2_decap_8 FILLER_32_1262 ();
 sg13g2_decap_8 FILLER_32_1269 ();
 sg13g2_decap_8 FILLER_32_1276 ();
 sg13g2_decap_8 FILLER_32_1283 ();
 sg13g2_decap_8 FILLER_32_1290 ();
 sg13g2_decap_8 FILLER_32_1297 ();
 sg13g2_decap_8 FILLER_32_1304 ();
 sg13g2_decap_4 FILLER_32_1311 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_37 ();
 sg13g2_fill_2 FILLER_33_43 ();
 sg13g2_fill_1 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_fill_2 FILLER_33_108 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_fill_2 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_146 ();
 sg13g2_fill_2 FILLER_33_225 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_decap_4 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_decap_8 FILLER_33_299 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_decap_4 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_317 ();
 sg13g2_fill_1 FILLER_33_323 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_fill_2 FILLER_33_395 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_decap_4 FILLER_33_407 ();
 sg13g2_decap_4 FILLER_33_448 ();
 sg13g2_fill_2 FILLER_33_458 ();
 sg13g2_fill_1 FILLER_33_492 ();
 sg13g2_decap_8 FILLER_33_509 ();
 sg13g2_fill_2 FILLER_33_516 ();
 sg13g2_fill_1 FILLER_33_518 ();
 sg13g2_fill_1 FILLER_33_525 ();
 sg13g2_decap_4 FILLER_33_546 ();
 sg13g2_fill_2 FILLER_33_561 ();
 sg13g2_fill_1 FILLER_33_563 ();
 sg13g2_fill_2 FILLER_33_582 ();
 sg13g2_fill_2 FILLER_33_590 ();
 sg13g2_fill_2 FILLER_33_601 ();
 sg13g2_fill_1 FILLER_33_603 ();
 sg13g2_fill_1 FILLER_33_613 ();
 sg13g2_decap_4 FILLER_33_622 ();
 sg13g2_fill_1 FILLER_33_631 ();
 sg13g2_decap_4 FILLER_33_635 ();
 sg13g2_decap_8 FILLER_33_643 ();
 sg13g2_fill_2 FILLER_33_659 ();
 sg13g2_decap_4 FILLER_33_665 ();
 sg13g2_fill_1 FILLER_33_669 ();
 sg13g2_fill_2 FILLER_33_684 ();
 sg13g2_fill_2 FILLER_33_701 ();
 sg13g2_fill_2 FILLER_33_711 ();
 sg13g2_fill_1 FILLER_33_713 ();
 sg13g2_decap_4 FILLER_33_729 ();
 sg13g2_fill_1 FILLER_33_733 ();
 sg13g2_fill_2 FILLER_33_750 ();
 sg13g2_decap_4 FILLER_33_781 ();
 sg13g2_fill_2 FILLER_33_823 ();
 sg13g2_fill_1 FILLER_33_825 ();
 sg13g2_decap_8 FILLER_33_850 ();
 sg13g2_decap_8 FILLER_33_870 ();
 sg13g2_decap_4 FILLER_33_877 ();
 sg13g2_fill_2 FILLER_33_922 ();
 sg13g2_fill_1 FILLER_33_924 ();
 sg13g2_fill_2 FILLER_33_943 ();
 sg13g2_fill_1 FILLER_33_945 ();
 sg13g2_decap_4 FILLER_33_972 ();
 sg13g2_fill_2 FILLER_33_976 ();
 sg13g2_fill_1 FILLER_33_986 ();
 sg13g2_fill_1 FILLER_33_1040 ();
 sg13g2_fill_2 FILLER_33_1064 ();
 sg13g2_fill_1 FILLER_33_1066 ();
 sg13g2_fill_1 FILLER_33_1092 ();
 sg13g2_fill_1 FILLER_33_1106 ();
 sg13g2_decap_8 FILLER_33_1142 ();
 sg13g2_decap_8 FILLER_33_1149 ();
 sg13g2_decap_8 FILLER_33_1156 ();
 sg13g2_decap_8 FILLER_33_1163 ();
 sg13g2_decap_8 FILLER_33_1170 ();
 sg13g2_decap_8 FILLER_33_1177 ();
 sg13g2_decap_8 FILLER_33_1184 ();
 sg13g2_decap_8 FILLER_33_1191 ();
 sg13g2_decap_8 FILLER_33_1198 ();
 sg13g2_decap_8 FILLER_33_1205 ();
 sg13g2_decap_8 FILLER_33_1212 ();
 sg13g2_decap_8 FILLER_33_1219 ();
 sg13g2_decap_8 FILLER_33_1226 ();
 sg13g2_decap_8 FILLER_33_1233 ();
 sg13g2_decap_8 FILLER_33_1240 ();
 sg13g2_decap_8 FILLER_33_1247 ();
 sg13g2_decap_8 FILLER_33_1254 ();
 sg13g2_decap_8 FILLER_33_1261 ();
 sg13g2_decap_8 FILLER_33_1268 ();
 sg13g2_decap_8 FILLER_33_1275 ();
 sg13g2_decap_8 FILLER_33_1282 ();
 sg13g2_decap_8 FILLER_33_1289 ();
 sg13g2_decap_8 FILLER_33_1296 ();
 sg13g2_decap_8 FILLER_33_1303 ();
 sg13g2_decap_4 FILLER_33_1310 ();
 sg13g2_fill_1 FILLER_33_1314 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_27 ();
 sg13g2_fill_1 FILLER_34_29 ();
 sg13g2_fill_2 FILLER_34_44 ();
 sg13g2_fill_1 FILLER_34_46 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_decap_4 FILLER_34_235 ();
 sg13g2_fill_2 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_fill_2 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_4 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_fill_2 FILLER_34_352 ();
 sg13g2_fill_2 FILLER_34_363 ();
 sg13g2_fill_1 FILLER_34_365 ();
 sg13g2_fill_2 FILLER_34_388 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_1 FILLER_34_451 ();
 sg13g2_fill_1 FILLER_34_475 ();
 sg13g2_fill_1 FILLER_34_486 ();
 sg13g2_fill_1 FILLER_34_495 ();
 sg13g2_fill_2 FILLER_34_506 ();
 sg13g2_fill_1 FILLER_34_508 ();
 sg13g2_decap_4 FILLER_34_523 ();
 sg13g2_fill_2 FILLER_34_548 ();
 sg13g2_fill_1 FILLER_34_550 ();
 sg13g2_decap_8 FILLER_34_557 ();
 sg13g2_fill_2 FILLER_34_564 ();
 sg13g2_fill_1 FILLER_34_589 ();
 sg13g2_fill_2 FILLER_34_616 ();
 sg13g2_fill_1 FILLER_34_645 ();
 sg13g2_fill_1 FILLER_34_651 ();
 sg13g2_decap_4 FILLER_34_658 ();
 sg13g2_fill_2 FILLER_34_662 ();
 sg13g2_fill_2 FILLER_34_676 ();
 sg13g2_fill_2 FILLER_34_696 ();
 sg13g2_decap_8 FILLER_34_705 ();
 sg13g2_fill_2 FILLER_34_712 ();
 sg13g2_fill_1 FILLER_34_749 ();
 sg13g2_decap_4 FILLER_34_766 ();
 sg13g2_fill_2 FILLER_34_776 ();
 sg13g2_fill_1 FILLER_34_786 ();
 sg13g2_fill_1 FILLER_34_792 ();
 sg13g2_fill_1 FILLER_34_798 ();
 sg13g2_fill_1 FILLER_34_816 ();
 sg13g2_fill_2 FILLER_34_831 ();
 sg13g2_fill_1 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_decap_8 FILLER_34_860 ();
 sg13g2_fill_2 FILLER_34_867 ();
 sg13g2_fill_1 FILLER_34_869 ();
 sg13g2_fill_1 FILLER_34_874 ();
 sg13g2_fill_2 FILLER_34_905 ();
 sg13g2_fill_1 FILLER_34_907 ();
 sg13g2_fill_1 FILLER_34_960 ();
 sg13g2_fill_2 FILLER_34_974 ();
 sg13g2_fill_1 FILLER_34_981 ();
 sg13g2_fill_2 FILLER_34_1013 ();
 sg13g2_decap_8 FILLER_34_1136 ();
 sg13g2_decap_8 FILLER_34_1143 ();
 sg13g2_decap_8 FILLER_34_1150 ();
 sg13g2_decap_8 FILLER_34_1157 ();
 sg13g2_decap_8 FILLER_34_1164 ();
 sg13g2_decap_8 FILLER_34_1171 ();
 sg13g2_decap_8 FILLER_34_1178 ();
 sg13g2_decap_8 FILLER_34_1185 ();
 sg13g2_decap_8 FILLER_34_1192 ();
 sg13g2_decap_8 FILLER_34_1199 ();
 sg13g2_decap_8 FILLER_34_1206 ();
 sg13g2_decap_8 FILLER_34_1213 ();
 sg13g2_decap_8 FILLER_34_1220 ();
 sg13g2_decap_8 FILLER_34_1227 ();
 sg13g2_decap_8 FILLER_34_1234 ();
 sg13g2_decap_8 FILLER_34_1241 ();
 sg13g2_decap_8 FILLER_34_1248 ();
 sg13g2_decap_8 FILLER_34_1255 ();
 sg13g2_decap_8 FILLER_34_1262 ();
 sg13g2_decap_8 FILLER_34_1269 ();
 sg13g2_decap_8 FILLER_34_1276 ();
 sg13g2_decap_8 FILLER_34_1283 ();
 sg13g2_decap_8 FILLER_34_1290 ();
 sg13g2_decap_8 FILLER_34_1297 ();
 sg13g2_decap_8 FILLER_34_1304 ();
 sg13g2_decap_4 FILLER_34_1311 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_32 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_fill_2 FILLER_35_92 ();
 sg13g2_fill_2 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_109 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_decap_4 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_141 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_2 FILLER_35_252 ();
 sg13g2_decap_4 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_fill_1 FILLER_35_311 ();
 sg13g2_decap_8 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_339 ();
 sg13g2_decap_8 FILLER_35_346 ();
 sg13g2_fill_1 FILLER_35_353 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_fill_2 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_2 FILLER_35_413 ();
 sg13g2_fill_1 FILLER_35_415 ();
 sg13g2_fill_2 FILLER_35_450 ();
 sg13g2_decap_8 FILLER_35_464 ();
 sg13g2_fill_1 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_487 ();
 sg13g2_fill_2 FILLER_35_494 ();
 sg13g2_fill_1 FILLER_35_496 ();
 sg13g2_fill_2 FILLER_35_502 ();
 sg13g2_fill_1 FILLER_35_554 ();
 sg13g2_decap_8 FILLER_35_579 ();
 sg13g2_fill_1 FILLER_35_586 ();
 sg13g2_fill_1 FILLER_35_605 ();
 sg13g2_decap_4 FILLER_35_612 ();
 sg13g2_fill_1 FILLER_35_624 ();
 sg13g2_fill_2 FILLER_35_663 ();
 sg13g2_fill_1 FILLER_35_665 ();
 sg13g2_fill_2 FILLER_35_671 ();
 sg13g2_fill_1 FILLER_35_678 ();
 sg13g2_decap_4 FILLER_35_687 ();
 sg13g2_fill_1 FILLER_35_691 ();
 sg13g2_decap_8 FILLER_35_718 ();
 sg13g2_fill_2 FILLER_35_725 ();
 sg13g2_decap_8 FILLER_35_731 ();
 sg13g2_decap_8 FILLER_35_738 ();
 sg13g2_decap_4 FILLER_35_745 ();
 sg13g2_decap_8 FILLER_35_753 ();
 sg13g2_decap_8 FILLER_35_760 ();
 sg13g2_fill_1 FILLER_35_767 ();
 sg13g2_fill_2 FILLER_35_781 ();
 sg13g2_fill_1 FILLER_35_819 ();
 sg13g2_fill_2 FILLER_35_835 ();
 sg13g2_fill_1 FILLER_35_837 ();
 sg13g2_fill_1 FILLER_35_916 ();
 sg13g2_fill_1 FILLER_35_964 ();
 sg13g2_fill_2 FILLER_35_999 ();
 sg13g2_fill_1 FILLER_35_1001 ();
 sg13g2_fill_1 FILLER_35_1028 ();
 sg13g2_fill_1 FILLER_35_1080 ();
 sg13g2_fill_2 FILLER_35_1094 ();
 sg13g2_decap_8 FILLER_35_1148 ();
 sg13g2_decap_8 FILLER_35_1155 ();
 sg13g2_decap_8 FILLER_35_1162 ();
 sg13g2_decap_8 FILLER_35_1169 ();
 sg13g2_decap_8 FILLER_35_1176 ();
 sg13g2_decap_8 FILLER_35_1183 ();
 sg13g2_decap_8 FILLER_35_1190 ();
 sg13g2_decap_8 FILLER_35_1197 ();
 sg13g2_decap_8 FILLER_35_1204 ();
 sg13g2_decap_8 FILLER_35_1211 ();
 sg13g2_decap_8 FILLER_35_1218 ();
 sg13g2_decap_8 FILLER_35_1225 ();
 sg13g2_decap_8 FILLER_35_1232 ();
 sg13g2_decap_8 FILLER_35_1239 ();
 sg13g2_decap_8 FILLER_35_1246 ();
 sg13g2_decap_8 FILLER_35_1253 ();
 sg13g2_decap_8 FILLER_35_1260 ();
 sg13g2_decap_8 FILLER_35_1267 ();
 sg13g2_decap_8 FILLER_35_1274 ();
 sg13g2_decap_8 FILLER_35_1281 ();
 sg13g2_decap_8 FILLER_35_1288 ();
 sg13g2_decap_8 FILLER_35_1295 ();
 sg13g2_decap_8 FILLER_35_1302 ();
 sg13g2_decap_4 FILLER_35_1309 ();
 sg13g2_fill_2 FILLER_35_1313 ();
 sg13g2_fill_2 FILLER_36_45 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_decap_4 FILLER_36_120 ();
 sg13g2_decap_8 FILLER_36_128 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_decap_4 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_decap_8 FILLER_36_265 ();
 sg13g2_fill_1 FILLER_36_272 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_327 ();
 sg13g2_decap_4 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_378 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_392 ();
 sg13g2_decap_4 FILLER_36_412 ();
 sg13g2_fill_1 FILLER_36_422 ();
 sg13g2_fill_1 FILLER_36_428 ();
 sg13g2_fill_2 FILLER_36_434 ();
 sg13g2_fill_1 FILLER_36_436 ();
 sg13g2_decap_4 FILLER_36_441 ();
 sg13g2_fill_1 FILLER_36_445 ();
 sg13g2_fill_1 FILLER_36_463 ();
 sg13g2_decap_8 FILLER_36_472 ();
 sg13g2_fill_2 FILLER_36_479 ();
 sg13g2_fill_1 FILLER_36_481 ();
 sg13g2_decap_4 FILLER_36_495 ();
 sg13g2_fill_2 FILLER_36_499 ();
 sg13g2_decap_4 FILLER_36_514 ();
 sg13g2_fill_2 FILLER_36_518 ();
 sg13g2_fill_2 FILLER_36_554 ();
 sg13g2_fill_1 FILLER_36_556 ();
 sg13g2_decap_8 FILLER_36_573 ();
 sg13g2_decap_4 FILLER_36_580 ();
 sg13g2_fill_2 FILLER_36_584 ();
 sg13g2_decap_8 FILLER_36_612 ();
 sg13g2_decap_8 FILLER_36_619 ();
 sg13g2_decap_8 FILLER_36_626 ();
 sg13g2_fill_1 FILLER_36_633 ();
 sg13g2_decap_4 FILLER_36_699 ();
 sg13g2_fill_1 FILLER_36_703 ();
 sg13g2_fill_1 FILLER_36_715 ();
 sg13g2_fill_1 FILLER_36_787 ();
 sg13g2_fill_2 FILLER_36_854 ();
 sg13g2_fill_2 FILLER_36_888 ();
 sg13g2_fill_1 FILLER_36_899 ();
 sg13g2_fill_2 FILLER_36_914 ();
 sg13g2_fill_1 FILLER_36_916 ();
 sg13g2_fill_2 FILLER_36_995 ();
 sg13g2_fill_1 FILLER_36_997 ();
 sg13g2_fill_1 FILLER_36_1121 ();
 sg13g2_decap_8 FILLER_36_1135 ();
 sg13g2_decap_8 FILLER_36_1142 ();
 sg13g2_decap_8 FILLER_36_1149 ();
 sg13g2_decap_8 FILLER_36_1156 ();
 sg13g2_decap_8 FILLER_36_1163 ();
 sg13g2_decap_8 FILLER_36_1170 ();
 sg13g2_decap_8 FILLER_36_1177 ();
 sg13g2_decap_8 FILLER_36_1184 ();
 sg13g2_decap_8 FILLER_36_1191 ();
 sg13g2_decap_8 FILLER_36_1198 ();
 sg13g2_decap_8 FILLER_36_1205 ();
 sg13g2_decap_8 FILLER_36_1212 ();
 sg13g2_decap_8 FILLER_36_1219 ();
 sg13g2_decap_8 FILLER_36_1226 ();
 sg13g2_decap_8 FILLER_36_1233 ();
 sg13g2_decap_8 FILLER_36_1240 ();
 sg13g2_decap_8 FILLER_36_1247 ();
 sg13g2_decap_8 FILLER_36_1254 ();
 sg13g2_decap_8 FILLER_36_1261 ();
 sg13g2_decap_8 FILLER_36_1268 ();
 sg13g2_decap_8 FILLER_36_1275 ();
 sg13g2_decap_8 FILLER_36_1282 ();
 sg13g2_decap_8 FILLER_36_1289 ();
 sg13g2_decap_8 FILLER_36_1296 ();
 sg13g2_decap_8 FILLER_36_1303 ();
 sg13g2_decap_4 FILLER_36_1310 ();
 sg13g2_fill_1 FILLER_36_1314 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_25 ();
 sg13g2_fill_1 FILLER_37_40 ();
 sg13g2_fill_2 FILLER_37_51 ();
 sg13g2_fill_1 FILLER_37_53 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_2 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_139 ();
 sg13g2_fill_2 FILLER_37_156 ();
 sg13g2_fill_2 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_204 ();
 sg13g2_fill_2 FILLER_37_215 ();
 sg13g2_fill_2 FILLER_37_225 ();
 sg13g2_decap_4 FILLER_37_234 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_2 FILLER_37_277 ();
 sg13g2_decap_8 FILLER_37_307 ();
 sg13g2_decap_4 FILLER_37_314 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_decap_4 FILLER_37_325 ();
 sg13g2_fill_1 FILLER_37_329 ();
 sg13g2_fill_1 FILLER_37_336 ();
 sg13g2_fill_1 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_fill_2 FILLER_37_386 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_fill_2 FILLER_37_434 ();
 sg13g2_decap_4 FILLER_37_460 ();
 sg13g2_fill_2 FILLER_37_464 ();
 sg13g2_fill_2 FILLER_37_484 ();
 sg13g2_decap_4 FILLER_37_555 ();
 sg13g2_fill_2 FILLER_37_559 ();
 sg13g2_decap_8 FILLER_37_580 ();
 sg13g2_decap_8 FILLER_37_587 ();
 sg13g2_fill_1 FILLER_37_594 ();
 sg13g2_decap_8 FILLER_37_599 ();
 sg13g2_fill_1 FILLER_37_606 ();
 sg13g2_decap_4 FILLER_37_631 ();
 sg13g2_fill_2 FILLER_37_660 ();
 sg13g2_fill_1 FILLER_37_662 ();
 sg13g2_decap_4 FILLER_37_677 ();
 sg13g2_fill_1 FILLER_37_681 ();
 sg13g2_decap_4 FILLER_37_688 ();
 sg13g2_fill_1 FILLER_37_692 ();
 sg13g2_decap_8 FILLER_37_712 ();
 sg13g2_decap_4 FILLER_37_719 ();
 sg13g2_fill_1 FILLER_37_723 ();
 sg13g2_fill_2 FILLER_37_728 ();
 sg13g2_fill_1 FILLER_37_730 ();
 sg13g2_fill_1 FILLER_37_736 ();
 sg13g2_fill_1 FILLER_37_750 ();
 sg13g2_fill_2 FILLER_37_777 ();
 sg13g2_decap_4 FILLER_37_805 ();
 sg13g2_fill_1 FILLER_37_809 ();
 sg13g2_fill_1 FILLER_37_836 ();
 sg13g2_fill_2 FILLER_37_889 ();
 sg13g2_fill_2 FILLER_37_947 ();
 sg13g2_fill_1 FILLER_37_949 ();
 sg13g2_fill_1 FILLER_37_985 ();
 sg13g2_fill_2 FILLER_37_1030 ();
 sg13g2_fill_1 FILLER_37_1032 ();
 sg13g2_fill_2 FILLER_37_1038 ();
 sg13g2_fill_1 FILLER_37_1040 ();
 sg13g2_decap_4 FILLER_37_1062 ();
 sg13g2_fill_1 FILLER_37_1066 ();
 sg13g2_decap_4 FILLER_37_1080 ();
 sg13g2_fill_1 FILLER_37_1084 ();
 sg13g2_fill_2 FILLER_37_1111 ();
 sg13g2_decap_8 FILLER_37_1117 ();
 sg13g2_decap_8 FILLER_37_1124 ();
 sg13g2_decap_8 FILLER_37_1131 ();
 sg13g2_decap_8 FILLER_37_1138 ();
 sg13g2_decap_8 FILLER_37_1145 ();
 sg13g2_decap_8 FILLER_37_1152 ();
 sg13g2_decap_8 FILLER_37_1159 ();
 sg13g2_decap_8 FILLER_37_1166 ();
 sg13g2_decap_8 FILLER_37_1173 ();
 sg13g2_decap_8 FILLER_37_1180 ();
 sg13g2_decap_8 FILLER_37_1187 ();
 sg13g2_decap_8 FILLER_37_1194 ();
 sg13g2_decap_8 FILLER_37_1201 ();
 sg13g2_decap_8 FILLER_37_1208 ();
 sg13g2_decap_8 FILLER_37_1215 ();
 sg13g2_decap_8 FILLER_37_1222 ();
 sg13g2_decap_8 FILLER_37_1229 ();
 sg13g2_decap_8 FILLER_37_1236 ();
 sg13g2_decap_8 FILLER_37_1243 ();
 sg13g2_decap_8 FILLER_37_1250 ();
 sg13g2_decap_8 FILLER_37_1257 ();
 sg13g2_decap_8 FILLER_37_1264 ();
 sg13g2_decap_8 FILLER_37_1271 ();
 sg13g2_decap_8 FILLER_37_1278 ();
 sg13g2_decap_8 FILLER_37_1285 ();
 sg13g2_decap_8 FILLER_37_1292 ();
 sg13g2_decap_8 FILLER_37_1299 ();
 sg13g2_decap_8 FILLER_37_1306 ();
 sg13g2_fill_2 FILLER_37_1313 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_48 ();
 sg13g2_fill_2 FILLER_38_81 ();
 sg13g2_decap_8 FILLER_38_88 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_162 ();
 sg13g2_fill_2 FILLER_38_178 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_fill_2 FILLER_38_227 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_decap_4 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_251 ();
 sg13g2_decap_4 FILLER_38_264 ();
 sg13g2_decap_4 FILLER_38_342 ();
 sg13g2_fill_2 FILLER_38_361 ();
 sg13g2_fill_1 FILLER_38_363 ();
 sg13g2_fill_2 FILLER_38_369 ();
 sg13g2_fill_2 FILLER_38_400 ();
 sg13g2_fill_1 FILLER_38_402 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_fill_1 FILLER_38_409 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_fill_2 FILLER_38_441 ();
 sg13g2_fill_1 FILLER_38_443 ();
 sg13g2_decap_4 FILLER_38_453 ();
 sg13g2_fill_1 FILLER_38_457 ();
 sg13g2_decap_8 FILLER_38_465 ();
 sg13g2_fill_2 FILLER_38_483 ();
 sg13g2_decap_4 FILLER_38_495 ();
 sg13g2_fill_2 FILLER_38_499 ();
 sg13g2_decap_4 FILLER_38_505 ();
 sg13g2_fill_2 FILLER_38_514 ();
 sg13g2_fill_2 FILLER_38_526 ();
 sg13g2_fill_1 FILLER_38_545 ();
 sg13g2_fill_1 FILLER_38_560 ();
 sg13g2_decap_4 FILLER_38_615 ();
 sg13g2_fill_2 FILLER_38_657 ();
 sg13g2_fill_1 FILLER_38_659 ();
 sg13g2_fill_1 FILLER_38_672 ();
 sg13g2_decap_4 FILLER_38_677 ();
 sg13g2_fill_1 FILLER_38_681 ();
 sg13g2_decap_4 FILLER_38_691 ();
 sg13g2_fill_2 FILLER_38_710 ();
 sg13g2_fill_1 FILLER_38_712 ();
 sg13g2_decap_4 FILLER_38_779 ();
 sg13g2_decap_8 FILLER_38_787 ();
 sg13g2_decap_4 FILLER_38_794 ();
 sg13g2_decap_8 FILLER_38_807 ();
 sg13g2_fill_1 FILLER_38_814 ();
 sg13g2_fill_2 FILLER_38_864 ();
 sg13g2_fill_1 FILLER_38_896 ();
 sg13g2_fill_2 FILLER_38_953 ();
 sg13g2_fill_1 FILLER_38_955 ();
 sg13g2_fill_2 FILLER_38_1013 ();
 sg13g2_fill_2 FILLER_38_1093 ();
 sg13g2_fill_1 FILLER_38_1095 ();
 sg13g2_fill_1 FILLER_38_1100 ();
 sg13g2_decap_8 FILLER_38_1110 ();
 sg13g2_decap_8 FILLER_38_1117 ();
 sg13g2_decap_8 FILLER_38_1124 ();
 sg13g2_decap_8 FILLER_38_1131 ();
 sg13g2_decap_8 FILLER_38_1138 ();
 sg13g2_decap_8 FILLER_38_1145 ();
 sg13g2_decap_8 FILLER_38_1152 ();
 sg13g2_decap_8 FILLER_38_1159 ();
 sg13g2_decap_8 FILLER_38_1166 ();
 sg13g2_decap_8 FILLER_38_1173 ();
 sg13g2_decap_8 FILLER_38_1180 ();
 sg13g2_decap_8 FILLER_38_1187 ();
 sg13g2_decap_8 FILLER_38_1194 ();
 sg13g2_decap_8 FILLER_38_1201 ();
 sg13g2_decap_8 FILLER_38_1208 ();
 sg13g2_decap_8 FILLER_38_1215 ();
 sg13g2_decap_8 FILLER_38_1222 ();
 sg13g2_decap_8 FILLER_38_1229 ();
 sg13g2_decap_8 FILLER_38_1236 ();
 sg13g2_decap_8 FILLER_38_1243 ();
 sg13g2_decap_8 FILLER_38_1250 ();
 sg13g2_decap_8 FILLER_38_1257 ();
 sg13g2_decap_8 FILLER_38_1264 ();
 sg13g2_decap_8 FILLER_38_1271 ();
 sg13g2_decap_8 FILLER_38_1278 ();
 sg13g2_decap_8 FILLER_38_1285 ();
 sg13g2_decap_8 FILLER_38_1292 ();
 sg13g2_decap_8 FILLER_38_1299 ();
 sg13g2_decap_8 FILLER_38_1306 ();
 sg13g2_fill_2 FILLER_38_1313 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_2 ();
 sg13g2_decap_4 FILLER_39_84 ();
 sg13g2_decap_4 FILLER_39_114 ();
 sg13g2_fill_1 FILLER_39_118 ();
 sg13g2_decap_4 FILLER_39_143 ();
 sg13g2_fill_1 FILLER_39_151 ();
 sg13g2_fill_2 FILLER_39_190 ();
 sg13g2_decap_4 FILLER_39_235 ();
 sg13g2_fill_1 FILLER_39_239 ();
 sg13g2_decap_4 FILLER_39_256 ();
 sg13g2_decap_4 FILLER_39_306 ();
 sg13g2_fill_1 FILLER_39_310 ();
 sg13g2_fill_2 FILLER_39_331 ();
 sg13g2_fill_1 FILLER_39_333 ();
 sg13g2_fill_2 FILLER_39_348 ();
 sg13g2_fill_1 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_360 ();
 sg13g2_fill_2 FILLER_39_367 ();
 sg13g2_fill_1 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_378 ();
 sg13g2_fill_1 FILLER_39_419 ();
 sg13g2_decap_8 FILLER_39_424 ();
 sg13g2_fill_2 FILLER_39_440 ();
 sg13g2_fill_1 FILLER_39_442 ();
 sg13g2_decap_8 FILLER_39_459 ();
 sg13g2_fill_1 FILLER_39_466 ();
 sg13g2_fill_2 FILLER_39_483 ();
 sg13g2_fill_2 FILLER_39_525 ();
 sg13g2_fill_1 FILLER_39_535 ();
 sg13g2_fill_2 FILLER_39_541 ();
 sg13g2_fill_1 FILLER_39_543 ();
 sg13g2_fill_1 FILLER_39_559 ();
 sg13g2_fill_1 FILLER_39_585 ();
 sg13g2_fill_1 FILLER_39_595 ();
 sg13g2_fill_2 FILLER_39_621 ();
 sg13g2_fill_1 FILLER_39_623 ();
 sg13g2_decap_4 FILLER_39_641 ();
 sg13g2_fill_1 FILLER_39_645 ();
 sg13g2_decap_4 FILLER_39_661 ();
 sg13g2_fill_2 FILLER_39_665 ();
 sg13g2_fill_2 FILLER_39_677 ();
 sg13g2_fill_2 FILLER_39_690 ();
 sg13g2_fill_2 FILLER_39_697 ();
 sg13g2_fill_1 FILLER_39_704 ();
 sg13g2_decap_4 FILLER_39_718 ();
 sg13g2_fill_1 FILLER_39_722 ();
 sg13g2_fill_2 FILLER_39_746 ();
 sg13g2_decap_8 FILLER_39_755 ();
 sg13g2_decap_4 FILLER_39_766 ();
 sg13g2_fill_2 FILLER_39_770 ();
 sg13g2_decap_8 FILLER_39_823 ();
 sg13g2_fill_1 FILLER_39_843 ();
 sg13g2_fill_2 FILLER_39_857 ();
 sg13g2_fill_1 FILLER_39_859 ();
 sg13g2_fill_2 FILLER_39_922 ();
 sg13g2_fill_1 FILLER_39_924 ();
 sg13g2_fill_2 FILLER_39_957 ();
 sg13g2_fill_2 FILLER_39_1024 ();
 sg13g2_fill_1 FILLER_39_1026 ();
 sg13g2_decap_8 FILLER_39_1053 ();
 sg13g2_decap_8 FILLER_39_1060 ();
 sg13g2_decap_8 FILLER_39_1067 ();
 sg13g2_decap_8 FILLER_39_1074 ();
 sg13g2_decap_8 FILLER_39_1081 ();
 sg13g2_decap_8 FILLER_39_1088 ();
 sg13g2_decap_8 FILLER_39_1095 ();
 sg13g2_decap_8 FILLER_39_1102 ();
 sg13g2_decap_8 FILLER_39_1109 ();
 sg13g2_decap_8 FILLER_39_1116 ();
 sg13g2_decap_8 FILLER_39_1123 ();
 sg13g2_decap_8 FILLER_39_1130 ();
 sg13g2_decap_8 FILLER_39_1137 ();
 sg13g2_decap_8 FILLER_39_1144 ();
 sg13g2_decap_8 FILLER_39_1151 ();
 sg13g2_decap_8 FILLER_39_1158 ();
 sg13g2_decap_8 FILLER_39_1165 ();
 sg13g2_decap_8 FILLER_39_1172 ();
 sg13g2_decap_8 FILLER_39_1179 ();
 sg13g2_decap_8 FILLER_39_1186 ();
 sg13g2_decap_8 FILLER_39_1193 ();
 sg13g2_decap_8 FILLER_39_1200 ();
 sg13g2_decap_8 FILLER_39_1207 ();
 sg13g2_decap_8 FILLER_39_1214 ();
 sg13g2_decap_8 FILLER_39_1221 ();
 sg13g2_decap_8 FILLER_39_1228 ();
 sg13g2_decap_8 FILLER_39_1235 ();
 sg13g2_decap_8 FILLER_39_1242 ();
 sg13g2_decap_8 FILLER_39_1249 ();
 sg13g2_decap_8 FILLER_39_1256 ();
 sg13g2_decap_8 FILLER_39_1263 ();
 sg13g2_decap_8 FILLER_39_1270 ();
 sg13g2_decap_8 FILLER_39_1277 ();
 sg13g2_decap_8 FILLER_39_1284 ();
 sg13g2_decap_8 FILLER_39_1291 ();
 sg13g2_decap_8 FILLER_39_1298 ();
 sg13g2_decap_8 FILLER_39_1305 ();
 sg13g2_fill_2 FILLER_39_1312 ();
 sg13g2_fill_1 FILLER_39_1314 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_1 FILLER_40_24 ();
 sg13g2_decap_4 FILLER_40_75 ();
 sg13g2_decap_8 FILLER_40_94 ();
 sg13g2_fill_2 FILLER_40_101 ();
 sg13g2_fill_1 FILLER_40_108 ();
 sg13g2_decap_8 FILLER_40_115 ();
 sg13g2_decap_4 FILLER_40_122 ();
 sg13g2_fill_1 FILLER_40_126 ();
 sg13g2_decap_4 FILLER_40_143 ();
 sg13g2_fill_1 FILLER_40_176 ();
 sg13g2_fill_2 FILLER_40_216 ();
 sg13g2_decap_4 FILLER_40_223 ();
 sg13g2_decap_8 FILLER_40_240 ();
 sg13g2_fill_1 FILLER_40_247 ();
 sg13g2_fill_1 FILLER_40_261 ();
 sg13g2_decap_8 FILLER_40_267 ();
 sg13g2_decap_8 FILLER_40_278 ();
 sg13g2_decap_8 FILLER_40_285 ();
 sg13g2_fill_2 FILLER_40_298 ();
 sg13g2_fill_1 FILLER_40_300 ();
 sg13g2_fill_1 FILLER_40_333 ();
 sg13g2_decap_8 FILLER_40_373 ();
 sg13g2_decap_8 FILLER_40_380 ();
 sg13g2_decap_4 FILLER_40_387 ();
 sg13g2_fill_1 FILLER_40_391 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_40_435 ();
 sg13g2_decap_4 FILLER_40_441 ();
 sg13g2_fill_1 FILLER_40_445 ();
 sg13g2_fill_2 FILLER_40_456 ();
 sg13g2_fill_1 FILLER_40_458 ();
 sg13g2_decap_8 FILLER_40_464 ();
 sg13g2_fill_1 FILLER_40_471 ();
 sg13g2_decap_8 FILLER_40_484 ();
 sg13g2_decap_8 FILLER_40_496 ();
 sg13g2_fill_2 FILLER_40_503 ();
 sg13g2_decap_8 FILLER_40_509 ();
 sg13g2_fill_2 FILLER_40_516 ();
 sg13g2_fill_1 FILLER_40_518 ();
 sg13g2_decap_4 FILLER_40_534 ();
 sg13g2_fill_1 FILLER_40_544 ();
 sg13g2_fill_1 FILLER_40_554 ();
 sg13g2_fill_1 FILLER_40_566 ();
 sg13g2_fill_2 FILLER_40_633 ();
 sg13g2_fill_2 FILLER_40_640 ();
 sg13g2_fill_1 FILLER_40_655 ();
 sg13g2_fill_2 FILLER_40_665 ();
 sg13g2_fill_1 FILLER_40_691 ();
 sg13g2_fill_1 FILLER_40_768 ();
 sg13g2_fill_1 FILLER_40_886 ();
 sg13g2_fill_2 FILLER_40_1004 ();
 sg13g2_decap_4 FILLER_40_1032 ();
 sg13g2_fill_1 FILLER_40_1036 ();
 sg13g2_decap_8 FILLER_40_1050 ();
 sg13g2_decap_8 FILLER_40_1057 ();
 sg13g2_decap_8 FILLER_40_1064 ();
 sg13g2_decap_8 FILLER_40_1071 ();
 sg13g2_decap_8 FILLER_40_1078 ();
 sg13g2_decap_8 FILLER_40_1085 ();
 sg13g2_decap_8 FILLER_40_1092 ();
 sg13g2_decap_8 FILLER_40_1099 ();
 sg13g2_decap_8 FILLER_40_1106 ();
 sg13g2_decap_8 FILLER_40_1113 ();
 sg13g2_decap_8 FILLER_40_1120 ();
 sg13g2_decap_8 FILLER_40_1127 ();
 sg13g2_decap_8 FILLER_40_1134 ();
 sg13g2_decap_8 FILLER_40_1141 ();
 sg13g2_decap_8 FILLER_40_1148 ();
 sg13g2_decap_8 FILLER_40_1155 ();
 sg13g2_decap_8 FILLER_40_1162 ();
 sg13g2_decap_8 FILLER_40_1169 ();
 sg13g2_decap_8 FILLER_40_1176 ();
 sg13g2_decap_8 FILLER_40_1183 ();
 sg13g2_decap_8 FILLER_40_1190 ();
 sg13g2_decap_8 FILLER_40_1197 ();
 sg13g2_decap_8 FILLER_40_1204 ();
 sg13g2_decap_8 FILLER_40_1211 ();
 sg13g2_decap_8 FILLER_40_1218 ();
 sg13g2_decap_8 FILLER_40_1225 ();
 sg13g2_decap_8 FILLER_40_1232 ();
 sg13g2_decap_8 FILLER_40_1239 ();
 sg13g2_decap_8 FILLER_40_1246 ();
 sg13g2_decap_8 FILLER_40_1253 ();
 sg13g2_decap_8 FILLER_40_1260 ();
 sg13g2_decap_8 FILLER_40_1267 ();
 sg13g2_decap_8 FILLER_40_1274 ();
 sg13g2_decap_8 FILLER_40_1281 ();
 sg13g2_decap_8 FILLER_40_1288 ();
 sg13g2_decap_8 FILLER_40_1295 ();
 sg13g2_decap_8 FILLER_40_1302 ();
 sg13g2_decap_4 FILLER_40_1309 ();
 sg13g2_fill_2 FILLER_40_1313 ();
 sg13g2_fill_2 FILLER_41_26 ();
 sg13g2_fill_1 FILLER_41_28 ();
 sg13g2_fill_2 FILLER_41_54 ();
 sg13g2_fill_1 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_66 ();
 sg13g2_fill_1 FILLER_41_78 ();
 sg13g2_fill_1 FILLER_41_82 ();
 sg13g2_fill_1 FILLER_41_93 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_fill_1 FILLER_41_175 ();
 sg13g2_decap_4 FILLER_41_195 ();
 sg13g2_fill_1 FILLER_41_199 ();
 sg13g2_decap_8 FILLER_41_214 ();
 sg13g2_fill_2 FILLER_41_221 ();
 sg13g2_fill_2 FILLER_41_252 ();
 sg13g2_fill_2 FILLER_41_300 ();
 sg13g2_fill_2 FILLER_41_311 ();
 sg13g2_decap_4 FILLER_41_367 ();
 sg13g2_decap_4 FILLER_41_376 ();
 sg13g2_decap_8 FILLER_41_384 ();
 sg13g2_fill_1 FILLER_41_391 ();
 sg13g2_fill_1 FILLER_41_437 ();
 sg13g2_fill_1 FILLER_41_443 ();
 sg13g2_fill_1 FILLER_41_448 ();
 sg13g2_decap_4 FILLER_41_463 ();
 sg13g2_fill_2 FILLER_41_467 ();
 sg13g2_fill_2 FILLER_41_474 ();
 sg13g2_fill_2 FILLER_41_533 ();
 sg13g2_fill_1 FILLER_41_535 ();
 sg13g2_decap_4 FILLER_41_546 ();
 sg13g2_fill_2 FILLER_41_584 ();
 sg13g2_fill_1 FILLER_41_586 ();
 sg13g2_decap_8 FILLER_41_591 ();
 sg13g2_fill_2 FILLER_41_602 ();
 sg13g2_fill_1 FILLER_41_604 ();
 sg13g2_fill_2 FILLER_41_628 ();
 sg13g2_fill_1 FILLER_41_630 ();
 sg13g2_fill_1 FILLER_41_636 ();
 sg13g2_fill_2 FILLER_41_642 ();
 sg13g2_fill_1 FILLER_41_649 ();
 sg13g2_fill_2 FILLER_41_661 ();
 sg13g2_fill_2 FILLER_41_689 ();
 sg13g2_decap_4 FILLER_41_717 ();
 sg13g2_decap_8 FILLER_41_729 ();
 sg13g2_decap_4 FILLER_41_736 ();
 sg13g2_fill_1 FILLER_41_740 ();
 sg13g2_fill_2 FILLER_41_750 ();
 sg13g2_decap_4 FILLER_41_756 ();
 sg13g2_fill_1 FILLER_41_799 ();
 sg13g2_decap_8 FILLER_41_810 ();
 sg13g2_fill_1 FILLER_41_821 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_fill_2 FILLER_41_849 ();
 sg13g2_fill_1 FILLER_41_851 ();
 sg13g2_fill_1 FILLER_41_864 ();
 sg13g2_fill_2 FILLER_41_910 ();
 sg13g2_fill_1 FILLER_41_912 ();
 sg13g2_fill_2 FILLER_41_947 ();
 sg13g2_fill_2 FILLER_41_962 ();
 sg13g2_fill_1 FILLER_41_964 ();
 sg13g2_fill_1 FILLER_41_978 ();
 sg13g2_decap_8 FILLER_41_1026 ();
 sg13g2_decap_8 FILLER_41_1033 ();
 sg13g2_decap_8 FILLER_41_1040 ();
 sg13g2_decap_8 FILLER_41_1047 ();
 sg13g2_decap_8 FILLER_41_1054 ();
 sg13g2_decap_8 FILLER_41_1061 ();
 sg13g2_decap_8 FILLER_41_1068 ();
 sg13g2_decap_8 FILLER_41_1075 ();
 sg13g2_decap_8 FILLER_41_1082 ();
 sg13g2_decap_8 FILLER_41_1089 ();
 sg13g2_decap_8 FILLER_41_1096 ();
 sg13g2_decap_8 FILLER_41_1103 ();
 sg13g2_decap_8 FILLER_41_1110 ();
 sg13g2_decap_8 FILLER_41_1117 ();
 sg13g2_decap_8 FILLER_41_1124 ();
 sg13g2_decap_8 FILLER_41_1131 ();
 sg13g2_decap_8 FILLER_41_1138 ();
 sg13g2_decap_8 FILLER_41_1145 ();
 sg13g2_decap_8 FILLER_41_1152 ();
 sg13g2_decap_8 FILLER_41_1159 ();
 sg13g2_decap_8 FILLER_41_1166 ();
 sg13g2_decap_8 FILLER_41_1173 ();
 sg13g2_decap_8 FILLER_41_1180 ();
 sg13g2_decap_8 FILLER_41_1187 ();
 sg13g2_decap_8 FILLER_41_1194 ();
 sg13g2_decap_8 FILLER_41_1201 ();
 sg13g2_decap_8 FILLER_41_1208 ();
 sg13g2_decap_8 FILLER_41_1215 ();
 sg13g2_decap_8 FILLER_41_1222 ();
 sg13g2_decap_8 FILLER_41_1229 ();
 sg13g2_decap_8 FILLER_41_1236 ();
 sg13g2_decap_8 FILLER_41_1243 ();
 sg13g2_decap_8 FILLER_41_1250 ();
 sg13g2_decap_8 FILLER_41_1257 ();
 sg13g2_decap_8 FILLER_41_1264 ();
 sg13g2_decap_8 FILLER_41_1271 ();
 sg13g2_decap_8 FILLER_41_1278 ();
 sg13g2_decap_8 FILLER_41_1285 ();
 sg13g2_decap_8 FILLER_41_1292 ();
 sg13g2_decap_8 FILLER_41_1299 ();
 sg13g2_decap_8 FILLER_41_1306 ();
 sg13g2_fill_2 FILLER_41_1313 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_75 ();
 sg13g2_fill_2 FILLER_42_82 ();
 sg13g2_decap_4 FILLER_42_95 ();
 sg13g2_decap_8 FILLER_42_104 ();
 sg13g2_decap_4 FILLER_42_115 ();
 sg13g2_fill_1 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_4 FILLER_42_140 ();
 sg13g2_fill_2 FILLER_42_144 ();
 sg13g2_decap_8 FILLER_42_150 ();
 sg13g2_fill_2 FILLER_42_157 ();
 sg13g2_fill_2 FILLER_42_190 ();
 sg13g2_fill_1 FILLER_42_192 ();
 sg13g2_decap_8 FILLER_42_235 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_fill_2 FILLER_42_249 ();
 sg13g2_fill_1 FILLER_42_256 ();
 sg13g2_fill_2 FILLER_42_264 ();
 sg13g2_fill_2 FILLER_42_275 ();
 sg13g2_decap_8 FILLER_42_281 ();
 sg13g2_fill_2 FILLER_42_344 ();
 sg13g2_decap_4 FILLER_42_355 ();
 sg13g2_fill_1 FILLER_42_395 ();
 sg13g2_fill_2 FILLER_42_405 ();
 sg13g2_fill_1 FILLER_42_407 ();
 sg13g2_decap_4 FILLER_42_416 ();
 sg13g2_fill_1 FILLER_42_420 ();
 sg13g2_fill_1 FILLER_42_431 ();
 sg13g2_fill_2 FILLER_42_444 ();
 sg13g2_fill_2 FILLER_42_452 ();
 sg13g2_fill_1 FILLER_42_454 ();
 sg13g2_fill_2 FILLER_42_461 ();
 sg13g2_fill_1 FILLER_42_463 ();
 sg13g2_fill_1 FILLER_42_470 ();
 sg13g2_fill_2 FILLER_42_482 ();
 sg13g2_fill_2 FILLER_42_493 ();
 sg13g2_fill_1 FILLER_42_495 ();
 sg13g2_decap_4 FILLER_42_513 ();
 sg13g2_fill_2 FILLER_42_517 ();
 sg13g2_decap_4 FILLER_42_527 ();
 sg13g2_decap_8 FILLER_42_579 ();
 sg13g2_fill_1 FILLER_42_586 ();
 sg13g2_decap_4 FILLER_42_601 ();
 sg13g2_fill_1 FILLER_42_605 ();
 sg13g2_decap_8 FILLER_42_616 ();
 sg13g2_fill_1 FILLER_42_623 ();
 sg13g2_fill_2 FILLER_42_634 ();
 sg13g2_fill_2 FILLER_42_643 ();
 sg13g2_fill_1 FILLER_42_657 ();
 sg13g2_decap_8 FILLER_42_670 ();
 sg13g2_fill_1 FILLER_42_677 ();
 sg13g2_decap_4 FILLER_42_687 ();
 sg13g2_fill_1 FILLER_42_691 ();
 sg13g2_decap_8 FILLER_42_712 ();
 sg13g2_fill_2 FILLER_42_719 ();
 sg13g2_fill_2 FILLER_42_747 ();
 sg13g2_fill_1 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_754 ();
 sg13g2_decap_8 FILLER_42_761 ();
 sg13g2_fill_2 FILLER_42_768 ();
 sg13g2_fill_1 FILLER_42_770 ();
 sg13g2_fill_1 FILLER_42_811 ();
 sg13g2_fill_2 FILLER_42_838 ();
 sg13g2_fill_1 FILLER_42_840 ();
 sg13g2_fill_2 FILLER_42_897 ();
 sg13g2_fill_1 FILLER_42_925 ();
 sg13g2_fill_1 FILLER_42_952 ();
 sg13g2_fill_2 FILLER_42_1005 ();
 sg13g2_fill_1 FILLER_42_1011 ();
 sg13g2_decap_8 FILLER_42_1021 ();
 sg13g2_decap_8 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_42_1035 ();
 sg13g2_decap_8 FILLER_42_1042 ();
 sg13g2_decap_8 FILLER_42_1049 ();
 sg13g2_decap_8 FILLER_42_1056 ();
 sg13g2_decap_8 FILLER_42_1063 ();
 sg13g2_decap_8 FILLER_42_1070 ();
 sg13g2_decap_8 FILLER_42_1077 ();
 sg13g2_decap_8 FILLER_42_1084 ();
 sg13g2_decap_8 FILLER_42_1091 ();
 sg13g2_decap_8 FILLER_42_1098 ();
 sg13g2_decap_8 FILLER_42_1105 ();
 sg13g2_decap_8 FILLER_42_1112 ();
 sg13g2_decap_8 FILLER_42_1119 ();
 sg13g2_decap_8 FILLER_42_1126 ();
 sg13g2_decap_8 FILLER_42_1133 ();
 sg13g2_decap_8 FILLER_42_1140 ();
 sg13g2_decap_8 FILLER_42_1147 ();
 sg13g2_decap_8 FILLER_42_1154 ();
 sg13g2_decap_8 FILLER_42_1161 ();
 sg13g2_decap_8 FILLER_42_1168 ();
 sg13g2_decap_8 FILLER_42_1175 ();
 sg13g2_decap_8 FILLER_42_1182 ();
 sg13g2_decap_8 FILLER_42_1189 ();
 sg13g2_decap_8 FILLER_42_1196 ();
 sg13g2_decap_8 FILLER_42_1203 ();
 sg13g2_decap_8 FILLER_42_1210 ();
 sg13g2_decap_8 FILLER_42_1217 ();
 sg13g2_decap_8 FILLER_42_1224 ();
 sg13g2_decap_8 FILLER_42_1231 ();
 sg13g2_decap_8 FILLER_42_1238 ();
 sg13g2_decap_8 FILLER_42_1245 ();
 sg13g2_decap_8 FILLER_42_1252 ();
 sg13g2_decap_8 FILLER_42_1259 ();
 sg13g2_decap_8 FILLER_42_1266 ();
 sg13g2_decap_8 FILLER_42_1273 ();
 sg13g2_decap_8 FILLER_42_1280 ();
 sg13g2_decap_8 FILLER_42_1287 ();
 sg13g2_decap_8 FILLER_42_1294 ();
 sg13g2_decap_8 FILLER_42_1301 ();
 sg13g2_decap_8 FILLER_42_1308 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_24 ();
 sg13g2_fill_1 FILLER_43_35 ();
 sg13g2_fill_2 FILLER_43_44 ();
 sg13g2_fill_1 FILLER_43_46 ();
 sg13g2_fill_2 FILLER_43_86 ();
 sg13g2_fill_1 FILLER_43_88 ();
 sg13g2_fill_2 FILLER_43_109 ();
 sg13g2_fill_1 FILLER_43_111 ();
 sg13g2_fill_2 FILLER_43_186 ();
 sg13g2_fill_1 FILLER_43_188 ();
 sg13g2_decap_4 FILLER_43_236 ();
 sg13g2_fill_1 FILLER_43_240 ();
 sg13g2_fill_2 FILLER_43_267 ();
 sg13g2_fill_2 FILLER_43_283 ();
 sg13g2_fill_2 FILLER_43_297 ();
 sg13g2_decap_4 FILLER_43_303 ();
 sg13g2_decap_8 FILLER_43_319 ();
 sg13g2_fill_2 FILLER_43_326 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_fill_2 FILLER_43_343 ();
 sg13g2_decap_4 FILLER_43_367 ();
 sg13g2_decap_4 FILLER_43_376 ();
 sg13g2_fill_1 FILLER_43_380 ();
 sg13g2_fill_2 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_434 ();
 sg13g2_decap_4 FILLER_43_449 ();
 sg13g2_fill_2 FILLER_43_453 ();
 sg13g2_fill_2 FILLER_43_485 ();
 sg13g2_decap_8 FILLER_43_495 ();
 sg13g2_decap_4 FILLER_43_527 ();
 sg13g2_fill_1 FILLER_43_531 ();
 sg13g2_decap_8 FILLER_43_537 ();
 sg13g2_decap_4 FILLER_43_544 ();
 sg13g2_decap_8 FILLER_43_556 ();
 sg13g2_decap_4 FILLER_43_563 ();
 sg13g2_fill_1 FILLER_43_574 ();
 sg13g2_fill_2 FILLER_43_580 ();
 sg13g2_fill_2 FILLER_43_597 ();
 sg13g2_decap_4 FILLER_43_609 ();
 sg13g2_fill_1 FILLER_43_651 ();
 sg13g2_fill_1 FILLER_43_666 ();
 sg13g2_fill_1 FILLER_43_680 ();
 sg13g2_fill_1 FILLER_43_689 ();
 sg13g2_fill_2 FILLER_43_699 ();
 sg13g2_fill_1 FILLER_43_701 ();
 sg13g2_decap_8 FILLER_43_712 ();
 sg13g2_fill_2 FILLER_43_719 ();
 sg13g2_fill_1 FILLER_43_738 ();
 sg13g2_fill_2 FILLER_43_795 ();
 sg13g2_fill_1 FILLER_43_821 ();
 sg13g2_fill_2 FILLER_43_848 ();
 sg13g2_fill_2 FILLER_43_876 ();
 sg13g2_decap_8 FILLER_43_908 ();
 sg13g2_fill_2 FILLER_43_915 ();
 sg13g2_fill_1 FILLER_43_917 ();
 sg13g2_fill_1 FILLER_43_961 ();
 sg13g2_decap_8 FILLER_43_1040 ();
 sg13g2_decap_8 FILLER_43_1047 ();
 sg13g2_decap_8 FILLER_43_1054 ();
 sg13g2_decap_8 FILLER_43_1061 ();
 sg13g2_decap_8 FILLER_43_1068 ();
 sg13g2_decap_8 FILLER_43_1075 ();
 sg13g2_decap_8 FILLER_43_1082 ();
 sg13g2_decap_8 FILLER_43_1089 ();
 sg13g2_decap_8 FILLER_43_1096 ();
 sg13g2_decap_8 FILLER_43_1103 ();
 sg13g2_decap_8 FILLER_43_1110 ();
 sg13g2_decap_8 FILLER_43_1117 ();
 sg13g2_decap_8 FILLER_43_1124 ();
 sg13g2_decap_8 FILLER_43_1131 ();
 sg13g2_decap_8 FILLER_43_1138 ();
 sg13g2_decap_8 FILLER_43_1145 ();
 sg13g2_decap_8 FILLER_43_1152 ();
 sg13g2_decap_8 FILLER_43_1159 ();
 sg13g2_decap_8 FILLER_43_1166 ();
 sg13g2_decap_8 FILLER_43_1173 ();
 sg13g2_decap_8 FILLER_43_1180 ();
 sg13g2_decap_8 FILLER_43_1187 ();
 sg13g2_decap_8 FILLER_43_1194 ();
 sg13g2_decap_8 FILLER_43_1201 ();
 sg13g2_decap_8 FILLER_43_1208 ();
 sg13g2_decap_8 FILLER_43_1215 ();
 sg13g2_decap_8 FILLER_43_1222 ();
 sg13g2_decap_8 FILLER_43_1229 ();
 sg13g2_decap_8 FILLER_43_1236 ();
 sg13g2_decap_8 FILLER_43_1243 ();
 sg13g2_decap_8 FILLER_43_1250 ();
 sg13g2_decap_8 FILLER_43_1257 ();
 sg13g2_decap_8 FILLER_43_1264 ();
 sg13g2_decap_8 FILLER_43_1271 ();
 sg13g2_decap_8 FILLER_43_1278 ();
 sg13g2_decap_8 FILLER_43_1285 ();
 sg13g2_decap_8 FILLER_43_1292 ();
 sg13g2_decap_8 FILLER_43_1299 ();
 sg13g2_decap_8 FILLER_43_1306 ();
 sg13g2_fill_2 FILLER_43_1313 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_57 ();
 sg13g2_fill_2 FILLER_44_77 ();
 sg13g2_fill_2 FILLER_44_98 ();
 sg13g2_fill_1 FILLER_44_100 ();
 sg13g2_decap_4 FILLER_44_110 ();
 sg13g2_fill_2 FILLER_44_114 ();
 sg13g2_fill_1 FILLER_44_125 ();
 sg13g2_decap_8 FILLER_44_130 ();
 sg13g2_decap_4 FILLER_44_137 ();
 sg13g2_fill_1 FILLER_44_141 ();
 sg13g2_fill_2 FILLER_44_166 ();
 sg13g2_fill_2 FILLER_44_190 ();
 sg13g2_fill_1 FILLER_44_192 ();
 sg13g2_fill_2 FILLER_44_218 ();
 sg13g2_fill_1 FILLER_44_220 ();
 sg13g2_fill_1 FILLER_44_233 ();
 sg13g2_fill_2 FILLER_44_269 ();
 sg13g2_fill_1 FILLER_44_307 ();
 sg13g2_fill_2 FILLER_44_322 ();
 sg13g2_fill_1 FILLER_44_324 ();
 sg13g2_fill_2 FILLER_44_338 ();
 sg13g2_fill_2 FILLER_44_353 ();
 sg13g2_fill_1 FILLER_44_368 ();
 sg13g2_fill_2 FILLER_44_389 ();
 sg13g2_fill_1 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_420 ();
 sg13g2_decap_4 FILLER_44_445 ();
 sg13g2_fill_1 FILLER_44_449 ();
 sg13g2_fill_2 FILLER_44_455 ();
 sg13g2_decap_4 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_483 ();
 sg13g2_fill_1 FILLER_44_490 ();
 sg13g2_decap_8 FILLER_44_503 ();
 sg13g2_fill_1 FILLER_44_510 ();
 sg13g2_fill_2 FILLER_44_519 ();
 sg13g2_fill_1 FILLER_44_542 ();
 sg13g2_fill_2 FILLER_44_565 ();
 sg13g2_fill_2 FILLER_44_583 ();
 sg13g2_decap_8 FILLER_44_595 ();
 sg13g2_fill_1 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_620 ();
 sg13g2_decap_8 FILLER_44_627 ();
 sg13g2_fill_1 FILLER_44_634 ();
 sg13g2_fill_1 FILLER_44_650 ();
 sg13g2_fill_2 FILLER_44_656 ();
 sg13g2_fill_1 FILLER_44_658 ();
 sg13g2_decap_4 FILLER_44_685 ();
 sg13g2_fill_1 FILLER_44_694 ();
 sg13g2_decap_4 FILLER_44_700 ();
 sg13g2_decap_4 FILLER_44_720 ();
 sg13g2_fill_1 FILLER_44_732 ();
 sg13g2_decap_4 FILLER_44_737 ();
 sg13g2_fill_2 FILLER_44_741 ();
 sg13g2_decap_8 FILLER_44_756 ();
 sg13g2_fill_2 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_778 ();
 sg13g2_decap_8 FILLER_44_785 ();
 sg13g2_fill_1 FILLER_44_848 ();
 sg13g2_fill_2 FILLER_44_907 ();
 sg13g2_fill_2 FILLER_44_918 ();
 sg13g2_fill_1 FILLER_44_980 ();
 sg13g2_fill_1 FILLER_44_1020 ();
 sg13g2_decap_8 FILLER_44_1025 ();
 sg13g2_decap_8 FILLER_44_1032 ();
 sg13g2_decap_8 FILLER_44_1039 ();
 sg13g2_decap_8 FILLER_44_1046 ();
 sg13g2_decap_8 FILLER_44_1053 ();
 sg13g2_decap_8 FILLER_44_1060 ();
 sg13g2_decap_8 FILLER_44_1067 ();
 sg13g2_decap_8 FILLER_44_1074 ();
 sg13g2_decap_8 FILLER_44_1081 ();
 sg13g2_decap_8 FILLER_44_1088 ();
 sg13g2_decap_8 FILLER_44_1095 ();
 sg13g2_decap_8 FILLER_44_1102 ();
 sg13g2_decap_8 FILLER_44_1109 ();
 sg13g2_decap_8 FILLER_44_1116 ();
 sg13g2_decap_8 FILLER_44_1123 ();
 sg13g2_decap_8 FILLER_44_1130 ();
 sg13g2_decap_8 FILLER_44_1137 ();
 sg13g2_decap_8 FILLER_44_1144 ();
 sg13g2_decap_8 FILLER_44_1151 ();
 sg13g2_decap_8 FILLER_44_1158 ();
 sg13g2_decap_8 FILLER_44_1165 ();
 sg13g2_decap_8 FILLER_44_1172 ();
 sg13g2_decap_8 FILLER_44_1179 ();
 sg13g2_decap_8 FILLER_44_1186 ();
 sg13g2_decap_8 FILLER_44_1193 ();
 sg13g2_decap_8 FILLER_44_1200 ();
 sg13g2_decap_8 FILLER_44_1207 ();
 sg13g2_decap_8 FILLER_44_1214 ();
 sg13g2_decap_8 FILLER_44_1221 ();
 sg13g2_decap_8 FILLER_44_1228 ();
 sg13g2_decap_8 FILLER_44_1235 ();
 sg13g2_decap_8 FILLER_44_1242 ();
 sg13g2_decap_8 FILLER_44_1249 ();
 sg13g2_decap_8 FILLER_44_1256 ();
 sg13g2_decap_8 FILLER_44_1263 ();
 sg13g2_decap_8 FILLER_44_1270 ();
 sg13g2_decap_8 FILLER_44_1277 ();
 sg13g2_decap_8 FILLER_44_1284 ();
 sg13g2_decap_8 FILLER_44_1291 ();
 sg13g2_decap_8 FILLER_44_1298 ();
 sg13g2_decap_8 FILLER_44_1305 ();
 sg13g2_fill_2 FILLER_44_1312 ();
 sg13g2_fill_1 FILLER_44_1314 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_11 ();
 sg13g2_decap_8 FILLER_45_31 ();
 sg13g2_fill_2 FILLER_45_60 ();
 sg13g2_fill_1 FILLER_45_62 ();
 sg13g2_fill_1 FILLER_45_68 ();
 sg13g2_fill_2 FILLER_45_100 ();
 sg13g2_fill_1 FILLER_45_102 ();
 sg13g2_fill_2 FILLER_45_155 ();
 sg13g2_fill_1 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_199 ();
 sg13g2_fill_2 FILLER_45_209 ();
 sg13g2_fill_1 FILLER_45_211 ();
 sg13g2_fill_2 FILLER_45_221 ();
 sg13g2_fill_1 FILLER_45_223 ();
 sg13g2_fill_2 FILLER_45_232 ();
 sg13g2_fill_2 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_244 ();
 sg13g2_fill_1 FILLER_45_258 ();
 sg13g2_fill_2 FILLER_45_286 ();
 sg13g2_fill_1 FILLER_45_288 ();
 sg13g2_fill_1 FILLER_45_298 ();
 sg13g2_fill_1 FILLER_45_339 ();
 sg13g2_fill_2 FILLER_45_348 ();
 sg13g2_fill_1 FILLER_45_365 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_fill_1 FILLER_45_378 ();
 sg13g2_decap_4 FILLER_45_387 ();
 sg13g2_fill_2 FILLER_45_391 ();
 sg13g2_decap_8 FILLER_45_410 ();
 sg13g2_fill_2 FILLER_45_417 ();
 sg13g2_fill_1 FILLER_45_419 ();
 sg13g2_decap_4 FILLER_45_425 ();
 sg13g2_fill_2 FILLER_45_439 ();
 sg13g2_fill_2 FILLER_45_465 ();
 sg13g2_fill_2 FILLER_45_483 ();
 sg13g2_fill_1 FILLER_45_485 ();
 sg13g2_fill_1 FILLER_45_529 ();
 sg13g2_decap_4 FILLER_45_535 ();
 sg13g2_decap_8 FILLER_45_560 ();
 sg13g2_decap_8 FILLER_45_567 ();
 sg13g2_decap_4 FILLER_45_574 ();
 sg13g2_fill_1 FILLER_45_591 ();
 sg13g2_fill_2 FILLER_45_601 ();
 sg13g2_fill_1 FILLER_45_603 ();
 sg13g2_decap_4 FILLER_45_613 ();
 sg13g2_decap_4 FILLER_45_643 ();
 sg13g2_fill_2 FILLER_45_679 ();
 sg13g2_fill_1 FILLER_45_681 ();
 sg13g2_fill_2 FILLER_45_690 ();
 sg13g2_fill_1 FILLER_45_692 ();
 sg13g2_decap_8 FILLER_45_698 ();
 sg13g2_fill_2 FILLER_45_720 ();
 sg13g2_fill_1 FILLER_45_722 ();
 sg13g2_fill_2 FILLER_45_756 ();
 sg13g2_fill_1 FILLER_45_758 ();
 sg13g2_decap_8 FILLER_45_785 ();
 sg13g2_decap_4 FILLER_45_792 ();
 sg13g2_fill_1 FILLER_45_810 ();
 sg13g2_fill_2 FILLER_45_830 ();
 sg13g2_fill_1 FILLER_45_832 ();
 sg13g2_fill_2 FILLER_45_894 ();
 sg13g2_fill_1 FILLER_45_896 ();
 sg13g2_fill_2 FILLER_45_1005 ();
 sg13g2_fill_1 FILLER_45_1007 ();
 sg13g2_fill_2 FILLER_45_1034 ();
 sg13g2_decap_8 FILLER_45_1045 ();
 sg13g2_decap_8 FILLER_45_1052 ();
 sg13g2_decap_8 FILLER_45_1059 ();
 sg13g2_decap_8 FILLER_45_1066 ();
 sg13g2_decap_8 FILLER_45_1073 ();
 sg13g2_decap_8 FILLER_45_1080 ();
 sg13g2_decap_8 FILLER_45_1087 ();
 sg13g2_decap_8 FILLER_45_1094 ();
 sg13g2_decap_8 FILLER_45_1101 ();
 sg13g2_decap_8 FILLER_45_1108 ();
 sg13g2_decap_8 FILLER_45_1115 ();
 sg13g2_decap_8 FILLER_45_1122 ();
 sg13g2_decap_8 FILLER_45_1129 ();
 sg13g2_decap_8 FILLER_45_1136 ();
 sg13g2_decap_8 FILLER_45_1143 ();
 sg13g2_decap_8 FILLER_45_1150 ();
 sg13g2_decap_8 FILLER_45_1157 ();
 sg13g2_decap_8 FILLER_45_1164 ();
 sg13g2_decap_8 FILLER_45_1171 ();
 sg13g2_decap_8 FILLER_45_1178 ();
 sg13g2_decap_8 FILLER_45_1185 ();
 sg13g2_decap_8 FILLER_45_1192 ();
 sg13g2_decap_8 FILLER_45_1199 ();
 sg13g2_decap_8 FILLER_45_1206 ();
 sg13g2_decap_8 FILLER_45_1213 ();
 sg13g2_decap_8 FILLER_45_1220 ();
 sg13g2_decap_8 FILLER_45_1227 ();
 sg13g2_decap_8 FILLER_45_1234 ();
 sg13g2_decap_8 FILLER_45_1241 ();
 sg13g2_decap_8 FILLER_45_1248 ();
 sg13g2_decap_8 FILLER_45_1255 ();
 sg13g2_decap_8 FILLER_45_1262 ();
 sg13g2_decap_8 FILLER_45_1269 ();
 sg13g2_decap_8 FILLER_45_1276 ();
 sg13g2_decap_8 FILLER_45_1283 ();
 sg13g2_decap_8 FILLER_45_1290 ();
 sg13g2_decap_8 FILLER_45_1297 ();
 sg13g2_decap_8 FILLER_45_1304 ();
 sg13g2_decap_4 FILLER_45_1311 ();
 sg13g2_fill_1 FILLER_46_50 ();
 sg13g2_decap_4 FILLER_46_83 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_decap_4 FILLER_46_96 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_fill_1 FILLER_46_106 ();
 sg13g2_fill_1 FILLER_46_150 ();
 sg13g2_fill_1 FILLER_46_194 ();
 sg13g2_decap_8 FILLER_46_230 ();
 sg13g2_fill_1 FILLER_46_237 ();
 sg13g2_fill_2 FILLER_46_287 ();
 sg13g2_fill_1 FILLER_46_298 ();
 sg13g2_fill_1 FILLER_46_318 ();
 sg13g2_fill_2 FILLER_46_348 ();
 sg13g2_fill_2 FILLER_46_389 ();
 sg13g2_decap_4 FILLER_46_401 ();
 sg13g2_fill_2 FILLER_46_435 ();
 sg13g2_decap_4 FILLER_46_445 ();
 sg13g2_decap_8 FILLER_46_465 ();
 sg13g2_decap_4 FILLER_46_484 ();
 sg13g2_fill_2 FILLER_46_488 ();
 sg13g2_fill_1 FILLER_46_495 ();
 sg13g2_decap_4 FILLER_46_506 ();
 sg13g2_fill_2 FILLER_46_510 ();
 sg13g2_fill_2 FILLER_46_522 ();
 sg13g2_fill_2 FILLER_46_532 ();
 sg13g2_decap_4 FILLER_46_538 ();
 sg13g2_fill_1 FILLER_46_577 ();
 sg13g2_fill_1 FILLER_46_619 ();
 sg13g2_decap_4 FILLER_46_632 ();
 sg13g2_fill_2 FILLER_46_658 ();
 sg13g2_fill_1 FILLER_46_660 ();
 sg13g2_fill_2 FILLER_46_675 ();
 sg13g2_fill_1 FILLER_46_677 ();
 sg13g2_fill_2 FILLER_46_683 ();
 sg13g2_fill_1 FILLER_46_685 ();
 sg13g2_fill_2 FILLER_46_699 ();
 sg13g2_decap_4 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_fill_1 FILLER_46_742 ();
 sg13g2_fill_1 FILLER_46_758 ();
 sg13g2_fill_2 FILLER_46_836 ();
 sg13g2_fill_1 FILLER_46_838 ();
 sg13g2_fill_1 FILLER_46_858 ();
 sg13g2_fill_2 FILLER_46_868 ();
 sg13g2_fill_1 FILLER_46_870 ();
 sg13g2_fill_2 FILLER_46_932 ();
 sg13g2_fill_1 FILLER_46_939 ();
 sg13g2_fill_2 FILLER_46_1005 ();
 sg13g2_decap_8 FILLER_46_1025 ();
 sg13g2_decap_8 FILLER_46_1032 ();
 sg13g2_decap_8 FILLER_46_1039 ();
 sg13g2_decap_8 FILLER_46_1046 ();
 sg13g2_decap_8 FILLER_46_1053 ();
 sg13g2_decap_8 FILLER_46_1060 ();
 sg13g2_decap_8 FILLER_46_1067 ();
 sg13g2_decap_8 FILLER_46_1074 ();
 sg13g2_decap_8 FILLER_46_1081 ();
 sg13g2_decap_8 FILLER_46_1088 ();
 sg13g2_decap_8 FILLER_46_1095 ();
 sg13g2_decap_8 FILLER_46_1102 ();
 sg13g2_decap_8 FILLER_46_1109 ();
 sg13g2_decap_8 FILLER_46_1116 ();
 sg13g2_decap_8 FILLER_46_1123 ();
 sg13g2_decap_8 FILLER_46_1130 ();
 sg13g2_decap_8 FILLER_46_1137 ();
 sg13g2_decap_8 FILLER_46_1144 ();
 sg13g2_decap_8 FILLER_46_1151 ();
 sg13g2_decap_8 FILLER_46_1158 ();
 sg13g2_decap_8 FILLER_46_1165 ();
 sg13g2_decap_8 FILLER_46_1172 ();
 sg13g2_decap_8 FILLER_46_1179 ();
 sg13g2_decap_8 FILLER_46_1186 ();
 sg13g2_decap_8 FILLER_46_1193 ();
 sg13g2_decap_8 FILLER_46_1200 ();
 sg13g2_decap_8 FILLER_46_1207 ();
 sg13g2_decap_8 FILLER_46_1214 ();
 sg13g2_decap_8 FILLER_46_1221 ();
 sg13g2_decap_8 FILLER_46_1228 ();
 sg13g2_decap_8 FILLER_46_1235 ();
 sg13g2_decap_8 FILLER_46_1242 ();
 sg13g2_decap_8 FILLER_46_1249 ();
 sg13g2_decap_8 FILLER_46_1256 ();
 sg13g2_decap_8 FILLER_46_1263 ();
 sg13g2_decap_8 FILLER_46_1270 ();
 sg13g2_decap_8 FILLER_46_1277 ();
 sg13g2_decap_8 FILLER_46_1284 ();
 sg13g2_decap_8 FILLER_46_1291 ();
 sg13g2_decap_8 FILLER_46_1298 ();
 sg13g2_decap_8 FILLER_46_1305 ();
 sg13g2_fill_2 FILLER_46_1312 ();
 sg13g2_fill_1 FILLER_46_1314 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_37 ();
 sg13g2_fill_1 FILLER_47_78 ();
 sg13g2_fill_1 FILLER_47_90 ();
 sg13g2_fill_2 FILLER_47_114 ();
 sg13g2_fill_1 FILLER_47_116 ();
 sg13g2_fill_2 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_172 ();
 sg13g2_fill_1 FILLER_47_189 ();
 sg13g2_fill_2 FILLER_47_196 ();
 sg13g2_fill_2 FILLER_47_207 ();
 sg13g2_fill_2 FILLER_47_228 ();
 sg13g2_decap_4 FILLER_47_237 ();
 sg13g2_fill_1 FILLER_47_261 ();
 sg13g2_fill_1 FILLER_47_292 ();
 sg13g2_fill_2 FILLER_47_354 ();
 sg13g2_fill_1 FILLER_47_356 ();
 sg13g2_fill_1 FILLER_47_368 ();
 sg13g2_decap_8 FILLER_47_373 ();
 sg13g2_decap_8 FILLER_47_380 ();
 sg13g2_fill_2 FILLER_47_387 ();
 sg13g2_fill_1 FILLER_47_389 ();
 sg13g2_fill_1 FILLER_47_393 ();
 sg13g2_decap_4 FILLER_47_408 ();
 sg13g2_decap_4 FILLER_47_438 ();
 sg13g2_decap_8 FILLER_47_445 ();
 sg13g2_fill_1 FILLER_47_452 ();
 sg13g2_fill_2 FILLER_47_480 ();
 sg13g2_decap_8 FILLER_47_499 ();
 sg13g2_fill_2 FILLER_47_541 ();
 sg13g2_fill_1 FILLER_47_543 ();
 sg13g2_fill_2 FILLER_47_560 ();
 sg13g2_decap_4 FILLER_47_566 ();
 sg13g2_fill_1 FILLER_47_570 ();
 sg13g2_fill_1 FILLER_47_580 ();
 sg13g2_decap_4 FILLER_47_616 ();
 sg13g2_fill_1 FILLER_47_620 ();
 sg13g2_fill_1 FILLER_47_639 ();
 sg13g2_fill_1 FILLER_47_688 ();
 sg13g2_decap_8 FILLER_47_732 ();
 sg13g2_decap_8 FILLER_47_757 ();
 sg13g2_decap_4 FILLER_47_764 ();
 sg13g2_fill_1 FILLER_47_768 ();
 sg13g2_fill_2 FILLER_47_807 ();
 sg13g2_fill_1 FILLER_47_809 ();
 sg13g2_fill_2 FILLER_47_820 ();
 sg13g2_fill_1 FILLER_47_848 ();
 sg13g2_fill_2 FILLER_47_875 ();
 sg13g2_fill_1 FILLER_47_877 ();
 sg13g2_fill_2 FILLER_47_887 ();
 sg13g2_fill_1 FILLER_47_907 ();
 sg13g2_fill_1 FILLER_47_948 ();
 sg13g2_fill_2 FILLER_47_967 ();
 sg13g2_fill_1 FILLER_47_969 ();
 sg13g2_decap_8 FILLER_47_1026 ();
 sg13g2_decap_8 FILLER_47_1033 ();
 sg13g2_decap_8 FILLER_47_1040 ();
 sg13g2_decap_8 FILLER_47_1047 ();
 sg13g2_decap_8 FILLER_47_1054 ();
 sg13g2_decap_8 FILLER_47_1061 ();
 sg13g2_decap_8 FILLER_47_1068 ();
 sg13g2_decap_8 FILLER_47_1075 ();
 sg13g2_decap_8 FILLER_47_1082 ();
 sg13g2_decap_8 FILLER_47_1089 ();
 sg13g2_decap_8 FILLER_47_1096 ();
 sg13g2_decap_8 FILLER_47_1103 ();
 sg13g2_decap_8 FILLER_47_1110 ();
 sg13g2_decap_8 FILLER_47_1117 ();
 sg13g2_decap_8 FILLER_47_1124 ();
 sg13g2_decap_8 FILLER_47_1131 ();
 sg13g2_decap_8 FILLER_47_1138 ();
 sg13g2_decap_8 FILLER_47_1145 ();
 sg13g2_decap_8 FILLER_47_1152 ();
 sg13g2_decap_8 FILLER_47_1159 ();
 sg13g2_decap_8 FILLER_47_1166 ();
 sg13g2_decap_8 FILLER_47_1173 ();
 sg13g2_decap_8 FILLER_47_1180 ();
 sg13g2_decap_8 FILLER_47_1187 ();
 sg13g2_decap_8 FILLER_47_1194 ();
 sg13g2_decap_8 FILLER_47_1201 ();
 sg13g2_decap_8 FILLER_47_1208 ();
 sg13g2_decap_8 FILLER_47_1215 ();
 sg13g2_decap_8 FILLER_47_1222 ();
 sg13g2_decap_8 FILLER_47_1229 ();
 sg13g2_decap_8 FILLER_47_1236 ();
 sg13g2_decap_8 FILLER_47_1243 ();
 sg13g2_decap_8 FILLER_47_1250 ();
 sg13g2_decap_8 FILLER_47_1257 ();
 sg13g2_decap_8 FILLER_47_1264 ();
 sg13g2_decap_8 FILLER_47_1271 ();
 sg13g2_decap_8 FILLER_47_1278 ();
 sg13g2_decap_8 FILLER_47_1285 ();
 sg13g2_decap_8 FILLER_47_1292 ();
 sg13g2_decap_8 FILLER_47_1299 ();
 sg13g2_decap_8 FILLER_47_1306 ();
 sg13g2_fill_2 FILLER_47_1313 ();
 sg13g2_fill_2 FILLER_48_31 ();
 sg13g2_fill_2 FILLER_48_48 ();
 sg13g2_decap_4 FILLER_48_70 ();
 sg13g2_fill_1 FILLER_48_74 ();
 sg13g2_fill_2 FILLER_48_80 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_fill_2 FILLER_48_103 ();
 sg13g2_fill_1 FILLER_48_105 ();
 sg13g2_fill_1 FILLER_48_154 ();
 sg13g2_fill_1 FILLER_48_244 ();
 sg13g2_fill_2 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_265 ();
 sg13g2_fill_2 FILLER_48_284 ();
 sg13g2_fill_2 FILLER_48_312 ();
 sg13g2_decap_4 FILLER_48_318 ();
 sg13g2_fill_2 FILLER_48_322 ();
 sg13g2_fill_1 FILLER_48_350 ();
 sg13g2_fill_1 FILLER_48_380 ();
 sg13g2_decap_8 FILLER_48_389 ();
 sg13g2_decap_8 FILLER_48_396 ();
 sg13g2_decap_4 FILLER_48_403 ();
 sg13g2_fill_2 FILLER_48_419 ();
 sg13g2_fill_1 FILLER_48_421 ();
 sg13g2_fill_1 FILLER_48_453 ();
 sg13g2_fill_1 FILLER_48_462 ();
 sg13g2_fill_2 FILLER_48_485 ();
 sg13g2_fill_1 FILLER_48_487 ();
 sg13g2_decap_4 FILLER_48_503 ();
 sg13g2_fill_2 FILLER_48_507 ();
 sg13g2_fill_1 FILLER_48_525 ();
 sg13g2_decap_4 FILLER_48_534 ();
 sg13g2_decap_4 FILLER_48_567 ();
 sg13g2_fill_1 FILLER_48_571 ();
 sg13g2_decap_4 FILLER_48_576 ();
 sg13g2_fill_2 FILLER_48_580 ();
 sg13g2_decap_8 FILLER_48_590 ();
 sg13g2_decap_8 FILLER_48_597 ();
 sg13g2_decap_4 FILLER_48_613 ();
 sg13g2_fill_2 FILLER_48_617 ();
 sg13g2_fill_1 FILLER_48_628 ();
 sg13g2_fill_1 FILLER_48_655 ();
 sg13g2_fill_1 FILLER_48_704 ();
 sg13g2_fill_2 FILLER_48_714 ();
 sg13g2_fill_1 FILLER_48_716 ();
 sg13g2_decap_4 FILLER_48_722 ();
 sg13g2_decap_4 FILLER_48_730 ();
 sg13g2_fill_1 FILLER_48_734 ();
 sg13g2_fill_2 FILLER_48_744 ();
 sg13g2_fill_1 FILLER_48_746 ();
 sg13g2_fill_1 FILLER_48_752 ();
 sg13g2_fill_1 FILLER_48_757 ();
 sg13g2_fill_1 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_797 ();
 sg13g2_fill_2 FILLER_48_804 ();
 sg13g2_fill_1 FILLER_48_806 ();
 sg13g2_decap_4 FILLER_48_816 ();
 sg13g2_fill_2 FILLER_48_820 ();
 sg13g2_fill_2 FILLER_48_856 ();
 sg13g2_fill_1 FILLER_48_858 ();
 sg13g2_fill_2 FILLER_48_994 ();
 sg13g2_fill_2 FILLER_48_1013 ();
 sg13g2_fill_1 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1042 ();
 sg13g2_decap_8 FILLER_48_1049 ();
 sg13g2_decap_8 FILLER_48_1056 ();
 sg13g2_decap_8 FILLER_48_1063 ();
 sg13g2_decap_8 FILLER_48_1070 ();
 sg13g2_decap_8 FILLER_48_1077 ();
 sg13g2_decap_8 FILLER_48_1084 ();
 sg13g2_decap_8 FILLER_48_1091 ();
 sg13g2_decap_8 FILLER_48_1098 ();
 sg13g2_decap_8 FILLER_48_1105 ();
 sg13g2_decap_8 FILLER_48_1112 ();
 sg13g2_decap_8 FILLER_48_1119 ();
 sg13g2_decap_8 FILLER_48_1126 ();
 sg13g2_decap_8 FILLER_48_1133 ();
 sg13g2_decap_8 FILLER_48_1140 ();
 sg13g2_decap_8 FILLER_48_1147 ();
 sg13g2_decap_8 FILLER_48_1154 ();
 sg13g2_decap_8 FILLER_48_1161 ();
 sg13g2_decap_8 FILLER_48_1168 ();
 sg13g2_decap_8 FILLER_48_1175 ();
 sg13g2_decap_8 FILLER_48_1182 ();
 sg13g2_decap_8 FILLER_48_1189 ();
 sg13g2_decap_8 FILLER_48_1196 ();
 sg13g2_decap_8 FILLER_48_1203 ();
 sg13g2_decap_8 FILLER_48_1210 ();
 sg13g2_decap_8 FILLER_48_1217 ();
 sg13g2_decap_8 FILLER_48_1224 ();
 sg13g2_decap_8 FILLER_48_1231 ();
 sg13g2_decap_8 FILLER_48_1238 ();
 sg13g2_decap_8 FILLER_48_1245 ();
 sg13g2_decap_8 FILLER_48_1252 ();
 sg13g2_decap_8 FILLER_48_1259 ();
 sg13g2_decap_8 FILLER_48_1266 ();
 sg13g2_decap_8 FILLER_48_1273 ();
 sg13g2_decap_8 FILLER_48_1280 ();
 sg13g2_decap_8 FILLER_48_1287 ();
 sg13g2_decap_8 FILLER_48_1294 ();
 sg13g2_decap_8 FILLER_48_1301 ();
 sg13g2_decap_8 FILLER_48_1308 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_26 ();
 sg13g2_fill_2 FILLER_49_35 ();
 sg13g2_decap_4 FILLER_49_47 ();
 sg13g2_fill_1 FILLER_49_51 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_decap_4 FILLER_49_83 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_fill_2 FILLER_49_160 ();
 sg13g2_fill_1 FILLER_49_162 ();
 sg13g2_fill_2 FILLER_49_168 ();
 sg13g2_decap_4 FILLER_49_174 ();
 sg13g2_fill_2 FILLER_49_178 ();
 sg13g2_decap_4 FILLER_49_240 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_decap_4 FILLER_49_297 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_fill_2 FILLER_49_334 ();
 sg13g2_decap_4 FILLER_49_367 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_386 ();
 sg13g2_decap_4 FILLER_49_393 ();
 sg13g2_fill_2 FILLER_49_401 ();
 sg13g2_decap_4 FILLER_49_424 ();
 sg13g2_fill_1 FILLER_49_428 ();
 sg13g2_decap_8 FILLER_49_447 ();
 sg13g2_decap_8 FILLER_49_485 ();
 sg13g2_decap_4 FILLER_49_492 ();
 sg13g2_fill_1 FILLER_49_496 ();
 sg13g2_fill_2 FILLER_49_501 ();
 sg13g2_fill_1 FILLER_49_529 ();
 sg13g2_decap_4 FILLER_49_587 ();
 sg13g2_fill_1 FILLER_49_591 ();
 sg13g2_fill_2 FILLER_49_621 ();
 sg13g2_fill_1 FILLER_49_623 ();
 sg13g2_fill_2 FILLER_49_650 ();
 sg13g2_fill_1 FILLER_49_652 ();
 sg13g2_decap_4 FILLER_49_679 ();
 sg13g2_fill_2 FILLER_49_683 ();
 sg13g2_decap_8 FILLER_49_706 ();
 sg13g2_decap_8 FILLER_49_713 ();
 sg13g2_decap_4 FILLER_49_720 ();
 sg13g2_fill_2 FILLER_49_724 ();
 sg13g2_fill_2 FILLER_49_739 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_4 FILLER_49_763 ();
 sg13g2_fill_2 FILLER_49_767 ();
 sg13g2_fill_2 FILLER_49_777 ();
 sg13g2_fill_1 FILLER_49_779 ();
 sg13g2_fill_2 FILLER_49_789 ();
 sg13g2_fill_2 FILLER_49_799 ();
 sg13g2_fill_2 FILLER_49_923 ();
 sg13g2_fill_2 FILLER_49_974 ();
 sg13g2_fill_1 FILLER_49_976 ();
 sg13g2_fill_1 FILLER_49_1033 ();
 sg13g2_decap_8 FILLER_49_1043 ();
 sg13g2_decap_8 FILLER_49_1050 ();
 sg13g2_decap_8 FILLER_49_1057 ();
 sg13g2_decap_8 FILLER_49_1064 ();
 sg13g2_decap_8 FILLER_49_1071 ();
 sg13g2_decap_8 FILLER_49_1078 ();
 sg13g2_decap_8 FILLER_49_1085 ();
 sg13g2_decap_8 FILLER_49_1092 ();
 sg13g2_decap_8 FILLER_49_1099 ();
 sg13g2_decap_8 FILLER_49_1106 ();
 sg13g2_decap_8 FILLER_49_1113 ();
 sg13g2_decap_8 FILLER_49_1120 ();
 sg13g2_decap_8 FILLER_49_1127 ();
 sg13g2_decap_8 FILLER_49_1134 ();
 sg13g2_decap_8 FILLER_49_1141 ();
 sg13g2_decap_8 FILLER_49_1148 ();
 sg13g2_decap_8 FILLER_49_1155 ();
 sg13g2_decap_8 FILLER_49_1162 ();
 sg13g2_decap_8 FILLER_49_1169 ();
 sg13g2_decap_8 FILLER_49_1176 ();
 sg13g2_decap_8 FILLER_49_1183 ();
 sg13g2_decap_8 FILLER_49_1190 ();
 sg13g2_decap_8 FILLER_49_1197 ();
 sg13g2_decap_8 FILLER_49_1204 ();
 sg13g2_decap_8 FILLER_49_1211 ();
 sg13g2_decap_8 FILLER_49_1218 ();
 sg13g2_decap_8 FILLER_49_1225 ();
 sg13g2_decap_8 FILLER_49_1232 ();
 sg13g2_decap_8 FILLER_49_1239 ();
 sg13g2_decap_8 FILLER_49_1246 ();
 sg13g2_decap_8 FILLER_49_1253 ();
 sg13g2_decap_8 FILLER_49_1260 ();
 sg13g2_decap_8 FILLER_49_1267 ();
 sg13g2_decap_8 FILLER_49_1274 ();
 sg13g2_decap_8 FILLER_49_1281 ();
 sg13g2_decap_8 FILLER_49_1288 ();
 sg13g2_decap_8 FILLER_49_1295 ();
 sg13g2_decap_8 FILLER_49_1302 ();
 sg13g2_decap_4 FILLER_49_1309 ();
 sg13g2_fill_2 FILLER_49_1313 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_36 ();
 sg13g2_fill_2 FILLER_50_43 ();
 sg13g2_fill_2 FILLER_50_53 ();
 sg13g2_decap_8 FILLER_50_65 ();
 sg13g2_fill_1 FILLER_50_72 ();
 sg13g2_decap_8 FILLER_50_78 ();
 sg13g2_fill_1 FILLER_50_95 ();
 sg13g2_decap_8 FILLER_50_101 ();
 sg13g2_fill_1 FILLER_50_108 ();
 sg13g2_fill_2 FILLER_50_152 ();
 sg13g2_fill_1 FILLER_50_215 ();
 sg13g2_fill_2 FILLER_50_231 ();
 sg13g2_fill_2 FILLER_50_241 ();
 sg13g2_fill_1 FILLER_50_258 ();
 sg13g2_fill_2 FILLER_50_274 ();
 sg13g2_decap_8 FILLER_50_280 ();
 sg13g2_fill_2 FILLER_50_291 ();
 sg13g2_fill_1 FILLER_50_293 ();
 sg13g2_fill_1 FILLER_50_315 ();
 sg13g2_fill_2 FILLER_50_320 ();
 sg13g2_fill_1 FILLER_50_322 ();
 sg13g2_fill_1 FILLER_50_340 ();
 sg13g2_decap_4 FILLER_50_354 ();
 sg13g2_fill_2 FILLER_50_361 ();
 sg13g2_fill_1 FILLER_50_363 ();
 sg13g2_fill_2 FILLER_50_373 ();
 sg13g2_fill_1 FILLER_50_375 ();
 sg13g2_decap_4 FILLER_50_381 ();
 sg13g2_fill_1 FILLER_50_385 ();
 sg13g2_decap_4 FILLER_50_429 ();
 sg13g2_fill_1 FILLER_50_438 ();
 sg13g2_decap_4 FILLER_50_448 ();
 sg13g2_fill_2 FILLER_50_462 ();
 sg13g2_fill_1 FILLER_50_464 ();
 sg13g2_decap_4 FILLER_50_469 ();
 sg13g2_fill_1 FILLER_50_473 ();
 sg13g2_fill_1 FILLER_50_487 ();
 sg13g2_fill_2 FILLER_50_508 ();
 sg13g2_fill_1 FILLER_50_523 ();
 sg13g2_fill_2 FILLER_50_544 ();
 sg13g2_fill_2 FILLER_50_576 ();
 sg13g2_fill_1 FILLER_50_582 ();
 sg13g2_decap_4 FILLER_50_616 ();
 sg13g2_fill_2 FILLER_50_635 ();
 sg13g2_decap_8 FILLER_50_650 ();
 sg13g2_decap_4 FILLER_50_657 ();
 sg13g2_fill_1 FILLER_50_661 ();
 sg13g2_decap_4 FILLER_50_685 ();
 sg13g2_decap_8 FILLER_50_693 ();
 sg13g2_decap_8 FILLER_50_700 ();
 sg13g2_fill_2 FILLER_50_717 ();
 sg13g2_fill_1 FILLER_50_719 ();
 sg13g2_fill_2 FILLER_50_730 ();
 sg13g2_fill_1 FILLER_50_745 ();
 sg13g2_fill_2 FILLER_50_772 ();
 sg13g2_decap_4 FILLER_50_778 ();
 sg13g2_fill_2 FILLER_50_808 ();
 sg13g2_fill_2 FILLER_50_827 ();
 sg13g2_fill_1 FILLER_50_829 ();
 sg13g2_fill_1 FILLER_50_834 ();
 sg13g2_fill_1 FILLER_50_878 ();
 sg13g2_fill_1 FILLER_50_901 ();
 sg13g2_fill_2 FILLER_50_928 ();
 sg13g2_decap_8 FILLER_50_1020 ();
 sg13g2_decap_8 FILLER_50_1027 ();
 sg13g2_decap_8 FILLER_50_1034 ();
 sg13g2_decap_8 FILLER_50_1041 ();
 sg13g2_decap_8 FILLER_50_1048 ();
 sg13g2_decap_8 FILLER_50_1055 ();
 sg13g2_decap_8 FILLER_50_1062 ();
 sg13g2_decap_8 FILLER_50_1069 ();
 sg13g2_decap_8 FILLER_50_1076 ();
 sg13g2_decap_8 FILLER_50_1083 ();
 sg13g2_decap_8 FILLER_50_1090 ();
 sg13g2_decap_8 FILLER_50_1097 ();
 sg13g2_decap_8 FILLER_50_1104 ();
 sg13g2_decap_8 FILLER_50_1111 ();
 sg13g2_decap_8 FILLER_50_1118 ();
 sg13g2_decap_8 FILLER_50_1125 ();
 sg13g2_decap_8 FILLER_50_1132 ();
 sg13g2_decap_8 FILLER_50_1139 ();
 sg13g2_decap_8 FILLER_50_1146 ();
 sg13g2_decap_8 FILLER_50_1153 ();
 sg13g2_decap_8 FILLER_50_1160 ();
 sg13g2_decap_8 FILLER_50_1167 ();
 sg13g2_decap_8 FILLER_50_1174 ();
 sg13g2_decap_8 FILLER_50_1181 ();
 sg13g2_decap_8 FILLER_50_1188 ();
 sg13g2_decap_8 FILLER_50_1195 ();
 sg13g2_decap_8 FILLER_50_1202 ();
 sg13g2_decap_8 FILLER_50_1209 ();
 sg13g2_decap_8 FILLER_50_1216 ();
 sg13g2_decap_8 FILLER_50_1223 ();
 sg13g2_decap_8 FILLER_50_1230 ();
 sg13g2_decap_8 FILLER_50_1237 ();
 sg13g2_decap_8 FILLER_50_1244 ();
 sg13g2_decap_8 FILLER_50_1251 ();
 sg13g2_decap_8 FILLER_50_1258 ();
 sg13g2_decap_8 FILLER_50_1265 ();
 sg13g2_decap_8 FILLER_50_1272 ();
 sg13g2_decap_8 FILLER_50_1279 ();
 sg13g2_decap_8 FILLER_50_1286 ();
 sg13g2_decap_8 FILLER_50_1293 ();
 sg13g2_decap_8 FILLER_50_1300 ();
 sg13g2_decap_8 FILLER_50_1307 ();
 sg13g2_fill_1 FILLER_50_1314 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_fill_1 FILLER_51_11 ();
 sg13g2_fill_1 FILLER_51_63 ();
 sg13g2_fill_1 FILLER_51_112 ();
 sg13g2_fill_1 FILLER_51_128 ();
 sg13g2_fill_1 FILLER_51_235 ();
 sg13g2_fill_2 FILLER_51_272 ();
 sg13g2_fill_1 FILLER_51_274 ();
 sg13g2_fill_2 FILLER_51_285 ();
 sg13g2_decap_8 FILLER_51_292 ();
 sg13g2_decap_4 FILLER_51_299 ();
 sg13g2_fill_2 FILLER_51_303 ();
 sg13g2_fill_2 FILLER_51_331 ();
 sg13g2_fill_1 FILLER_51_333 ();
 sg13g2_fill_2 FILLER_51_339 ();
 sg13g2_fill_1 FILLER_51_341 ();
 sg13g2_decap_4 FILLER_51_354 ();
 sg13g2_fill_2 FILLER_51_378 ();
 sg13g2_decap_8 FILLER_51_388 ();
 sg13g2_decap_4 FILLER_51_395 ();
 sg13g2_fill_2 FILLER_51_399 ();
 sg13g2_fill_1 FILLER_51_411 ();
 sg13g2_fill_1 FILLER_51_431 ();
 sg13g2_fill_2 FILLER_51_451 ();
 sg13g2_fill_1 FILLER_51_453 ();
 sg13g2_fill_2 FILLER_51_467 ();
 sg13g2_fill_1 FILLER_51_469 ();
 sg13g2_decap_8 FILLER_51_486 ();
 sg13g2_decap_8 FILLER_51_502 ();
 sg13g2_fill_2 FILLER_51_509 ();
 sg13g2_fill_1 FILLER_51_525 ();
 sg13g2_fill_1 FILLER_51_603 ();
 sg13g2_decap_8 FILLER_51_613 ();
 sg13g2_fill_2 FILLER_51_620 ();
 sg13g2_fill_1 FILLER_51_622 ();
 sg13g2_fill_2 FILLER_51_667 ();
 sg13g2_fill_2 FILLER_51_674 ();
 sg13g2_fill_1 FILLER_51_697 ();
 sg13g2_decap_4 FILLER_51_755 ();
 sg13g2_fill_1 FILLER_51_777 ();
 sg13g2_fill_2 FILLER_51_799 ();
 sg13g2_fill_1 FILLER_51_801 ();
 sg13g2_decap_8 FILLER_51_806 ();
 sg13g2_decap_4 FILLER_51_813 ();
 sg13g2_fill_1 FILLER_51_817 ();
 sg13g2_fill_1 FILLER_51_828 ();
 sg13g2_fill_1 FILLER_51_859 ();
 sg13g2_fill_2 FILLER_51_972 ();
 sg13g2_fill_1 FILLER_51_974 ();
 sg13g2_decap_8 FILLER_51_1001 ();
 sg13g2_decap_8 FILLER_51_1008 ();
 sg13g2_decap_8 FILLER_51_1015 ();
 sg13g2_decap_8 FILLER_51_1022 ();
 sg13g2_decap_8 FILLER_51_1029 ();
 sg13g2_decap_8 FILLER_51_1036 ();
 sg13g2_decap_8 FILLER_51_1043 ();
 sg13g2_decap_8 FILLER_51_1050 ();
 sg13g2_decap_8 FILLER_51_1057 ();
 sg13g2_decap_8 FILLER_51_1064 ();
 sg13g2_decap_8 FILLER_51_1071 ();
 sg13g2_decap_8 FILLER_51_1078 ();
 sg13g2_decap_8 FILLER_51_1085 ();
 sg13g2_decap_8 FILLER_51_1092 ();
 sg13g2_decap_8 FILLER_51_1099 ();
 sg13g2_decap_8 FILLER_51_1106 ();
 sg13g2_decap_8 FILLER_51_1113 ();
 sg13g2_decap_8 FILLER_51_1120 ();
 sg13g2_decap_8 FILLER_51_1127 ();
 sg13g2_decap_8 FILLER_51_1134 ();
 sg13g2_decap_8 FILLER_51_1141 ();
 sg13g2_decap_8 FILLER_51_1148 ();
 sg13g2_decap_8 FILLER_51_1155 ();
 sg13g2_decap_8 FILLER_51_1162 ();
 sg13g2_decap_8 FILLER_51_1169 ();
 sg13g2_decap_8 FILLER_51_1176 ();
 sg13g2_decap_8 FILLER_51_1183 ();
 sg13g2_decap_8 FILLER_51_1190 ();
 sg13g2_decap_8 FILLER_51_1197 ();
 sg13g2_decap_8 FILLER_51_1204 ();
 sg13g2_decap_8 FILLER_51_1211 ();
 sg13g2_decap_8 FILLER_51_1218 ();
 sg13g2_decap_8 FILLER_51_1225 ();
 sg13g2_decap_8 FILLER_51_1232 ();
 sg13g2_decap_8 FILLER_51_1239 ();
 sg13g2_decap_8 FILLER_51_1246 ();
 sg13g2_decap_8 FILLER_51_1253 ();
 sg13g2_decap_8 FILLER_51_1260 ();
 sg13g2_decap_8 FILLER_51_1267 ();
 sg13g2_decap_8 FILLER_51_1274 ();
 sg13g2_decap_8 FILLER_51_1281 ();
 sg13g2_decap_8 FILLER_51_1288 ();
 sg13g2_decap_8 FILLER_51_1295 ();
 sg13g2_decap_8 FILLER_51_1302 ();
 sg13g2_decap_4 FILLER_51_1309 ();
 sg13g2_fill_2 FILLER_51_1313 ();
 sg13g2_fill_1 FILLER_52_39 ();
 sg13g2_fill_2 FILLER_52_64 ();
 sg13g2_fill_1 FILLER_52_66 ();
 sg13g2_fill_1 FILLER_52_74 ();
 sg13g2_decap_4 FILLER_52_81 ();
 sg13g2_decap_4 FILLER_52_96 ();
 sg13g2_fill_2 FILLER_52_110 ();
 sg13g2_fill_2 FILLER_52_131 ();
 sg13g2_fill_1 FILLER_52_150 ();
 sg13g2_decap_4 FILLER_52_174 ();
 sg13g2_fill_1 FILLER_52_257 ();
 sg13g2_decap_4 FILLER_52_289 ();
 sg13g2_fill_1 FILLER_52_293 ();
 sg13g2_decap_4 FILLER_52_304 ();
 sg13g2_decap_4 FILLER_52_331 ();
 sg13g2_decap_4 FILLER_52_340 ();
 sg13g2_fill_1 FILLER_52_354 ();
 sg13g2_fill_2 FILLER_52_362 ();
 sg13g2_fill_1 FILLER_52_364 ();
 sg13g2_fill_2 FILLER_52_397 ();
 sg13g2_fill_2 FILLER_52_417 ();
 sg13g2_fill_1 FILLER_52_419 ();
 sg13g2_decap_8 FILLER_52_425 ();
 sg13g2_fill_1 FILLER_52_432 ();
 sg13g2_decap_4 FILLER_52_449 ();
 sg13g2_fill_2 FILLER_52_460 ();
 sg13g2_fill_1 FILLER_52_462 ();
 sg13g2_decap_4 FILLER_52_468 ();
 sg13g2_fill_1 FILLER_52_472 ();
 sg13g2_decap_4 FILLER_52_488 ();
 sg13g2_fill_1 FILLER_52_492 ();
 sg13g2_fill_2 FILLER_52_507 ();
 sg13g2_fill_1 FILLER_52_509 ();
 sg13g2_fill_2 FILLER_52_528 ();
 sg13g2_fill_1 FILLER_52_534 ();
 sg13g2_decap_4 FILLER_52_557 ();
 sg13g2_decap_8 FILLER_52_565 ();
 sg13g2_fill_2 FILLER_52_572 ();
 sg13g2_fill_1 FILLER_52_574 ();
 sg13g2_decap_8 FILLER_52_579 ();
 sg13g2_fill_1 FILLER_52_609 ();
 sg13g2_decap_4 FILLER_52_636 ();
 sg13g2_fill_1 FILLER_52_640 ();
 sg13g2_fill_2 FILLER_52_672 ();
 sg13g2_fill_2 FILLER_52_679 ();
 sg13g2_decap_8 FILLER_52_695 ();
 sg13g2_fill_1 FILLER_52_702 ();
 sg13g2_decap_8 FILLER_52_716 ();
 sg13g2_decap_4 FILLER_52_723 ();
 sg13g2_fill_2 FILLER_52_727 ();
 sg13g2_fill_1 FILLER_52_745 ();
 sg13g2_fill_1 FILLER_52_765 ();
 sg13g2_decap_8 FILLER_52_778 ();
 sg13g2_fill_2 FILLER_52_785 ();
 sg13g2_fill_1 FILLER_52_790 ();
 sg13g2_fill_2 FILLER_52_861 ();
 sg13g2_fill_1 FILLER_52_876 ();
 sg13g2_fill_2 FILLER_52_952 ();
 sg13g2_fill_1 FILLER_52_954 ();
 sg13g2_decap_4 FILLER_52_981 ();
 sg13g2_fill_1 FILLER_52_985 ();
 sg13g2_decap_8 FILLER_52_999 ();
 sg13g2_decap_8 FILLER_52_1006 ();
 sg13g2_decap_8 FILLER_52_1013 ();
 sg13g2_decap_8 FILLER_52_1020 ();
 sg13g2_decap_8 FILLER_52_1027 ();
 sg13g2_decap_8 FILLER_52_1034 ();
 sg13g2_decap_8 FILLER_52_1041 ();
 sg13g2_decap_8 FILLER_52_1048 ();
 sg13g2_decap_8 FILLER_52_1055 ();
 sg13g2_decap_8 FILLER_52_1062 ();
 sg13g2_decap_8 FILLER_52_1069 ();
 sg13g2_decap_8 FILLER_52_1076 ();
 sg13g2_decap_8 FILLER_52_1083 ();
 sg13g2_decap_8 FILLER_52_1090 ();
 sg13g2_decap_8 FILLER_52_1097 ();
 sg13g2_decap_8 FILLER_52_1104 ();
 sg13g2_decap_8 FILLER_52_1111 ();
 sg13g2_decap_8 FILLER_52_1118 ();
 sg13g2_decap_8 FILLER_52_1125 ();
 sg13g2_decap_8 FILLER_52_1132 ();
 sg13g2_decap_8 FILLER_52_1139 ();
 sg13g2_decap_8 FILLER_52_1146 ();
 sg13g2_decap_8 FILLER_52_1153 ();
 sg13g2_decap_8 FILLER_52_1160 ();
 sg13g2_decap_8 FILLER_52_1167 ();
 sg13g2_decap_8 FILLER_52_1174 ();
 sg13g2_decap_8 FILLER_52_1181 ();
 sg13g2_decap_8 FILLER_52_1188 ();
 sg13g2_decap_8 FILLER_52_1195 ();
 sg13g2_decap_8 FILLER_52_1202 ();
 sg13g2_decap_8 FILLER_52_1209 ();
 sg13g2_decap_8 FILLER_52_1216 ();
 sg13g2_decap_8 FILLER_52_1223 ();
 sg13g2_decap_8 FILLER_52_1230 ();
 sg13g2_decap_8 FILLER_52_1237 ();
 sg13g2_decap_8 FILLER_52_1244 ();
 sg13g2_decap_8 FILLER_52_1251 ();
 sg13g2_decap_8 FILLER_52_1258 ();
 sg13g2_decap_8 FILLER_52_1265 ();
 sg13g2_decap_8 FILLER_52_1272 ();
 sg13g2_decap_8 FILLER_52_1279 ();
 sg13g2_decap_8 FILLER_52_1286 ();
 sg13g2_decap_8 FILLER_52_1293 ();
 sg13g2_decap_8 FILLER_52_1300 ();
 sg13g2_decap_8 FILLER_52_1307 ();
 sg13g2_fill_1 FILLER_52_1314 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_15 ();
 sg13g2_fill_1 FILLER_53_17 ();
 sg13g2_fill_2 FILLER_53_48 ();
 sg13g2_fill_1 FILLER_53_50 ();
 sg13g2_fill_2 FILLER_53_59 ();
 sg13g2_fill_1 FILLER_53_61 ();
 sg13g2_decap_4 FILLER_53_67 ();
 sg13g2_fill_1 FILLER_53_71 ();
 sg13g2_fill_2 FILLER_53_77 ();
 sg13g2_fill_1 FILLER_53_79 ();
 sg13g2_fill_2 FILLER_53_122 ();
 sg13g2_fill_2 FILLER_53_150 ();
 sg13g2_fill_1 FILLER_53_152 ();
 sg13g2_fill_2 FILLER_53_161 ();
 sg13g2_fill_2 FILLER_53_178 ();
 sg13g2_fill_1 FILLER_53_180 ();
 sg13g2_fill_2 FILLER_53_210 ();
 sg13g2_fill_1 FILLER_53_212 ();
 sg13g2_fill_2 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_224 ();
 sg13g2_fill_1 FILLER_53_252 ();
 sg13g2_decap_8 FILLER_53_277 ();
 sg13g2_decap_4 FILLER_53_284 ();
 sg13g2_fill_1 FILLER_53_288 ();
 sg13g2_fill_1 FILLER_53_337 ();
 sg13g2_decap_4 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_354 ();
 sg13g2_fill_2 FILLER_53_367 ();
 sg13g2_decap_8 FILLER_53_383 ();
 sg13g2_fill_2 FILLER_53_390 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_fill_1 FILLER_53_409 ();
 sg13g2_fill_1 FILLER_53_415 ();
 sg13g2_decap_4 FILLER_53_433 ();
 sg13g2_decap_4 FILLER_53_466 ();
 sg13g2_decap_4 FILLER_53_487 ();
 sg13g2_fill_2 FILLER_53_508 ();
 sg13g2_fill_1 FILLER_53_522 ();
 sg13g2_fill_1 FILLER_53_616 ();
 sg13g2_decap_8 FILLER_53_646 ();
 sg13g2_fill_1 FILLER_53_674 ();
 sg13g2_fill_2 FILLER_53_701 ();
 sg13g2_fill_1 FILLER_53_703 ();
 sg13g2_decap_4 FILLER_53_746 ();
 sg13g2_fill_2 FILLER_53_766 ();
 sg13g2_fill_1 FILLER_53_776 ();
 sg13g2_decap_4 FILLER_53_800 ();
 sg13g2_fill_2 FILLER_53_804 ();
 sg13g2_decap_4 FILLER_53_832 ();
 sg13g2_fill_2 FILLER_53_844 ();
 sg13g2_fill_1 FILLER_53_959 ();
 sg13g2_decap_8 FILLER_53_973 ();
 sg13g2_decap_8 FILLER_53_980 ();
 sg13g2_decap_8 FILLER_53_987 ();
 sg13g2_decap_8 FILLER_53_994 ();
 sg13g2_decap_8 FILLER_53_1001 ();
 sg13g2_decap_8 FILLER_53_1008 ();
 sg13g2_decap_8 FILLER_53_1015 ();
 sg13g2_decap_8 FILLER_53_1022 ();
 sg13g2_decap_8 FILLER_53_1029 ();
 sg13g2_decap_8 FILLER_53_1036 ();
 sg13g2_decap_8 FILLER_53_1043 ();
 sg13g2_decap_8 FILLER_53_1050 ();
 sg13g2_decap_8 FILLER_53_1057 ();
 sg13g2_decap_8 FILLER_53_1064 ();
 sg13g2_decap_8 FILLER_53_1071 ();
 sg13g2_decap_8 FILLER_53_1078 ();
 sg13g2_decap_8 FILLER_53_1085 ();
 sg13g2_decap_8 FILLER_53_1092 ();
 sg13g2_decap_8 FILLER_53_1099 ();
 sg13g2_decap_8 FILLER_53_1106 ();
 sg13g2_decap_8 FILLER_53_1113 ();
 sg13g2_decap_8 FILLER_53_1120 ();
 sg13g2_decap_8 FILLER_53_1127 ();
 sg13g2_decap_8 FILLER_53_1134 ();
 sg13g2_decap_8 FILLER_53_1141 ();
 sg13g2_decap_8 FILLER_53_1148 ();
 sg13g2_decap_8 FILLER_53_1155 ();
 sg13g2_decap_8 FILLER_53_1162 ();
 sg13g2_decap_8 FILLER_53_1169 ();
 sg13g2_decap_8 FILLER_53_1176 ();
 sg13g2_decap_8 FILLER_53_1183 ();
 sg13g2_decap_8 FILLER_53_1190 ();
 sg13g2_decap_8 FILLER_53_1197 ();
 sg13g2_decap_8 FILLER_53_1204 ();
 sg13g2_decap_8 FILLER_53_1211 ();
 sg13g2_decap_8 FILLER_53_1218 ();
 sg13g2_decap_8 FILLER_53_1225 ();
 sg13g2_decap_8 FILLER_53_1232 ();
 sg13g2_decap_8 FILLER_53_1239 ();
 sg13g2_decap_8 FILLER_53_1246 ();
 sg13g2_decap_8 FILLER_53_1253 ();
 sg13g2_decap_8 FILLER_53_1260 ();
 sg13g2_decap_8 FILLER_53_1267 ();
 sg13g2_decap_8 FILLER_53_1274 ();
 sg13g2_decap_8 FILLER_53_1281 ();
 sg13g2_decap_8 FILLER_53_1288 ();
 sg13g2_decap_8 FILLER_53_1295 ();
 sg13g2_decap_8 FILLER_53_1302 ();
 sg13g2_decap_4 FILLER_53_1309 ();
 sg13g2_fill_2 FILLER_53_1313 ();
 sg13g2_fill_2 FILLER_54_31 ();
 sg13g2_decap_4 FILLER_54_56 ();
 sg13g2_fill_2 FILLER_54_65 ();
 sg13g2_fill_2 FILLER_54_83 ();
 sg13g2_decap_8 FILLER_54_97 ();
 sg13g2_fill_2 FILLER_54_111 ();
 sg13g2_decap_4 FILLER_54_118 ();
 sg13g2_decap_8 FILLER_54_189 ();
 sg13g2_fill_2 FILLER_54_196 ();
 sg13g2_fill_1 FILLER_54_198 ();
 sg13g2_fill_1 FILLER_54_203 ();
 sg13g2_fill_2 FILLER_54_231 ();
 sg13g2_fill_1 FILLER_54_271 ();
 sg13g2_fill_2 FILLER_54_298 ();
 sg13g2_decap_8 FILLER_54_304 ();
 sg13g2_fill_2 FILLER_54_311 ();
 sg13g2_fill_1 FILLER_54_313 ();
 sg13g2_decap_4 FILLER_54_361 ();
 sg13g2_fill_1 FILLER_54_365 ();
 sg13g2_fill_1 FILLER_54_376 ();
 sg13g2_fill_2 FILLER_54_390 ();
 sg13g2_fill_1 FILLER_54_397 ();
 sg13g2_fill_2 FILLER_54_403 ();
 sg13g2_decap_4 FILLER_54_410 ();
 sg13g2_fill_2 FILLER_54_414 ();
 sg13g2_decap_4 FILLER_54_426 ();
 sg13g2_decap_4 FILLER_54_435 ();
 sg13g2_fill_2 FILLER_54_447 ();
 sg13g2_fill_1 FILLER_54_449 ();
 sg13g2_fill_2 FILLER_54_458 ();
 sg13g2_fill_2 FILLER_54_472 ();
 sg13g2_fill_1 FILLER_54_474 ();
 sg13g2_decap_8 FILLER_54_482 ();
 sg13g2_decap_4 FILLER_54_489 ();
 sg13g2_fill_1 FILLER_54_509 ();
 sg13g2_fill_1 FILLER_54_513 ();
 sg13g2_fill_1 FILLER_54_524 ();
 sg13g2_fill_2 FILLER_54_540 ();
 sg13g2_fill_1 FILLER_54_542 ();
 sg13g2_fill_2 FILLER_54_589 ();
 sg13g2_fill_1 FILLER_54_591 ();
 sg13g2_fill_1 FILLER_54_613 ();
 sg13g2_decap_8 FILLER_54_657 ();
 sg13g2_decap_8 FILLER_54_664 ();
 sg13g2_fill_2 FILLER_54_671 ();
 sg13g2_fill_1 FILLER_54_673 ();
 sg13g2_decap_8 FILLER_54_682 ();
 sg13g2_fill_1 FILLER_54_694 ();
 sg13g2_decap_4 FILLER_54_703 ();
 sg13g2_fill_1 FILLER_54_707 ();
 sg13g2_fill_2 FILLER_54_718 ();
 sg13g2_fill_1 FILLER_54_720 ();
 sg13g2_decap_4 FILLER_54_730 ();
 sg13g2_fill_1 FILLER_54_734 ();
 sg13g2_fill_2 FILLER_54_739 ();
 sg13g2_decap_4 FILLER_54_751 ();
 sg13g2_decap_4 FILLER_54_763 ();
 sg13g2_fill_1 FILLER_54_767 ();
 sg13g2_decap_8 FILLER_54_778 ();
 sg13g2_fill_2 FILLER_54_785 ();
 sg13g2_fill_1 FILLER_54_787 ();
 sg13g2_fill_2 FILLER_54_793 ();
 sg13g2_fill_1 FILLER_54_821 ();
 sg13g2_fill_1 FILLER_54_919 ();
 sg13g2_fill_2 FILLER_54_967 ();
 sg13g2_decap_8 FILLER_54_978 ();
 sg13g2_decap_8 FILLER_54_985 ();
 sg13g2_decap_8 FILLER_54_992 ();
 sg13g2_decap_8 FILLER_54_999 ();
 sg13g2_decap_8 FILLER_54_1006 ();
 sg13g2_decap_8 FILLER_54_1013 ();
 sg13g2_decap_8 FILLER_54_1020 ();
 sg13g2_decap_8 FILLER_54_1027 ();
 sg13g2_decap_8 FILLER_54_1034 ();
 sg13g2_decap_8 FILLER_54_1041 ();
 sg13g2_decap_8 FILLER_54_1048 ();
 sg13g2_decap_8 FILLER_54_1055 ();
 sg13g2_decap_8 FILLER_54_1062 ();
 sg13g2_decap_8 FILLER_54_1069 ();
 sg13g2_decap_8 FILLER_54_1076 ();
 sg13g2_decap_8 FILLER_54_1083 ();
 sg13g2_decap_8 FILLER_54_1090 ();
 sg13g2_decap_8 FILLER_54_1097 ();
 sg13g2_decap_8 FILLER_54_1104 ();
 sg13g2_decap_8 FILLER_54_1111 ();
 sg13g2_decap_8 FILLER_54_1118 ();
 sg13g2_decap_8 FILLER_54_1125 ();
 sg13g2_decap_8 FILLER_54_1132 ();
 sg13g2_decap_8 FILLER_54_1139 ();
 sg13g2_decap_8 FILLER_54_1146 ();
 sg13g2_decap_8 FILLER_54_1153 ();
 sg13g2_decap_8 FILLER_54_1160 ();
 sg13g2_decap_8 FILLER_54_1167 ();
 sg13g2_decap_8 FILLER_54_1174 ();
 sg13g2_decap_8 FILLER_54_1181 ();
 sg13g2_decap_8 FILLER_54_1188 ();
 sg13g2_decap_8 FILLER_54_1195 ();
 sg13g2_decap_8 FILLER_54_1202 ();
 sg13g2_decap_8 FILLER_54_1209 ();
 sg13g2_decap_8 FILLER_54_1216 ();
 sg13g2_decap_8 FILLER_54_1223 ();
 sg13g2_decap_8 FILLER_54_1230 ();
 sg13g2_decap_8 FILLER_54_1237 ();
 sg13g2_decap_8 FILLER_54_1244 ();
 sg13g2_decap_8 FILLER_54_1251 ();
 sg13g2_decap_8 FILLER_54_1258 ();
 sg13g2_decap_8 FILLER_54_1265 ();
 sg13g2_decap_8 FILLER_54_1272 ();
 sg13g2_decap_8 FILLER_54_1279 ();
 sg13g2_decap_8 FILLER_54_1286 ();
 sg13g2_decap_8 FILLER_54_1293 ();
 sg13g2_decap_8 FILLER_54_1300 ();
 sg13g2_decap_8 FILLER_54_1307 ();
 sg13g2_fill_1 FILLER_54_1314 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_fill_2 FILLER_55_60 ();
 sg13g2_fill_2 FILLER_55_90 ();
 sg13g2_decap_4 FILLER_55_122 ();
 sg13g2_fill_1 FILLER_55_126 ();
 sg13g2_fill_2 FILLER_55_132 ();
 sg13g2_fill_1 FILLER_55_134 ();
 sg13g2_fill_2 FILLER_55_139 ();
 sg13g2_fill_1 FILLER_55_159 ();
 sg13g2_fill_1 FILLER_55_166 ();
 sg13g2_fill_1 FILLER_55_188 ();
 sg13g2_fill_2 FILLER_55_220 ();
 sg13g2_fill_1 FILLER_55_222 ();
 sg13g2_decap_8 FILLER_55_227 ();
 sg13g2_fill_2 FILLER_55_276 ();
 sg13g2_fill_1 FILLER_55_278 ();
 sg13g2_fill_2 FILLER_55_289 ();
 sg13g2_fill_1 FILLER_55_291 ();
 sg13g2_fill_1 FILLER_55_318 ();
 sg13g2_fill_1 FILLER_55_324 ();
 sg13g2_fill_2 FILLER_55_344 ();
 sg13g2_decap_4 FILLER_55_350 ();
 sg13g2_fill_2 FILLER_55_379 ();
 sg13g2_fill_1 FILLER_55_421 ();
 sg13g2_fill_2 FILLER_55_438 ();
 sg13g2_fill_1 FILLER_55_468 ();
 sg13g2_fill_2 FILLER_55_493 ();
 sg13g2_fill_2 FILLER_55_514 ();
 sg13g2_fill_1 FILLER_55_586 ();
 sg13g2_decap_4 FILLER_55_622 ();
 sg13g2_fill_1 FILLER_55_626 ();
 sg13g2_fill_2 FILLER_55_635 ();
 sg13g2_fill_1 FILLER_55_637 ();
 sg13g2_fill_2 FILLER_55_651 ();
 sg13g2_fill_1 FILLER_55_653 ();
 sg13g2_fill_2 FILLER_55_664 ();
 sg13g2_fill_1 FILLER_55_666 ();
 sg13g2_decap_4 FILLER_55_686 ();
 sg13g2_fill_1 FILLER_55_690 ();
 sg13g2_fill_1 FILLER_55_706 ();
 sg13g2_fill_2 FILLER_55_716 ();
 sg13g2_fill_2 FILLER_55_726 ();
 sg13g2_fill_1 FILLER_55_728 ();
 sg13g2_fill_1 FILLER_55_737 ();
 sg13g2_decap_4 FILLER_55_754 ();
 sg13g2_fill_1 FILLER_55_758 ();
 sg13g2_fill_2 FILLER_55_763 ();
 sg13g2_fill_1 FILLER_55_791 ();
 sg13g2_decap_8 FILLER_55_796 ();
 sg13g2_fill_2 FILLER_55_803 ();
 sg13g2_fill_1 FILLER_55_805 ();
 sg13g2_decap_4 FILLER_55_810 ();
 sg13g2_fill_2 FILLER_55_814 ();
 sg13g2_fill_2 FILLER_55_819 ();
 sg13g2_decap_4 FILLER_55_825 ();
 sg13g2_fill_1 FILLER_55_829 ();
 sg13g2_fill_2 FILLER_55_843 ();
 sg13g2_fill_2 FILLER_55_935 ();
 sg13g2_decap_8 FILLER_55_958 ();
 sg13g2_decap_8 FILLER_55_965 ();
 sg13g2_decap_8 FILLER_55_972 ();
 sg13g2_decap_8 FILLER_55_979 ();
 sg13g2_decap_8 FILLER_55_986 ();
 sg13g2_decap_8 FILLER_55_993 ();
 sg13g2_decap_8 FILLER_55_1000 ();
 sg13g2_decap_8 FILLER_55_1007 ();
 sg13g2_decap_8 FILLER_55_1014 ();
 sg13g2_decap_8 FILLER_55_1021 ();
 sg13g2_decap_8 FILLER_55_1028 ();
 sg13g2_decap_8 FILLER_55_1035 ();
 sg13g2_decap_8 FILLER_55_1042 ();
 sg13g2_decap_8 FILLER_55_1049 ();
 sg13g2_decap_8 FILLER_55_1056 ();
 sg13g2_decap_8 FILLER_55_1063 ();
 sg13g2_decap_8 FILLER_55_1070 ();
 sg13g2_decap_8 FILLER_55_1077 ();
 sg13g2_decap_8 FILLER_55_1084 ();
 sg13g2_decap_8 FILLER_55_1091 ();
 sg13g2_decap_8 FILLER_55_1098 ();
 sg13g2_decap_8 FILLER_55_1105 ();
 sg13g2_decap_8 FILLER_55_1112 ();
 sg13g2_decap_8 FILLER_55_1119 ();
 sg13g2_decap_8 FILLER_55_1126 ();
 sg13g2_decap_8 FILLER_55_1133 ();
 sg13g2_decap_8 FILLER_55_1140 ();
 sg13g2_decap_8 FILLER_55_1147 ();
 sg13g2_decap_8 FILLER_55_1154 ();
 sg13g2_decap_8 FILLER_55_1161 ();
 sg13g2_decap_8 FILLER_55_1168 ();
 sg13g2_decap_8 FILLER_55_1175 ();
 sg13g2_decap_8 FILLER_55_1182 ();
 sg13g2_decap_8 FILLER_55_1189 ();
 sg13g2_decap_8 FILLER_55_1196 ();
 sg13g2_decap_8 FILLER_55_1203 ();
 sg13g2_decap_8 FILLER_55_1210 ();
 sg13g2_decap_8 FILLER_55_1217 ();
 sg13g2_decap_8 FILLER_55_1224 ();
 sg13g2_decap_8 FILLER_55_1231 ();
 sg13g2_decap_8 FILLER_55_1238 ();
 sg13g2_decap_8 FILLER_55_1245 ();
 sg13g2_decap_8 FILLER_55_1252 ();
 sg13g2_decap_8 FILLER_55_1259 ();
 sg13g2_decap_8 FILLER_55_1266 ();
 sg13g2_decap_8 FILLER_55_1273 ();
 sg13g2_decap_8 FILLER_55_1280 ();
 sg13g2_decap_8 FILLER_55_1287 ();
 sg13g2_decap_8 FILLER_55_1294 ();
 sg13g2_decap_8 FILLER_55_1301 ();
 sg13g2_decap_8 FILLER_55_1308 ();
 sg13g2_fill_1 FILLER_56_72 ();
 sg13g2_decap_4 FILLER_56_82 ();
 sg13g2_fill_1 FILLER_56_108 ();
 sg13g2_fill_2 FILLER_56_169 ();
 sg13g2_fill_2 FILLER_56_180 ();
 sg13g2_fill_2 FILLER_56_200 ();
 sg13g2_fill_1 FILLER_56_202 ();
 sg13g2_decap_4 FILLER_56_299 ();
 sg13g2_fill_1 FILLER_56_307 ();
 sg13g2_fill_1 FILLER_56_320 ();
 sg13g2_decap_4 FILLER_56_326 ();
 sg13g2_fill_2 FILLER_56_330 ();
 sg13g2_decap_8 FILLER_56_358 ();
 sg13g2_fill_1 FILLER_56_365 ();
 sg13g2_fill_2 FILLER_56_381 ();
 sg13g2_decap_8 FILLER_56_418 ();
 sg13g2_fill_1 FILLER_56_430 ();
 sg13g2_decap_4 FILLER_56_447 ();
 sg13g2_fill_2 FILLER_56_463 ();
 sg13g2_fill_2 FILLER_56_511 ();
 sg13g2_fill_2 FILLER_56_565 ();
 sg13g2_fill_2 FILLER_56_617 ();
 sg13g2_fill_2 FILLER_56_653 ();
 sg13g2_fill_1 FILLER_56_655 ();
 sg13g2_decap_8 FILLER_56_682 ();
 sg13g2_fill_2 FILLER_56_689 ();
 sg13g2_fill_1 FILLER_56_691 ();
 sg13g2_fill_1 FILLER_56_734 ();
 sg13g2_fill_2 FILLER_56_741 ();
 sg13g2_fill_1 FILLER_56_785 ();
 sg13g2_fill_1 FILLER_56_791 ();
 sg13g2_decap_8 FILLER_56_805 ();
 sg13g2_fill_2 FILLER_56_812 ();
 sg13g2_fill_2 FILLER_56_843 ();
 sg13g2_fill_2 FILLER_56_858 ();
 sg13g2_fill_1 FILLER_56_860 ();
 sg13g2_fill_2 FILLER_56_932 ();
 sg13g2_fill_1 FILLER_56_934 ();
 sg13g2_decap_8 FILLER_56_961 ();
 sg13g2_decap_8 FILLER_56_968 ();
 sg13g2_decap_8 FILLER_56_975 ();
 sg13g2_decap_8 FILLER_56_982 ();
 sg13g2_decap_8 FILLER_56_989 ();
 sg13g2_decap_8 FILLER_56_996 ();
 sg13g2_decap_8 FILLER_56_1003 ();
 sg13g2_decap_8 FILLER_56_1010 ();
 sg13g2_decap_8 FILLER_56_1017 ();
 sg13g2_decap_8 FILLER_56_1024 ();
 sg13g2_decap_8 FILLER_56_1031 ();
 sg13g2_decap_8 FILLER_56_1038 ();
 sg13g2_decap_8 FILLER_56_1045 ();
 sg13g2_decap_8 FILLER_56_1052 ();
 sg13g2_decap_8 FILLER_56_1059 ();
 sg13g2_decap_8 FILLER_56_1066 ();
 sg13g2_decap_8 FILLER_56_1073 ();
 sg13g2_decap_8 FILLER_56_1080 ();
 sg13g2_decap_8 FILLER_56_1087 ();
 sg13g2_decap_8 FILLER_56_1094 ();
 sg13g2_decap_8 FILLER_56_1101 ();
 sg13g2_decap_8 FILLER_56_1108 ();
 sg13g2_decap_8 FILLER_56_1115 ();
 sg13g2_decap_8 FILLER_56_1122 ();
 sg13g2_decap_8 FILLER_56_1129 ();
 sg13g2_decap_8 FILLER_56_1136 ();
 sg13g2_decap_8 FILLER_56_1143 ();
 sg13g2_decap_8 FILLER_56_1150 ();
 sg13g2_decap_8 FILLER_56_1157 ();
 sg13g2_decap_8 FILLER_56_1164 ();
 sg13g2_decap_8 FILLER_56_1171 ();
 sg13g2_decap_8 FILLER_56_1178 ();
 sg13g2_decap_8 FILLER_56_1185 ();
 sg13g2_decap_8 FILLER_56_1192 ();
 sg13g2_decap_8 FILLER_56_1199 ();
 sg13g2_decap_8 FILLER_56_1206 ();
 sg13g2_decap_8 FILLER_56_1213 ();
 sg13g2_decap_8 FILLER_56_1220 ();
 sg13g2_decap_8 FILLER_56_1227 ();
 sg13g2_decap_8 FILLER_56_1234 ();
 sg13g2_decap_8 FILLER_56_1241 ();
 sg13g2_decap_8 FILLER_56_1248 ();
 sg13g2_decap_8 FILLER_56_1255 ();
 sg13g2_decap_8 FILLER_56_1262 ();
 sg13g2_decap_8 FILLER_56_1269 ();
 sg13g2_decap_8 FILLER_56_1276 ();
 sg13g2_decap_8 FILLER_56_1283 ();
 sg13g2_decap_8 FILLER_56_1290 ();
 sg13g2_decap_8 FILLER_56_1297 ();
 sg13g2_decap_8 FILLER_56_1304 ();
 sg13g2_decap_4 FILLER_56_1311 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_1 FILLER_57_47 ();
 sg13g2_fill_2 FILLER_57_78 ();
 sg13g2_fill_2 FILLER_57_141 ();
 sg13g2_fill_1 FILLER_57_143 ();
 sg13g2_fill_1 FILLER_57_229 ();
 sg13g2_decap_8 FILLER_57_284 ();
 sg13g2_fill_2 FILLER_57_317 ();
 sg13g2_fill_1 FILLER_57_319 ();
 sg13g2_decap_8 FILLER_57_333 ();
 sg13g2_fill_2 FILLER_57_340 ();
 sg13g2_decap_4 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_fill_2 FILLER_57_506 ();
 sg13g2_fill_1 FILLER_57_508 ();
 sg13g2_fill_1 FILLER_57_555 ();
 sg13g2_fill_2 FILLER_57_561 ();
 sg13g2_fill_1 FILLER_57_563 ();
 sg13g2_fill_2 FILLER_57_635 ();
 sg13g2_fill_1 FILLER_57_637 ();
 sg13g2_fill_2 FILLER_57_643 ();
 sg13g2_decap_8 FILLER_57_657 ();
 sg13g2_decap_4 FILLER_57_664 ();
 sg13g2_fill_1 FILLER_57_668 ();
 sg13g2_fill_2 FILLER_57_701 ();
 sg13g2_fill_1 FILLER_57_703 ();
 sg13g2_fill_2 FILLER_57_723 ();
 sg13g2_fill_1 FILLER_57_725 ();
 sg13g2_fill_2 FILLER_57_735 ();
 sg13g2_fill_1 FILLER_57_748 ();
 sg13g2_decap_4 FILLER_57_765 ();
 sg13g2_fill_2 FILLER_57_774 ();
 sg13g2_fill_1 FILLER_57_776 ();
 sg13g2_decap_8 FILLER_57_782 ();
 sg13g2_decap_4 FILLER_57_789 ();
 sg13g2_fill_2 FILLER_57_797 ();
 sg13g2_fill_1 FILLER_57_799 ();
 sg13g2_fill_2 FILLER_57_826 ();
 sg13g2_decap_4 FILLER_57_832 ();
 sg13g2_fill_1 FILLER_57_836 ();
 sg13g2_fill_1 FILLER_57_889 ();
 sg13g2_fill_2 FILLER_57_950 ();
 sg13g2_decap_8 FILLER_57_961 ();
 sg13g2_decap_8 FILLER_57_968 ();
 sg13g2_decap_8 FILLER_57_975 ();
 sg13g2_decap_8 FILLER_57_982 ();
 sg13g2_decap_8 FILLER_57_989 ();
 sg13g2_decap_8 FILLER_57_996 ();
 sg13g2_decap_8 FILLER_57_1003 ();
 sg13g2_decap_8 FILLER_57_1010 ();
 sg13g2_decap_8 FILLER_57_1017 ();
 sg13g2_decap_8 FILLER_57_1024 ();
 sg13g2_decap_8 FILLER_57_1031 ();
 sg13g2_decap_8 FILLER_57_1038 ();
 sg13g2_decap_8 FILLER_57_1045 ();
 sg13g2_decap_8 FILLER_57_1052 ();
 sg13g2_decap_8 FILLER_57_1059 ();
 sg13g2_decap_8 FILLER_57_1066 ();
 sg13g2_decap_8 FILLER_57_1073 ();
 sg13g2_decap_8 FILLER_57_1080 ();
 sg13g2_decap_8 FILLER_57_1087 ();
 sg13g2_decap_8 FILLER_57_1094 ();
 sg13g2_decap_8 FILLER_57_1101 ();
 sg13g2_decap_8 FILLER_57_1108 ();
 sg13g2_decap_8 FILLER_57_1115 ();
 sg13g2_decap_8 FILLER_57_1122 ();
 sg13g2_decap_8 FILLER_57_1129 ();
 sg13g2_decap_8 FILLER_57_1136 ();
 sg13g2_decap_8 FILLER_57_1143 ();
 sg13g2_decap_8 FILLER_57_1150 ();
 sg13g2_decap_8 FILLER_57_1157 ();
 sg13g2_decap_8 FILLER_57_1164 ();
 sg13g2_decap_8 FILLER_57_1171 ();
 sg13g2_decap_8 FILLER_57_1178 ();
 sg13g2_decap_8 FILLER_57_1185 ();
 sg13g2_decap_8 FILLER_57_1192 ();
 sg13g2_decap_8 FILLER_57_1199 ();
 sg13g2_decap_8 FILLER_57_1206 ();
 sg13g2_decap_8 FILLER_57_1213 ();
 sg13g2_decap_8 FILLER_57_1220 ();
 sg13g2_decap_8 FILLER_57_1227 ();
 sg13g2_decap_8 FILLER_57_1234 ();
 sg13g2_decap_8 FILLER_57_1241 ();
 sg13g2_decap_8 FILLER_57_1248 ();
 sg13g2_decap_8 FILLER_57_1255 ();
 sg13g2_decap_8 FILLER_57_1262 ();
 sg13g2_decap_8 FILLER_57_1269 ();
 sg13g2_decap_8 FILLER_57_1276 ();
 sg13g2_decap_8 FILLER_57_1283 ();
 sg13g2_decap_8 FILLER_57_1290 ();
 sg13g2_decap_8 FILLER_57_1297 ();
 sg13g2_decap_8 FILLER_57_1304 ();
 sg13g2_decap_4 FILLER_57_1311 ();
 sg13g2_fill_2 FILLER_58_69 ();
 sg13g2_fill_1 FILLER_58_71 ();
 sg13g2_fill_1 FILLER_58_85 ();
 sg13g2_decap_4 FILLER_58_90 ();
 sg13g2_fill_1 FILLER_58_110 ();
 sg13g2_fill_1 FILLER_58_127 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_fill_2 FILLER_58_178 ();
 sg13g2_fill_2 FILLER_58_210 ();
 sg13g2_fill_2 FILLER_58_255 ();
 sg13g2_decap_4 FILLER_58_272 ();
 sg13g2_fill_1 FILLER_58_276 ();
 sg13g2_fill_2 FILLER_58_281 ();
 sg13g2_fill_1 FILLER_58_283 ();
 sg13g2_fill_2 FILLER_58_288 ();
 sg13g2_fill_1 FILLER_58_290 ();
 sg13g2_decap_4 FILLER_58_295 ();
 sg13g2_fill_1 FILLER_58_299 ();
 sg13g2_fill_2 FILLER_58_326 ();
 sg13g2_fill_1 FILLER_58_328 ();
 sg13g2_fill_1 FILLER_58_364 ();
 sg13g2_decap_4 FILLER_58_373 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_decap_8 FILLER_58_409 ();
 sg13g2_fill_2 FILLER_58_416 ();
 sg13g2_fill_1 FILLER_58_418 ();
 sg13g2_fill_1 FILLER_58_428 ();
 sg13g2_decap_4 FILLER_58_438 ();
 sg13g2_fill_1 FILLER_58_442 ();
 sg13g2_fill_2 FILLER_58_447 ();
 sg13g2_fill_1 FILLER_58_449 ();
 sg13g2_decap_4 FILLER_58_454 ();
 sg13g2_fill_1 FILLER_58_458 ();
 sg13g2_fill_1 FILLER_58_463 ();
 sg13g2_fill_2 FILLER_58_468 ();
 sg13g2_fill_1 FILLER_58_470 ();
 sg13g2_decap_8 FILLER_58_475 ();
 sg13g2_fill_1 FILLER_58_482 ();
 sg13g2_fill_2 FILLER_58_532 ();
 sg13g2_fill_1 FILLER_58_534 ();
 sg13g2_fill_1 FILLER_58_561 ();
 sg13g2_fill_2 FILLER_58_600 ();
 sg13g2_fill_2 FILLER_58_607 ();
 sg13g2_decap_4 FILLER_58_618 ();
 sg13g2_fill_1 FILLER_58_622 ();
 sg13g2_decap_4 FILLER_58_654 ();
 sg13g2_fill_2 FILLER_58_688 ();
 sg13g2_fill_2 FILLER_58_712 ();
 sg13g2_fill_1 FILLER_58_714 ();
 sg13g2_fill_2 FILLER_58_741 ();
 sg13g2_fill_1 FILLER_58_743 ();
 sg13g2_fill_1 FILLER_58_749 ();
 sg13g2_fill_2 FILLER_58_755 ();
 sg13g2_fill_1 FILLER_58_757 ();
 sg13g2_fill_1 FILLER_58_766 ();
 sg13g2_decap_4 FILLER_58_815 ();
 sg13g2_fill_2 FILLER_58_819 ();
 sg13g2_decap_8 FILLER_58_856 ();
 sg13g2_fill_1 FILLER_58_919 ();
 sg13g2_decap_8 FILLER_58_963 ();
 sg13g2_decap_8 FILLER_58_970 ();
 sg13g2_decap_8 FILLER_58_977 ();
 sg13g2_decap_8 FILLER_58_984 ();
 sg13g2_decap_8 FILLER_58_991 ();
 sg13g2_decap_8 FILLER_58_998 ();
 sg13g2_decap_8 FILLER_58_1005 ();
 sg13g2_decap_8 FILLER_58_1012 ();
 sg13g2_decap_8 FILLER_58_1019 ();
 sg13g2_decap_8 FILLER_58_1026 ();
 sg13g2_decap_8 FILLER_58_1033 ();
 sg13g2_decap_8 FILLER_58_1040 ();
 sg13g2_decap_8 FILLER_58_1047 ();
 sg13g2_decap_8 FILLER_58_1054 ();
 sg13g2_decap_8 FILLER_58_1061 ();
 sg13g2_decap_8 FILLER_58_1068 ();
 sg13g2_decap_8 FILLER_58_1075 ();
 sg13g2_decap_8 FILLER_58_1082 ();
 sg13g2_decap_8 FILLER_58_1089 ();
 sg13g2_decap_8 FILLER_58_1096 ();
 sg13g2_decap_8 FILLER_58_1103 ();
 sg13g2_decap_8 FILLER_58_1110 ();
 sg13g2_decap_8 FILLER_58_1117 ();
 sg13g2_decap_8 FILLER_58_1124 ();
 sg13g2_decap_8 FILLER_58_1131 ();
 sg13g2_decap_8 FILLER_58_1138 ();
 sg13g2_decap_8 FILLER_58_1145 ();
 sg13g2_decap_8 FILLER_58_1152 ();
 sg13g2_decap_8 FILLER_58_1159 ();
 sg13g2_decap_8 FILLER_58_1166 ();
 sg13g2_decap_8 FILLER_58_1173 ();
 sg13g2_decap_8 FILLER_58_1180 ();
 sg13g2_decap_8 FILLER_58_1187 ();
 sg13g2_decap_8 FILLER_58_1194 ();
 sg13g2_decap_8 FILLER_58_1201 ();
 sg13g2_decap_8 FILLER_58_1208 ();
 sg13g2_decap_8 FILLER_58_1215 ();
 sg13g2_decap_8 FILLER_58_1222 ();
 sg13g2_decap_8 FILLER_58_1229 ();
 sg13g2_decap_8 FILLER_58_1236 ();
 sg13g2_decap_8 FILLER_58_1243 ();
 sg13g2_decap_8 FILLER_58_1250 ();
 sg13g2_decap_8 FILLER_58_1257 ();
 sg13g2_decap_8 FILLER_58_1264 ();
 sg13g2_decap_8 FILLER_58_1271 ();
 sg13g2_decap_8 FILLER_58_1278 ();
 sg13g2_decap_8 FILLER_58_1285 ();
 sg13g2_decap_8 FILLER_58_1292 ();
 sg13g2_decap_8 FILLER_58_1299 ();
 sg13g2_decap_8 FILLER_58_1306 ();
 sg13g2_fill_2 FILLER_58_1313 ();
 sg13g2_fill_2 FILLER_59_46 ();
 sg13g2_fill_1 FILLER_59_48 ();
 sg13g2_fill_1 FILLER_59_108 ();
 sg13g2_fill_1 FILLER_59_129 ();
 sg13g2_fill_1 FILLER_59_159 ();
 sg13g2_fill_2 FILLER_59_197 ();
 sg13g2_fill_2 FILLER_59_240 ();
 sg13g2_fill_1 FILLER_59_242 ();
 sg13g2_fill_1 FILLER_59_259 ();
 sg13g2_decap_4 FILLER_59_266 ();
 sg13g2_fill_2 FILLER_59_270 ();
 sg13g2_fill_1 FILLER_59_277 ();
 sg13g2_fill_1 FILLER_59_295 ();
 sg13g2_decap_4 FILLER_59_336 ();
 sg13g2_decap_4 FILLER_59_348 ();
 sg13g2_fill_2 FILLER_59_352 ();
 sg13g2_fill_2 FILLER_59_380 ();
 sg13g2_fill_1 FILLER_59_382 ();
 sg13g2_decap_4 FILLER_59_444 ();
 sg13g2_decap_4 FILLER_59_474 ();
 sg13g2_fill_2 FILLER_59_478 ();
 sg13g2_fill_2 FILLER_59_514 ();
 sg13g2_fill_2 FILLER_59_542 ();
 sg13g2_fill_1 FILLER_59_544 ();
 sg13g2_decap_8 FILLER_59_549 ();
 sg13g2_fill_1 FILLER_59_569 ();
 sg13g2_fill_2 FILLER_59_578 ();
 sg13g2_fill_2 FILLER_59_585 ();
 sg13g2_fill_2 FILLER_59_595 ();
 sg13g2_fill_1 FILLER_59_597 ();
 sg13g2_fill_1 FILLER_59_634 ();
 sg13g2_fill_2 FILLER_59_656 ();
 sg13g2_fill_1 FILLER_59_658 ();
 sg13g2_decap_8 FILLER_59_679 ();
 sg13g2_fill_1 FILLER_59_686 ();
 sg13g2_fill_2 FILLER_59_705 ();
 sg13g2_fill_1 FILLER_59_715 ();
 sg13g2_fill_1 FILLER_59_730 ();
 sg13g2_fill_2 FILLER_59_746 ();
 sg13g2_fill_1 FILLER_59_748 ();
 sg13g2_decap_8 FILLER_59_758 ();
 sg13g2_fill_2 FILLER_59_765 ();
 sg13g2_fill_1 FILLER_59_767 ();
 sg13g2_decap_8 FILLER_59_772 ();
 sg13g2_fill_1 FILLER_59_779 ();
 sg13g2_decap_8 FILLER_59_785 ();
 sg13g2_fill_2 FILLER_59_792 ();
 sg13g2_decap_8 FILLER_59_803 ();
 sg13g2_fill_1 FILLER_59_840 ();
 sg13g2_fill_2 FILLER_59_898 ();
 sg13g2_decap_8 FILLER_59_965 ();
 sg13g2_decap_8 FILLER_59_972 ();
 sg13g2_decap_8 FILLER_59_979 ();
 sg13g2_decap_8 FILLER_59_986 ();
 sg13g2_decap_8 FILLER_59_993 ();
 sg13g2_decap_8 FILLER_59_1000 ();
 sg13g2_decap_8 FILLER_59_1007 ();
 sg13g2_decap_8 FILLER_59_1014 ();
 sg13g2_decap_8 FILLER_59_1021 ();
 sg13g2_decap_8 FILLER_59_1028 ();
 sg13g2_decap_8 FILLER_59_1035 ();
 sg13g2_decap_8 FILLER_59_1042 ();
 sg13g2_decap_8 FILLER_59_1049 ();
 sg13g2_decap_8 FILLER_59_1056 ();
 sg13g2_decap_8 FILLER_59_1063 ();
 sg13g2_decap_8 FILLER_59_1070 ();
 sg13g2_decap_8 FILLER_59_1077 ();
 sg13g2_decap_8 FILLER_59_1084 ();
 sg13g2_decap_8 FILLER_59_1091 ();
 sg13g2_decap_8 FILLER_59_1098 ();
 sg13g2_decap_8 FILLER_59_1105 ();
 sg13g2_decap_8 FILLER_59_1112 ();
 sg13g2_decap_8 FILLER_59_1119 ();
 sg13g2_decap_8 FILLER_59_1126 ();
 sg13g2_decap_8 FILLER_59_1133 ();
 sg13g2_decap_8 FILLER_59_1140 ();
 sg13g2_decap_8 FILLER_59_1147 ();
 sg13g2_decap_8 FILLER_59_1154 ();
 sg13g2_decap_8 FILLER_59_1161 ();
 sg13g2_decap_8 FILLER_59_1168 ();
 sg13g2_decap_8 FILLER_59_1175 ();
 sg13g2_decap_8 FILLER_59_1182 ();
 sg13g2_decap_8 FILLER_59_1189 ();
 sg13g2_decap_8 FILLER_59_1196 ();
 sg13g2_decap_8 FILLER_59_1203 ();
 sg13g2_decap_8 FILLER_59_1210 ();
 sg13g2_decap_8 FILLER_59_1217 ();
 sg13g2_decap_8 FILLER_59_1224 ();
 sg13g2_decap_8 FILLER_59_1231 ();
 sg13g2_decap_8 FILLER_59_1238 ();
 sg13g2_decap_8 FILLER_59_1245 ();
 sg13g2_decap_8 FILLER_59_1252 ();
 sg13g2_decap_8 FILLER_59_1259 ();
 sg13g2_decap_8 FILLER_59_1266 ();
 sg13g2_decap_8 FILLER_59_1273 ();
 sg13g2_decap_8 FILLER_59_1280 ();
 sg13g2_decap_8 FILLER_59_1287 ();
 sg13g2_decap_8 FILLER_59_1294 ();
 sg13g2_decap_8 FILLER_59_1301 ();
 sg13g2_decap_8 FILLER_59_1308 ();
 sg13g2_fill_1 FILLER_60_35 ();
 sg13g2_fill_1 FILLER_60_68 ();
 sg13g2_fill_1 FILLER_60_92 ();
 sg13g2_fill_2 FILLER_60_155 ();
 sg13g2_fill_2 FILLER_60_162 ();
 sg13g2_fill_1 FILLER_60_164 ();
 sg13g2_fill_2 FILLER_60_169 ();
 sg13g2_fill_2 FILLER_60_184 ();
 sg13g2_fill_1 FILLER_60_186 ();
 sg13g2_fill_1 FILLER_60_236 ();
 sg13g2_fill_1 FILLER_60_243 ();
 sg13g2_fill_2 FILLER_60_255 ();
 sg13g2_fill_1 FILLER_60_257 ();
 sg13g2_fill_2 FILLER_60_267 ();
 sg13g2_fill_1 FILLER_60_269 ();
 sg13g2_fill_2 FILLER_60_306 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_2 FILLER_60_417 ();
 sg13g2_fill_1 FILLER_60_454 ();
 sg13g2_fill_2 FILLER_60_525 ();
 sg13g2_decap_8 FILLER_60_534 ();
 sg13g2_fill_2 FILLER_60_541 ();
 sg13g2_decap_4 FILLER_60_547 ();
 sg13g2_fill_1 FILLER_60_551 ();
 sg13g2_fill_1 FILLER_60_578 ();
 sg13g2_decap_8 FILLER_60_608 ();
 sg13g2_fill_2 FILLER_60_615 ();
 sg13g2_fill_1 FILLER_60_617 ();
 sg13g2_fill_1 FILLER_60_631 ();
 sg13g2_fill_2 FILLER_60_698 ();
 sg13g2_decap_4 FILLER_60_733 ();
 sg13g2_fill_2 FILLER_60_737 ();
 sg13g2_decap_4 FILLER_60_763 ();
 sg13g2_fill_1 FILLER_60_771 ();
 sg13g2_fill_2 FILLER_60_780 ();
 sg13g2_decap_4 FILLER_60_825 ();
 sg13g2_decap_8 FILLER_60_832 ();
 sg13g2_decap_4 FILLER_60_839 ();
 sg13g2_fill_1 FILLER_60_843 ();
 sg13g2_decap_8 FILLER_60_857 ();
 sg13g2_fill_2 FILLER_60_864 ();
 sg13g2_fill_1 FILLER_60_866 ();
 sg13g2_fill_2 FILLER_60_880 ();
 sg13g2_fill_2 FILLER_60_900 ();
 sg13g2_fill_1 FILLER_60_902 ();
 sg13g2_decap_4 FILLER_60_920 ();
 sg13g2_fill_2 FILLER_60_924 ();
 sg13g2_decap_8 FILLER_60_935 ();
 sg13g2_decap_8 FILLER_60_942 ();
 sg13g2_decap_8 FILLER_60_949 ();
 sg13g2_decap_8 FILLER_60_956 ();
 sg13g2_decap_8 FILLER_60_963 ();
 sg13g2_decap_8 FILLER_60_970 ();
 sg13g2_decap_8 FILLER_60_977 ();
 sg13g2_decap_8 FILLER_60_984 ();
 sg13g2_decap_8 FILLER_60_991 ();
 sg13g2_decap_8 FILLER_60_998 ();
 sg13g2_decap_8 FILLER_60_1005 ();
 sg13g2_decap_8 FILLER_60_1012 ();
 sg13g2_decap_8 FILLER_60_1019 ();
 sg13g2_decap_8 FILLER_60_1026 ();
 sg13g2_decap_8 FILLER_60_1033 ();
 sg13g2_decap_8 FILLER_60_1040 ();
 sg13g2_decap_8 FILLER_60_1047 ();
 sg13g2_decap_8 FILLER_60_1054 ();
 sg13g2_decap_8 FILLER_60_1061 ();
 sg13g2_decap_8 FILLER_60_1068 ();
 sg13g2_decap_8 FILLER_60_1075 ();
 sg13g2_decap_8 FILLER_60_1082 ();
 sg13g2_decap_8 FILLER_60_1089 ();
 sg13g2_decap_8 FILLER_60_1096 ();
 sg13g2_decap_8 FILLER_60_1103 ();
 sg13g2_decap_8 FILLER_60_1110 ();
 sg13g2_decap_8 FILLER_60_1117 ();
 sg13g2_decap_8 FILLER_60_1124 ();
 sg13g2_decap_8 FILLER_60_1131 ();
 sg13g2_decap_8 FILLER_60_1138 ();
 sg13g2_decap_8 FILLER_60_1145 ();
 sg13g2_decap_8 FILLER_60_1152 ();
 sg13g2_decap_8 FILLER_60_1159 ();
 sg13g2_decap_8 FILLER_60_1166 ();
 sg13g2_decap_8 FILLER_60_1173 ();
 sg13g2_decap_8 FILLER_60_1180 ();
 sg13g2_decap_8 FILLER_60_1187 ();
 sg13g2_decap_8 FILLER_60_1194 ();
 sg13g2_decap_8 FILLER_60_1201 ();
 sg13g2_decap_8 FILLER_60_1208 ();
 sg13g2_decap_8 FILLER_60_1215 ();
 sg13g2_decap_8 FILLER_60_1222 ();
 sg13g2_decap_8 FILLER_60_1229 ();
 sg13g2_decap_8 FILLER_60_1236 ();
 sg13g2_decap_8 FILLER_60_1243 ();
 sg13g2_decap_8 FILLER_60_1250 ();
 sg13g2_decap_8 FILLER_60_1257 ();
 sg13g2_decap_8 FILLER_60_1264 ();
 sg13g2_decap_8 FILLER_60_1271 ();
 sg13g2_decap_8 FILLER_60_1278 ();
 sg13g2_decap_8 FILLER_60_1285 ();
 sg13g2_decap_8 FILLER_60_1292 ();
 sg13g2_decap_8 FILLER_60_1299 ();
 sg13g2_decap_8 FILLER_60_1306 ();
 sg13g2_fill_2 FILLER_60_1313 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_29 ();
 sg13g2_fill_1 FILLER_61_85 ();
 sg13g2_fill_1 FILLER_61_118 ();
 sg13g2_fill_1 FILLER_61_129 ();
 sg13g2_fill_2 FILLER_61_133 ();
 sg13g2_fill_1 FILLER_61_244 ();
 sg13g2_fill_2 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_262 ();
 sg13g2_fill_2 FILLER_61_280 ();
 sg13g2_fill_1 FILLER_61_282 ();
 sg13g2_fill_1 FILLER_61_345 ();
 sg13g2_fill_2 FILLER_61_363 ();
 sg13g2_fill_2 FILLER_61_374 ();
 sg13g2_fill_1 FILLER_61_376 ();
 sg13g2_fill_1 FILLER_61_386 ();
 sg13g2_fill_1 FILLER_61_402 ();
 sg13g2_fill_2 FILLER_61_416 ();
 sg13g2_fill_1 FILLER_61_418 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_fill_1 FILLER_61_442 ();
 sg13g2_fill_1 FILLER_61_498 ();
 sg13g2_fill_2 FILLER_61_521 ();
 sg13g2_fill_2 FILLER_61_564 ();
 sg13g2_fill_1 FILLER_61_566 ();
 sg13g2_fill_2 FILLER_61_575 ();
 sg13g2_decap_4 FILLER_61_585 ();
 sg13g2_decap_8 FILLER_61_633 ();
 sg13g2_decap_8 FILLER_61_640 ();
 sg13g2_decap_8 FILLER_61_647 ();
 sg13g2_fill_2 FILLER_61_654 ();
 sg13g2_fill_2 FILLER_61_672 ();
 sg13g2_decap_8 FILLER_61_678 ();
 sg13g2_decap_4 FILLER_61_685 ();
 sg13g2_fill_2 FILLER_61_689 ();
 sg13g2_decap_4 FILLER_61_742 ();
 sg13g2_fill_2 FILLER_61_746 ();
 sg13g2_fill_2 FILLER_61_753 ();
 sg13g2_fill_1 FILLER_61_755 ();
 sg13g2_fill_2 FILLER_61_772 ();
 sg13g2_decap_8 FILLER_61_804 ();
 sg13g2_fill_1 FILLER_61_811 ();
 sg13g2_decap_8 FILLER_61_820 ();
 sg13g2_fill_1 FILLER_61_827 ();
 sg13g2_decap_4 FILLER_61_832 ();
 sg13g2_fill_1 FILLER_61_836 ();
 sg13g2_decap_8 FILLER_61_840 ();
 sg13g2_decap_8 FILLER_61_847 ();
 sg13g2_decap_8 FILLER_61_854 ();
 sg13g2_decap_8 FILLER_61_861 ();
 sg13g2_fill_2 FILLER_61_868 ();
 sg13g2_fill_1 FILLER_61_870 ();
 sg13g2_decap_8 FILLER_61_875 ();
 sg13g2_decap_8 FILLER_61_882 ();
 sg13g2_fill_2 FILLER_61_889 ();
 sg13g2_decap_8 FILLER_61_895 ();
 sg13g2_decap_8 FILLER_61_902 ();
 sg13g2_decap_8 FILLER_61_909 ();
 sg13g2_decap_8 FILLER_61_916 ();
 sg13g2_decap_8 FILLER_61_923 ();
 sg13g2_decap_8 FILLER_61_930 ();
 sg13g2_decap_8 FILLER_61_937 ();
 sg13g2_decap_8 FILLER_61_944 ();
 sg13g2_decap_8 FILLER_61_951 ();
 sg13g2_decap_8 FILLER_61_958 ();
 sg13g2_decap_8 FILLER_61_965 ();
 sg13g2_decap_8 FILLER_61_972 ();
 sg13g2_decap_8 FILLER_61_979 ();
 sg13g2_decap_8 FILLER_61_986 ();
 sg13g2_decap_8 FILLER_61_993 ();
 sg13g2_decap_8 FILLER_61_1000 ();
 sg13g2_decap_8 FILLER_61_1007 ();
 sg13g2_decap_8 FILLER_61_1014 ();
 sg13g2_decap_8 FILLER_61_1021 ();
 sg13g2_decap_8 FILLER_61_1028 ();
 sg13g2_decap_8 FILLER_61_1035 ();
 sg13g2_decap_8 FILLER_61_1042 ();
 sg13g2_decap_8 FILLER_61_1049 ();
 sg13g2_decap_8 FILLER_61_1056 ();
 sg13g2_decap_8 FILLER_61_1063 ();
 sg13g2_decap_8 FILLER_61_1070 ();
 sg13g2_decap_8 FILLER_61_1077 ();
 sg13g2_decap_8 FILLER_61_1084 ();
 sg13g2_decap_8 FILLER_61_1091 ();
 sg13g2_decap_8 FILLER_61_1098 ();
 sg13g2_decap_8 FILLER_61_1105 ();
 sg13g2_decap_8 FILLER_61_1112 ();
 sg13g2_decap_8 FILLER_61_1119 ();
 sg13g2_decap_8 FILLER_61_1126 ();
 sg13g2_decap_8 FILLER_61_1133 ();
 sg13g2_decap_8 FILLER_61_1140 ();
 sg13g2_decap_8 FILLER_61_1147 ();
 sg13g2_decap_8 FILLER_61_1154 ();
 sg13g2_decap_8 FILLER_61_1161 ();
 sg13g2_decap_8 FILLER_61_1168 ();
 sg13g2_decap_8 FILLER_61_1175 ();
 sg13g2_decap_8 FILLER_61_1182 ();
 sg13g2_decap_8 FILLER_61_1189 ();
 sg13g2_decap_8 FILLER_61_1196 ();
 sg13g2_decap_8 FILLER_61_1203 ();
 sg13g2_decap_8 FILLER_61_1210 ();
 sg13g2_decap_8 FILLER_61_1217 ();
 sg13g2_decap_8 FILLER_61_1224 ();
 sg13g2_decap_8 FILLER_61_1231 ();
 sg13g2_decap_8 FILLER_61_1238 ();
 sg13g2_decap_8 FILLER_61_1245 ();
 sg13g2_decap_8 FILLER_61_1252 ();
 sg13g2_decap_8 FILLER_61_1259 ();
 sg13g2_decap_8 FILLER_61_1266 ();
 sg13g2_decap_8 FILLER_61_1273 ();
 sg13g2_decap_8 FILLER_61_1280 ();
 sg13g2_decap_8 FILLER_61_1287 ();
 sg13g2_decap_8 FILLER_61_1294 ();
 sg13g2_decap_8 FILLER_61_1301 ();
 sg13g2_decap_8 FILLER_61_1308 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_2 FILLER_62_27 ();
 sg13g2_fill_1 FILLER_62_29 ();
 sg13g2_fill_2 FILLER_62_38 ();
 sg13g2_fill_1 FILLER_62_40 ();
 sg13g2_fill_1 FILLER_62_53 ();
 sg13g2_fill_2 FILLER_62_68 ();
 sg13g2_fill_1 FILLER_62_70 ();
 sg13g2_fill_2 FILLER_62_103 ();
 sg13g2_fill_2 FILLER_62_115 ();
 sg13g2_fill_2 FILLER_62_192 ();
 sg13g2_fill_2 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_210 ();
 sg13g2_fill_2 FILLER_62_233 ();
 sg13g2_fill_1 FILLER_62_235 ();
 sg13g2_fill_2 FILLER_62_241 ();
 sg13g2_fill_2 FILLER_62_259 ();
 sg13g2_decap_8 FILLER_62_274 ();
 sg13g2_fill_1 FILLER_62_286 ();
 sg13g2_decap_4 FILLER_62_293 ();
 sg13g2_fill_1 FILLER_62_297 ();
 sg13g2_decap_8 FILLER_62_302 ();
 sg13g2_decap_4 FILLER_62_309 ();
 sg13g2_fill_1 FILLER_62_313 ();
 sg13g2_fill_2 FILLER_62_381 ();
 sg13g2_fill_1 FILLER_62_383 ();
 sg13g2_fill_1 FILLER_62_483 ();
 sg13g2_fill_2 FILLER_62_516 ();
 sg13g2_decap_8 FILLER_62_566 ();
 sg13g2_fill_2 FILLER_62_573 ();
 sg13g2_fill_1 FILLER_62_575 ();
 sg13g2_fill_2 FILLER_62_631 ();
 sg13g2_fill_1 FILLER_62_633 ();
 sg13g2_decap_8 FILLER_62_655 ();
 sg13g2_fill_2 FILLER_62_662 ();
 sg13g2_fill_2 FILLER_62_678 ();
 sg13g2_fill_1 FILLER_62_680 ();
 sg13g2_fill_2 FILLER_62_686 ();
 sg13g2_fill_2 FILLER_62_701 ();
 sg13g2_fill_1 FILLER_62_744 ();
 sg13g2_fill_1 FILLER_62_749 ();
 sg13g2_fill_2 FILLER_62_763 ();
 sg13g2_fill_1 FILLER_62_765 ();
 sg13g2_fill_2 FILLER_62_780 ();
 sg13g2_fill_1 FILLER_62_782 ();
 sg13g2_fill_2 FILLER_62_788 ();
 sg13g2_fill_1 FILLER_62_790 ();
 sg13g2_fill_2 FILLER_62_799 ();
 sg13g2_fill_1 FILLER_62_801 ();
 sg13g2_decap_8 FILLER_62_810 ();
 sg13g2_decap_8 FILLER_62_843 ();
 sg13g2_decap_8 FILLER_62_850 ();
 sg13g2_decap_8 FILLER_62_857 ();
 sg13g2_decap_8 FILLER_62_864 ();
 sg13g2_decap_8 FILLER_62_871 ();
 sg13g2_decap_8 FILLER_62_878 ();
 sg13g2_decap_8 FILLER_62_885 ();
 sg13g2_decap_8 FILLER_62_892 ();
 sg13g2_decap_8 FILLER_62_899 ();
 sg13g2_decap_8 FILLER_62_906 ();
 sg13g2_decap_8 FILLER_62_913 ();
 sg13g2_decap_8 FILLER_62_920 ();
 sg13g2_decap_8 FILLER_62_927 ();
 sg13g2_decap_8 FILLER_62_934 ();
 sg13g2_decap_8 FILLER_62_941 ();
 sg13g2_decap_8 FILLER_62_948 ();
 sg13g2_decap_8 FILLER_62_955 ();
 sg13g2_decap_8 FILLER_62_962 ();
 sg13g2_decap_8 FILLER_62_969 ();
 sg13g2_decap_8 FILLER_62_976 ();
 sg13g2_decap_8 FILLER_62_983 ();
 sg13g2_decap_8 FILLER_62_990 ();
 sg13g2_decap_8 FILLER_62_997 ();
 sg13g2_decap_8 FILLER_62_1004 ();
 sg13g2_decap_8 FILLER_62_1011 ();
 sg13g2_decap_8 FILLER_62_1018 ();
 sg13g2_decap_8 FILLER_62_1025 ();
 sg13g2_decap_8 FILLER_62_1032 ();
 sg13g2_decap_8 FILLER_62_1039 ();
 sg13g2_decap_8 FILLER_62_1046 ();
 sg13g2_decap_8 FILLER_62_1053 ();
 sg13g2_decap_8 FILLER_62_1060 ();
 sg13g2_decap_8 FILLER_62_1067 ();
 sg13g2_decap_8 FILLER_62_1074 ();
 sg13g2_decap_8 FILLER_62_1081 ();
 sg13g2_decap_8 FILLER_62_1088 ();
 sg13g2_decap_8 FILLER_62_1095 ();
 sg13g2_decap_8 FILLER_62_1102 ();
 sg13g2_decap_8 FILLER_62_1109 ();
 sg13g2_decap_8 FILLER_62_1116 ();
 sg13g2_decap_8 FILLER_62_1123 ();
 sg13g2_decap_8 FILLER_62_1130 ();
 sg13g2_decap_8 FILLER_62_1137 ();
 sg13g2_decap_8 FILLER_62_1144 ();
 sg13g2_decap_8 FILLER_62_1151 ();
 sg13g2_decap_8 FILLER_62_1158 ();
 sg13g2_decap_8 FILLER_62_1165 ();
 sg13g2_decap_8 FILLER_62_1172 ();
 sg13g2_decap_8 FILLER_62_1179 ();
 sg13g2_decap_8 FILLER_62_1186 ();
 sg13g2_decap_8 FILLER_62_1193 ();
 sg13g2_decap_8 FILLER_62_1200 ();
 sg13g2_decap_8 FILLER_62_1207 ();
 sg13g2_decap_8 FILLER_62_1214 ();
 sg13g2_decap_8 FILLER_62_1221 ();
 sg13g2_decap_8 FILLER_62_1228 ();
 sg13g2_decap_8 FILLER_62_1235 ();
 sg13g2_decap_8 FILLER_62_1242 ();
 sg13g2_decap_8 FILLER_62_1249 ();
 sg13g2_decap_8 FILLER_62_1256 ();
 sg13g2_decap_8 FILLER_62_1263 ();
 sg13g2_decap_8 FILLER_62_1270 ();
 sg13g2_decap_8 FILLER_62_1277 ();
 sg13g2_decap_8 FILLER_62_1284 ();
 sg13g2_decap_8 FILLER_62_1291 ();
 sg13g2_decap_8 FILLER_62_1298 ();
 sg13g2_decap_8 FILLER_62_1305 ();
 sg13g2_fill_2 FILLER_62_1312 ();
 sg13g2_fill_1 FILLER_62_1314 ();
 sg13g2_fill_1 FILLER_63_41 ();
 sg13g2_fill_1 FILLER_63_50 ();
 sg13g2_fill_1 FILLER_63_96 ();
 sg13g2_fill_2 FILLER_63_102 ();
 sg13g2_fill_2 FILLER_63_128 ();
 sg13g2_fill_1 FILLER_63_135 ();
 sg13g2_fill_2 FILLER_63_197 ();
 sg13g2_fill_1 FILLER_63_199 ();
 sg13g2_decap_4 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_263 ();
 sg13g2_decap_4 FILLER_63_270 ();
 sg13g2_fill_2 FILLER_63_274 ();
 sg13g2_fill_1 FILLER_63_285 ();
 sg13g2_fill_1 FILLER_63_291 ();
 sg13g2_fill_2 FILLER_63_361 ();
 sg13g2_fill_2 FILLER_63_375 ();
 sg13g2_fill_1 FILLER_63_432 ();
 sg13g2_fill_2 FILLER_63_463 ();
 sg13g2_fill_1 FILLER_63_534 ();
 sg13g2_decap_4 FILLER_63_545 ();
 sg13g2_decap_4 FILLER_63_562 ();
 sg13g2_decap_4 FILLER_63_582 ();
 sg13g2_decap_4 FILLER_63_630 ();
 sg13g2_fill_2 FILLER_63_655 ();
 sg13g2_fill_1 FILLER_63_657 ();
 sg13g2_decap_4 FILLER_63_661 ();
 sg13g2_fill_1 FILLER_63_665 ();
 sg13g2_decap_8 FILLER_63_696 ();
 sg13g2_decap_8 FILLER_63_703 ();
 sg13g2_fill_2 FILLER_63_710 ();
 sg13g2_fill_2 FILLER_63_748 ();
 sg13g2_fill_1 FILLER_63_750 ();
 sg13g2_fill_1 FILLER_63_755 ();
 sg13g2_fill_1 FILLER_63_760 ();
 sg13g2_fill_1 FILLER_63_773 ();
 sg13g2_fill_2 FILLER_63_808 ();
 sg13g2_fill_1 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_825 ();
 sg13g2_decap_8 FILLER_63_832 ();
 sg13g2_fill_2 FILLER_63_839 ();
 sg13g2_fill_1 FILLER_63_841 ();
 sg13g2_decap_8 FILLER_63_845 ();
 sg13g2_decap_8 FILLER_63_852 ();
 sg13g2_decap_8 FILLER_63_859 ();
 sg13g2_decap_8 FILLER_63_866 ();
 sg13g2_decap_8 FILLER_63_873 ();
 sg13g2_decap_8 FILLER_63_880 ();
 sg13g2_decap_8 FILLER_63_887 ();
 sg13g2_decap_8 FILLER_63_894 ();
 sg13g2_decap_8 FILLER_63_901 ();
 sg13g2_decap_8 FILLER_63_908 ();
 sg13g2_decap_8 FILLER_63_915 ();
 sg13g2_decap_8 FILLER_63_922 ();
 sg13g2_decap_8 FILLER_63_929 ();
 sg13g2_decap_8 FILLER_63_936 ();
 sg13g2_decap_8 FILLER_63_943 ();
 sg13g2_decap_8 FILLER_63_950 ();
 sg13g2_decap_8 FILLER_63_957 ();
 sg13g2_decap_8 FILLER_63_964 ();
 sg13g2_decap_8 FILLER_63_971 ();
 sg13g2_decap_8 FILLER_63_978 ();
 sg13g2_decap_8 FILLER_63_985 ();
 sg13g2_decap_8 FILLER_63_992 ();
 sg13g2_decap_8 FILLER_63_999 ();
 sg13g2_decap_8 FILLER_63_1006 ();
 sg13g2_decap_8 FILLER_63_1013 ();
 sg13g2_decap_8 FILLER_63_1020 ();
 sg13g2_decap_8 FILLER_63_1027 ();
 sg13g2_decap_8 FILLER_63_1034 ();
 sg13g2_decap_8 FILLER_63_1041 ();
 sg13g2_decap_8 FILLER_63_1048 ();
 sg13g2_decap_8 FILLER_63_1055 ();
 sg13g2_decap_8 FILLER_63_1062 ();
 sg13g2_decap_8 FILLER_63_1069 ();
 sg13g2_decap_8 FILLER_63_1076 ();
 sg13g2_decap_8 FILLER_63_1083 ();
 sg13g2_decap_8 FILLER_63_1090 ();
 sg13g2_decap_8 FILLER_63_1097 ();
 sg13g2_decap_8 FILLER_63_1104 ();
 sg13g2_decap_8 FILLER_63_1111 ();
 sg13g2_decap_8 FILLER_63_1118 ();
 sg13g2_decap_8 FILLER_63_1125 ();
 sg13g2_decap_8 FILLER_63_1132 ();
 sg13g2_decap_8 FILLER_63_1139 ();
 sg13g2_decap_8 FILLER_63_1146 ();
 sg13g2_decap_8 FILLER_63_1153 ();
 sg13g2_decap_8 FILLER_63_1160 ();
 sg13g2_decap_8 FILLER_63_1167 ();
 sg13g2_decap_8 FILLER_63_1174 ();
 sg13g2_decap_8 FILLER_63_1181 ();
 sg13g2_decap_8 FILLER_63_1188 ();
 sg13g2_decap_8 FILLER_63_1195 ();
 sg13g2_decap_8 FILLER_63_1202 ();
 sg13g2_decap_8 FILLER_63_1209 ();
 sg13g2_decap_8 FILLER_63_1216 ();
 sg13g2_decap_8 FILLER_63_1223 ();
 sg13g2_decap_8 FILLER_63_1230 ();
 sg13g2_decap_8 FILLER_63_1237 ();
 sg13g2_decap_8 FILLER_63_1244 ();
 sg13g2_decap_8 FILLER_63_1251 ();
 sg13g2_decap_8 FILLER_63_1258 ();
 sg13g2_decap_8 FILLER_63_1265 ();
 sg13g2_decap_8 FILLER_63_1272 ();
 sg13g2_decap_8 FILLER_63_1279 ();
 sg13g2_decap_8 FILLER_63_1286 ();
 sg13g2_decap_8 FILLER_63_1293 ();
 sg13g2_decap_8 FILLER_63_1300 ();
 sg13g2_decap_8 FILLER_63_1307 ();
 sg13g2_fill_1 FILLER_63_1314 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_45 ();
 sg13g2_fill_1 FILLER_64_47 ();
 sg13g2_fill_1 FILLER_64_63 ();
 sg13g2_fill_2 FILLER_64_112 ();
 sg13g2_fill_1 FILLER_64_145 ();
 sg13g2_fill_1 FILLER_64_155 ();
 sg13g2_fill_2 FILLER_64_165 ();
 sg13g2_fill_1 FILLER_64_167 ();
 sg13g2_decap_4 FILLER_64_234 ();
 sg13g2_fill_2 FILLER_64_238 ();
 sg13g2_fill_1 FILLER_64_261 ();
 sg13g2_fill_1 FILLER_64_286 ();
 sg13g2_fill_1 FILLER_64_306 ();
 sg13g2_decap_8 FILLER_64_359 ();
 sg13g2_fill_1 FILLER_64_384 ();
 sg13g2_fill_2 FILLER_64_417 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_fill_1 FILLER_64_470 ();
 sg13g2_fill_1 FILLER_64_508 ();
 sg13g2_fill_1 FILLER_64_522 ();
 sg13g2_fill_2 FILLER_64_531 ();
 sg13g2_fill_1 FILLER_64_569 ();
 sg13g2_fill_2 FILLER_64_575 ();
 sg13g2_decap_8 FILLER_64_597 ();
 sg13g2_decap_8 FILLER_64_604 ();
 sg13g2_decap_4 FILLER_64_611 ();
 sg13g2_decap_8 FILLER_64_619 ();
 sg13g2_decap_4 FILLER_64_626 ();
 sg13g2_fill_2 FILLER_64_651 ();
 sg13g2_fill_1 FILLER_64_653 ();
 sg13g2_fill_2 FILLER_64_662 ();
 sg13g2_fill_1 FILLER_64_664 ();
 sg13g2_fill_1 FILLER_64_674 ();
 sg13g2_decap_4 FILLER_64_679 ();
 sg13g2_fill_1 FILLER_64_683 ();
 sg13g2_decap_4 FILLER_64_702 ();
 sg13g2_fill_1 FILLER_64_706 ();
 sg13g2_fill_2 FILLER_64_717 ();
 sg13g2_fill_1 FILLER_64_719 ();
 sg13g2_fill_1 FILLER_64_733 ();
 sg13g2_fill_1 FILLER_64_743 ();
 sg13g2_fill_2 FILLER_64_757 ();
 sg13g2_fill_1 FILLER_64_759 ();
 sg13g2_fill_2 FILLER_64_783 ();
 sg13g2_fill_2 FILLER_64_803 ();
 sg13g2_fill_1 FILLER_64_821 ();
 sg13g2_decap_8 FILLER_64_848 ();
 sg13g2_decap_8 FILLER_64_855 ();
 sg13g2_decap_8 FILLER_64_862 ();
 sg13g2_decap_8 FILLER_64_869 ();
 sg13g2_decap_8 FILLER_64_876 ();
 sg13g2_decap_8 FILLER_64_883 ();
 sg13g2_decap_8 FILLER_64_890 ();
 sg13g2_decap_8 FILLER_64_897 ();
 sg13g2_decap_8 FILLER_64_904 ();
 sg13g2_decap_8 FILLER_64_911 ();
 sg13g2_decap_8 FILLER_64_918 ();
 sg13g2_decap_8 FILLER_64_925 ();
 sg13g2_decap_8 FILLER_64_932 ();
 sg13g2_decap_8 FILLER_64_939 ();
 sg13g2_decap_8 FILLER_64_946 ();
 sg13g2_decap_8 FILLER_64_953 ();
 sg13g2_decap_8 FILLER_64_960 ();
 sg13g2_decap_8 FILLER_64_967 ();
 sg13g2_decap_8 FILLER_64_974 ();
 sg13g2_decap_8 FILLER_64_981 ();
 sg13g2_decap_8 FILLER_64_988 ();
 sg13g2_decap_8 FILLER_64_995 ();
 sg13g2_decap_8 FILLER_64_1002 ();
 sg13g2_decap_8 FILLER_64_1009 ();
 sg13g2_decap_8 FILLER_64_1016 ();
 sg13g2_decap_8 FILLER_64_1023 ();
 sg13g2_decap_8 FILLER_64_1030 ();
 sg13g2_decap_8 FILLER_64_1037 ();
 sg13g2_decap_8 FILLER_64_1044 ();
 sg13g2_decap_8 FILLER_64_1051 ();
 sg13g2_decap_8 FILLER_64_1058 ();
 sg13g2_decap_8 FILLER_64_1065 ();
 sg13g2_decap_8 FILLER_64_1072 ();
 sg13g2_decap_8 FILLER_64_1079 ();
 sg13g2_decap_8 FILLER_64_1086 ();
 sg13g2_decap_8 FILLER_64_1093 ();
 sg13g2_decap_8 FILLER_64_1100 ();
 sg13g2_decap_8 FILLER_64_1107 ();
 sg13g2_decap_8 FILLER_64_1114 ();
 sg13g2_decap_8 FILLER_64_1121 ();
 sg13g2_decap_8 FILLER_64_1128 ();
 sg13g2_decap_8 FILLER_64_1135 ();
 sg13g2_decap_8 FILLER_64_1142 ();
 sg13g2_decap_8 FILLER_64_1149 ();
 sg13g2_decap_8 FILLER_64_1156 ();
 sg13g2_decap_8 FILLER_64_1163 ();
 sg13g2_decap_8 FILLER_64_1170 ();
 sg13g2_decap_8 FILLER_64_1177 ();
 sg13g2_decap_8 FILLER_64_1184 ();
 sg13g2_decap_8 FILLER_64_1191 ();
 sg13g2_decap_8 FILLER_64_1198 ();
 sg13g2_decap_8 FILLER_64_1205 ();
 sg13g2_decap_8 FILLER_64_1212 ();
 sg13g2_decap_8 FILLER_64_1219 ();
 sg13g2_decap_8 FILLER_64_1226 ();
 sg13g2_decap_8 FILLER_64_1233 ();
 sg13g2_decap_8 FILLER_64_1240 ();
 sg13g2_decap_8 FILLER_64_1247 ();
 sg13g2_decap_8 FILLER_64_1254 ();
 sg13g2_decap_8 FILLER_64_1261 ();
 sg13g2_decap_8 FILLER_64_1268 ();
 sg13g2_decap_8 FILLER_64_1275 ();
 sg13g2_decap_8 FILLER_64_1282 ();
 sg13g2_decap_8 FILLER_64_1289 ();
 sg13g2_decap_8 FILLER_64_1296 ();
 sg13g2_decap_8 FILLER_64_1303 ();
 sg13g2_decap_4 FILLER_64_1310 ();
 sg13g2_fill_1 FILLER_64_1314 ();
 sg13g2_fill_1 FILLER_65_26 ();
 sg13g2_fill_2 FILLER_65_36 ();
 sg13g2_fill_1 FILLER_65_38 ();
 sg13g2_fill_1 FILLER_65_46 ();
 sg13g2_fill_1 FILLER_65_73 ();
 sg13g2_fill_2 FILLER_65_79 ();
 sg13g2_fill_1 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_117 ();
 sg13g2_fill_2 FILLER_65_128 ();
 sg13g2_fill_1 FILLER_65_183 ();
 sg13g2_fill_2 FILLER_65_215 ();
 sg13g2_fill_1 FILLER_65_217 ();
 sg13g2_fill_1 FILLER_65_243 ();
 sg13g2_decap_4 FILLER_65_264 ();
 sg13g2_fill_1 FILLER_65_268 ();
 sg13g2_fill_2 FILLER_65_277 ();
 sg13g2_decap_4 FILLER_65_285 ();
 sg13g2_fill_1 FILLER_65_289 ();
 sg13g2_decap_4 FILLER_65_298 ();
 sg13g2_fill_1 FILLER_65_302 ();
 sg13g2_fill_2 FILLER_65_334 ();
 sg13g2_fill_2 FILLER_65_341 ();
 sg13g2_fill_2 FILLER_65_571 ();
 sg13g2_fill_1 FILLER_65_573 ();
 sg13g2_fill_2 FILLER_65_584 ();
 sg13g2_fill_1 FILLER_65_591 ();
 sg13g2_decap_4 FILLER_65_596 ();
 sg13g2_fill_2 FILLER_65_600 ();
 sg13g2_decap_4 FILLER_65_628 ();
 sg13g2_fill_1 FILLER_65_632 ();
 sg13g2_fill_2 FILLER_65_659 ();
 sg13g2_fill_2 FILLER_65_666 ();
 sg13g2_decap_4 FILLER_65_681 ();
 sg13g2_fill_1 FILLER_65_685 ();
 sg13g2_fill_2 FILLER_65_696 ();
 sg13g2_fill_2 FILLER_65_715 ();
 sg13g2_fill_2 FILLER_65_722 ();
 sg13g2_fill_1 FILLER_65_724 ();
 sg13g2_fill_1 FILLER_65_764 ();
 sg13g2_fill_2 FILLER_65_774 ();
 sg13g2_fill_1 FILLER_65_792 ();
 sg13g2_decap_8 FILLER_65_823 ();
 sg13g2_fill_2 FILLER_65_830 ();
 sg13g2_fill_1 FILLER_65_832 ();
 sg13g2_decap_8 FILLER_65_837 ();
 sg13g2_decap_8 FILLER_65_844 ();
 sg13g2_decap_8 FILLER_65_851 ();
 sg13g2_decap_8 FILLER_65_858 ();
 sg13g2_decap_8 FILLER_65_865 ();
 sg13g2_decap_8 FILLER_65_872 ();
 sg13g2_decap_8 FILLER_65_879 ();
 sg13g2_decap_8 FILLER_65_886 ();
 sg13g2_decap_8 FILLER_65_893 ();
 sg13g2_decap_8 FILLER_65_900 ();
 sg13g2_decap_8 FILLER_65_907 ();
 sg13g2_decap_8 FILLER_65_914 ();
 sg13g2_decap_8 FILLER_65_921 ();
 sg13g2_decap_8 FILLER_65_928 ();
 sg13g2_decap_8 FILLER_65_935 ();
 sg13g2_decap_8 FILLER_65_942 ();
 sg13g2_decap_8 FILLER_65_949 ();
 sg13g2_decap_8 FILLER_65_956 ();
 sg13g2_decap_8 FILLER_65_963 ();
 sg13g2_decap_8 FILLER_65_970 ();
 sg13g2_decap_8 FILLER_65_977 ();
 sg13g2_decap_8 FILLER_65_984 ();
 sg13g2_decap_8 FILLER_65_991 ();
 sg13g2_decap_8 FILLER_65_998 ();
 sg13g2_decap_8 FILLER_65_1005 ();
 sg13g2_decap_8 FILLER_65_1012 ();
 sg13g2_decap_8 FILLER_65_1019 ();
 sg13g2_decap_8 FILLER_65_1026 ();
 sg13g2_decap_8 FILLER_65_1033 ();
 sg13g2_decap_8 FILLER_65_1040 ();
 sg13g2_decap_8 FILLER_65_1047 ();
 sg13g2_decap_8 FILLER_65_1054 ();
 sg13g2_decap_8 FILLER_65_1061 ();
 sg13g2_decap_8 FILLER_65_1068 ();
 sg13g2_decap_8 FILLER_65_1075 ();
 sg13g2_decap_8 FILLER_65_1082 ();
 sg13g2_decap_8 FILLER_65_1089 ();
 sg13g2_decap_8 FILLER_65_1096 ();
 sg13g2_decap_8 FILLER_65_1103 ();
 sg13g2_decap_8 FILLER_65_1110 ();
 sg13g2_decap_8 FILLER_65_1117 ();
 sg13g2_decap_8 FILLER_65_1124 ();
 sg13g2_decap_8 FILLER_65_1131 ();
 sg13g2_decap_8 FILLER_65_1138 ();
 sg13g2_decap_8 FILLER_65_1145 ();
 sg13g2_decap_8 FILLER_65_1152 ();
 sg13g2_decap_8 FILLER_65_1159 ();
 sg13g2_decap_8 FILLER_65_1166 ();
 sg13g2_decap_8 FILLER_65_1173 ();
 sg13g2_decap_8 FILLER_65_1180 ();
 sg13g2_decap_8 FILLER_65_1187 ();
 sg13g2_decap_8 FILLER_65_1194 ();
 sg13g2_decap_8 FILLER_65_1201 ();
 sg13g2_decap_8 FILLER_65_1208 ();
 sg13g2_decap_8 FILLER_65_1215 ();
 sg13g2_decap_8 FILLER_65_1222 ();
 sg13g2_decap_8 FILLER_65_1229 ();
 sg13g2_decap_8 FILLER_65_1236 ();
 sg13g2_decap_8 FILLER_65_1243 ();
 sg13g2_decap_8 FILLER_65_1250 ();
 sg13g2_decap_8 FILLER_65_1257 ();
 sg13g2_decap_8 FILLER_65_1264 ();
 sg13g2_decap_8 FILLER_65_1271 ();
 sg13g2_decap_8 FILLER_65_1278 ();
 sg13g2_decap_8 FILLER_65_1285 ();
 sg13g2_decap_8 FILLER_65_1292 ();
 sg13g2_decap_8 FILLER_65_1299 ();
 sg13g2_decap_8 FILLER_65_1306 ();
 sg13g2_fill_2 FILLER_65_1313 ();
 sg13g2_fill_2 FILLER_66_26 ();
 sg13g2_fill_1 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_48 ();
 sg13g2_fill_2 FILLER_66_105 ();
 sg13g2_fill_1 FILLER_66_107 ();
 sg13g2_fill_1 FILLER_66_141 ();
 sg13g2_decap_4 FILLER_66_249 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_fill_2 FILLER_66_266 ();
 sg13g2_decap_4 FILLER_66_274 ();
 sg13g2_fill_2 FILLER_66_285 ();
 sg13g2_fill_1 FILLER_66_287 ();
 sg13g2_decap_4 FILLER_66_307 ();
 sg13g2_fill_2 FILLER_66_351 ();
 sg13g2_fill_1 FILLER_66_367 ();
 sg13g2_fill_2 FILLER_66_383 ();
 sg13g2_fill_1 FILLER_66_391 ();
 sg13g2_fill_2 FILLER_66_401 ();
 sg13g2_fill_2 FILLER_66_408 ();
 sg13g2_fill_1 FILLER_66_410 ();
 sg13g2_fill_2 FILLER_66_469 ();
 sg13g2_fill_1 FILLER_66_502 ();
 sg13g2_fill_1 FILLER_66_516 ();
 sg13g2_fill_1 FILLER_66_521 ();
 sg13g2_fill_1 FILLER_66_540 ();
 sg13g2_decap_4 FILLER_66_577 ();
 sg13g2_fill_2 FILLER_66_607 ();
 sg13g2_fill_1 FILLER_66_631 ();
 sg13g2_decap_8 FILLER_66_653 ();
 sg13g2_decap_8 FILLER_66_660 ();
 sg13g2_decap_4 FILLER_66_693 ();
 sg13g2_fill_1 FILLER_66_705 ();
 sg13g2_fill_1 FILLER_66_714 ();
 sg13g2_fill_1 FILLER_66_720 ();
 sg13g2_fill_2 FILLER_66_744 ();
 sg13g2_fill_1 FILLER_66_746 ();
 sg13g2_fill_2 FILLER_66_759 ();
 sg13g2_decap_8 FILLER_66_785 ();
 sg13g2_decap_8 FILLER_66_792 ();
 sg13g2_decap_4 FILLER_66_799 ();
 sg13g2_fill_2 FILLER_66_803 ();
 sg13g2_fill_2 FILLER_66_809 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_decap_8 FILLER_66_857 ();
 sg13g2_decap_8 FILLER_66_864 ();
 sg13g2_decap_8 FILLER_66_871 ();
 sg13g2_decap_8 FILLER_66_878 ();
 sg13g2_decap_8 FILLER_66_885 ();
 sg13g2_decap_8 FILLER_66_892 ();
 sg13g2_decap_8 FILLER_66_899 ();
 sg13g2_decap_8 FILLER_66_906 ();
 sg13g2_decap_8 FILLER_66_913 ();
 sg13g2_decap_8 FILLER_66_920 ();
 sg13g2_decap_8 FILLER_66_927 ();
 sg13g2_decap_8 FILLER_66_934 ();
 sg13g2_decap_8 FILLER_66_941 ();
 sg13g2_decap_8 FILLER_66_948 ();
 sg13g2_decap_8 FILLER_66_955 ();
 sg13g2_decap_8 FILLER_66_962 ();
 sg13g2_decap_8 FILLER_66_969 ();
 sg13g2_decap_8 FILLER_66_976 ();
 sg13g2_decap_8 FILLER_66_983 ();
 sg13g2_decap_8 FILLER_66_990 ();
 sg13g2_decap_8 FILLER_66_997 ();
 sg13g2_decap_8 FILLER_66_1004 ();
 sg13g2_decap_8 FILLER_66_1011 ();
 sg13g2_decap_8 FILLER_66_1018 ();
 sg13g2_decap_8 FILLER_66_1025 ();
 sg13g2_decap_8 FILLER_66_1032 ();
 sg13g2_decap_8 FILLER_66_1039 ();
 sg13g2_decap_8 FILLER_66_1046 ();
 sg13g2_decap_8 FILLER_66_1053 ();
 sg13g2_decap_8 FILLER_66_1060 ();
 sg13g2_decap_8 FILLER_66_1067 ();
 sg13g2_decap_8 FILLER_66_1074 ();
 sg13g2_decap_8 FILLER_66_1081 ();
 sg13g2_decap_8 FILLER_66_1088 ();
 sg13g2_decap_8 FILLER_66_1095 ();
 sg13g2_decap_8 FILLER_66_1102 ();
 sg13g2_decap_8 FILLER_66_1109 ();
 sg13g2_decap_8 FILLER_66_1116 ();
 sg13g2_decap_8 FILLER_66_1123 ();
 sg13g2_decap_8 FILLER_66_1130 ();
 sg13g2_decap_8 FILLER_66_1137 ();
 sg13g2_decap_8 FILLER_66_1144 ();
 sg13g2_decap_8 FILLER_66_1151 ();
 sg13g2_decap_8 FILLER_66_1158 ();
 sg13g2_decap_8 FILLER_66_1165 ();
 sg13g2_decap_8 FILLER_66_1172 ();
 sg13g2_decap_8 FILLER_66_1179 ();
 sg13g2_decap_8 FILLER_66_1186 ();
 sg13g2_decap_8 FILLER_66_1193 ();
 sg13g2_decap_8 FILLER_66_1200 ();
 sg13g2_decap_8 FILLER_66_1207 ();
 sg13g2_decap_8 FILLER_66_1214 ();
 sg13g2_decap_8 FILLER_66_1221 ();
 sg13g2_decap_8 FILLER_66_1228 ();
 sg13g2_decap_8 FILLER_66_1235 ();
 sg13g2_decap_8 FILLER_66_1242 ();
 sg13g2_decap_8 FILLER_66_1249 ();
 sg13g2_decap_8 FILLER_66_1256 ();
 sg13g2_decap_8 FILLER_66_1263 ();
 sg13g2_decap_8 FILLER_66_1270 ();
 sg13g2_decap_8 FILLER_66_1277 ();
 sg13g2_decap_8 FILLER_66_1284 ();
 sg13g2_decap_8 FILLER_66_1291 ();
 sg13g2_decap_8 FILLER_66_1298 ();
 sg13g2_decap_8 FILLER_66_1305 ();
 sg13g2_fill_2 FILLER_66_1312 ();
 sg13g2_fill_1 FILLER_66_1314 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_86 ();
 sg13g2_fill_1 FILLER_67_88 ();
 sg13g2_fill_2 FILLER_67_156 ();
 sg13g2_fill_2 FILLER_67_163 ();
 sg13g2_fill_1 FILLER_67_165 ();
 sg13g2_fill_2 FILLER_67_197 ();
 sg13g2_fill_1 FILLER_67_199 ();
 sg13g2_fill_2 FILLER_67_205 ();
 sg13g2_fill_2 FILLER_67_216 ();
 sg13g2_fill_1 FILLER_67_218 ();
 sg13g2_fill_2 FILLER_67_285 ();
 sg13g2_fill_1 FILLER_67_287 ();
 sg13g2_fill_1 FILLER_67_311 ();
 sg13g2_fill_1 FILLER_67_349 ();
 sg13g2_fill_2 FILLER_67_438 ();
 sg13g2_fill_2 FILLER_67_475 ();
 sg13g2_fill_1 FILLER_67_485 ();
 sg13g2_fill_1 FILLER_67_491 ();
 sg13g2_fill_1 FILLER_67_537 ();
 sg13g2_fill_2 FILLER_67_555 ();
 sg13g2_fill_2 FILLER_67_580 ();
 sg13g2_fill_1 FILLER_67_582 ();
 sg13g2_fill_1 FILLER_67_596 ();
 sg13g2_fill_2 FILLER_67_654 ();
 sg13g2_fill_1 FILLER_67_656 ();
 sg13g2_decap_8 FILLER_67_661 ();
 sg13g2_decap_4 FILLER_67_668 ();
 sg13g2_fill_2 FILLER_67_672 ();
 sg13g2_fill_1 FILLER_67_687 ();
 sg13g2_fill_1 FILLER_67_701 ();
 sg13g2_fill_2 FILLER_67_712 ();
 sg13g2_decap_4 FILLER_67_733 ();
 sg13g2_fill_2 FILLER_67_737 ();
 sg13g2_fill_2 FILLER_67_743 ();
 sg13g2_decap_4 FILLER_67_754 ();
 sg13g2_fill_1 FILLER_67_758 ();
 sg13g2_fill_1 FILLER_67_764 ();
 sg13g2_fill_2 FILLER_67_774 ();
 sg13g2_fill_1 FILLER_67_776 ();
 sg13g2_fill_2 FILLER_67_785 ();
 sg13g2_fill_2 FILLER_67_808 ();
 sg13g2_fill_1 FILLER_67_831 ();
 sg13g2_decap_8 FILLER_67_836 ();
 sg13g2_decap_8 FILLER_67_843 ();
 sg13g2_decap_8 FILLER_67_850 ();
 sg13g2_decap_8 FILLER_67_857 ();
 sg13g2_decap_8 FILLER_67_864 ();
 sg13g2_decap_8 FILLER_67_871 ();
 sg13g2_decap_8 FILLER_67_878 ();
 sg13g2_decap_8 FILLER_67_885 ();
 sg13g2_decap_8 FILLER_67_892 ();
 sg13g2_decap_8 FILLER_67_899 ();
 sg13g2_decap_8 FILLER_67_906 ();
 sg13g2_decap_8 FILLER_67_913 ();
 sg13g2_decap_8 FILLER_67_920 ();
 sg13g2_decap_8 FILLER_67_927 ();
 sg13g2_decap_8 FILLER_67_934 ();
 sg13g2_decap_8 FILLER_67_941 ();
 sg13g2_decap_8 FILLER_67_948 ();
 sg13g2_decap_8 FILLER_67_955 ();
 sg13g2_decap_8 FILLER_67_962 ();
 sg13g2_decap_8 FILLER_67_969 ();
 sg13g2_decap_8 FILLER_67_976 ();
 sg13g2_decap_8 FILLER_67_983 ();
 sg13g2_decap_8 FILLER_67_990 ();
 sg13g2_decap_8 FILLER_67_997 ();
 sg13g2_decap_8 FILLER_67_1004 ();
 sg13g2_decap_8 FILLER_67_1011 ();
 sg13g2_decap_8 FILLER_67_1018 ();
 sg13g2_decap_8 FILLER_67_1025 ();
 sg13g2_decap_8 FILLER_67_1032 ();
 sg13g2_decap_8 FILLER_67_1039 ();
 sg13g2_decap_8 FILLER_67_1046 ();
 sg13g2_decap_8 FILLER_67_1053 ();
 sg13g2_decap_8 FILLER_67_1060 ();
 sg13g2_decap_8 FILLER_67_1067 ();
 sg13g2_decap_8 FILLER_67_1074 ();
 sg13g2_decap_8 FILLER_67_1081 ();
 sg13g2_decap_8 FILLER_67_1088 ();
 sg13g2_decap_8 FILLER_67_1095 ();
 sg13g2_decap_8 FILLER_67_1102 ();
 sg13g2_decap_8 FILLER_67_1109 ();
 sg13g2_decap_8 FILLER_67_1116 ();
 sg13g2_decap_8 FILLER_67_1123 ();
 sg13g2_decap_8 FILLER_67_1130 ();
 sg13g2_decap_8 FILLER_67_1137 ();
 sg13g2_decap_8 FILLER_67_1144 ();
 sg13g2_decap_8 FILLER_67_1151 ();
 sg13g2_decap_8 FILLER_67_1158 ();
 sg13g2_decap_8 FILLER_67_1165 ();
 sg13g2_decap_8 FILLER_67_1172 ();
 sg13g2_decap_8 FILLER_67_1179 ();
 sg13g2_decap_8 FILLER_67_1186 ();
 sg13g2_decap_8 FILLER_67_1193 ();
 sg13g2_decap_8 FILLER_67_1200 ();
 sg13g2_decap_8 FILLER_67_1207 ();
 sg13g2_decap_8 FILLER_67_1214 ();
 sg13g2_decap_8 FILLER_67_1221 ();
 sg13g2_decap_8 FILLER_67_1228 ();
 sg13g2_decap_8 FILLER_67_1235 ();
 sg13g2_decap_8 FILLER_67_1242 ();
 sg13g2_decap_8 FILLER_67_1249 ();
 sg13g2_decap_8 FILLER_67_1256 ();
 sg13g2_decap_8 FILLER_67_1263 ();
 sg13g2_decap_8 FILLER_67_1270 ();
 sg13g2_decap_8 FILLER_67_1277 ();
 sg13g2_decap_8 FILLER_67_1284 ();
 sg13g2_decap_8 FILLER_67_1291 ();
 sg13g2_decap_8 FILLER_67_1298 ();
 sg13g2_decap_8 FILLER_67_1305 ();
 sg13g2_fill_2 FILLER_67_1312 ();
 sg13g2_fill_1 FILLER_67_1314 ();
 sg13g2_fill_2 FILLER_68_40 ();
 sg13g2_fill_2 FILLER_68_51 ();
 sg13g2_fill_2 FILLER_68_70 ();
 sg13g2_fill_1 FILLER_68_72 ();
 sg13g2_fill_2 FILLER_68_83 ();
 sg13g2_fill_1 FILLER_68_85 ();
 sg13g2_fill_1 FILLER_68_135 ();
 sg13g2_fill_2 FILLER_68_166 ();
 sg13g2_fill_1 FILLER_68_168 ();
 sg13g2_fill_2 FILLER_68_207 ();
 sg13g2_fill_1 FILLER_68_209 ();
 sg13g2_fill_2 FILLER_68_258 ();
 sg13g2_fill_2 FILLER_68_272 ();
 sg13g2_fill_1 FILLER_68_274 ();
 sg13g2_fill_2 FILLER_68_281 ();
 sg13g2_fill_1 FILLER_68_283 ();
 sg13g2_fill_2 FILLER_68_384 ();
 sg13g2_fill_1 FILLER_68_386 ();
 sg13g2_fill_1 FILLER_68_416 ();
 sg13g2_fill_1 FILLER_68_432 ();
 sg13g2_fill_1 FILLER_68_448 ();
 sg13g2_fill_2 FILLER_68_471 ();
 sg13g2_fill_1 FILLER_68_473 ();
 sg13g2_fill_2 FILLER_68_505 ();
 sg13g2_fill_2 FILLER_68_533 ();
 sg13g2_fill_1 FILLER_68_573 ();
 sg13g2_decap_8 FILLER_68_635 ();
 sg13g2_decap_8 FILLER_68_642 ();
 sg13g2_fill_1 FILLER_68_649 ();
 sg13g2_fill_2 FILLER_68_671 ();
 sg13g2_fill_1 FILLER_68_673 ();
 sg13g2_fill_1 FILLER_68_708 ();
 sg13g2_decap_4 FILLER_68_724 ();
 sg13g2_fill_2 FILLER_68_728 ();
 sg13g2_fill_1 FILLER_68_740 ();
 sg13g2_fill_2 FILLER_68_761 ();
 sg13g2_decap_8 FILLER_68_767 ();
 sg13g2_decap_4 FILLER_68_774 ();
 sg13g2_fill_1 FILLER_68_778 ();
 sg13g2_fill_1 FILLER_68_787 ();
 sg13g2_fill_2 FILLER_68_793 ();
 sg13g2_decap_4 FILLER_68_808 ();
 sg13g2_fill_2 FILLER_68_812 ();
 sg13g2_fill_1 FILLER_68_817 ();
 sg13g2_decap_8 FILLER_68_821 ();
 sg13g2_decap_8 FILLER_68_828 ();
 sg13g2_fill_1 FILLER_68_835 ();
 sg13g2_decap_8 FILLER_68_839 ();
 sg13g2_decap_8 FILLER_68_846 ();
 sg13g2_decap_8 FILLER_68_853 ();
 sg13g2_decap_8 FILLER_68_860 ();
 sg13g2_decap_8 FILLER_68_867 ();
 sg13g2_decap_8 FILLER_68_874 ();
 sg13g2_decap_8 FILLER_68_881 ();
 sg13g2_decap_8 FILLER_68_888 ();
 sg13g2_decap_8 FILLER_68_895 ();
 sg13g2_decap_8 FILLER_68_902 ();
 sg13g2_decap_8 FILLER_68_909 ();
 sg13g2_decap_8 FILLER_68_916 ();
 sg13g2_decap_8 FILLER_68_923 ();
 sg13g2_decap_8 FILLER_68_930 ();
 sg13g2_decap_8 FILLER_68_937 ();
 sg13g2_decap_8 FILLER_68_944 ();
 sg13g2_decap_8 FILLER_68_951 ();
 sg13g2_decap_8 FILLER_68_958 ();
 sg13g2_decap_8 FILLER_68_965 ();
 sg13g2_decap_8 FILLER_68_972 ();
 sg13g2_decap_8 FILLER_68_979 ();
 sg13g2_decap_8 FILLER_68_986 ();
 sg13g2_decap_8 FILLER_68_993 ();
 sg13g2_decap_8 FILLER_68_1000 ();
 sg13g2_decap_8 FILLER_68_1007 ();
 sg13g2_decap_8 FILLER_68_1014 ();
 sg13g2_decap_8 FILLER_68_1021 ();
 sg13g2_decap_8 FILLER_68_1028 ();
 sg13g2_decap_8 FILLER_68_1035 ();
 sg13g2_decap_8 FILLER_68_1042 ();
 sg13g2_decap_8 FILLER_68_1049 ();
 sg13g2_decap_8 FILLER_68_1056 ();
 sg13g2_decap_8 FILLER_68_1063 ();
 sg13g2_decap_8 FILLER_68_1070 ();
 sg13g2_decap_8 FILLER_68_1077 ();
 sg13g2_decap_8 FILLER_68_1084 ();
 sg13g2_decap_8 FILLER_68_1091 ();
 sg13g2_decap_8 FILLER_68_1098 ();
 sg13g2_decap_8 FILLER_68_1105 ();
 sg13g2_decap_8 FILLER_68_1112 ();
 sg13g2_decap_8 FILLER_68_1119 ();
 sg13g2_decap_8 FILLER_68_1126 ();
 sg13g2_decap_8 FILLER_68_1133 ();
 sg13g2_decap_8 FILLER_68_1140 ();
 sg13g2_decap_8 FILLER_68_1147 ();
 sg13g2_decap_8 FILLER_68_1154 ();
 sg13g2_decap_8 FILLER_68_1161 ();
 sg13g2_decap_8 FILLER_68_1168 ();
 sg13g2_decap_8 FILLER_68_1175 ();
 sg13g2_decap_8 FILLER_68_1182 ();
 sg13g2_decap_8 FILLER_68_1189 ();
 sg13g2_decap_8 FILLER_68_1196 ();
 sg13g2_decap_8 FILLER_68_1203 ();
 sg13g2_decap_8 FILLER_68_1210 ();
 sg13g2_decap_8 FILLER_68_1217 ();
 sg13g2_decap_8 FILLER_68_1224 ();
 sg13g2_decap_8 FILLER_68_1231 ();
 sg13g2_decap_8 FILLER_68_1238 ();
 sg13g2_decap_8 FILLER_68_1245 ();
 sg13g2_decap_8 FILLER_68_1252 ();
 sg13g2_decap_8 FILLER_68_1259 ();
 sg13g2_decap_8 FILLER_68_1266 ();
 sg13g2_decap_8 FILLER_68_1273 ();
 sg13g2_decap_8 FILLER_68_1280 ();
 sg13g2_decap_8 FILLER_68_1287 ();
 sg13g2_decap_8 FILLER_68_1294 ();
 sg13g2_decap_8 FILLER_68_1301 ();
 sg13g2_decap_8 FILLER_68_1308 ();
 sg13g2_fill_1 FILLER_69_83 ();
 sg13g2_fill_1 FILLER_69_99 ();
 sg13g2_fill_1 FILLER_69_109 ();
 sg13g2_fill_2 FILLER_69_151 ();
 sg13g2_fill_1 FILLER_69_153 ();
 sg13g2_fill_2 FILLER_69_180 ();
 sg13g2_fill_1 FILLER_69_182 ();
 sg13g2_fill_1 FILLER_69_227 ();
 sg13g2_fill_2 FILLER_69_240 ();
 sg13g2_fill_1 FILLER_69_242 ();
 sg13g2_decap_8 FILLER_69_249 ();
 sg13g2_fill_1 FILLER_69_256 ();
 sg13g2_fill_2 FILLER_69_269 ();
 sg13g2_fill_1 FILLER_69_271 ();
 sg13g2_decap_4 FILLER_69_316 ();
 sg13g2_fill_2 FILLER_69_320 ();
 sg13g2_fill_2 FILLER_69_332 ();
 sg13g2_fill_2 FILLER_69_369 ();
 sg13g2_fill_1 FILLER_69_414 ();
 sg13g2_fill_2 FILLER_69_543 ();
 sg13g2_fill_2 FILLER_69_559 ();
 sg13g2_fill_2 FILLER_69_566 ();
 sg13g2_decap_4 FILLER_69_602 ();
 sg13g2_fill_1 FILLER_69_606 ();
 sg13g2_fill_1 FILLER_69_620 ();
 sg13g2_decap_8 FILLER_69_668 ();
 sg13g2_decap_4 FILLER_69_675 ();
 sg13g2_fill_1 FILLER_69_684 ();
 sg13g2_decap_8 FILLER_69_690 ();
 sg13g2_decap_8 FILLER_69_718 ();
 sg13g2_decap_8 FILLER_69_725 ();
 sg13g2_decap_8 FILLER_69_732 ();
 sg13g2_decap_4 FILLER_69_739 ();
 sg13g2_fill_2 FILLER_69_743 ();
 sg13g2_decap_8 FILLER_69_750 ();
 sg13g2_fill_1 FILLER_69_757 ();
 sg13g2_fill_2 FILLER_69_762 ();
 sg13g2_fill_2 FILLER_69_788 ();
 sg13g2_fill_1 FILLER_69_790 ();
 sg13g2_fill_1 FILLER_69_816 ();
 sg13g2_decap_8 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_69_850 ();
 sg13g2_decap_8 FILLER_69_857 ();
 sg13g2_decap_8 FILLER_69_864 ();
 sg13g2_decap_8 FILLER_69_871 ();
 sg13g2_decap_8 FILLER_69_878 ();
 sg13g2_decap_8 FILLER_69_885 ();
 sg13g2_decap_8 FILLER_69_892 ();
 sg13g2_decap_8 FILLER_69_899 ();
 sg13g2_decap_8 FILLER_69_906 ();
 sg13g2_decap_8 FILLER_69_913 ();
 sg13g2_decap_8 FILLER_69_920 ();
 sg13g2_decap_8 FILLER_69_927 ();
 sg13g2_decap_8 FILLER_69_934 ();
 sg13g2_decap_8 FILLER_69_941 ();
 sg13g2_decap_8 FILLER_69_948 ();
 sg13g2_decap_8 FILLER_69_955 ();
 sg13g2_decap_8 FILLER_69_962 ();
 sg13g2_decap_8 FILLER_69_969 ();
 sg13g2_decap_8 FILLER_69_976 ();
 sg13g2_decap_8 FILLER_69_983 ();
 sg13g2_decap_8 FILLER_69_990 ();
 sg13g2_decap_8 FILLER_69_997 ();
 sg13g2_decap_8 FILLER_69_1004 ();
 sg13g2_decap_8 FILLER_69_1011 ();
 sg13g2_decap_8 FILLER_69_1018 ();
 sg13g2_decap_8 FILLER_69_1025 ();
 sg13g2_decap_8 FILLER_69_1032 ();
 sg13g2_decap_8 FILLER_69_1039 ();
 sg13g2_decap_8 FILLER_69_1046 ();
 sg13g2_decap_8 FILLER_69_1053 ();
 sg13g2_decap_8 FILLER_69_1060 ();
 sg13g2_decap_8 FILLER_69_1067 ();
 sg13g2_decap_8 FILLER_69_1074 ();
 sg13g2_decap_8 FILLER_69_1081 ();
 sg13g2_decap_8 FILLER_69_1088 ();
 sg13g2_decap_8 FILLER_69_1095 ();
 sg13g2_decap_8 FILLER_69_1102 ();
 sg13g2_decap_8 FILLER_69_1109 ();
 sg13g2_decap_8 FILLER_69_1116 ();
 sg13g2_decap_8 FILLER_69_1123 ();
 sg13g2_decap_8 FILLER_69_1130 ();
 sg13g2_decap_8 FILLER_69_1137 ();
 sg13g2_decap_8 FILLER_69_1144 ();
 sg13g2_decap_8 FILLER_69_1151 ();
 sg13g2_decap_8 FILLER_69_1158 ();
 sg13g2_decap_8 FILLER_69_1165 ();
 sg13g2_decap_8 FILLER_69_1172 ();
 sg13g2_decap_8 FILLER_69_1179 ();
 sg13g2_decap_8 FILLER_69_1186 ();
 sg13g2_decap_8 FILLER_69_1193 ();
 sg13g2_decap_8 FILLER_69_1200 ();
 sg13g2_decap_8 FILLER_69_1207 ();
 sg13g2_decap_8 FILLER_69_1214 ();
 sg13g2_decap_8 FILLER_69_1221 ();
 sg13g2_decap_8 FILLER_69_1228 ();
 sg13g2_decap_8 FILLER_69_1235 ();
 sg13g2_decap_8 FILLER_69_1242 ();
 sg13g2_decap_8 FILLER_69_1249 ();
 sg13g2_decap_8 FILLER_69_1256 ();
 sg13g2_decap_8 FILLER_69_1263 ();
 sg13g2_decap_8 FILLER_69_1270 ();
 sg13g2_decap_8 FILLER_69_1277 ();
 sg13g2_decap_8 FILLER_69_1284 ();
 sg13g2_decap_8 FILLER_69_1291 ();
 sg13g2_decap_8 FILLER_69_1298 ();
 sg13g2_decap_8 FILLER_69_1305 ();
 sg13g2_fill_2 FILLER_69_1312 ();
 sg13g2_fill_1 FILLER_69_1314 ();
 sg13g2_fill_1 FILLER_70_45 ();
 sg13g2_fill_2 FILLER_70_55 ();
 sg13g2_fill_1 FILLER_70_95 ();
 sg13g2_fill_2 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_135 ();
 sg13g2_fill_2 FILLER_70_150 ();
 sg13g2_fill_1 FILLER_70_152 ();
 sg13g2_fill_2 FILLER_70_162 ();
 sg13g2_fill_2 FILLER_70_215 ();
 sg13g2_fill_1 FILLER_70_226 ();
 sg13g2_fill_2 FILLER_70_245 ();
 sg13g2_fill_1 FILLER_70_252 ();
 sg13g2_fill_1 FILLER_70_276 ();
 sg13g2_fill_2 FILLER_70_285 ();
 sg13g2_fill_1 FILLER_70_287 ();
 sg13g2_fill_1 FILLER_70_297 ();
 sg13g2_fill_2 FILLER_70_311 ();
 sg13g2_fill_1 FILLER_70_313 ();
 sg13g2_fill_2 FILLER_70_333 ();
 sg13g2_fill_1 FILLER_70_344 ();
 sg13g2_fill_2 FILLER_70_349 ();
 sg13g2_fill_2 FILLER_70_377 ();
 sg13g2_fill_2 FILLER_70_405 ();
 sg13g2_fill_1 FILLER_70_407 ();
 sg13g2_fill_2 FILLER_70_430 ();
 sg13g2_fill_2 FILLER_70_465 ();
 sg13g2_fill_1 FILLER_70_467 ();
 sg13g2_fill_1 FILLER_70_560 ();
 sg13g2_fill_1 FILLER_70_584 ();
 sg13g2_fill_1 FILLER_70_631 ();
 sg13g2_fill_2 FILLER_70_658 ();
 sg13g2_fill_2 FILLER_70_681 ();
 sg13g2_fill_1 FILLER_70_683 ();
 sg13g2_decap_8 FILLER_70_715 ();
 sg13g2_decap_4 FILLER_70_748 ();
 sg13g2_fill_1 FILLER_70_752 ();
 sg13g2_fill_2 FILLER_70_758 ();
 sg13g2_fill_1 FILLER_70_760 ();
 sg13g2_decap_8 FILLER_70_779 ();
 sg13g2_decap_4 FILLER_70_786 ();
 sg13g2_fill_2 FILLER_70_790 ();
 sg13g2_fill_1 FILLER_70_797 ();
 sg13g2_decap_4 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_818 ();
 sg13g2_fill_2 FILLER_70_825 ();
 sg13g2_fill_1 FILLER_70_827 ();
 sg13g2_decap_8 FILLER_70_835 ();
 sg13g2_decap_8 FILLER_70_842 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_8 FILLER_70_856 ();
 sg13g2_decap_8 FILLER_70_863 ();
 sg13g2_decap_8 FILLER_70_870 ();
 sg13g2_decap_8 FILLER_70_877 ();
 sg13g2_decap_8 FILLER_70_884 ();
 sg13g2_decap_8 FILLER_70_891 ();
 sg13g2_decap_8 FILLER_70_898 ();
 sg13g2_decap_8 FILLER_70_905 ();
 sg13g2_decap_8 FILLER_70_912 ();
 sg13g2_decap_8 FILLER_70_919 ();
 sg13g2_decap_8 FILLER_70_926 ();
 sg13g2_decap_8 FILLER_70_933 ();
 sg13g2_decap_8 FILLER_70_940 ();
 sg13g2_decap_8 FILLER_70_947 ();
 sg13g2_decap_8 FILLER_70_954 ();
 sg13g2_decap_8 FILLER_70_961 ();
 sg13g2_decap_8 FILLER_70_968 ();
 sg13g2_decap_8 FILLER_70_975 ();
 sg13g2_decap_8 FILLER_70_982 ();
 sg13g2_decap_8 FILLER_70_989 ();
 sg13g2_decap_8 FILLER_70_996 ();
 sg13g2_decap_8 FILLER_70_1003 ();
 sg13g2_decap_8 FILLER_70_1010 ();
 sg13g2_decap_8 FILLER_70_1017 ();
 sg13g2_decap_8 FILLER_70_1024 ();
 sg13g2_decap_8 FILLER_70_1031 ();
 sg13g2_decap_8 FILLER_70_1038 ();
 sg13g2_decap_8 FILLER_70_1045 ();
 sg13g2_decap_8 FILLER_70_1052 ();
 sg13g2_decap_8 FILLER_70_1059 ();
 sg13g2_decap_8 FILLER_70_1066 ();
 sg13g2_decap_8 FILLER_70_1073 ();
 sg13g2_decap_8 FILLER_70_1080 ();
 sg13g2_decap_8 FILLER_70_1087 ();
 sg13g2_decap_8 FILLER_70_1094 ();
 sg13g2_decap_8 FILLER_70_1101 ();
 sg13g2_decap_8 FILLER_70_1108 ();
 sg13g2_decap_8 FILLER_70_1115 ();
 sg13g2_decap_8 FILLER_70_1122 ();
 sg13g2_decap_8 FILLER_70_1129 ();
 sg13g2_decap_8 FILLER_70_1136 ();
 sg13g2_decap_8 FILLER_70_1143 ();
 sg13g2_decap_8 FILLER_70_1150 ();
 sg13g2_decap_8 FILLER_70_1157 ();
 sg13g2_decap_8 FILLER_70_1164 ();
 sg13g2_decap_8 FILLER_70_1171 ();
 sg13g2_decap_8 FILLER_70_1178 ();
 sg13g2_decap_8 FILLER_70_1185 ();
 sg13g2_decap_8 FILLER_70_1192 ();
 sg13g2_decap_8 FILLER_70_1199 ();
 sg13g2_decap_8 FILLER_70_1206 ();
 sg13g2_decap_8 FILLER_70_1213 ();
 sg13g2_decap_8 FILLER_70_1220 ();
 sg13g2_decap_8 FILLER_70_1227 ();
 sg13g2_decap_8 FILLER_70_1234 ();
 sg13g2_decap_8 FILLER_70_1241 ();
 sg13g2_decap_8 FILLER_70_1248 ();
 sg13g2_decap_8 FILLER_70_1255 ();
 sg13g2_decap_8 FILLER_70_1262 ();
 sg13g2_decap_8 FILLER_70_1269 ();
 sg13g2_decap_8 FILLER_70_1276 ();
 sg13g2_decap_8 FILLER_70_1283 ();
 sg13g2_decap_8 FILLER_70_1290 ();
 sg13g2_decap_8 FILLER_70_1297 ();
 sg13g2_decap_8 FILLER_70_1304 ();
 sg13g2_decap_4 FILLER_70_1311 ();
 sg13g2_fill_1 FILLER_71_26 ();
 sg13g2_fill_1 FILLER_71_120 ();
 sg13g2_fill_1 FILLER_71_147 ();
 sg13g2_fill_2 FILLER_71_161 ();
 sg13g2_fill_1 FILLER_71_270 ();
 sg13g2_fill_2 FILLER_71_302 ();
 sg13g2_fill_1 FILLER_71_304 ();
 sg13g2_fill_2 FILLER_71_404 ();
 sg13g2_fill_2 FILLER_71_437 ();
 sg13g2_fill_2 FILLER_71_465 ();
 sg13g2_fill_2 FILLER_71_571 ();
 sg13g2_fill_1 FILLER_71_605 ();
 sg13g2_decap_4 FILLER_71_625 ();
 sg13g2_fill_1 FILLER_71_629 ();
 sg13g2_fill_2 FILLER_71_643 ();
 sg13g2_fill_1 FILLER_71_645 ();
 sg13g2_fill_2 FILLER_71_654 ();
 sg13g2_decap_4 FILLER_71_677 ();
 sg13g2_fill_1 FILLER_71_681 ();
 sg13g2_decap_8 FILLER_71_700 ();
 sg13g2_decap_8 FILLER_71_707 ();
 sg13g2_decap_4 FILLER_71_714 ();
 sg13g2_decap_4 FILLER_71_769 ();
 sg13g2_fill_2 FILLER_71_773 ();
 sg13g2_fill_1 FILLER_71_810 ();
 sg13g2_decap_8 FILLER_71_820 ();
 sg13g2_decap_8 FILLER_71_827 ();
 sg13g2_decap_8 FILLER_71_834 ();
 sg13g2_decap_8 FILLER_71_841 ();
 sg13g2_decap_8 FILLER_71_848 ();
 sg13g2_decap_8 FILLER_71_855 ();
 sg13g2_decap_8 FILLER_71_862 ();
 sg13g2_decap_8 FILLER_71_869 ();
 sg13g2_decap_8 FILLER_71_876 ();
 sg13g2_decap_8 FILLER_71_883 ();
 sg13g2_decap_8 FILLER_71_890 ();
 sg13g2_decap_8 FILLER_71_897 ();
 sg13g2_decap_8 FILLER_71_904 ();
 sg13g2_decap_8 FILLER_71_911 ();
 sg13g2_decap_8 FILLER_71_918 ();
 sg13g2_decap_8 FILLER_71_925 ();
 sg13g2_decap_8 FILLER_71_932 ();
 sg13g2_decap_8 FILLER_71_939 ();
 sg13g2_decap_8 FILLER_71_946 ();
 sg13g2_decap_8 FILLER_71_953 ();
 sg13g2_decap_8 FILLER_71_960 ();
 sg13g2_decap_8 FILLER_71_967 ();
 sg13g2_decap_8 FILLER_71_974 ();
 sg13g2_decap_8 FILLER_71_981 ();
 sg13g2_decap_8 FILLER_71_988 ();
 sg13g2_decap_8 FILLER_71_995 ();
 sg13g2_decap_8 FILLER_71_1002 ();
 sg13g2_decap_8 FILLER_71_1009 ();
 sg13g2_decap_8 FILLER_71_1016 ();
 sg13g2_decap_8 FILLER_71_1023 ();
 sg13g2_decap_8 FILLER_71_1030 ();
 sg13g2_decap_8 FILLER_71_1037 ();
 sg13g2_decap_8 FILLER_71_1044 ();
 sg13g2_decap_8 FILLER_71_1051 ();
 sg13g2_decap_8 FILLER_71_1058 ();
 sg13g2_decap_8 FILLER_71_1065 ();
 sg13g2_decap_8 FILLER_71_1072 ();
 sg13g2_decap_8 FILLER_71_1079 ();
 sg13g2_decap_8 FILLER_71_1086 ();
 sg13g2_decap_8 FILLER_71_1093 ();
 sg13g2_decap_8 FILLER_71_1100 ();
 sg13g2_decap_8 FILLER_71_1107 ();
 sg13g2_decap_8 FILLER_71_1114 ();
 sg13g2_decap_8 FILLER_71_1121 ();
 sg13g2_decap_8 FILLER_71_1128 ();
 sg13g2_decap_8 FILLER_71_1135 ();
 sg13g2_decap_8 FILLER_71_1142 ();
 sg13g2_decap_8 FILLER_71_1149 ();
 sg13g2_decap_8 FILLER_71_1156 ();
 sg13g2_decap_8 FILLER_71_1163 ();
 sg13g2_decap_8 FILLER_71_1170 ();
 sg13g2_decap_8 FILLER_71_1177 ();
 sg13g2_decap_8 FILLER_71_1184 ();
 sg13g2_decap_8 FILLER_71_1191 ();
 sg13g2_decap_8 FILLER_71_1198 ();
 sg13g2_decap_8 FILLER_71_1205 ();
 sg13g2_decap_8 FILLER_71_1212 ();
 sg13g2_decap_8 FILLER_71_1219 ();
 sg13g2_decap_8 FILLER_71_1226 ();
 sg13g2_decap_8 FILLER_71_1233 ();
 sg13g2_decap_8 FILLER_71_1240 ();
 sg13g2_decap_8 FILLER_71_1247 ();
 sg13g2_decap_8 FILLER_71_1254 ();
 sg13g2_decap_8 FILLER_71_1261 ();
 sg13g2_decap_8 FILLER_71_1268 ();
 sg13g2_decap_8 FILLER_71_1275 ();
 sg13g2_decap_8 FILLER_71_1282 ();
 sg13g2_decap_8 FILLER_71_1289 ();
 sg13g2_decap_8 FILLER_71_1296 ();
 sg13g2_decap_8 FILLER_71_1303 ();
 sg13g2_decap_4 FILLER_71_1310 ();
 sg13g2_fill_1 FILLER_71_1314 ();
 sg13g2_fill_2 FILLER_72_83 ();
 sg13g2_fill_1 FILLER_72_114 ();
 sg13g2_fill_2 FILLER_72_135 ();
 sg13g2_fill_1 FILLER_72_137 ();
 sg13g2_fill_2 FILLER_72_169 ();
 sg13g2_fill_2 FILLER_72_179 ();
 sg13g2_fill_2 FILLER_72_186 ();
 sg13g2_fill_1 FILLER_72_197 ();
 sg13g2_fill_1 FILLER_72_233 ();
 sg13g2_fill_2 FILLER_72_255 ();
 sg13g2_fill_1 FILLER_72_257 ();
 sg13g2_fill_2 FILLER_72_275 ();
 sg13g2_fill_1 FILLER_72_326 ();
 sg13g2_fill_1 FILLER_72_340 ();
 sg13g2_fill_2 FILLER_72_375 ();
 sg13g2_fill_2 FILLER_72_463 ();
 sg13g2_fill_1 FILLER_72_465 ();
 sg13g2_fill_2 FILLER_72_472 ();
 sg13g2_fill_1 FILLER_72_474 ();
 sg13g2_fill_2 FILLER_72_518 ();
 sg13g2_fill_1 FILLER_72_557 ();
 sg13g2_fill_2 FILLER_72_603 ();
 sg13g2_fill_1 FILLER_72_605 ();
 sg13g2_fill_1 FILLER_72_623 ();
 sg13g2_fill_2 FILLER_72_650 ();
 sg13g2_decap_8 FILLER_72_661 ();
 sg13g2_decap_4 FILLER_72_668 ();
 sg13g2_fill_2 FILLER_72_672 ();
 sg13g2_decap_4 FILLER_72_687 ();
 sg13g2_fill_1 FILLER_72_714 ();
 sg13g2_decap_8 FILLER_72_745 ();
 sg13g2_fill_1 FILLER_72_752 ();
 sg13g2_fill_2 FILLER_72_766 ();
 sg13g2_decap_4 FILLER_72_777 ();
 sg13g2_fill_1 FILLER_72_790 ();
 sg13g2_fill_2 FILLER_72_812 ();
 sg13g2_decap_8 FILLER_72_827 ();
 sg13g2_decap_8 FILLER_72_834 ();
 sg13g2_decap_8 FILLER_72_841 ();
 sg13g2_decap_8 FILLER_72_848 ();
 sg13g2_decap_8 FILLER_72_855 ();
 sg13g2_decap_8 FILLER_72_862 ();
 sg13g2_decap_8 FILLER_72_869 ();
 sg13g2_decap_8 FILLER_72_876 ();
 sg13g2_decap_8 FILLER_72_883 ();
 sg13g2_decap_8 FILLER_72_890 ();
 sg13g2_decap_8 FILLER_72_897 ();
 sg13g2_decap_8 FILLER_72_904 ();
 sg13g2_decap_8 FILLER_72_911 ();
 sg13g2_decap_8 FILLER_72_918 ();
 sg13g2_decap_8 FILLER_72_925 ();
 sg13g2_decap_8 FILLER_72_932 ();
 sg13g2_decap_8 FILLER_72_939 ();
 sg13g2_decap_8 FILLER_72_946 ();
 sg13g2_decap_8 FILLER_72_953 ();
 sg13g2_decap_8 FILLER_72_960 ();
 sg13g2_decap_8 FILLER_72_967 ();
 sg13g2_decap_8 FILLER_72_974 ();
 sg13g2_decap_8 FILLER_72_981 ();
 sg13g2_decap_8 FILLER_72_988 ();
 sg13g2_decap_8 FILLER_72_995 ();
 sg13g2_decap_8 FILLER_72_1002 ();
 sg13g2_decap_8 FILLER_72_1009 ();
 sg13g2_decap_8 FILLER_72_1016 ();
 sg13g2_decap_8 FILLER_72_1023 ();
 sg13g2_decap_8 FILLER_72_1030 ();
 sg13g2_decap_8 FILLER_72_1037 ();
 sg13g2_decap_8 FILLER_72_1044 ();
 sg13g2_decap_8 FILLER_72_1051 ();
 sg13g2_decap_8 FILLER_72_1058 ();
 sg13g2_decap_8 FILLER_72_1065 ();
 sg13g2_decap_8 FILLER_72_1072 ();
 sg13g2_decap_8 FILLER_72_1079 ();
 sg13g2_decap_8 FILLER_72_1086 ();
 sg13g2_decap_8 FILLER_72_1093 ();
 sg13g2_decap_8 FILLER_72_1100 ();
 sg13g2_decap_8 FILLER_72_1107 ();
 sg13g2_decap_8 FILLER_72_1114 ();
 sg13g2_decap_8 FILLER_72_1121 ();
 sg13g2_decap_8 FILLER_72_1128 ();
 sg13g2_decap_8 FILLER_72_1135 ();
 sg13g2_decap_8 FILLER_72_1142 ();
 sg13g2_decap_8 FILLER_72_1149 ();
 sg13g2_decap_8 FILLER_72_1156 ();
 sg13g2_decap_8 FILLER_72_1163 ();
 sg13g2_decap_8 FILLER_72_1170 ();
 sg13g2_decap_8 FILLER_72_1177 ();
 sg13g2_decap_8 FILLER_72_1184 ();
 sg13g2_decap_8 FILLER_72_1191 ();
 sg13g2_decap_8 FILLER_72_1198 ();
 sg13g2_decap_8 FILLER_72_1205 ();
 sg13g2_decap_8 FILLER_72_1212 ();
 sg13g2_decap_8 FILLER_72_1219 ();
 sg13g2_decap_8 FILLER_72_1226 ();
 sg13g2_decap_8 FILLER_72_1233 ();
 sg13g2_decap_8 FILLER_72_1240 ();
 sg13g2_decap_8 FILLER_72_1247 ();
 sg13g2_decap_8 FILLER_72_1254 ();
 sg13g2_decap_8 FILLER_72_1261 ();
 sg13g2_decap_8 FILLER_72_1268 ();
 sg13g2_decap_8 FILLER_72_1275 ();
 sg13g2_decap_8 FILLER_72_1282 ();
 sg13g2_decap_8 FILLER_72_1289 ();
 sg13g2_decap_8 FILLER_72_1296 ();
 sg13g2_decap_8 FILLER_72_1303 ();
 sg13g2_decap_4 FILLER_72_1310 ();
 sg13g2_fill_1 FILLER_72_1314 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_2 ();
 sg13g2_fill_1 FILLER_73_25 ();
 sg13g2_fill_1 FILLER_73_48 ();
 sg13g2_fill_1 FILLER_73_55 ();
 sg13g2_fill_2 FILLER_73_62 ();
 sg13g2_fill_2 FILLER_73_87 ();
 sg13g2_fill_1 FILLER_73_89 ();
 sg13g2_fill_2 FILLER_73_108 ();
 sg13g2_fill_2 FILLER_73_129 ();
 sg13g2_fill_1 FILLER_73_131 ();
 sg13g2_fill_2 FILLER_73_141 ();
 sg13g2_fill_1 FILLER_73_143 ();
 sg13g2_fill_2 FILLER_73_152 ();
 sg13g2_fill_1 FILLER_73_190 ();
 sg13g2_fill_2 FILLER_73_222 ();
 sg13g2_fill_2 FILLER_73_280 ();
 sg13g2_fill_1 FILLER_73_282 ();
 sg13g2_fill_1 FILLER_73_314 ();
 sg13g2_fill_2 FILLER_73_338 ();
 sg13g2_fill_2 FILLER_73_477 ();
 sg13g2_fill_2 FILLER_73_484 ();
 sg13g2_fill_1 FILLER_73_556 ();
 sg13g2_fill_1 FILLER_73_576 ();
 sg13g2_fill_2 FILLER_73_661 ();
 sg13g2_fill_1 FILLER_73_663 ();
 sg13g2_fill_1 FILLER_73_693 ();
 sg13g2_decap_8 FILLER_73_698 ();
 sg13g2_fill_2 FILLER_73_705 ();
 sg13g2_fill_2 FILLER_73_717 ();
 sg13g2_fill_1 FILLER_73_719 ();
 sg13g2_fill_2 FILLER_73_724 ();
 sg13g2_fill_2 FILLER_73_744 ();
 sg13g2_fill_1 FILLER_73_746 ();
 sg13g2_fill_2 FILLER_73_756 ();
 sg13g2_decap_8 FILLER_73_795 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_8 FILLER_73_857 ();
 sg13g2_decap_8 FILLER_73_864 ();
 sg13g2_decap_8 FILLER_73_871 ();
 sg13g2_decap_8 FILLER_73_878 ();
 sg13g2_decap_8 FILLER_73_885 ();
 sg13g2_decap_8 FILLER_73_892 ();
 sg13g2_decap_8 FILLER_73_899 ();
 sg13g2_decap_8 FILLER_73_906 ();
 sg13g2_decap_8 FILLER_73_913 ();
 sg13g2_decap_8 FILLER_73_920 ();
 sg13g2_decap_8 FILLER_73_927 ();
 sg13g2_decap_8 FILLER_73_934 ();
 sg13g2_decap_8 FILLER_73_941 ();
 sg13g2_decap_8 FILLER_73_948 ();
 sg13g2_decap_8 FILLER_73_955 ();
 sg13g2_decap_8 FILLER_73_962 ();
 sg13g2_decap_8 FILLER_73_969 ();
 sg13g2_decap_8 FILLER_73_976 ();
 sg13g2_decap_8 FILLER_73_983 ();
 sg13g2_decap_8 FILLER_73_990 ();
 sg13g2_decap_8 FILLER_73_997 ();
 sg13g2_decap_8 FILLER_73_1004 ();
 sg13g2_decap_8 FILLER_73_1011 ();
 sg13g2_decap_8 FILLER_73_1018 ();
 sg13g2_decap_8 FILLER_73_1025 ();
 sg13g2_decap_8 FILLER_73_1032 ();
 sg13g2_decap_8 FILLER_73_1039 ();
 sg13g2_decap_8 FILLER_73_1046 ();
 sg13g2_decap_8 FILLER_73_1053 ();
 sg13g2_decap_8 FILLER_73_1060 ();
 sg13g2_decap_8 FILLER_73_1067 ();
 sg13g2_decap_8 FILLER_73_1074 ();
 sg13g2_decap_8 FILLER_73_1081 ();
 sg13g2_decap_8 FILLER_73_1088 ();
 sg13g2_decap_8 FILLER_73_1095 ();
 sg13g2_decap_8 FILLER_73_1102 ();
 sg13g2_decap_8 FILLER_73_1109 ();
 sg13g2_decap_8 FILLER_73_1116 ();
 sg13g2_decap_8 FILLER_73_1123 ();
 sg13g2_decap_8 FILLER_73_1130 ();
 sg13g2_decap_8 FILLER_73_1137 ();
 sg13g2_decap_8 FILLER_73_1144 ();
 sg13g2_decap_8 FILLER_73_1151 ();
 sg13g2_decap_8 FILLER_73_1158 ();
 sg13g2_decap_8 FILLER_73_1165 ();
 sg13g2_decap_8 FILLER_73_1172 ();
 sg13g2_decap_8 FILLER_73_1179 ();
 sg13g2_decap_8 FILLER_73_1186 ();
 sg13g2_decap_8 FILLER_73_1193 ();
 sg13g2_decap_8 FILLER_73_1200 ();
 sg13g2_decap_8 FILLER_73_1207 ();
 sg13g2_decap_8 FILLER_73_1214 ();
 sg13g2_decap_8 FILLER_73_1221 ();
 sg13g2_decap_8 FILLER_73_1228 ();
 sg13g2_decap_8 FILLER_73_1235 ();
 sg13g2_decap_8 FILLER_73_1242 ();
 sg13g2_decap_8 FILLER_73_1249 ();
 sg13g2_decap_8 FILLER_73_1256 ();
 sg13g2_decap_8 FILLER_73_1263 ();
 sg13g2_decap_8 FILLER_73_1270 ();
 sg13g2_decap_8 FILLER_73_1277 ();
 sg13g2_decap_8 FILLER_73_1284 ();
 sg13g2_decap_8 FILLER_73_1291 ();
 sg13g2_decap_8 FILLER_73_1298 ();
 sg13g2_decap_8 FILLER_73_1305 ();
 sg13g2_fill_2 FILLER_73_1312 ();
 sg13g2_fill_1 FILLER_73_1314 ();
 sg13g2_fill_2 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_49 ();
 sg13g2_fill_1 FILLER_74_51 ();
 sg13g2_fill_1 FILLER_74_92 ();
 sg13g2_fill_2 FILLER_74_121 ();
 sg13g2_fill_2 FILLER_74_149 ();
 sg13g2_fill_2 FILLER_74_198 ();
 sg13g2_fill_1 FILLER_74_208 ();
 sg13g2_fill_2 FILLER_74_254 ();
 sg13g2_fill_1 FILLER_74_305 ();
 sg13g2_fill_2 FILLER_74_320 ();
 sg13g2_fill_1 FILLER_74_411 ();
 sg13g2_fill_1 FILLER_74_517 ();
 sg13g2_fill_2 FILLER_74_523 ();
 sg13g2_fill_2 FILLER_74_534 ();
 sg13g2_fill_1 FILLER_74_536 ();
 sg13g2_fill_2 FILLER_74_583 ();
 sg13g2_fill_1 FILLER_74_585 ();
 sg13g2_fill_2 FILLER_74_615 ();
 sg13g2_fill_1 FILLER_74_663 ();
 sg13g2_fill_2 FILLER_74_673 ();
 sg13g2_fill_1 FILLER_74_675 ();
 sg13g2_fill_2 FILLER_74_710 ();
 sg13g2_fill_1 FILLER_74_737 ();
 sg13g2_fill_2 FILLER_74_763 ();
 sg13g2_fill_1 FILLER_74_765 ();
 sg13g2_decap_8 FILLER_74_779 ();
 sg13g2_decap_8 FILLER_74_786 ();
 sg13g2_fill_1 FILLER_74_801 ();
 sg13g2_fill_1 FILLER_74_811 ();
 sg13g2_decap_8 FILLER_74_838 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_decap_8 FILLER_74_852 ();
 sg13g2_decap_8 FILLER_74_859 ();
 sg13g2_decap_8 FILLER_74_866 ();
 sg13g2_decap_8 FILLER_74_873 ();
 sg13g2_decap_8 FILLER_74_880 ();
 sg13g2_decap_8 FILLER_74_887 ();
 sg13g2_decap_8 FILLER_74_894 ();
 sg13g2_decap_8 FILLER_74_901 ();
 sg13g2_decap_8 FILLER_74_908 ();
 sg13g2_decap_8 FILLER_74_915 ();
 sg13g2_decap_8 FILLER_74_922 ();
 sg13g2_decap_8 FILLER_74_929 ();
 sg13g2_decap_8 FILLER_74_936 ();
 sg13g2_decap_8 FILLER_74_943 ();
 sg13g2_decap_8 FILLER_74_950 ();
 sg13g2_decap_8 FILLER_74_957 ();
 sg13g2_decap_8 FILLER_74_964 ();
 sg13g2_decap_8 FILLER_74_971 ();
 sg13g2_decap_8 FILLER_74_978 ();
 sg13g2_decap_8 FILLER_74_985 ();
 sg13g2_decap_8 FILLER_74_992 ();
 sg13g2_decap_8 FILLER_74_999 ();
 sg13g2_decap_8 FILLER_74_1006 ();
 sg13g2_decap_8 FILLER_74_1013 ();
 sg13g2_decap_8 FILLER_74_1020 ();
 sg13g2_decap_8 FILLER_74_1027 ();
 sg13g2_decap_8 FILLER_74_1034 ();
 sg13g2_decap_8 FILLER_74_1041 ();
 sg13g2_decap_8 FILLER_74_1048 ();
 sg13g2_decap_8 FILLER_74_1055 ();
 sg13g2_decap_8 FILLER_74_1062 ();
 sg13g2_decap_8 FILLER_74_1069 ();
 sg13g2_decap_8 FILLER_74_1076 ();
 sg13g2_decap_8 FILLER_74_1083 ();
 sg13g2_decap_8 FILLER_74_1090 ();
 sg13g2_decap_8 FILLER_74_1097 ();
 sg13g2_decap_8 FILLER_74_1104 ();
 sg13g2_decap_8 FILLER_74_1111 ();
 sg13g2_decap_8 FILLER_74_1118 ();
 sg13g2_decap_8 FILLER_74_1125 ();
 sg13g2_decap_8 FILLER_74_1132 ();
 sg13g2_decap_8 FILLER_74_1139 ();
 sg13g2_decap_8 FILLER_74_1146 ();
 sg13g2_decap_8 FILLER_74_1153 ();
 sg13g2_decap_8 FILLER_74_1160 ();
 sg13g2_decap_8 FILLER_74_1167 ();
 sg13g2_decap_8 FILLER_74_1174 ();
 sg13g2_decap_8 FILLER_74_1181 ();
 sg13g2_decap_8 FILLER_74_1188 ();
 sg13g2_decap_8 FILLER_74_1195 ();
 sg13g2_decap_8 FILLER_74_1202 ();
 sg13g2_decap_8 FILLER_74_1209 ();
 sg13g2_decap_8 FILLER_74_1216 ();
 sg13g2_decap_8 FILLER_74_1223 ();
 sg13g2_decap_8 FILLER_74_1230 ();
 sg13g2_decap_8 FILLER_74_1237 ();
 sg13g2_decap_8 FILLER_74_1244 ();
 sg13g2_decap_8 FILLER_74_1251 ();
 sg13g2_decap_8 FILLER_74_1258 ();
 sg13g2_decap_8 FILLER_74_1265 ();
 sg13g2_decap_8 FILLER_74_1272 ();
 sg13g2_decap_8 FILLER_74_1279 ();
 sg13g2_decap_8 FILLER_74_1286 ();
 sg13g2_decap_8 FILLER_74_1293 ();
 sg13g2_decap_8 FILLER_74_1300 ();
 sg13g2_decap_8 FILLER_74_1307 ();
 sg13g2_fill_1 FILLER_74_1314 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_45 ();
 sg13g2_fill_2 FILLER_75_66 ();
 sg13g2_fill_2 FILLER_75_93 ();
 sg13g2_fill_2 FILLER_75_105 ();
 sg13g2_fill_2 FILLER_75_115 ();
 sg13g2_fill_1 FILLER_75_117 ();
 sg13g2_fill_1 FILLER_75_128 ();
 sg13g2_fill_2 FILLER_75_161 ();
 sg13g2_fill_1 FILLER_75_163 ();
 sg13g2_fill_2 FILLER_75_227 ();
 sg13g2_fill_1 FILLER_75_229 ();
 sg13g2_fill_2 FILLER_75_282 ();
 sg13g2_fill_2 FILLER_75_310 ();
 sg13g2_fill_1 FILLER_75_319 ();
 sg13g2_fill_1 FILLER_75_325 ();
 sg13g2_fill_2 FILLER_75_460 ();
 sg13g2_fill_1 FILLER_75_462 ();
 sg13g2_fill_2 FILLER_75_472 ();
 sg13g2_fill_1 FILLER_75_474 ();
 sg13g2_fill_1 FILLER_75_497 ();
 sg13g2_fill_2 FILLER_75_548 ();
 sg13g2_fill_1 FILLER_75_622 ();
 sg13g2_fill_1 FILLER_75_650 ();
 sg13g2_fill_1 FILLER_75_661 ();
 sg13g2_decap_8 FILLER_75_695 ();
 sg13g2_decap_8 FILLER_75_702 ();
 sg13g2_decap_8 FILLER_75_709 ();
 sg13g2_decap_8 FILLER_75_733 ();
 sg13g2_decap_8 FILLER_75_740 ();
 sg13g2_decap_4 FILLER_75_752 ();
 sg13g2_fill_2 FILLER_75_756 ();
 sg13g2_fill_1 FILLER_75_804 ();
 sg13g2_decap_4 FILLER_75_817 ();
 sg13g2_fill_2 FILLER_75_821 ();
 sg13g2_decap_8 FILLER_75_827 ();
 sg13g2_decap_8 FILLER_75_834 ();
 sg13g2_decap_8 FILLER_75_841 ();
 sg13g2_decap_8 FILLER_75_848 ();
 sg13g2_decap_8 FILLER_75_855 ();
 sg13g2_decap_8 FILLER_75_862 ();
 sg13g2_decap_8 FILLER_75_869 ();
 sg13g2_decap_8 FILLER_75_876 ();
 sg13g2_decap_8 FILLER_75_883 ();
 sg13g2_decap_8 FILLER_75_890 ();
 sg13g2_decap_8 FILLER_75_897 ();
 sg13g2_decap_8 FILLER_75_904 ();
 sg13g2_decap_8 FILLER_75_911 ();
 sg13g2_decap_8 FILLER_75_918 ();
 sg13g2_decap_8 FILLER_75_925 ();
 sg13g2_decap_8 FILLER_75_932 ();
 sg13g2_decap_8 FILLER_75_939 ();
 sg13g2_decap_8 FILLER_75_946 ();
 sg13g2_decap_8 FILLER_75_953 ();
 sg13g2_decap_8 FILLER_75_960 ();
 sg13g2_decap_8 FILLER_75_967 ();
 sg13g2_decap_8 FILLER_75_974 ();
 sg13g2_decap_8 FILLER_75_981 ();
 sg13g2_decap_8 FILLER_75_988 ();
 sg13g2_decap_8 FILLER_75_995 ();
 sg13g2_decap_8 FILLER_75_1002 ();
 sg13g2_decap_8 FILLER_75_1009 ();
 sg13g2_decap_8 FILLER_75_1016 ();
 sg13g2_decap_8 FILLER_75_1023 ();
 sg13g2_decap_8 FILLER_75_1030 ();
 sg13g2_decap_8 FILLER_75_1037 ();
 sg13g2_decap_8 FILLER_75_1044 ();
 sg13g2_decap_8 FILLER_75_1051 ();
 sg13g2_decap_8 FILLER_75_1058 ();
 sg13g2_decap_8 FILLER_75_1065 ();
 sg13g2_decap_8 FILLER_75_1072 ();
 sg13g2_decap_8 FILLER_75_1079 ();
 sg13g2_decap_8 FILLER_75_1086 ();
 sg13g2_decap_8 FILLER_75_1093 ();
 sg13g2_decap_8 FILLER_75_1100 ();
 sg13g2_decap_8 FILLER_75_1107 ();
 sg13g2_decap_8 FILLER_75_1114 ();
 sg13g2_decap_8 FILLER_75_1121 ();
 sg13g2_decap_8 FILLER_75_1128 ();
 sg13g2_decap_8 FILLER_75_1135 ();
 sg13g2_decap_8 FILLER_75_1142 ();
 sg13g2_decap_8 FILLER_75_1149 ();
 sg13g2_decap_8 FILLER_75_1156 ();
 sg13g2_decap_8 FILLER_75_1163 ();
 sg13g2_decap_8 FILLER_75_1170 ();
 sg13g2_decap_8 FILLER_75_1177 ();
 sg13g2_decap_8 FILLER_75_1184 ();
 sg13g2_decap_8 FILLER_75_1191 ();
 sg13g2_decap_8 FILLER_75_1198 ();
 sg13g2_decap_8 FILLER_75_1205 ();
 sg13g2_decap_8 FILLER_75_1212 ();
 sg13g2_decap_8 FILLER_75_1219 ();
 sg13g2_decap_8 FILLER_75_1226 ();
 sg13g2_decap_8 FILLER_75_1233 ();
 sg13g2_decap_8 FILLER_75_1240 ();
 sg13g2_decap_8 FILLER_75_1247 ();
 sg13g2_decap_8 FILLER_75_1254 ();
 sg13g2_decap_8 FILLER_75_1261 ();
 sg13g2_decap_8 FILLER_75_1268 ();
 sg13g2_decap_8 FILLER_75_1275 ();
 sg13g2_decap_8 FILLER_75_1282 ();
 sg13g2_decap_8 FILLER_75_1289 ();
 sg13g2_decap_8 FILLER_75_1296 ();
 sg13g2_decap_8 FILLER_75_1303 ();
 sg13g2_decap_4 FILLER_75_1310 ();
 sg13g2_fill_1 FILLER_75_1314 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_2 ();
 sg13g2_fill_2 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_9 ();
 sg13g2_fill_1 FILLER_76_19 ();
 sg13g2_fill_2 FILLER_76_77 ();
 sg13g2_fill_1 FILLER_76_79 ();
 sg13g2_fill_2 FILLER_76_172 ();
 sg13g2_fill_1 FILLER_76_185 ();
 sg13g2_fill_1 FILLER_76_312 ();
 sg13g2_fill_1 FILLER_76_342 ();
 sg13g2_fill_1 FILLER_76_393 ();
 sg13g2_fill_2 FILLER_76_432 ();
 sg13g2_fill_2 FILLER_76_460 ();
 sg13g2_fill_2 FILLER_76_498 ();
 sg13g2_fill_1 FILLER_76_500 ();
 sg13g2_fill_1 FILLER_76_510 ();
 sg13g2_fill_2 FILLER_76_521 ();
 sg13g2_fill_1 FILLER_76_523 ();
 sg13g2_fill_1 FILLER_76_547 ();
 sg13g2_fill_2 FILLER_76_582 ();
 sg13g2_decap_4 FILLER_76_668 ();
 sg13g2_fill_2 FILLER_76_708 ();
 sg13g2_fill_1 FILLER_76_710 ();
 sg13g2_decap_8 FILLER_76_720 ();
 sg13g2_fill_1 FILLER_76_738 ();
 sg13g2_fill_2 FILLER_76_759 ();
 sg13g2_fill_2 FILLER_76_787 ();
 sg13g2_fill_1 FILLER_76_789 ();
 sg13g2_decap_8 FILLER_76_803 ();
 sg13g2_decap_4 FILLER_76_810 ();
 sg13g2_fill_2 FILLER_76_814 ();
 sg13g2_decap_8 FILLER_76_819 ();
 sg13g2_decap_8 FILLER_76_826 ();
 sg13g2_decap_8 FILLER_76_833 ();
 sg13g2_decap_8 FILLER_76_840 ();
 sg13g2_decap_8 FILLER_76_847 ();
 sg13g2_decap_8 FILLER_76_854 ();
 sg13g2_decap_8 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_76_868 ();
 sg13g2_decap_8 FILLER_76_875 ();
 sg13g2_decap_8 FILLER_76_882 ();
 sg13g2_decap_8 FILLER_76_889 ();
 sg13g2_decap_8 FILLER_76_896 ();
 sg13g2_decap_8 FILLER_76_903 ();
 sg13g2_decap_8 FILLER_76_910 ();
 sg13g2_decap_8 FILLER_76_917 ();
 sg13g2_decap_8 FILLER_76_924 ();
 sg13g2_decap_8 FILLER_76_931 ();
 sg13g2_decap_8 FILLER_76_938 ();
 sg13g2_decap_8 FILLER_76_945 ();
 sg13g2_decap_8 FILLER_76_952 ();
 sg13g2_decap_8 FILLER_76_959 ();
 sg13g2_decap_8 FILLER_76_966 ();
 sg13g2_decap_8 FILLER_76_973 ();
 sg13g2_decap_8 FILLER_76_980 ();
 sg13g2_decap_8 FILLER_76_987 ();
 sg13g2_decap_8 FILLER_76_994 ();
 sg13g2_decap_8 FILLER_76_1001 ();
 sg13g2_decap_8 FILLER_76_1008 ();
 sg13g2_decap_8 FILLER_76_1015 ();
 sg13g2_decap_8 FILLER_76_1022 ();
 sg13g2_decap_8 FILLER_76_1029 ();
 sg13g2_decap_8 FILLER_76_1036 ();
 sg13g2_decap_8 FILLER_76_1043 ();
 sg13g2_decap_8 FILLER_76_1050 ();
 sg13g2_decap_8 FILLER_76_1057 ();
 sg13g2_decap_8 FILLER_76_1064 ();
 sg13g2_decap_8 FILLER_76_1071 ();
 sg13g2_decap_8 FILLER_76_1078 ();
 sg13g2_decap_8 FILLER_76_1085 ();
 sg13g2_decap_8 FILLER_76_1092 ();
 sg13g2_decap_8 FILLER_76_1099 ();
 sg13g2_decap_8 FILLER_76_1106 ();
 sg13g2_decap_8 FILLER_76_1113 ();
 sg13g2_decap_8 FILLER_76_1120 ();
 sg13g2_decap_8 FILLER_76_1127 ();
 sg13g2_decap_8 FILLER_76_1134 ();
 sg13g2_decap_8 FILLER_76_1141 ();
 sg13g2_decap_8 FILLER_76_1148 ();
 sg13g2_decap_8 FILLER_76_1155 ();
 sg13g2_decap_8 FILLER_76_1162 ();
 sg13g2_decap_8 FILLER_76_1169 ();
 sg13g2_decap_8 FILLER_76_1176 ();
 sg13g2_decap_8 FILLER_76_1183 ();
 sg13g2_decap_8 FILLER_76_1190 ();
 sg13g2_decap_8 FILLER_76_1197 ();
 sg13g2_decap_8 FILLER_76_1204 ();
 sg13g2_decap_8 FILLER_76_1211 ();
 sg13g2_decap_8 FILLER_76_1218 ();
 sg13g2_decap_8 FILLER_76_1225 ();
 sg13g2_decap_8 FILLER_76_1232 ();
 sg13g2_decap_8 FILLER_76_1239 ();
 sg13g2_decap_8 FILLER_76_1246 ();
 sg13g2_decap_8 FILLER_76_1253 ();
 sg13g2_decap_8 FILLER_76_1260 ();
 sg13g2_decap_8 FILLER_76_1267 ();
 sg13g2_decap_8 FILLER_76_1274 ();
 sg13g2_decap_8 FILLER_76_1281 ();
 sg13g2_decap_8 FILLER_76_1288 ();
 sg13g2_decap_8 FILLER_76_1295 ();
 sg13g2_decap_8 FILLER_76_1302 ();
 sg13g2_decap_4 FILLER_76_1309 ();
 sg13g2_fill_2 FILLER_76_1313 ();
 sg13g2_fill_2 FILLER_77_90 ();
 sg13g2_fill_1 FILLER_77_136 ();
 sg13g2_fill_2 FILLER_77_145 ();
 sg13g2_fill_1 FILLER_77_156 ();
 sg13g2_fill_2 FILLER_77_163 ();
 sg13g2_fill_1 FILLER_77_165 ();
 sg13g2_fill_2 FILLER_77_220 ();
 sg13g2_fill_1 FILLER_77_222 ();
 sg13g2_fill_2 FILLER_77_231 ();
 sg13g2_fill_1 FILLER_77_252 ();
 sg13g2_fill_2 FILLER_77_347 ();
 sg13g2_fill_1 FILLER_77_400 ();
 sg13g2_fill_2 FILLER_77_442 ();
 sg13g2_fill_2 FILLER_77_448 ();
 sg13g2_fill_1 FILLER_77_476 ();
 sg13g2_fill_2 FILLER_77_525 ();
 sg13g2_fill_1 FILLER_77_527 ();
 sg13g2_fill_2 FILLER_77_562 ();
 sg13g2_fill_1 FILLER_77_590 ();
 sg13g2_fill_2 FILLER_77_617 ();
 sg13g2_fill_1 FILLER_77_619 ();
 sg13g2_fill_1 FILLER_77_642 ();
 sg13g2_decap_8 FILLER_77_679 ();
 sg13g2_fill_2 FILLER_77_686 ();
 sg13g2_decap_4 FILLER_77_701 ();
 sg13g2_fill_1 FILLER_77_722 ();
 sg13g2_decap_4 FILLER_77_744 ();
 sg13g2_fill_1 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_757 ();
 sg13g2_decap_4 FILLER_77_768 ();
 sg13g2_fill_1 FILLER_77_772 ();
 sg13g2_decap_4 FILLER_77_781 ();
 sg13g2_fill_1 FILLER_77_785 ();
 sg13g2_decap_8 FILLER_77_824 ();
 sg13g2_decap_8 FILLER_77_831 ();
 sg13g2_decap_8 FILLER_77_838 ();
 sg13g2_decap_8 FILLER_77_845 ();
 sg13g2_decap_8 FILLER_77_852 ();
 sg13g2_decap_8 FILLER_77_859 ();
 sg13g2_decap_8 FILLER_77_866 ();
 sg13g2_decap_8 FILLER_77_873 ();
 sg13g2_decap_8 FILLER_77_880 ();
 sg13g2_decap_8 FILLER_77_887 ();
 sg13g2_decap_8 FILLER_77_894 ();
 sg13g2_decap_8 FILLER_77_901 ();
 sg13g2_decap_8 FILLER_77_908 ();
 sg13g2_decap_8 FILLER_77_915 ();
 sg13g2_decap_8 FILLER_77_922 ();
 sg13g2_decap_8 FILLER_77_929 ();
 sg13g2_decap_8 FILLER_77_936 ();
 sg13g2_decap_8 FILLER_77_943 ();
 sg13g2_decap_8 FILLER_77_950 ();
 sg13g2_decap_8 FILLER_77_957 ();
 sg13g2_decap_8 FILLER_77_964 ();
 sg13g2_decap_8 FILLER_77_971 ();
 sg13g2_decap_8 FILLER_77_978 ();
 sg13g2_decap_8 FILLER_77_985 ();
 sg13g2_decap_8 FILLER_77_992 ();
 sg13g2_decap_8 FILLER_77_999 ();
 sg13g2_decap_8 FILLER_77_1006 ();
 sg13g2_decap_8 FILLER_77_1013 ();
 sg13g2_decap_8 FILLER_77_1020 ();
 sg13g2_decap_8 FILLER_77_1027 ();
 sg13g2_decap_8 FILLER_77_1034 ();
 sg13g2_decap_8 FILLER_77_1041 ();
 sg13g2_decap_8 FILLER_77_1048 ();
 sg13g2_decap_8 FILLER_77_1055 ();
 sg13g2_decap_8 FILLER_77_1062 ();
 sg13g2_decap_8 FILLER_77_1069 ();
 sg13g2_decap_8 FILLER_77_1076 ();
 sg13g2_decap_8 FILLER_77_1083 ();
 sg13g2_decap_8 FILLER_77_1090 ();
 sg13g2_decap_8 FILLER_77_1097 ();
 sg13g2_decap_8 FILLER_77_1104 ();
 sg13g2_decap_8 FILLER_77_1111 ();
 sg13g2_decap_8 FILLER_77_1118 ();
 sg13g2_decap_8 FILLER_77_1125 ();
 sg13g2_decap_8 FILLER_77_1132 ();
 sg13g2_decap_8 FILLER_77_1139 ();
 sg13g2_decap_8 FILLER_77_1146 ();
 sg13g2_decap_8 FILLER_77_1153 ();
 sg13g2_decap_8 FILLER_77_1160 ();
 sg13g2_decap_8 FILLER_77_1167 ();
 sg13g2_decap_8 FILLER_77_1174 ();
 sg13g2_decap_8 FILLER_77_1181 ();
 sg13g2_decap_8 FILLER_77_1188 ();
 sg13g2_decap_8 FILLER_77_1195 ();
 sg13g2_decap_8 FILLER_77_1202 ();
 sg13g2_decap_8 FILLER_77_1209 ();
 sg13g2_decap_8 FILLER_77_1216 ();
 sg13g2_decap_8 FILLER_77_1223 ();
 sg13g2_decap_8 FILLER_77_1230 ();
 sg13g2_decap_8 FILLER_77_1237 ();
 sg13g2_decap_8 FILLER_77_1244 ();
 sg13g2_decap_8 FILLER_77_1251 ();
 sg13g2_decap_8 FILLER_77_1258 ();
 sg13g2_decap_8 FILLER_77_1265 ();
 sg13g2_decap_8 FILLER_77_1272 ();
 sg13g2_decap_8 FILLER_77_1279 ();
 sg13g2_decap_8 FILLER_77_1286 ();
 sg13g2_decap_8 FILLER_77_1293 ();
 sg13g2_decap_8 FILLER_77_1300 ();
 sg13g2_decap_8 FILLER_77_1307 ();
 sg13g2_fill_1 FILLER_77_1314 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_23 ();
 sg13g2_fill_1 FILLER_78_25 ();
 sg13g2_fill_2 FILLER_78_66 ();
 sg13g2_fill_1 FILLER_78_68 ();
 sg13g2_fill_1 FILLER_78_78 ();
 sg13g2_fill_1 FILLER_78_158 ();
 sg13g2_fill_2 FILLER_78_168 ();
 sg13g2_fill_1 FILLER_78_170 ();
 sg13g2_fill_1 FILLER_78_180 ();
 sg13g2_fill_2 FILLER_78_232 ();
 sg13g2_fill_1 FILLER_78_234 ();
 sg13g2_fill_2 FILLER_78_334 ();
 sg13g2_fill_1 FILLER_78_379 ();
 sg13g2_fill_1 FILLER_78_433 ();
 sg13g2_fill_1 FILLER_78_442 ();
 sg13g2_fill_1 FILLER_78_455 ();
 sg13g2_fill_1 FILLER_78_470 ();
 sg13g2_fill_2 FILLER_78_505 ();
 sg13g2_fill_1 FILLER_78_507 ();
 sg13g2_fill_2 FILLER_78_518 ();
 sg13g2_fill_2 FILLER_78_581 ();
 sg13g2_fill_1 FILLER_78_587 ();
 sg13g2_fill_1 FILLER_78_607 ();
 sg13g2_fill_2 FILLER_78_617 ();
 sg13g2_decap_4 FILLER_78_704 ();
 sg13g2_fill_1 FILLER_78_708 ();
 sg13g2_fill_1 FILLER_78_728 ();
 sg13g2_decap_4 FILLER_78_744 ();
 sg13g2_decap_4 FILLER_78_760 ();
 sg13g2_fill_1 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_779 ();
 sg13g2_decap_8 FILLER_78_786 ();
 sg13g2_fill_1 FILLER_78_793 ();
 sg13g2_decap_8 FILLER_78_799 ();
 sg13g2_fill_2 FILLER_78_806 ();
 sg13g2_fill_1 FILLER_78_808 ();
 sg13g2_decap_8 FILLER_78_813 ();
 sg13g2_decap_8 FILLER_78_820 ();
 sg13g2_decap_8 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_834 ();
 sg13g2_decap_8 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_848 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_decap_8 FILLER_78_862 ();
 sg13g2_decap_8 FILLER_78_869 ();
 sg13g2_decap_8 FILLER_78_876 ();
 sg13g2_decap_8 FILLER_78_883 ();
 sg13g2_decap_8 FILLER_78_890 ();
 sg13g2_decap_8 FILLER_78_897 ();
 sg13g2_decap_8 FILLER_78_904 ();
 sg13g2_decap_8 FILLER_78_911 ();
 sg13g2_decap_8 FILLER_78_918 ();
 sg13g2_decap_8 FILLER_78_925 ();
 sg13g2_decap_8 FILLER_78_932 ();
 sg13g2_decap_8 FILLER_78_939 ();
 sg13g2_decap_8 FILLER_78_946 ();
 sg13g2_decap_8 FILLER_78_953 ();
 sg13g2_decap_8 FILLER_78_960 ();
 sg13g2_decap_8 FILLER_78_967 ();
 sg13g2_decap_8 FILLER_78_974 ();
 sg13g2_decap_8 FILLER_78_981 ();
 sg13g2_decap_8 FILLER_78_988 ();
 sg13g2_decap_8 FILLER_78_995 ();
 sg13g2_decap_8 FILLER_78_1002 ();
 sg13g2_decap_8 FILLER_78_1009 ();
 sg13g2_decap_8 FILLER_78_1016 ();
 sg13g2_decap_8 FILLER_78_1023 ();
 sg13g2_decap_8 FILLER_78_1030 ();
 sg13g2_decap_8 FILLER_78_1037 ();
 sg13g2_decap_8 FILLER_78_1044 ();
 sg13g2_decap_8 FILLER_78_1051 ();
 sg13g2_decap_8 FILLER_78_1058 ();
 sg13g2_decap_8 FILLER_78_1065 ();
 sg13g2_decap_8 FILLER_78_1072 ();
 sg13g2_decap_8 FILLER_78_1079 ();
 sg13g2_decap_8 FILLER_78_1086 ();
 sg13g2_decap_8 FILLER_78_1093 ();
 sg13g2_decap_8 FILLER_78_1100 ();
 sg13g2_decap_8 FILLER_78_1107 ();
 sg13g2_decap_8 FILLER_78_1114 ();
 sg13g2_decap_8 FILLER_78_1121 ();
 sg13g2_decap_8 FILLER_78_1128 ();
 sg13g2_decap_8 FILLER_78_1135 ();
 sg13g2_decap_8 FILLER_78_1142 ();
 sg13g2_decap_8 FILLER_78_1149 ();
 sg13g2_decap_8 FILLER_78_1156 ();
 sg13g2_decap_8 FILLER_78_1163 ();
 sg13g2_decap_8 FILLER_78_1170 ();
 sg13g2_decap_8 FILLER_78_1177 ();
 sg13g2_decap_8 FILLER_78_1184 ();
 sg13g2_decap_8 FILLER_78_1191 ();
 sg13g2_decap_8 FILLER_78_1198 ();
 sg13g2_decap_8 FILLER_78_1205 ();
 sg13g2_decap_8 FILLER_78_1212 ();
 sg13g2_decap_8 FILLER_78_1219 ();
 sg13g2_decap_8 FILLER_78_1226 ();
 sg13g2_decap_8 FILLER_78_1233 ();
 sg13g2_decap_8 FILLER_78_1240 ();
 sg13g2_decap_8 FILLER_78_1247 ();
 sg13g2_decap_8 FILLER_78_1254 ();
 sg13g2_decap_8 FILLER_78_1261 ();
 sg13g2_decap_8 FILLER_78_1268 ();
 sg13g2_decap_8 FILLER_78_1275 ();
 sg13g2_decap_8 FILLER_78_1282 ();
 sg13g2_decap_8 FILLER_78_1289 ();
 sg13g2_decap_8 FILLER_78_1296 ();
 sg13g2_decap_8 FILLER_78_1303 ();
 sg13g2_decap_4 FILLER_78_1310 ();
 sg13g2_fill_1 FILLER_78_1314 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_2 FILLER_79_15 ();
 sg13g2_fill_1 FILLER_79_17 ();
 sg13g2_decap_8 FILLER_79_22 ();
 sg13g2_fill_1 FILLER_79_29 ();
 sg13g2_decap_8 FILLER_79_34 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_4 FILLER_79_56 ();
 sg13g2_decap_4 FILLER_79_68 ();
 sg13g2_fill_2 FILLER_79_72 ();
 sg13g2_fill_2 FILLER_79_86 ();
 sg13g2_fill_1 FILLER_79_88 ();
 sg13g2_fill_1 FILLER_79_94 ();
 sg13g2_fill_2 FILLER_79_103 ();
 sg13g2_fill_2 FILLER_79_114 ();
 sg13g2_fill_2 FILLER_79_125 ();
 sg13g2_fill_1 FILLER_79_127 ();
 sg13g2_fill_2 FILLER_79_136 ();
 sg13g2_fill_1 FILLER_79_138 ();
 sg13g2_fill_1 FILLER_79_147 ();
 sg13g2_fill_1 FILLER_79_152 ();
 sg13g2_fill_1 FILLER_79_179 ();
 sg13g2_fill_2 FILLER_79_189 ();
 sg13g2_fill_2 FILLER_79_217 ();
 sg13g2_fill_1 FILLER_79_219 ();
 sg13g2_fill_1 FILLER_79_229 ();
 sg13g2_fill_1 FILLER_79_244 ();
 sg13g2_fill_2 FILLER_79_258 ();
 sg13g2_fill_2 FILLER_79_340 ();
 sg13g2_fill_2 FILLER_79_356 ();
 sg13g2_fill_1 FILLER_79_404 ();
 sg13g2_decap_8 FILLER_79_453 ();
 sg13g2_fill_1 FILLER_79_460 ();
 sg13g2_decap_4 FILLER_79_465 ();
 sg13g2_decap_4 FILLER_79_473 ();
 sg13g2_fill_2 FILLER_79_477 ();
 sg13g2_fill_2 FILLER_79_522 ();
 sg13g2_fill_1 FILLER_79_524 ();
 sg13g2_fill_2 FILLER_79_559 ();
 sg13g2_fill_1 FILLER_79_561 ();
 sg13g2_fill_1 FILLER_79_571 ();
 sg13g2_fill_1 FILLER_79_657 ();
 sg13g2_fill_2 FILLER_79_676 ();
 sg13g2_decap_8 FILLER_79_695 ();
 sg13g2_decap_8 FILLER_79_702 ();
 sg13g2_fill_1 FILLER_79_709 ();
 sg13g2_fill_2 FILLER_79_727 ();
 sg13g2_fill_1 FILLER_79_732 ();
 sg13g2_fill_1 FILLER_79_740 ();
 sg13g2_fill_2 FILLER_79_760 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_decap_8 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_827 ();
 sg13g2_decap_8 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_decap_8 FILLER_79_862 ();
 sg13g2_decap_8 FILLER_79_869 ();
 sg13g2_decap_8 FILLER_79_876 ();
 sg13g2_decap_8 FILLER_79_883 ();
 sg13g2_decap_8 FILLER_79_890 ();
 sg13g2_decap_8 FILLER_79_897 ();
 sg13g2_decap_8 FILLER_79_904 ();
 sg13g2_decap_8 FILLER_79_911 ();
 sg13g2_decap_8 FILLER_79_918 ();
 sg13g2_decap_8 FILLER_79_925 ();
 sg13g2_decap_8 FILLER_79_932 ();
 sg13g2_decap_8 FILLER_79_939 ();
 sg13g2_decap_8 FILLER_79_946 ();
 sg13g2_decap_8 FILLER_79_953 ();
 sg13g2_decap_8 FILLER_79_960 ();
 sg13g2_decap_8 FILLER_79_967 ();
 sg13g2_decap_8 FILLER_79_974 ();
 sg13g2_decap_8 FILLER_79_981 ();
 sg13g2_decap_8 FILLER_79_988 ();
 sg13g2_decap_8 FILLER_79_995 ();
 sg13g2_decap_8 FILLER_79_1002 ();
 sg13g2_decap_8 FILLER_79_1009 ();
 sg13g2_decap_8 FILLER_79_1016 ();
 sg13g2_decap_8 FILLER_79_1023 ();
 sg13g2_decap_8 FILLER_79_1030 ();
 sg13g2_decap_8 FILLER_79_1037 ();
 sg13g2_decap_8 FILLER_79_1044 ();
 sg13g2_decap_8 FILLER_79_1051 ();
 sg13g2_decap_8 FILLER_79_1058 ();
 sg13g2_decap_8 FILLER_79_1065 ();
 sg13g2_decap_8 FILLER_79_1072 ();
 sg13g2_decap_8 FILLER_79_1079 ();
 sg13g2_decap_8 FILLER_79_1086 ();
 sg13g2_decap_8 FILLER_79_1093 ();
 sg13g2_decap_8 FILLER_79_1100 ();
 sg13g2_decap_8 FILLER_79_1107 ();
 sg13g2_decap_8 FILLER_79_1114 ();
 sg13g2_decap_8 FILLER_79_1121 ();
 sg13g2_decap_8 FILLER_79_1128 ();
 sg13g2_decap_8 FILLER_79_1135 ();
 sg13g2_decap_8 FILLER_79_1142 ();
 sg13g2_decap_8 FILLER_79_1149 ();
 sg13g2_decap_8 FILLER_79_1156 ();
 sg13g2_decap_8 FILLER_79_1163 ();
 sg13g2_decap_8 FILLER_79_1170 ();
 sg13g2_decap_8 FILLER_79_1177 ();
 sg13g2_decap_8 FILLER_79_1184 ();
 sg13g2_decap_8 FILLER_79_1191 ();
 sg13g2_decap_8 FILLER_79_1198 ();
 sg13g2_decap_8 FILLER_79_1205 ();
 sg13g2_decap_8 FILLER_79_1212 ();
 sg13g2_decap_8 FILLER_79_1219 ();
 sg13g2_decap_8 FILLER_79_1226 ();
 sg13g2_decap_8 FILLER_79_1233 ();
 sg13g2_decap_8 FILLER_79_1240 ();
 sg13g2_decap_8 FILLER_79_1247 ();
 sg13g2_decap_8 FILLER_79_1254 ();
 sg13g2_decap_8 FILLER_79_1261 ();
 sg13g2_decap_8 FILLER_79_1268 ();
 sg13g2_decap_8 FILLER_79_1275 ();
 sg13g2_decap_8 FILLER_79_1282 ();
 sg13g2_decap_8 FILLER_79_1289 ();
 sg13g2_decap_8 FILLER_79_1296 ();
 sg13g2_decap_8 FILLER_79_1303 ();
 sg13g2_decap_4 FILLER_79_1310 ();
 sg13g2_fill_1 FILLER_79_1314 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_4 FILLER_80_77 ();
 sg13g2_fill_1 FILLER_80_81 ();
 sg13g2_decap_8 FILLER_80_133 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_fill_1 FILLER_80_144 ();
 sg13g2_fill_2 FILLER_80_174 ();
 sg13g2_fill_2 FILLER_80_199 ();
 sg13g2_fill_1 FILLER_80_244 ();
 sg13g2_fill_1 FILLER_80_275 ();
 sg13g2_fill_2 FILLER_80_386 ();
 sg13g2_fill_1 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_454 ();
 sg13g2_decap_8 FILLER_80_461 ();
 sg13g2_decap_8 FILLER_80_468 ();
 sg13g2_decap_8 FILLER_80_475 ();
 sg13g2_fill_2 FILLER_80_482 ();
 sg13g2_fill_1 FILLER_80_520 ();
 sg13g2_fill_2 FILLER_80_561 ();
 sg13g2_fill_2 FILLER_80_586 ();
 sg13g2_fill_1 FILLER_80_588 ();
 sg13g2_fill_2 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_624 ();
 sg13g2_fill_1 FILLER_80_631 ();
 sg13g2_fill_2 FILLER_80_666 ();
 sg13g2_fill_1 FILLER_80_668 ();
 sg13g2_decap_4 FILLER_80_695 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_fill_2 FILLER_80_739 ();
 sg13g2_fill_1 FILLER_80_741 ();
 sg13g2_decap_8 FILLER_80_768 ();
 sg13g2_decap_4 FILLER_80_775 ();
 sg13g2_fill_1 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_833 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_decap_8 FILLER_80_861 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_decap_8 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_889 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_decap_8 FILLER_80_903 ();
 sg13g2_decap_8 FILLER_80_910 ();
 sg13g2_decap_8 FILLER_80_917 ();
 sg13g2_decap_8 FILLER_80_924 ();
 sg13g2_decap_8 FILLER_80_931 ();
 sg13g2_decap_8 FILLER_80_938 ();
 sg13g2_decap_8 FILLER_80_945 ();
 sg13g2_decap_8 FILLER_80_952 ();
 sg13g2_decap_8 FILLER_80_959 ();
 sg13g2_decap_8 FILLER_80_966 ();
 sg13g2_decap_8 FILLER_80_973 ();
 sg13g2_decap_8 FILLER_80_980 ();
 sg13g2_decap_8 FILLER_80_987 ();
 sg13g2_decap_8 FILLER_80_994 ();
 sg13g2_decap_8 FILLER_80_1001 ();
 sg13g2_decap_8 FILLER_80_1008 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_decap_8 FILLER_80_1022 ();
 sg13g2_decap_8 FILLER_80_1029 ();
 sg13g2_decap_8 FILLER_80_1036 ();
 sg13g2_decap_8 FILLER_80_1043 ();
 sg13g2_decap_8 FILLER_80_1050 ();
 sg13g2_decap_8 FILLER_80_1057 ();
 sg13g2_decap_8 FILLER_80_1064 ();
 sg13g2_decap_8 FILLER_80_1071 ();
 sg13g2_decap_8 FILLER_80_1078 ();
 sg13g2_decap_8 FILLER_80_1085 ();
 sg13g2_decap_8 FILLER_80_1092 ();
 sg13g2_decap_8 FILLER_80_1099 ();
 sg13g2_decap_8 FILLER_80_1106 ();
 sg13g2_decap_8 FILLER_80_1113 ();
 sg13g2_decap_8 FILLER_80_1120 ();
 sg13g2_decap_8 FILLER_80_1127 ();
 sg13g2_decap_8 FILLER_80_1134 ();
 sg13g2_decap_8 FILLER_80_1141 ();
 sg13g2_decap_8 FILLER_80_1148 ();
 sg13g2_decap_8 FILLER_80_1155 ();
 sg13g2_decap_8 FILLER_80_1162 ();
 sg13g2_decap_8 FILLER_80_1169 ();
 sg13g2_decap_8 FILLER_80_1176 ();
 sg13g2_decap_8 FILLER_80_1183 ();
 sg13g2_decap_8 FILLER_80_1190 ();
 sg13g2_decap_8 FILLER_80_1197 ();
 sg13g2_decap_8 FILLER_80_1204 ();
 sg13g2_decap_8 FILLER_80_1211 ();
 sg13g2_decap_8 FILLER_80_1218 ();
 sg13g2_decap_8 FILLER_80_1225 ();
 sg13g2_decap_8 FILLER_80_1232 ();
 sg13g2_decap_8 FILLER_80_1239 ();
 sg13g2_decap_8 FILLER_80_1246 ();
 sg13g2_decap_8 FILLER_80_1253 ();
 sg13g2_decap_8 FILLER_80_1260 ();
 sg13g2_decap_8 FILLER_80_1267 ();
 sg13g2_decap_8 FILLER_80_1274 ();
 sg13g2_decap_8 FILLER_80_1281 ();
 sg13g2_decap_8 FILLER_80_1288 ();
 sg13g2_decap_8 FILLER_80_1295 ();
 sg13g2_decap_8 FILLER_80_1302 ();
 sg13g2_decap_4 FILLER_80_1309 ();
 sg13g2_fill_2 FILLER_80_1313 ();
endmodule
